**************************************************
* OpenRAM generated memory.
* Words: 64
* Data bits: 256
* Banks: 1
* Column mux: 1:1
**************************************************
* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
*
.subckt dff D Q clk vdd gnd
*
MM21 Q a_66_6# gnd gnd NMOS_VTG L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd NMOS_VTG L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd PMOS_VTG L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd PMOS_VTG L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd PMOS_VTG L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd PMOS_VTG L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.SUBCKT row_addr_dff din_0 din_1 din_2 din_3 din_4 din_5 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 6 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r1_c0 din_1 dout_1 clk vdd gnd dff
Xdff_r2_c0 din_2 dout_2 clk vdd gnd dff
Xdff_r3_c0 din_3 dout_3 clk vdd gnd dff
Xdff_r4_c0 din_4 dout_4 clk vdd gnd dff
Xdff_r5_c0 din_5 dout_5 clk vdd gnd dff
.ENDS row_addr_dff

.SUBCKT data_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 din_128 din_129 din_130 din_131 din_132 din_133 din_134 din_135 din_136 din_137 din_138 din_139 din_140 din_141 din_142 din_143 din_144 din_145 din_146 din_147 din_148 din_149 din_150 din_151 din_152 din_153 din_154 din_155 din_156 din_157 din_158 din_159 din_160 din_161 din_162 din_163 din_164 din_165 din_166 din_167 din_168 din_169 din_170 din_171 din_172 din_173 din_174 din_175 din_176 din_177 din_178 din_179 din_180 din_181 din_182 din_183 din_184 din_185 din_186 din_187 din_188 din_189 din_190 din_191 din_192 din_193 din_194 din_195 din_196 din_197 din_198 din_199 din_200 din_201 din_202 din_203 din_204 din_205 din_206 din_207 din_208 din_209 din_210 din_211 din_212 din_213 din_214 din_215 din_216 din_217 din_218 din_219 din_220 din_221 din_222 din_223 din_224 din_225 din_226 din_227 din_228 din_229 din_230 din_231 din_232 din_233 din_234 din_235 din_236 din_237 din_238 din_239 din_240 din_241 din_242 din_243 din_244 din_245 din_246 din_247 din_248 din_249 din_250 din_251 din_252 din_253 din_254 din_255 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38 dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46 dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54 dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62 dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70 dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78 dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86 dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94 dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102 dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109 dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116 dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123 dout_124 dout_125 dout_126 dout_127 dout_128 dout_129 dout_130 dout_131 dout_132 dout_133 dout_134 dout_135 dout_136 dout_137 dout_138 dout_139 dout_140 dout_141 dout_142 dout_143 dout_144 dout_145 dout_146 dout_147 dout_148 dout_149 dout_150 dout_151 dout_152 dout_153 dout_154 dout_155 dout_156 dout_157 dout_158 dout_159 dout_160 dout_161 dout_162 dout_163 dout_164 dout_165 dout_166 dout_167 dout_168 dout_169 dout_170 dout_171 dout_172 dout_173 dout_174 dout_175 dout_176 dout_177 dout_178 dout_179 dout_180 dout_181 dout_182 dout_183 dout_184 dout_185 dout_186 dout_187 dout_188 dout_189 dout_190 dout_191 dout_192 dout_193 dout_194 dout_195 dout_196 dout_197 dout_198 dout_199 dout_200 dout_201 dout_202 dout_203 dout_204 dout_205 dout_206 dout_207 dout_208 dout_209 dout_210 dout_211 dout_212 dout_213 dout_214 dout_215 dout_216 dout_217 dout_218 dout_219 dout_220 dout_221 dout_222 dout_223 dout_224 dout_225 dout_226 dout_227 dout_228 dout_229 dout_230 dout_231 dout_232 dout_233 dout_234 dout_235 dout_236 dout_237 dout_238 dout_239 dout_240 dout_241 dout_242 dout_243 dout_244 dout_245 dout_246 dout_247 dout_248 dout_249 dout_250 dout_251 dout_252 dout_253 dout_254 dout_255 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* INPUT : din_128 
* INPUT : din_129 
* INPUT : din_130 
* INPUT : din_131 
* INPUT : din_132 
* INPUT : din_133 
* INPUT : din_134 
* INPUT : din_135 
* INPUT : din_136 
* INPUT : din_137 
* INPUT : din_138 
* INPUT : din_139 
* INPUT : din_140 
* INPUT : din_141 
* INPUT : din_142 
* INPUT : din_143 
* INPUT : din_144 
* INPUT : din_145 
* INPUT : din_146 
* INPUT : din_147 
* INPUT : din_148 
* INPUT : din_149 
* INPUT : din_150 
* INPUT : din_151 
* INPUT : din_152 
* INPUT : din_153 
* INPUT : din_154 
* INPUT : din_155 
* INPUT : din_156 
* INPUT : din_157 
* INPUT : din_158 
* INPUT : din_159 
* INPUT : din_160 
* INPUT : din_161 
* INPUT : din_162 
* INPUT : din_163 
* INPUT : din_164 
* INPUT : din_165 
* INPUT : din_166 
* INPUT : din_167 
* INPUT : din_168 
* INPUT : din_169 
* INPUT : din_170 
* INPUT : din_171 
* INPUT : din_172 
* INPUT : din_173 
* INPUT : din_174 
* INPUT : din_175 
* INPUT : din_176 
* INPUT : din_177 
* INPUT : din_178 
* INPUT : din_179 
* INPUT : din_180 
* INPUT : din_181 
* INPUT : din_182 
* INPUT : din_183 
* INPUT : din_184 
* INPUT : din_185 
* INPUT : din_186 
* INPUT : din_187 
* INPUT : din_188 
* INPUT : din_189 
* INPUT : din_190 
* INPUT : din_191 
* INPUT : din_192 
* INPUT : din_193 
* INPUT : din_194 
* INPUT : din_195 
* INPUT : din_196 
* INPUT : din_197 
* INPUT : din_198 
* INPUT : din_199 
* INPUT : din_200 
* INPUT : din_201 
* INPUT : din_202 
* INPUT : din_203 
* INPUT : din_204 
* INPUT : din_205 
* INPUT : din_206 
* INPUT : din_207 
* INPUT : din_208 
* INPUT : din_209 
* INPUT : din_210 
* INPUT : din_211 
* INPUT : din_212 
* INPUT : din_213 
* INPUT : din_214 
* INPUT : din_215 
* INPUT : din_216 
* INPUT : din_217 
* INPUT : din_218 
* INPUT : din_219 
* INPUT : din_220 
* INPUT : din_221 
* INPUT : din_222 
* INPUT : din_223 
* INPUT : din_224 
* INPUT : din_225 
* INPUT : din_226 
* INPUT : din_227 
* INPUT : din_228 
* INPUT : din_229 
* INPUT : din_230 
* INPUT : din_231 
* INPUT : din_232 
* INPUT : din_233 
* INPUT : din_234 
* INPUT : din_235 
* INPUT : din_236 
* INPUT : din_237 
* INPUT : din_238 
* INPUT : din_239 
* INPUT : din_240 
* INPUT : din_241 
* INPUT : din_242 
* INPUT : din_243 
* INPUT : din_244 
* INPUT : din_245 
* INPUT : din_246 
* INPUT : din_247 
* INPUT : din_248 
* INPUT : din_249 
* INPUT : din_250 
* INPUT : din_251 
* INPUT : din_252 
* INPUT : din_253 
* INPUT : din_254 
* INPUT : din_255 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* OUTPUT: dout_128 
* OUTPUT: dout_129 
* OUTPUT: dout_130 
* OUTPUT: dout_131 
* OUTPUT: dout_132 
* OUTPUT: dout_133 
* OUTPUT: dout_134 
* OUTPUT: dout_135 
* OUTPUT: dout_136 
* OUTPUT: dout_137 
* OUTPUT: dout_138 
* OUTPUT: dout_139 
* OUTPUT: dout_140 
* OUTPUT: dout_141 
* OUTPUT: dout_142 
* OUTPUT: dout_143 
* OUTPUT: dout_144 
* OUTPUT: dout_145 
* OUTPUT: dout_146 
* OUTPUT: dout_147 
* OUTPUT: dout_148 
* OUTPUT: dout_149 
* OUTPUT: dout_150 
* OUTPUT: dout_151 
* OUTPUT: dout_152 
* OUTPUT: dout_153 
* OUTPUT: dout_154 
* OUTPUT: dout_155 
* OUTPUT: dout_156 
* OUTPUT: dout_157 
* OUTPUT: dout_158 
* OUTPUT: dout_159 
* OUTPUT: dout_160 
* OUTPUT: dout_161 
* OUTPUT: dout_162 
* OUTPUT: dout_163 
* OUTPUT: dout_164 
* OUTPUT: dout_165 
* OUTPUT: dout_166 
* OUTPUT: dout_167 
* OUTPUT: dout_168 
* OUTPUT: dout_169 
* OUTPUT: dout_170 
* OUTPUT: dout_171 
* OUTPUT: dout_172 
* OUTPUT: dout_173 
* OUTPUT: dout_174 
* OUTPUT: dout_175 
* OUTPUT: dout_176 
* OUTPUT: dout_177 
* OUTPUT: dout_178 
* OUTPUT: dout_179 
* OUTPUT: dout_180 
* OUTPUT: dout_181 
* OUTPUT: dout_182 
* OUTPUT: dout_183 
* OUTPUT: dout_184 
* OUTPUT: dout_185 
* OUTPUT: dout_186 
* OUTPUT: dout_187 
* OUTPUT: dout_188 
* OUTPUT: dout_189 
* OUTPUT: dout_190 
* OUTPUT: dout_191 
* OUTPUT: dout_192 
* OUTPUT: dout_193 
* OUTPUT: dout_194 
* OUTPUT: dout_195 
* OUTPUT: dout_196 
* OUTPUT: dout_197 
* OUTPUT: dout_198 
* OUTPUT: dout_199 
* OUTPUT: dout_200 
* OUTPUT: dout_201 
* OUTPUT: dout_202 
* OUTPUT: dout_203 
* OUTPUT: dout_204 
* OUTPUT: dout_205 
* OUTPUT: dout_206 
* OUTPUT: dout_207 
* OUTPUT: dout_208 
* OUTPUT: dout_209 
* OUTPUT: dout_210 
* OUTPUT: dout_211 
* OUTPUT: dout_212 
* OUTPUT: dout_213 
* OUTPUT: dout_214 
* OUTPUT: dout_215 
* OUTPUT: dout_216 
* OUTPUT: dout_217 
* OUTPUT: dout_218 
* OUTPUT: dout_219 
* OUTPUT: dout_220 
* OUTPUT: dout_221 
* OUTPUT: dout_222 
* OUTPUT: dout_223 
* OUTPUT: dout_224 
* OUTPUT: dout_225 
* OUTPUT: dout_226 
* OUTPUT: dout_227 
* OUTPUT: dout_228 
* OUTPUT: dout_229 
* OUTPUT: dout_230 
* OUTPUT: dout_231 
* OUTPUT: dout_232 
* OUTPUT: dout_233 
* OUTPUT: dout_234 
* OUTPUT: dout_235 
* OUTPUT: dout_236 
* OUTPUT: dout_237 
* OUTPUT: dout_238 
* OUTPUT: dout_239 
* OUTPUT: dout_240 
* OUTPUT: dout_241 
* OUTPUT: dout_242 
* OUTPUT: dout_243 
* OUTPUT: dout_244 
* OUTPUT: dout_245 
* OUTPUT: dout_246 
* OUTPUT: dout_247 
* OUTPUT: dout_248 
* OUTPUT: dout_249 
* OUTPUT: dout_250 
* OUTPUT: dout_251 
* OUTPUT: dout_252 
* OUTPUT: dout_253 
* OUTPUT: dout_254 
* OUTPUT: dout_255 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 256
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
Xdff_r0_c3 din_3 dout_3 clk vdd gnd dff
Xdff_r0_c4 din_4 dout_4 clk vdd gnd dff
Xdff_r0_c5 din_5 dout_5 clk vdd gnd dff
Xdff_r0_c6 din_6 dout_6 clk vdd gnd dff
Xdff_r0_c7 din_7 dout_7 clk vdd gnd dff
Xdff_r0_c8 din_8 dout_8 clk vdd gnd dff
Xdff_r0_c9 din_9 dout_9 clk vdd gnd dff
Xdff_r0_c10 din_10 dout_10 clk vdd gnd dff
Xdff_r0_c11 din_11 dout_11 clk vdd gnd dff
Xdff_r0_c12 din_12 dout_12 clk vdd gnd dff
Xdff_r0_c13 din_13 dout_13 clk vdd gnd dff
Xdff_r0_c14 din_14 dout_14 clk vdd gnd dff
Xdff_r0_c15 din_15 dout_15 clk vdd gnd dff
Xdff_r0_c16 din_16 dout_16 clk vdd gnd dff
Xdff_r0_c17 din_17 dout_17 clk vdd gnd dff
Xdff_r0_c18 din_18 dout_18 clk vdd gnd dff
Xdff_r0_c19 din_19 dout_19 clk vdd gnd dff
Xdff_r0_c20 din_20 dout_20 clk vdd gnd dff
Xdff_r0_c21 din_21 dout_21 clk vdd gnd dff
Xdff_r0_c22 din_22 dout_22 clk vdd gnd dff
Xdff_r0_c23 din_23 dout_23 clk vdd gnd dff
Xdff_r0_c24 din_24 dout_24 clk vdd gnd dff
Xdff_r0_c25 din_25 dout_25 clk vdd gnd dff
Xdff_r0_c26 din_26 dout_26 clk vdd gnd dff
Xdff_r0_c27 din_27 dout_27 clk vdd gnd dff
Xdff_r0_c28 din_28 dout_28 clk vdd gnd dff
Xdff_r0_c29 din_29 dout_29 clk vdd gnd dff
Xdff_r0_c30 din_30 dout_30 clk vdd gnd dff
Xdff_r0_c31 din_31 dout_31 clk vdd gnd dff
Xdff_r0_c32 din_32 dout_32 clk vdd gnd dff
Xdff_r0_c33 din_33 dout_33 clk vdd gnd dff
Xdff_r0_c34 din_34 dout_34 clk vdd gnd dff
Xdff_r0_c35 din_35 dout_35 clk vdd gnd dff
Xdff_r0_c36 din_36 dout_36 clk vdd gnd dff
Xdff_r0_c37 din_37 dout_37 clk vdd gnd dff
Xdff_r0_c38 din_38 dout_38 clk vdd gnd dff
Xdff_r0_c39 din_39 dout_39 clk vdd gnd dff
Xdff_r0_c40 din_40 dout_40 clk vdd gnd dff
Xdff_r0_c41 din_41 dout_41 clk vdd gnd dff
Xdff_r0_c42 din_42 dout_42 clk vdd gnd dff
Xdff_r0_c43 din_43 dout_43 clk vdd gnd dff
Xdff_r0_c44 din_44 dout_44 clk vdd gnd dff
Xdff_r0_c45 din_45 dout_45 clk vdd gnd dff
Xdff_r0_c46 din_46 dout_46 clk vdd gnd dff
Xdff_r0_c47 din_47 dout_47 clk vdd gnd dff
Xdff_r0_c48 din_48 dout_48 clk vdd gnd dff
Xdff_r0_c49 din_49 dout_49 clk vdd gnd dff
Xdff_r0_c50 din_50 dout_50 clk vdd gnd dff
Xdff_r0_c51 din_51 dout_51 clk vdd gnd dff
Xdff_r0_c52 din_52 dout_52 clk vdd gnd dff
Xdff_r0_c53 din_53 dout_53 clk vdd gnd dff
Xdff_r0_c54 din_54 dout_54 clk vdd gnd dff
Xdff_r0_c55 din_55 dout_55 clk vdd gnd dff
Xdff_r0_c56 din_56 dout_56 clk vdd gnd dff
Xdff_r0_c57 din_57 dout_57 clk vdd gnd dff
Xdff_r0_c58 din_58 dout_58 clk vdd gnd dff
Xdff_r0_c59 din_59 dout_59 clk vdd gnd dff
Xdff_r0_c60 din_60 dout_60 clk vdd gnd dff
Xdff_r0_c61 din_61 dout_61 clk vdd gnd dff
Xdff_r0_c62 din_62 dout_62 clk vdd gnd dff
Xdff_r0_c63 din_63 dout_63 clk vdd gnd dff
Xdff_r0_c64 din_64 dout_64 clk vdd gnd dff
Xdff_r0_c65 din_65 dout_65 clk vdd gnd dff
Xdff_r0_c66 din_66 dout_66 clk vdd gnd dff
Xdff_r0_c67 din_67 dout_67 clk vdd gnd dff
Xdff_r0_c68 din_68 dout_68 clk vdd gnd dff
Xdff_r0_c69 din_69 dout_69 clk vdd gnd dff
Xdff_r0_c70 din_70 dout_70 clk vdd gnd dff
Xdff_r0_c71 din_71 dout_71 clk vdd gnd dff
Xdff_r0_c72 din_72 dout_72 clk vdd gnd dff
Xdff_r0_c73 din_73 dout_73 clk vdd gnd dff
Xdff_r0_c74 din_74 dout_74 clk vdd gnd dff
Xdff_r0_c75 din_75 dout_75 clk vdd gnd dff
Xdff_r0_c76 din_76 dout_76 clk vdd gnd dff
Xdff_r0_c77 din_77 dout_77 clk vdd gnd dff
Xdff_r0_c78 din_78 dout_78 clk vdd gnd dff
Xdff_r0_c79 din_79 dout_79 clk vdd gnd dff
Xdff_r0_c80 din_80 dout_80 clk vdd gnd dff
Xdff_r0_c81 din_81 dout_81 clk vdd gnd dff
Xdff_r0_c82 din_82 dout_82 clk vdd gnd dff
Xdff_r0_c83 din_83 dout_83 clk vdd gnd dff
Xdff_r0_c84 din_84 dout_84 clk vdd gnd dff
Xdff_r0_c85 din_85 dout_85 clk vdd gnd dff
Xdff_r0_c86 din_86 dout_86 clk vdd gnd dff
Xdff_r0_c87 din_87 dout_87 clk vdd gnd dff
Xdff_r0_c88 din_88 dout_88 clk vdd gnd dff
Xdff_r0_c89 din_89 dout_89 clk vdd gnd dff
Xdff_r0_c90 din_90 dout_90 clk vdd gnd dff
Xdff_r0_c91 din_91 dout_91 clk vdd gnd dff
Xdff_r0_c92 din_92 dout_92 clk vdd gnd dff
Xdff_r0_c93 din_93 dout_93 clk vdd gnd dff
Xdff_r0_c94 din_94 dout_94 clk vdd gnd dff
Xdff_r0_c95 din_95 dout_95 clk vdd gnd dff
Xdff_r0_c96 din_96 dout_96 clk vdd gnd dff
Xdff_r0_c97 din_97 dout_97 clk vdd gnd dff
Xdff_r0_c98 din_98 dout_98 clk vdd gnd dff
Xdff_r0_c99 din_99 dout_99 clk vdd gnd dff
Xdff_r0_c100 din_100 dout_100 clk vdd gnd dff
Xdff_r0_c101 din_101 dout_101 clk vdd gnd dff
Xdff_r0_c102 din_102 dout_102 clk vdd gnd dff
Xdff_r0_c103 din_103 dout_103 clk vdd gnd dff
Xdff_r0_c104 din_104 dout_104 clk vdd gnd dff
Xdff_r0_c105 din_105 dout_105 clk vdd gnd dff
Xdff_r0_c106 din_106 dout_106 clk vdd gnd dff
Xdff_r0_c107 din_107 dout_107 clk vdd gnd dff
Xdff_r0_c108 din_108 dout_108 clk vdd gnd dff
Xdff_r0_c109 din_109 dout_109 clk vdd gnd dff
Xdff_r0_c110 din_110 dout_110 clk vdd gnd dff
Xdff_r0_c111 din_111 dout_111 clk vdd gnd dff
Xdff_r0_c112 din_112 dout_112 clk vdd gnd dff
Xdff_r0_c113 din_113 dout_113 clk vdd gnd dff
Xdff_r0_c114 din_114 dout_114 clk vdd gnd dff
Xdff_r0_c115 din_115 dout_115 clk vdd gnd dff
Xdff_r0_c116 din_116 dout_116 clk vdd gnd dff
Xdff_r0_c117 din_117 dout_117 clk vdd gnd dff
Xdff_r0_c118 din_118 dout_118 clk vdd gnd dff
Xdff_r0_c119 din_119 dout_119 clk vdd gnd dff
Xdff_r0_c120 din_120 dout_120 clk vdd gnd dff
Xdff_r0_c121 din_121 dout_121 clk vdd gnd dff
Xdff_r0_c122 din_122 dout_122 clk vdd gnd dff
Xdff_r0_c123 din_123 dout_123 clk vdd gnd dff
Xdff_r0_c124 din_124 dout_124 clk vdd gnd dff
Xdff_r0_c125 din_125 dout_125 clk vdd gnd dff
Xdff_r0_c126 din_126 dout_126 clk vdd gnd dff
Xdff_r0_c127 din_127 dout_127 clk vdd gnd dff
Xdff_r0_c128 din_128 dout_128 clk vdd gnd dff
Xdff_r0_c129 din_129 dout_129 clk vdd gnd dff
Xdff_r0_c130 din_130 dout_130 clk vdd gnd dff
Xdff_r0_c131 din_131 dout_131 clk vdd gnd dff
Xdff_r0_c132 din_132 dout_132 clk vdd gnd dff
Xdff_r0_c133 din_133 dout_133 clk vdd gnd dff
Xdff_r0_c134 din_134 dout_134 clk vdd gnd dff
Xdff_r0_c135 din_135 dout_135 clk vdd gnd dff
Xdff_r0_c136 din_136 dout_136 clk vdd gnd dff
Xdff_r0_c137 din_137 dout_137 clk vdd gnd dff
Xdff_r0_c138 din_138 dout_138 clk vdd gnd dff
Xdff_r0_c139 din_139 dout_139 clk vdd gnd dff
Xdff_r0_c140 din_140 dout_140 clk vdd gnd dff
Xdff_r0_c141 din_141 dout_141 clk vdd gnd dff
Xdff_r0_c142 din_142 dout_142 clk vdd gnd dff
Xdff_r0_c143 din_143 dout_143 clk vdd gnd dff
Xdff_r0_c144 din_144 dout_144 clk vdd gnd dff
Xdff_r0_c145 din_145 dout_145 clk vdd gnd dff
Xdff_r0_c146 din_146 dout_146 clk vdd gnd dff
Xdff_r0_c147 din_147 dout_147 clk vdd gnd dff
Xdff_r0_c148 din_148 dout_148 clk vdd gnd dff
Xdff_r0_c149 din_149 dout_149 clk vdd gnd dff
Xdff_r0_c150 din_150 dout_150 clk vdd gnd dff
Xdff_r0_c151 din_151 dout_151 clk vdd gnd dff
Xdff_r0_c152 din_152 dout_152 clk vdd gnd dff
Xdff_r0_c153 din_153 dout_153 clk vdd gnd dff
Xdff_r0_c154 din_154 dout_154 clk vdd gnd dff
Xdff_r0_c155 din_155 dout_155 clk vdd gnd dff
Xdff_r0_c156 din_156 dout_156 clk vdd gnd dff
Xdff_r0_c157 din_157 dout_157 clk vdd gnd dff
Xdff_r0_c158 din_158 dout_158 clk vdd gnd dff
Xdff_r0_c159 din_159 dout_159 clk vdd gnd dff
Xdff_r0_c160 din_160 dout_160 clk vdd gnd dff
Xdff_r0_c161 din_161 dout_161 clk vdd gnd dff
Xdff_r0_c162 din_162 dout_162 clk vdd gnd dff
Xdff_r0_c163 din_163 dout_163 clk vdd gnd dff
Xdff_r0_c164 din_164 dout_164 clk vdd gnd dff
Xdff_r0_c165 din_165 dout_165 clk vdd gnd dff
Xdff_r0_c166 din_166 dout_166 clk vdd gnd dff
Xdff_r0_c167 din_167 dout_167 clk vdd gnd dff
Xdff_r0_c168 din_168 dout_168 clk vdd gnd dff
Xdff_r0_c169 din_169 dout_169 clk vdd gnd dff
Xdff_r0_c170 din_170 dout_170 clk vdd gnd dff
Xdff_r0_c171 din_171 dout_171 clk vdd gnd dff
Xdff_r0_c172 din_172 dout_172 clk vdd gnd dff
Xdff_r0_c173 din_173 dout_173 clk vdd gnd dff
Xdff_r0_c174 din_174 dout_174 clk vdd gnd dff
Xdff_r0_c175 din_175 dout_175 clk vdd gnd dff
Xdff_r0_c176 din_176 dout_176 clk vdd gnd dff
Xdff_r0_c177 din_177 dout_177 clk vdd gnd dff
Xdff_r0_c178 din_178 dout_178 clk vdd gnd dff
Xdff_r0_c179 din_179 dout_179 clk vdd gnd dff
Xdff_r0_c180 din_180 dout_180 clk vdd gnd dff
Xdff_r0_c181 din_181 dout_181 clk vdd gnd dff
Xdff_r0_c182 din_182 dout_182 clk vdd gnd dff
Xdff_r0_c183 din_183 dout_183 clk vdd gnd dff
Xdff_r0_c184 din_184 dout_184 clk vdd gnd dff
Xdff_r0_c185 din_185 dout_185 clk vdd gnd dff
Xdff_r0_c186 din_186 dout_186 clk vdd gnd dff
Xdff_r0_c187 din_187 dout_187 clk vdd gnd dff
Xdff_r0_c188 din_188 dout_188 clk vdd gnd dff
Xdff_r0_c189 din_189 dout_189 clk vdd gnd dff
Xdff_r0_c190 din_190 dout_190 clk vdd gnd dff
Xdff_r0_c191 din_191 dout_191 clk vdd gnd dff
Xdff_r0_c192 din_192 dout_192 clk vdd gnd dff
Xdff_r0_c193 din_193 dout_193 clk vdd gnd dff
Xdff_r0_c194 din_194 dout_194 clk vdd gnd dff
Xdff_r0_c195 din_195 dout_195 clk vdd gnd dff
Xdff_r0_c196 din_196 dout_196 clk vdd gnd dff
Xdff_r0_c197 din_197 dout_197 clk vdd gnd dff
Xdff_r0_c198 din_198 dout_198 clk vdd gnd dff
Xdff_r0_c199 din_199 dout_199 clk vdd gnd dff
Xdff_r0_c200 din_200 dout_200 clk vdd gnd dff
Xdff_r0_c201 din_201 dout_201 clk vdd gnd dff
Xdff_r0_c202 din_202 dout_202 clk vdd gnd dff
Xdff_r0_c203 din_203 dout_203 clk vdd gnd dff
Xdff_r0_c204 din_204 dout_204 clk vdd gnd dff
Xdff_r0_c205 din_205 dout_205 clk vdd gnd dff
Xdff_r0_c206 din_206 dout_206 clk vdd gnd dff
Xdff_r0_c207 din_207 dout_207 clk vdd gnd dff
Xdff_r0_c208 din_208 dout_208 clk vdd gnd dff
Xdff_r0_c209 din_209 dout_209 clk vdd gnd dff
Xdff_r0_c210 din_210 dout_210 clk vdd gnd dff
Xdff_r0_c211 din_211 dout_211 clk vdd gnd dff
Xdff_r0_c212 din_212 dout_212 clk vdd gnd dff
Xdff_r0_c213 din_213 dout_213 clk vdd gnd dff
Xdff_r0_c214 din_214 dout_214 clk vdd gnd dff
Xdff_r0_c215 din_215 dout_215 clk vdd gnd dff
Xdff_r0_c216 din_216 dout_216 clk vdd gnd dff
Xdff_r0_c217 din_217 dout_217 clk vdd gnd dff
Xdff_r0_c218 din_218 dout_218 clk vdd gnd dff
Xdff_r0_c219 din_219 dout_219 clk vdd gnd dff
Xdff_r0_c220 din_220 dout_220 clk vdd gnd dff
Xdff_r0_c221 din_221 dout_221 clk vdd gnd dff
Xdff_r0_c222 din_222 dout_222 clk vdd gnd dff
Xdff_r0_c223 din_223 dout_223 clk vdd gnd dff
Xdff_r0_c224 din_224 dout_224 clk vdd gnd dff
Xdff_r0_c225 din_225 dout_225 clk vdd gnd dff
Xdff_r0_c226 din_226 dout_226 clk vdd gnd dff
Xdff_r0_c227 din_227 dout_227 clk vdd gnd dff
Xdff_r0_c228 din_228 dout_228 clk vdd gnd dff
Xdff_r0_c229 din_229 dout_229 clk vdd gnd dff
Xdff_r0_c230 din_230 dout_230 clk vdd gnd dff
Xdff_r0_c231 din_231 dout_231 clk vdd gnd dff
Xdff_r0_c232 din_232 dout_232 clk vdd gnd dff
Xdff_r0_c233 din_233 dout_233 clk vdd gnd dff
Xdff_r0_c234 din_234 dout_234 clk vdd gnd dff
Xdff_r0_c235 din_235 dout_235 clk vdd gnd dff
Xdff_r0_c236 din_236 dout_236 clk vdd gnd dff
Xdff_r0_c237 din_237 dout_237 clk vdd gnd dff
Xdff_r0_c238 din_238 dout_238 clk vdd gnd dff
Xdff_r0_c239 din_239 dout_239 clk vdd gnd dff
Xdff_r0_c240 din_240 dout_240 clk vdd gnd dff
Xdff_r0_c241 din_241 dout_241 clk vdd gnd dff
Xdff_r0_c242 din_242 dout_242 clk vdd gnd dff
Xdff_r0_c243 din_243 dout_243 clk vdd gnd dff
Xdff_r0_c244 din_244 dout_244 clk vdd gnd dff
Xdff_r0_c245 din_245 dout_245 clk vdd gnd dff
Xdff_r0_c246 din_246 dout_246 clk vdd gnd dff
Xdff_r0_c247 din_247 dout_247 clk vdd gnd dff
Xdff_r0_c248 din_248 dout_248 clk vdd gnd dff
Xdff_r0_c249 din_249 dout_249 clk vdd gnd dff
Xdff_r0_c250 din_250 dout_250 clk vdd gnd dff
Xdff_r0_c251 din_251 dout_251 clk vdd gnd dff
Xdff_r0_c252 din_252 dout_252 clk vdd gnd dff
Xdff_r0_c253 din_253 dout_253 clk vdd gnd dff
Xdff_r0_c254 din_254 dout_254 clk vdd gnd dff
Xdff_r0_c255 din_255 dout_255 clk vdd gnd dff
.ENDS data_dff

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT precharge_1 bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos1 bl en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos2 br en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS precharge_1

.SUBCKT precharge_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 bl_256 br_256 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* INPUT : en_bar 
* POWER : vdd 
* cols: 257 size: 1 bl: bl br: br
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_1
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_1
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_1
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_1
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_1
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_1
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_1
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_1
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_1
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_1
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_1
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_1
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_1
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_1
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_1
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_1
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_1
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_1
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_1
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_1
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_1
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_1
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_1
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_1
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_1
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_1
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_1
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_1
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_1
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_1
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_1
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_1
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_1
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_1
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_1
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_1
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_1
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_1
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_1
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_1
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_1
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_1
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_1
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_1
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_1
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_1
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_1
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_1
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_1
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_1
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_1
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_1
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_1
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_1
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_1
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_1
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_1
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_1
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_1
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_1
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_1
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_1
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_1
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_1
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_1
Xpre_column_65 bl_65 br_65 en_bar vdd precharge_1
Xpre_column_66 bl_66 br_66 en_bar vdd precharge_1
Xpre_column_67 bl_67 br_67 en_bar vdd precharge_1
Xpre_column_68 bl_68 br_68 en_bar vdd precharge_1
Xpre_column_69 bl_69 br_69 en_bar vdd precharge_1
Xpre_column_70 bl_70 br_70 en_bar vdd precharge_1
Xpre_column_71 bl_71 br_71 en_bar vdd precharge_1
Xpre_column_72 bl_72 br_72 en_bar vdd precharge_1
Xpre_column_73 bl_73 br_73 en_bar vdd precharge_1
Xpre_column_74 bl_74 br_74 en_bar vdd precharge_1
Xpre_column_75 bl_75 br_75 en_bar vdd precharge_1
Xpre_column_76 bl_76 br_76 en_bar vdd precharge_1
Xpre_column_77 bl_77 br_77 en_bar vdd precharge_1
Xpre_column_78 bl_78 br_78 en_bar vdd precharge_1
Xpre_column_79 bl_79 br_79 en_bar vdd precharge_1
Xpre_column_80 bl_80 br_80 en_bar vdd precharge_1
Xpre_column_81 bl_81 br_81 en_bar vdd precharge_1
Xpre_column_82 bl_82 br_82 en_bar vdd precharge_1
Xpre_column_83 bl_83 br_83 en_bar vdd precharge_1
Xpre_column_84 bl_84 br_84 en_bar vdd precharge_1
Xpre_column_85 bl_85 br_85 en_bar vdd precharge_1
Xpre_column_86 bl_86 br_86 en_bar vdd precharge_1
Xpre_column_87 bl_87 br_87 en_bar vdd precharge_1
Xpre_column_88 bl_88 br_88 en_bar vdd precharge_1
Xpre_column_89 bl_89 br_89 en_bar vdd precharge_1
Xpre_column_90 bl_90 br_90 en_bar vdd precharge_1
Xpre_column_91 bl_91 br_91 en_bar vdd precharge_1
Xpre_column_92 bl_92 br_92 en_bar vdd precharge_1
Xpre_column_93 bl_93 br_93 en_bar vdd precharge_1
Xpre_column_94 bl_94 br_94 en_bar vdd precharge_1
Xpre_column_95 bl_95 br_95 en_bar vdd precharge_1
Xpre_column_96 bl_96 br_96 en_bar vdd precharge_1
Xpre_column_97 bl_97 br_97 en_bar vdd precharge_1
Xpre_column_98 bl_98 br_98 en_bar vdd precharge_1
Xpre_column_99 bl_99 br_99 en_bar vdd precharge_1
Xpre_column_100 bl_100 br_100 en_bar vdd precharge_1
Xpre_column_101 bl_101 br_101 en_bar vdd precharge_1
Xpre_column_102 bl_102 br_102 en_bar vdd precharge_1
Xpre_column_103 bl_103 br_103 en_bar vdd precharge_1
Xpre_column_104 bl_104 br_104 en_bar vdd precharge_1
Xpre_column_105 bl_105 br_105 en_bar vdd precharge_1
Xpre_column_106 bl_106 br_106 en_bar vdd precharge_1
Xpre_column_107 bl_107 br_107 en_bar vdd precharge_1
Xpre_column_108 bl_108 br_108 en_bar vdd precharge_1
Xpre_column_109 bl_109 br_109 en_bar vdd precharge_1
Xpre_column_110 bl_110 br_110 en_bar vdd precharge_1
Xpre_column_111 bl_111 br_111 en_bar vdd precharge_1
Xpre_column_112 bl_112 br_112 en_bar vdd precharge_1
Xpre_column_113 bl_113 br_113 en_bar vdd precharge_1
Xpre_column_114 bl_114 br_114 en_bar vdd precharge_1
Xpre_column_115 bl_115 br_115 en_bar vdd precharge_1
Xpre_column_116 bl_116 br_116 en_bar vdd precharge_1
Xpre_column_117 bl_117 br_117 en_bar vdd precharge_1
Xpre_column_118 bl_118 br_118 en_bar vdd precharge_1
Xpre_column_119 bl_119 br_119 en_bar vdd precharge_1
Xpre_column_120 bl_120 br_120 en_bar vdd precharge_1
Xpre_column_121 bl_121 br_121 en_bar vdd precharge_1
Xpre_column_122 bl_122 br_122 en_bar vdd precharge_1
Xpre_column_123 bl_123 br_123 en_bar vdd precharge_1
Xpre_column_124 bl_124 br_124 en_bar vdd precharge_1
Xpre_column_125 bl_125 br_125 en_bar vdd precharge_1
Xpre_column_126 bl_126 br_126 en_bar vdd precharge_1
Xpre_column_127 bl_127 br_127 en_bar vdd precharge_1
Xpre_column_128 bl_128 br_128 en_bar vdd precharge_1
Xpre_column_129 bl_129 br_129 en_bar vdd precharge_1
Xpre_column_130 bl_130 br_130 en_bar vdd precharge_1
Xpre_column_131 bl_131 br_131 en_bar vdd precharge_1
Xpre_column_132 bl_132 br_132 en_bar vdd precharge_1
Xpre_column_133 bl_133 br_133 en_bar vdd precharge_1
Xpre_column_134 bl_134 br_134 en_bar vdd precharge_1
Xpre_column_135 bl_135 br_135 en_bar vdd precharge_1
Xpre_column_136 bl_136 br_136 en_bar vdd precharge_1
Xpre_column_137 bl_137 br_137 en_bar vdd precharge_1
Xpre_column_138 bl_138 br_138 en_bar vdd precharge_1
Xpre_column_139 bl_139 br_139 en_bar vdd precharge_1
Xpre_column_140 bl_140 br_140 en_bar vdd precharge_1
Xpre_column_141 bl_141 br_141 en_bar vdd precharge_1
Xpre_column_142 bl_142 br_142 en_bar vdd precharge_1
Xpre_column_143 bl_143 br_143 en_bar vdd precharge_1
Xpre_column_144 bl_144 br_144 en_bar vdd precharge_1
Xpre_column_145 bl_145 br_145 en_bar vdd precharge_1
Xpre_column_146 bl_146 br_146 en_bar vdd precharge_1
Xpre_column_147 bl_147 br_147 en_bar vdd precharge_1
Xpre_column_148 bl_148 br_148 en_bar vdd precharge_1
Xpre_column_149 bl_149 br_149 en_bar vdd precharge_1
Xpre_column_150 bl_150 br_150 en_bar vdd precharge_1
Xpre_column_151 bl_151 br_151 en_bar vdd precharge_1
Xpre_column_152 bl_152 br_152 en_bar vdd precharge_1
Xpre_column_153 bl_153 br_153 en_bar vdd precharge_1
Xpre_column_154 bl_154 br_154 en_bar vdd precharge_1
Xpre_column_155 bl_155 br_155 en_bar vdd precharge_1
Xpre_column_156 bl_156 br_156 en_bar vdd precharge_1
Xpre_column_157 bl_157 br_157 en_bar vdd precharge_1
Xpre_column_158 bl_158 br_158 en_bar vdd precharge_1
Xpre_column_159 bl_159 br_159 en_bar vdd precharge_1
Xpre_column_160 bl_160 br_160 en_bar vdd precharge_1
Xpre_column_161 bl_161 br_161 en_bar vdd precharge_1
Xpre_column_162 bl_162 br_162 en_bar vdd precharge_1
Xpre_column_163 bl_163 br_163 en_bar vdd precharge_1
Xpre_column_164 bl_164 br_164 en_bar vdd precharge_1
Xpre_column_165 bl_165 br_165 en_bar vdd precharge_1
Xpre_column_166 bl_166 br_166 en_bar vdd precharge_1
Xpre_column_167 bl_167 br_167 en_bar vdd precharge_1
Xpre_column_168 bl_168 br_168 en_bar vdd precharge_1
Xpre_column_169 bl_169 br_169 en_bar vdd precharge_1
Xpre_column_170 bl_170 br_170 en_bar vdd precharge_1
Xpre_column_171 bl_171 br_171 en_bar vdd precharge_1
Xpre_column_172 bl_172 br_172 en_bar vdd precharge_1
Xpre_column_173 bl_173 br_173 en_bar vdd precharge_1
Xpre_column_174 bl_174 br_174 en_bar vdd precharge_1
Xpre_column_175 bl_175 br_175 en_bar vdd precharge_1
Xpre_column_176 bl_176 br_176 en_bar vdd precharge_1
Xpre_column_177 bl_177 br_177 en_bar vdd precharge_1
Xpre_column_178 bl_178 br_178 en_bar vdd precharge_1
Xpre_column_179 bl_179 br_179 en_bar vdd precharge_1
Xpre_column_180 bl_180 br_180 en_bar vdd precharge_1
Xpre_column_181 bl_181 br_181 en_bar vdd precharge_1
Xpre_column_182 bl_182 br_182 en_bar vdd precharge_1
Xpre_column_183 bl_183 br_183 en_bar vdd precharge_1
Xpre_column_184 bl_184 br_184 en_bar vdd precharge_1
Xpre_column_185 bl_185 br_185 en_bar vdd precharge_1
Xpre_column_186 bl_186 br_186 en_bar vdd precharge_1
Xpre_column_187 bl_187 br_187 en_bar vdd precharge_1
Xpre_column_188 bl_188 br_188 en_bar vdd precharge_1
Xpre_column_189 bl_189 br_189 en_bar vdd precharge_1
Xpre_column_190 bl_190 br_190 en_bar vdd precharge_1
Xpre_column_191 bl_191 br_191 en_bar vdd precharge_1
Xpre_column_192 bl_192 br_192 en_bar vdd precharge_1
Xpre_column_193 bl_193 br_193 en_bar vdd precharge_1
Xpre_column_194 bl_194 br_194 en_bar vdd precharge_1
Xpre_column_195 bl_195 br_195 en_bar vdd precharge_1
Xpre_column_196 bl_196 br_196 en_bar vdd precharge_1
Xpre_column_197 bl_197 br_197 en_bar vdd precharge_1
Xpre_column_198 bl_198 br_198 en_bar vdd precharge_1
Xpre_column_199 bl_199 br_199 en_bar vdd precharge_1
Xpre_column_200 bl_200 br_200 en_bar vdd precharge_1
Xpre_column_201 bl_201 br_201 en_bar vdd precharge_1
Xpre_column_202 bl_202 br_202 en_bar vdd precharge_1
Xpre_column_203 bl_203 br_203 en_bar vdd precharge_1
Xpre_column_204 bl_204 br_204 en_bar vdd precharge_1
Xpre_column_205 bl_205 br_205 en_bar vdd precharge_1
Xpre_column_206 bl_206 br_206 en_bar vdd precharge_1
Xpre_column_207 bl_207 br_207 en_bar vdd precharge_1
Xpre_column_208 bl_208 br_208 en_bar vdd precharge_1
Xpre_column_209 bl_209 br_209 en_bar vdd precharge_1
Xpre_column_210 bl_210 br_210 en_bar vdd precharge_1
Xpre_column_211 bl_211 br_211 en_bar vdd precharge_1
Xpre_column_212 bl_212 br_212 en_bar vdd precharge_1
Xpre_column_213 bl_213 br_213 en_bar vdd precharge_1
Xpre_column_214 bl_214 br_214 en_bar vdd precharge_1
Xpre_column_215 bl_215 br_215 en_bar vdd precharge_1
Xpre_column_216 bl_216 br_216 en_bar vdd precharge_1
Xpre_column_217 bl_217 br_217 en_bar vdd precharge_1
Xpre_column_218 bl_218 br_218 en_bar vdd precharge_1
Xpre_column_219 bl_219 br_219 en_bar vdd precharge_1
Xpre_column_220 bl_220 br_220 en_bar vdd precharge_1
Xpre_column_221 bl_221 br_221 en_bar vdd precharge_1
Xpre_column_222 bl_222 br_222 en_bar vdd precharge_1
Xpre_column_223 bl_223 br_223 en_bar vdd precharge_1
Xpre_column_224 bl_224 br_224 en_bar vdd precharge_1
Xpre_column_225 bl_225 br_225 en_bar vdd precharge_1
Xpre_column_226 bl_226 br_226 en_bar vdd precharge_1
Xpre_column_227 bl_227 br_227 en_bar vdd precharge_1
Xpre_column_228 bl_228 br_228 en_bar vdd precharge_1
Xpre_column_229 bl_229 br_229 en_bar vdd precharge_1
Xpre_column_230 bl_230 br_230 en_bar vdd precharge_1
Xpre_column_231 bl_231 br_231 en_bar vdd precharge_1
Xpre_column_232 bl_232 br_232 en_bar vdd precharge_1
Xpre_column_233 bl_233 br_233 en_bar vdd precharge_1
Xpre_column_234 bl_234 br_234 en_bar vdd precharge_1
Xpre_column_235 bl_235 br_235 en_bar vdd precharge_1
Xpre_column_236 bl_236 br_236 en_bar vdd precharge_1
Xpre_column_237 bl_237 br_237 en_bar vdd precharge_1
Xpre_column_238 bl_238 br_238 en_bar vdd precharge_1
Xpre_column_239 bl_239 br_239 en_bar vdd precharge_1
Xpre_column_240 bl_240 br_240 en_bar vdd precharge_1
Xpre_column_241 bl_241 br_241 en_bar vdd precharge_1
Xpre_column_242 bl_242 br_242 en_bar vdd precharge_1
Xpre_column_243 bl_243 br_243 en_bar vdd precharge_1
Xpre_column_244 bl_244 br_244 en_bar vdd precharge_1
Xpre_column_245 bl_245 br_245 en_bar vdd precharge_1
Xpre_column_246 bl_246 br_246 en_bar vdd precharge_1
Xpre_column_247 bl_247 br_247 en_bar vdd precharge_1
Xpre_column_248 bl_248 br_248 en_bar vdd precharge_1
Xpre_column_249 bl_249 br_249 en_bar vdd precharge_1
Xpre_column_250 bl_250 br_250 en_bar vdd precharge_1
Xpre_column_251 bl_251 br_251 en_bar vdd precharge_1
Xpre_column_252 bl_252 br_252 en_bar vdd precharge_1
Xpre_column_253 bl_253 br_253 en_bar vdd precharge_1
Xpre_column_254 bl_254 br_254 en_bar vdd precharge_1
Xpre_column_255 bl_255 br_255 en_bar vdd precharge_1
Xpre_column_256 bl_256 br_256 en_bar vdd precharge_1
.ENDS precharge_array_0

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sense_amp_array_0 data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14 data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18 bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31 br_31 data_32 bl_32 br_32 data_33 bl_33 br_33 data_34 bl_34 br_34 data_35 bl_35 br_35 data_36 bl_36 br_36 data_37 bl_37 br_37 data_38 bl_38 br_38 data_39 bl_39 br_39 data_40 bl_40 br_40 data_41 bl_41 br_41 data_42 bl_42 br_42 data_43 bl_43 br_43 data_44 bl_44 br_44 data_45 bl_45 br_45 data_46 bl_46 br_46 data_47 bl_47 br_47 data_48 bl_48 br_48 data_49 bl_49 br_49 data_50 bl_50 br_50 data_51 bl_51 br_51 data_52 bl_52 br_52 data_53 bl_53 br_53 data_54 bl_54 br_54 data_55 bl_55 br_55 data_56 bl_56 br_56 data_57 bl_57 br_57 data_58 bl_58 br_58 data_59 bl_59 br_59 data_60 bl_60 br_60 data_61 bl_61 br_61 data_62 bl_62 br_62 data_63 bl_63 br_63 data_64 bl_64 br_64 data_65 bl_65 br_65 data_66 bl_66 br_66 data_67 bl_67 br_67 data_68 bl_68 br_68 data_69 bl_69 br_69 data_70 bl_70 br_70 data_71 bl_71 br_71 data_72 bl_72 br_72 data_73 bl_73 br_73 data_74 bl_74 br_74 data_75 bl_75 br_75 data_76 bl_76 br_76 data_77 bl_77 br_77 data_78 bl_78 br_78 data_79 bl_79 br_79 data_80 bl_80 br_80 data_81 bl_81 br_81 data_82 bl_82 br_82 data_83 bl_83 br_83 data_84 bl_84 br_84 data_85 bl_85 br_85 data_86 bl_86 br_86 data_87 bl_87 br_87 data_88 bl_88 br_88 data_89 bl_89 br_89 data_90 bl_90 br_90 data_91 bl_91 br_91 data_92 bl_92 br_92 data_93 bl_93 br_93 data_94 bl_94 br_94 data_95 bl_95 br_95 data_96 bl_96 br_96 data_97 bl_97 br_97 data_98 bl_98 br_98 data_99 bl_99 br_99 data_100 bl_100 br_100 data_101 bl_101 br_101 data_102 bl_102 br_102 data_103 bl_103 br_103 data_104 bl_104 br_104 data_105 bl_105 br_105 data_106 bl_106 br_106 data_107 bl_107 br_107 data_108 bl_108 br_108 data_109 bl_109 br_109 data_110 bl_110 br_110 data_111 bl_111 br_111 data_112 bl_112 br_112 data_113 bl_113 br_113 data_114 bl_114 br_114 data_115 bl_115 br_115 data_116 bl_116 br_116 data_117 bl_117 br_117 data_118 bl_118 br_118 data_119 bl_119 br_119 data_120 bl_120 br_120 data_121 bl_121 br_121 data_122 bl_122 br_122 data_123 bl_123 br_123 data_124 bl_124 br_124 data_125 bl_125 br_125 data_126 bl_126 br_126 data_127 bl_127 br_127 data_128 bl_128 br_128 data_129 bl_129 br_129 data_130 bl_130 br_130 data_131 bl_131 br_131 data_132 bl_132 br_132 data_133 bl_133 br_133 data_134 bl_134 br_134 data_135 bl_135 br_135 data_136 bl_136 br_136 data_137 bl_137 br_137 data_138 bl_138 br_138 data_139 bl_139 br_139 data_140 bl_140 br_140 data_141 bl_141 br_141 data_142 bl_142 br_142 data_143 bl_143 br_143 data_144 bl_144 br_144 data_145 bl_145 br_145 data_146 bl_146 br_146 data_147 bl_147 br_147 data_148 bl_148 br_148 data_149 bl_149 br_149 data_150 bl_150 br_150 data_151 bl_151 br_151 data_152 bl_152 br_152 data_153 bl_153 br_153 data_154 bl_154 br_154 data_155 bl_155 br_155 data_156 bl_156 br_156 data_157 bl_157 br_157 data_158 bl_158 br_158 data_159 bl_159 br_159 data_160 bl_160 br_160 data_161 bl_161 br_161 data_162 bl_162 br_162 data_163 bl_163 br_163 data_164 bl_164 br_164 data_165 bl_165 br_165 data_166 bl_166 br_166 data_167 bl_167 br_167 data_168 bl_168 br_168 data_169 bl_169 br_169 data_170 bl_170 br_170 data_171 bl_171 br_171 data_172 bl_172 br_172 data_173 bl_173 br_173 data_174 bl_174 br_174 data_175 bl_175 br_175 data_176 bl_176 br_176 data_177 bl_177 br_177 data_178 bl_178 br_178 data_179 bl_179 br_179 data_180 bl_180 br_180 data_181 bl_181 br_181 data_182 bl_182 br_182 data_183 bl_183 br_183 data_184 bl_184 br_184 data_185 bl_185 br_185 data_186 bl_186 br_186 data_187 bl_187 br_187 data_188 bl_188 br_188 data_189 bl_189 br_189 data_190 bl_190 br_190 data_191 bl_191 br_191 data_192 bl_192 br_192 data_193 bl_193 br_193 data_194 bl_194 br_194 data_195 bl_195 br_195 data_196 bl_196 br_196 data_197 bl_197 br_197 data_198 bl_198 br_198 data_199 bl_199 br_199 data_200 bl_200 br_200 data_201 bl_201 br_201 data_202 bl_202 br_202 data_203 bl_203 br_203 data_204 bl_204 br_204 data_205 bl_205 br_205 data_206 bl_206 br_206 data_207 bl_207 br_207 data_208 bl_208 br_208 data_209 bl_209 br_209 data_210 bl_210 br_210 data_211 bl_211 br_211 data_212 bl_212 br_212 data_213 bl_213 br_213 data_214 bl_214 br_214 data_215 bl_215 br_215 data_216 bl_216 br_216 data_217 bl_217 br_217 data_218 bl_218 br_218 data_219 bl_219 br_219 data_220 bl_220 br_220 data_221 bl_221 br_221 data_222 bl_222 br_222 data_223 bl_223 br_223 data_224 bl_224 br_224 data_225 bl_225 br_225 data_226 bl_226 br_226 data_227 bl_227 br_227 data_228 bl_228 br_228 data_229 bl_229 br_229 data_230 bl_230 br_230 data_231 bl_231 br_231 data_232 bl_232 br_232 data_233 bl_233 br_233 data_234 bl_234 br_234 data_235 bl_235 br_235 data_236 bl_236 br_236 data_237 bl_237 br_237 data_238 bl_238 br_238 data_239 bl_239 br_239 data_240 bl_240 br_240 data_241 bl_241 br_241 data_242 bl_242 br_242 data_243 bl_243 br_243 data_244 bl_244 br_244 data_245 bl_245 br_245 data_246 bl_246 br_246 data_247 bl_247 br_247 data_248 bl_248 br_248 data_249 bl_249 br_249 data_250 bl_250 br_250 data_251 bl_251 br_251 data_252 bl_252 br_252 data_253 bl_253 br_253 data_254 bl_254 br_254 data_255 bl_255 br_255 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* OUTPUT: data_32 
* INPUT : bl_32 
* INPUT : br_32 
* OUTPUT: data_33 
* INPUT : bl_33 
* INPUT : br_33 
* OUTPUT: data_34 
* INPUT : bl_34 
* INPUT : br_34 
* OUTPUT: data_35 
* INPUT : bl_35 
* INPUT : br_35 
* OUTPUT: data_36 
* INPUT : bl_36 
* INPUT : br_36 
* OUTPUT: data_37 
* INPUT : bl_37 
* INPUT : br_37 
* OUTPUT: data_38 
* INPUT : bl_38 
* INPUT : br_38 
* OUTPUT: data_39 
* INPUT : bl_39 
* INPUT : br_39 
* OUTPUT: data_40 
* INPUT : bl_40 
* INPUT : br_40 
* OUTPUT: data_41 
* INPUT : bl_41 
* INPUT : br_41 
* OUTPUT: data_42 
* INPUT : bl_42 
* INPUT : br_42 
* OUTPUT: data_43 
* INPUT : bl_43 
* INPUT : br_43 
* OUTPUT: data_44 
* INPUT : bl_44 
* INPUT : br_44 
* OUTPUT: data_45 
* INPUT : bl_45 
* INPUT : br_45 
* OUTPUT: data_46 
* INPUT : bl_46 
* INPUT : br_46 
* OUTPUT: data_47 
* INPUT : bl_47 
* INPUT : br_47 
* OUTPUT: data_48 
* INPUT : bl_48 
* INPUT : br_48 
* OUTPUT: data_49 
* INPUT : bl_49 
* INPUT : br_49 
* OUTPUT: data_50 
* INPUT : bl_50 
* INPUT : br_50 
* OUTPUT: data_51 
* INPUT : bl_51 
* INPUT : br_51 
* OUTPUT: data_52 
* INPUT : bl_52 
* INPUT : br_52 
* OUTPUT: data_53 
* INPUT : bl_53 
* INPUT : br_53 
* OUTPUT: data_54 
* INPUT : bl_54 
* INPUT : br_54 
* OUTPUT: data_55 
* INPUT : bl_55 
* INPUT : br_55 
* OUTPUT: data_56 
* INPUT : bl_56 
* INPUT : br_56 
* OUTPUT: data_57 
* INPUT : bl_57 
* INPUT : br_57 
* OUTPUT: data_58 
* INPUT : bl_58 
* INPUT : br_58 
* OUTPUT: data_59 
* INPUT : bl_59 
* INPUT : br_59 
* OUTPUT: data_60 
* INPUT : bl_60 
* INPUT : br_60 
* OUTPUT: data_61 
* INPUT : bl_61 
* INPUT : br_61 
* OUTPUT: data_62 
* INPUT : bl_62 
* INPUT : br_62 
* OUTPUT: data_63 
* INPUT : bl_63 
* INPUT : br_63 
* OUTPUT: data_64 
* INPUT : bl_64 
* INPUT : br_64 
* OUTPUT: data_65 
* INPUT : bl_65 
* INPUT : br_65 
* OUTPUT: data_66 
* INPUT : bl_66 
* INPUT : br_66 
* OUTPUT: data_67 
* INPUT : bl_67 
* INPUT : br_67 
* OUTPUT: data_68 
* INPUT : bl_68 
* INPUT : br_68 
* OUTPUT: data_69 
* INPUT : bl_69 
* INPUT : br_69 
* OUTPUT: data_70 
* INPUT : bl_70 
* INPUT : br_70 
* OUTPUT: data_71 
* INPUT : bl_71 
* INPUT : br_71 
* OUTPUT: data_72 
* INPUT : bl_72 
* INPUT : br_72 
* OUTPUT: data_73 
* INPUT : bl_73 
* INPUT : br_73 
* OUTPUT: data_74 
* INPUT : bl_74 
* INPUT : br_74 
* OUTPUT: data_75 
* INPUT : bl_75 
* INPUT : br_75 
* OUTPUT: data_76 
* INPUT : bl_76 
* INPUT : br_76 
* OUTPUT: data_77 
* INPUT : bl_77 
* INPUT : br_77 
* OUTPUT: data_78 
* INPUT : bl_78 
* INPUT : br_78 
* OUTPUT: data_79 
* INPUT : bl_79 
* INPUT : br_79 
* OUTPUT: data_80 
* INPUT : bl_80 
* INPUT : br_80 
* OUTPUT: data_81 
* INPUT : bl_81 
* INPUT : br_81 
* OUTPUT: data_82 
* INPUT : bl_82 
* INPUT : br_82 
* OUTPUT: data_83 
* INPUT : bl_83 
* INPUT : br_83 
* OUTPUT: data_84 
* INPUT : bl_84 
* INPUT : br_84 
* OUTPUT: data_85 
* INPUT : bl_85 
* INPUT : br_85 
* OUTPUT: data_86 
* INPUT : bl_86 
* INPUT : br_86 
* OUTPUT: data_87 
* INPUT : bl_87 
* INPUT : br_87 
* OUTPUT: data_88 
* INPUT : bl_88 
* INPUT : br_88 
* OUTPUT: data_89 
* INPUT : bl_89 
* INPUT : br_89 
* OUTPUT: data_90 
* INPUT : bl_90 
* INPUT : br_90 
* OUTPUT: data_91 
* INPUT : bl_91 
* INPUT : br_91 
* OUTPUT: data_92 
* INPUT : bl_92 
* INPUT : br_92 
* OUTPUT: data_93 
* INPUT : bl_93 
* INPUT : br_93 
* OUTPUT: data_94 
* INPUT : bl_94 
* INPUT : br_94 
* OUTPUT: data_95 
* INPUT : bl_95 
* INPUT : br_95 
* OUTPUT: data_96 
* INPUT : bl_96 
* INPUT : br_96 
* OUTPUT: data_97 
* INPUT : bl_97 
* INPUT : br_97 
* OUTPUT: data_98 
* INPUT : bl_98 
* INPUT : br_98 
* OUTPUT: data_99 
* INPUT : bl_99 
* INPUT : br_99 
* OUTPUT: data_100 
* INPUT : bl_100 
* INPUT : br_100 
* OUTPUT: data_101 
* INPUT : bl_101 
* INPUT : br_101 
* OUTPUT: data_102 
* INPUT : bl_102 
* INPUT : br_102 
* OUTPUT: data_103 
* INPUT : bl_103 
* INPUT : br_103 
* OUTPUT: data_104 
* INPUT : bl_104 
* INPUT : br_104 
* OUTPUT: data_105 
* INPUT : bl_105 
* INPUT : br_105 
* OUTPUT: data_106 
* INPUT : bl_106 
* INPUT : br_106 
* OUTPUT: data_107 
* INPUT : bl_107 
* INPUT : br_107 
* OUTPUT: data_108 
* INPUT : bl_108 
* INPUT : br_108 
* OUTPUT: data_109 
* INPUT : bl_109 
* INPUT : br_109 
* OUTPUT: data_110 
* INPUT : bl_110 
* INPUT : br_110 
* OUTPUT: data_111 
* INPUT : bl_111 
* INPUT : br_111 
* OUTPUT: data_112 
* INPUT : bl_112 
* INPUT : br_112 
* OUTPUT: data_113 
* INPUT : bl_113 
* INPUT : br_113 
* OUTPUT: data_114 
* INPUT : bl_114 
* INPUT : br_114 
* OUTPUT: data_115 
* INPUT : bl_115 
* INPUT : br_115 
* OUTPUT: data_116 
* INPUT : bl_116 
* INPUT : br_116 
* OUTPUT: data_117 
* INPUT : bl_117 
* INPUT : br_117 
* OUTPUT: data_118 
* INPUT : bl_118 
* INPUT : br_118 
* OUTPUT: data_119 
* INPUT : bl_119 
* INPUT : br_119 
* OUTPUT: data_120 
* INPUT : bl_120 
* INPUT : br_120 
* OUTPUT: data_121 
* INPUT : bl_121 
* INPUT : br_121 
* OUTPUT: data_122 
* INPUT : bl_122 
* INPUT : br_122 
* OUTPUT: data_123 
* INPUT : bl_123 
* INPUT : br_123 
* OUTPUT: data_124 
* INPUT : bl_124 
* INPUT : br_124 
* OUTPUT: data_125 
* INPUT : bl_125 
* INPUT : br_125 
* OUTPUT: data_126 
* INPUT : bl_126 
* INPUT : br_126 
* OUTPUT: data_127 
* INPUT : bl_127 
* INPUT : br_127 
* OUTPUT: data_128 
* INPUT : bl_128 
* INPUT : br_128 
* OUTPUT: data_129 
* INPUT : bl_129 
* INPUT : br_129 
* OUTPUT: data_130 
* INPUT : bl_130 
* INPUT : br_130 
* OUTPUT: data_131 
* INPUT : bl_131 
* INPUT : br_131 
* OUTPUT: data_132 
* INPUT : bl_132 
* INPUT : br_132 
* OUTPUT: data_133 
* INPUT : bl_133 
* INPUT : br_133 
* OUTPUT: data_134 
* INPUT : bl_134 
* INPUT : br_134 
* OUTPUT: data_135 
* INPUT : bl_135 
* INPUT : br_135 
* OUTPUT: data_136 
* INPUT : bl_136 
* INPUT : br_136 
* OUTPUT: data_137 
* INPUT : bl_137 
* INPUT : br_137 
* OUTPUT: data_138 
* INPUT : bl_138 
* INPUT : br_138 
* OUTPUT: data_139 
* INPUT : bl_139 
* INPUT : br_139 
* OUTPUT: data_140 
* INPUT : bl_140 
* INPUT : br_140 
* OUTPUT: data_141 
* INPUT : bl_141 
* INPUT : br_141 
* OUTPUT: data_142 
* INPUT : bl_142 
* INPUT : br_142 
* OUTPUT: data_143 
* INPUT : bl_143 
* INPUT : br_143 
* OUTPUT: data_144 
* INPUT : bl_144 
* INPUT : br_144 
* OUTPUT: data_145 
* INPUT : bl_145 
* INPUT : br_145 
* OUTPUT: data_146 
* INPUT : bl_146 
* INPUT : br_146 
* OUTPUT: data_147 
* INPUT : bl_147 
* INPUT : br_147 
* OUTPUT: data_148 
* INPUT : bl_148 
* INPUT : br_148 
* OUTPUT: data_149 
* INPUT : bl_149 
* INPUT : br_149 
* OUTPUT: data_150 
* INPUT : bl_150 
* INPUT : br_150 
* OUTPUT: data_151 
* INPUT : bl_151 
* INPUT : br_151 
* OUTPUT: data_152 
* INPUT : bl_152 
* INPUT : br_152 
* OUTPUT: data_153 
* INPUT : bl_153 
* INPUT : br_153 
* OUTPUT: data_154 
* INPUT : bl_154 
* INPUT : br_154 
* OUTPUT: data_155 
* INPUT : bl_155 
* INPUT : br_155 
* OUTPUT: data_156 
* INPUT : bl_156 
* INPUT : br_156 
* OUTPUT: data_157 
* INPUT : bl_157 
* INPUT : br_157 
* OUTPUT: data_158 
* INPUT : bl_158 
* INPUT : br_158 
* OUTPUT: data_159 
* INPUT : bl_159 
* INPUT : br_159 
* OUTPUT: data_160 
* INPUT : bl_160 
* INPUT : br_160 
* OUTPUT: data_161 
* INPUT : bl_161 
* INPUT : br_161 
* OUTPUT: data_162 
* INPUT : bl_162 
* INPUT : br_162 
* OUTPUT: data_163 
* INPUT : bl_163 
* INPUT : br_163 
* OUTPUT: data_164 
* INPUT : bl_164 
* INPUT : br_164 
* OUTPUT: data_165 
* INPUT : bl_165 
* INPUT : br_165 
* OUTPUT: data_166 
* INPUT : bl_166 
* INPUT : br_166 
* OUTPUT: data_167 
* INPUT : bl_167 
* INPUT : br_167 
* OUTPUT: data_168 
* INPUT : bl_168 
* INPUT : br_168 
* OUTPUT: data_169 
* INPUT : bl_169 
* INPUT : br_169 
* OUTPUT: data_170 
* INPUT : bl_170 
* INPUT : br_170 
* OUTPUT: data_171 
* INPUT : bl_171 
* INPUT : br_171 
* OUTPUT: data_172 
* INPUT : bl_172 
* INPUT : br_172 
* OUTPUT: data_173 
* INPUT : bl_173 
* INPUT : br_173 
* OUTPUT: data_174 
* INPUT : bl_174 
* INPUT : br_174 
* OUTPUT: data_175 
* INPUT : bl_175 
* INPUT : br_175 
* OUTPUT: data_176 
* INPUT : bl_176 
* INPUT : br_176 
* OUTPUT: data_177 
* INPUT : bl_177 
* INPUT : br_177 
* OUTPUT: data_178 
* INPUT : bl_178 
* INPUT : br_178 
* OUTPUT: data_179 
* INPUT : bl_179 
* INPUT : br_179 
* OUTPUT: data_180 
* INPUT : bl_180 
* INPUT : br_180 
* OUTPUT: data_181 
* INPUT : bl_181 
* INPUT : br_181 
* OUTPUT: data_182 
* INPUT : bl_182 
* INPUT : br_182 
* OUTPUT: data_183 
* INPUT : bl_183 
* INPUT : br_183 
* OUTPUT: data_184 
* INPUT : bl_184 
* INPUT : br_184 
* OUTPUT: data_185 
* INPUT : bl_185 
* INPUT : br_185 
* OUTPUT: data_186 
* INPUT : bl_186 
* INPUT : br_186 
* OUTPUT: data_187 
* INPUT : bl_187 
* INPUT : br_187 
* OUTPUT: data_188 
* INPUT : bl_188 
* INPUT : br_188 
* OUTPUT: data_189 
* INPUT : bl_189 
* INPUT : br_189 
* OUTPUT: data_190 
* INPUT : bl_190 
* INPUT : br_190 
* OUTPUT: data_191 
* INPUT : bl_191 
* INPUT : br_191 
* OUTPUT: data_192 
* INPUT : bl_192 
* INPUT : br_192 
* OUTPUT: data_193 
* INPUT : bl_193 
* INPUT : br_193 
* OUTPUT: data_194 
* INPUT : bl_194 
* INPUT : br_194 
* OUTPUT: data_195 
* INPUT : bl_195 
* INPUT : br_195 
* OUTPUT: data_196 
* INPUT : bl_196 
* INPUT : br_196 
* OUTPUT: data_197 
* INPUT : bl_197 
* INPUT : br_197 
* OUTPUT: data_198 
* INPUT : bl_198 
* INPUT : br_198 
* OUTPUT: data_199 
* INPUT : bl_199 
* INPUT : br_199 
* OUTPUT: data_200 
* INPUT : bl_200 
* INPUT : br_200 
* OUTPUT: data_201 
* INPUT : bl_201 
* INPUT : br_201 
* OUTPUT: data_202 
* INPUT : bl_202 
* INPUT : br_202 
* OUTPUT: data_203 
* INPUT : bl_203 
* INPUT : br_203 
* OUTPUT: data_204 
* INPUT : bl_204 
* INPUT : br_204 
* OUTPUT: data_205 
* INPUT : bl_205 
* INPUT : br_205 
* OUTPUT: data_206 
* INPUT : bl_206 
* INPUT : br_206 
* OUTPUT: data_207 
* INPUT : bl_207 
* INPUT : br_207 
* OUTPUT: data_208 
* INPUT : bl_208 
* INPUT : br_208 
* OUTPUT: data_209 
* INPUT : bl_209 
* INPUT : br_209 
* OUTPUT: data_210 
* INPUT : bl_210 
* INPUT : br_210 
* OUTPUT: data_211 
* INPUT : bl_211 
* INPUT : br_211 
* OUTPUT: data_212 
* INPUT : bl_212 
* INPUT : br_212 
* OUTPUT: data_213 
* INPUT : bl_213 
* INPUT : br_213 
* OUTPUT: data_214 
* INPUT : bl_214 
* INPUT : br_214 
* OUTPUT: data_215 
* INPUT : bl_215 
* INPUT : br_215 
* OUTPUT: data_216 
* INPUT : bl_216 
* INPUT : br_216 
* OUTPUT: data_217 
* INPUT : bl_217 
* INPUT : br_217 
* OUTPUT: data_218 
* INPUT : bl_218 
* INPUT : br_218 
* OUTPUT: data_219 
* INPUT : bl_219 
* INPUT : br_219 
* OUTPUT: data_220 
* INPUT : bl_220 
* INPUT : br_220 
* OUTPUT: data_221 
* INPUT : bl_221 
* INPUT : br_221 
* OUTPUT: data_222 
* INPUT : bl_222 
* INPUT : br_222 
* OUTPUT: data_223 
* INPUT : bl_223 
* INPUT : br_223 
* OUTPUT: data_224 
* INPUT : bl_224 
* INPUT : br_224 
* OUTPUT: data_225 
* INPUT : bl_225 
* INPUT : br_225 
* OUTPUT: data_226 
* INPUT : bl_226 
* INPUT : br_226 
* OUTPUT: data_227 
* INPUT : bl_227 
* INPUT : br_227 
* OUTPUT: data_228 
* INPUT : bl_228 
* INPUT : br_228 
* OUTPUT: data_229 
* INPUT : bl_229 
* INPUT : br_229 
* OUTPUT: data_230 
* INPUT : bl_230 
* INPUT : br_230 
* OUTPUT: data_231 
* INPUT : bl_231 
* INPUT : br_231 
* OUTPUT: data_232 
* INPUT : bl_232 
* INPUT : br_232 
* OUTPUT: data_233 
* INPUT : bl_233 
* INPUT : br_233 
* OUTPUT: data_234 
* INPUT : bl_234 
* INPUT : br_234 
* OUTPUT: data_235 
* INPUT : bl_235 
* INPUT : br_235 
* OUTPUT: data_236 
* INPUT : bl_236 
* INPUT : br_236 
* OUTPUT: data_237 
* INPUT : bl_237 
* INPUT : br_237 
* OUTPUT: data_238 
* INPUT : bl_238 
* INPUT : br_238 
* OUTPUT: data_239 
* INPUT : bl_239 
* INPUT : br_239 
* OUTPUT: data_240 
* INPUT : bl_240 
* INPUT : br_240 
* OUTPUT: data_241 
* INPUT : bl_241 
* INPUT : br_241 
* OUTPUT: data_242 
* INPUT : bl_242 
* INPUT : br_242 
* OUTPUT: data_243 
* INPUT : bl_243 
* INPUT : br_243 
* OUTPUT: data_244 
* INPUT : bl_244 
* INPUT : br_244 
* OUTPUT: data_245 
* INPUT : bl_245 
* INPUT : br_245 
* OUTPUT: data_246 
* INPUT : bl_246 
* INPUT : br_246 
* OUTPUT: data_247 
* INPUT : bl_247 
* INPUT : br_247 
* OUTPUT: data_248 
* INPUT : bl_248 
* INPUT : br_248 
* OUTPUT: data_249 
* INPUT : bl_249 
* INPUT : br_249 
* OUTPUT: data_250 
* INPUT : bl_250 
* INPUT : br_250 
* OUTPUT: data_251 
* INPUT : bl_251 
* INPUT : br_251 
* OUTPUT: data_252 
* INPUT : bl_252 
* INPUT : br_252 
* OUTPUT: data_253 
* INPUT : bl_253 
* INPUT : br_253 
* OUTPUT: data_254 
* INPUT : bl_254 
* INPUT : br_254 
* OUTPUT: data_255 
* INPUT : bl_255 
* INPUT : br_255 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 1
Xsa_d0 bl_0 br_0 data_0 en vdd gnd sense_amp
Xsa_d1 bl_1 br_1 data_1 en vdd gnd sense_amp
Xsa_d2 bl_2 br_2 data_2 en vdd gnd sense_amp
Xsa_d3 bl_3 br_3 data_3 en vdd gnd sense_amp
Xsa_d4 bl_4 br_4 data_4 en vdd gnd sense_amp
Xsa_d5 bl_5 br_5 data_5 en vdd gnd sense_amp
Xsa_d6 bl_6 br_6 data_6 en vdd gnd sense_amp
Xsa_d7 bl_7 br_7 data_7 en vdd gnd sense_amp
Xsa_d8 bl_8 br_8 data_8 en vdd gnd sense_amp
Xsa_d9 bl_9 br_9 data_9 en vdd gnd sense_amp
Xsa_d10 bl_10 br_10 data_10 en vdd gnd sense_amp
Xsa_d11 bl_11 br_11 data_11 en vdd gnd sense_amp
Xsa_d12 bl_12 br_12 data_12 en vdd gnd sense_amp
Xsa_d13 bl_13 br_13 data_13 en vdd gnd sense_amp
Xsa_d14 bl_14 br_14 data_14 en vdd gnd sense_amp
Xsa_d15 bl_15 br_15 data_15 en vdd gnd sense_amp
Xsa_d16 bl_16 br_16 data_16 en vdd gnd sense_amp
Xsa_d17 bl_17 br_17 data_17 en vdd gnd sense_amp
Xsa_d18 bl_18 br_18 data_18 en vdd gnd sense_amp
Xsa_d19 bl_19 br_19 data_19 en vdd gnd sense_amp
Xsa_d20 bl_20 br_20 data_20 en vdd gnd sense_amp
Xsa_d21 bl_21 br_21 data_21 en vdd gnd sense_amp
Xsa_d22 bl_22 br_22 data_22 en vdd gnd sense_amp
Xsa_d23 bl_23 br_23 data_23 en vdd gnd sense_amp
Xsa_d24 bl_24 br_24 data_24 en vdd gnd sense_amp
Xsa_d25 bl_25 br_25 data_25 en vdd gnd sense_amp
Xsa_d26 bl_26 br_26 data_26 en vdd gnd sense_amp
Xsa_d27 bl_27 br_27 data_27 en vdd gnd sense_amp
Xsa_d28 bl_28 br_28 data_28 en vdd gnd sense_amp
Xsa_d29 bl_29 br_29 data_29 en vdd gnd sense_amp
Xsa_d30 bl_30 br_30 data_30 en vdd gnd sense_amp
Xsa_d31 bl_31 br_31 data_31 en vdd gnd sense_amp
Xsa_d32 bl_32 br_32 data_32 en vdd gnd sense_amp
Xsa_d33 bl_33 br_33 data_33 en vdd gnd sense_amp
Xsa_d34 bl_34 br_34 data_34 en vdd gnd sense_amp
Xsa_d35 bl_35 br_35 data_35 en vdd gnd sense_amp
Xsa_d36 bl_36 br_36 data_36 en vdd gnd sense_amp
Xsa_d37 bl_37 br_37 data_37 en vdd gnd sense_amp
Xsa_d38 bl_38 br_38 data_38 en vdd gnd sense_amp
Xsa_d39 bl_39 br_39 data_39 en vdd gnd sense_amp
Xsa_d40 bl_40 br_40 data_40 en vdd gnd sense_amp
Xsa_d41 bl_41 br_41 data_41 en vdd gnd sense_amp
Xsa_d42 bl_42 br_42 data_42 en vdd gnd sense_amp
Xsa_d43 bl_43 br_43 data_43 en vdd gnd sense_amp
Xsa_d44 bl_44 br_44 data_44 en vdd gnd sense_amp
Xsa_d45 bl_45 br_45 data_45 en vdd gnd sense_amp
Xsa_d46 bl_46 br_46 data_46 en vdd gnd sense_amp
Xsa_d47 bl_47 br_47 data_47 en vdd gnd sense_amp
Xsa_d48 bl_48 br_48 data_48 en vdd gnd sense_amp
Xsa_d49 bl_49 br_49 data_49 en vdd gnd sense_amp
Xsa_d50 bl_50 br_50 data_50 en vdd gnd sense_amp
Xsa_d51 bl_51 br_51 data_51 en vdd gnd sense_amp
Xsa_d52 bl_52 br_52 data_52 en vdd gnd sense_amp
Xsa_d53 bl_53 br_53 data_53 en vdd gnd sense_amp
Xsa_d54 bl_54 br_54 data_54 en vdd gnd sense_amp
Xsa_d55 bl_55 br_55 data_55 en vdd gnd sense_amp
Xsa_d56 bl_56 br_56 data_56 en vdd gnd sense_amp
Xsa_d57 bl_57 br_57 data_57 en vdd gnd sense_amp
Xsa_d58 bl_58 br_58 data_58 en vdd gnd sense_amp
Xsa_d59 bl_59 br_59 data_59 en vdd gnd sense_amp
Xsa_d60 bl_60 br_60 data_60 en vdd gnd sense_amp
Xsa_d61 bl_61 br_61 data_61 en vdd gnd sense_amp
Xsa_d62 bl_62 br_62 data_62 en vdd gnd sense_amp
Xsa_d63 bl_63 br_63 data_63 en vdd gnd sense_amp
Xsa_d64 bl_64 br_64 data_64 en vdd gnd sense_amp
Xsa_d65 bl_65 br_65 data_65 en vdd gnd sense_amp
Xsa_d66 bl_66 br_66 data_66 en vdd gnd sense_amp
Xsa_d67 bl_67 br_67 data_67 en vdd gnd sense_amp
Xsa_d68 bl_68 br_68 data_68 en vdd gnd sense_amp
Xsa_d69 bl_69 br_69 data_69 en vdd gnd sense_amp
Xsa_d70 bl_70 br_70 data_70 en vdd gnd sense_amp
Xsa_d71 bl_71 br_71 data_71 en vdd gnd sense_amp
Xsa_d72 bl_72 br_72 data_72 en vdd gnd sense_amp
Xsa_d73 bl_73 br_73 data_73 en vdd gnd sense_amp
Xsa_d74 bl_74 br_74 data_74 en vdd gnd sense_amp
Xsa_d75 bl_75 br_75 data_75 en vdd gnd sense_amp
Xsa_d76 bl_76 br_76 data_76 en vdd gnd sense_amp
Xsa_d77 bl_77 br_77 data_77 en vdd gnd sense_amp
Xsa_d78 bl_78 br_78 data_78 en vdd gnd sense_amp
Xsa_d79 bl_79 br_79 data_79 en vdd gnd sense_amp
Xsa_d80 bl_80 br_80 data_80 en vdd gnd sense_amp
Xsa_d81 bl_81 br_81 data_81 en vdd gnd sense_amp
Xsa_d82 bl_82 br_82 data_82 en vdd gnd sense_amp
Xsa_d83 bl_83 br_83 data_83 en vdd gnd sense_amp
Xsa_d84 bl_84 br_84 data_84 en vdd gnd sense_amp
Xsa_d85 bl_85 br_85 data_85 en vdd gnd sense_amp
Xsa_d86 bl_86 br_86 data_86 en vdd gnd sense_amp
Xsa_d87 bl_87 br_87 data_87 en vdd gnd sense_amp
Xsa_d88 bl_88 br_88 data_88 en vdd gnd sense_amp
Xsa_d89 bl_89 br_89 data_89 en vdd gnd sense_amp
Xsa_d90 bl_90 br_90 data_90 en vdd gnd sense_amp
Xsa_d91 bl_91 br_91 data_91 en vdd gnd sense_amp
Xsa_d92 bl_92 br_92 data_92 en vdd gnd sense_amp
Xsa_d93 bl_93 br_93 data_93 en vdd gnd sense_amp
Xsa_d94 bl_94 br_94 data_94 en vdd gnd sense_amp
Xsa_d95 bl_95 br_95 data_95 en vdd gnd sense_amp
Xsa_d96 bl_96 br_96 data_96 en vdd gnd sense_amp
Xsa_d97 bl_97 br_97 data_97 en vdd gnd sense_amp
Xsa_d98 bl_98 br_98 data_98 en vdd gnd sense_amp
Xsa_d99 bl_99 br_99 data_99 en vdd gnd sense_amp
Xsa_d100 bl_100 br_100 data_100 en vdd gnd sense_amp
Xsa_d101 bl_101 br_101 data_101 en vdd gnd sense_amp
Xsa_d102 bl_102 br_102 data_102 en vdd gnd sense_amp
Xsa_d103 bl_103 br_103 data_103 en vdd gnd sense_amp
Xsa_d104 bl_104 br_104 data_104 en vdd gnd sense_amp
Xsa_d105 bl_105 br_105 data_105 en vdd gnd sense_amp
Xsa_d106 bl_106 br_106 data_106 en vdd gnd sense_amp
Xsa_d107 bl_107 br_107 data_107 en vdd gnd sense_amp
Xsa_d108 bl_108 br_108 data_108 en vdd gnd sense_amp
Xsa_d109 bl_109 br_109 data_109 en vdd gnd sense_amp
Xsa_d110 bl_110 br_110 data_110 en vdd gnd sense_amp
Xsa_d111 bl_111 br_111 data_111 en vdd gnd sense_amp
Xsa_d112 bl_112 br_112 data_112 en vdd gnd sense_amp
Xsa_d113 bl_113 br_113 data_113 en vdd gnd sense_amp
Xsa_d114 bl_114 br_114 data_114 en vdd gnd sense_amp
Xsa_d115 bl_115 br_115 data_115 en vdd gnd sense_amp
Xsa_d116 bl_116 br_116 data_116 en vdd gnd sense_amp
Xsa_d117 bl_117 br_117 data_117 en vdd gnd sense_amp
Xsa_d118 bl_118 br_118 data_118 en vdd gnd sense_amp
Xsa_d119 bl_119 br_119 data_119 en vdd gnd sense_amp
Xsa_d120 bl_120 br_120 data_120 en vdd gnd sense_amp
Xsa_d121 bl_121 br_121 data_121 en vdd gnd sense_amp
Xsa_d122 bl_122 br_122 data_122 en vdd gnd sense_amp
Xsa_d123 bl_123 br_123 data_123 en vdd gnd sense_amp
Xsa_d124 bl_124 br_124 data_124 en vdd gnd sense_amp
Xsa_d125 bl_125 br_125 data_125 en vdd gnd sense_amp
Xsa_d126 bl_126 br_126 data_126 en vdd gnd sense_amp
Xsa_d127 bl_127 br_127 data_127 en vdd gnd sense_amp
Xsa_d128 bl_128 br_128 data_128 en vdd gnd sense_amp
Xsa_d129 bl_129 br_129 data_129 en vdd gnd sense_amp
Xsa_d130 bl_130 br_130 data_130 en vdd gnd sense_amp
Xsa_d131 bl_131 br_131 data_131 en vdd gnd sense_amp
Xsa_d132 bl_132 br_132 data_132 en vdd gnd sense_amp
Xsa_d133 bl_133 br_133 data_133 en vdd gnd sense_amp
Xsa_d134 bl_134 br_134 data_134 en vdd gnd sense_amp
Xsa_d135 bl_135 br_135 data_135 en vdd gnd sense_amp
Xsa_d136 bl_136 br_136 data_136 en vdd gnd sense_amp
Xsa_d137 bl_137 br_137 data_137 en vdd gnd sense_amp
Xsa_d138 bl_138 br_138 data_138 en vdd gnd sense_amp
Xsa_d139 bl_139 br_139 data_139 en vdd gnd sense_amp
Xsa_d140 bl_140 br_140 data_140 en vdd gnd sense_amp
Xsa_d141 bl_141 br_141 data_141 en vdd gnd sense_amp
Xsa_d142 bl_142 br_142 data_142 en vdd gnd sense_amp
Xsa_d143 bl_143 br_143 data_143 en vdd gnd sense_amp
Xsa_d144 bl_144 br_144 data_144 en vdd gnd sense_amp
Xsa_d145 bl_145 br_145 data_145 en vdd gnd sense_amp
Xsa_d146 bl_146 br_146 data_146 en vdd gnd sense_amp
Xsa_d147 bl_147 br_147 data_147 en vdd gnd sense_amp
Xsa_d148 bl_148 br_148 data_148 en vdd gnd sense_amp
Xsa_d149 bl_149 br_149 data_149 en vdd gnd sense_amp
Xsa_d150 bl_150 br_150 data_150 en vdd gnd sense_amp
Xsa_d151 bl_151 br_151 data_151 en vdd gnd sense_amp
Xsa_d152 bl_152 br_152 data_152 en vdd gnd sense_amp
Xsa_d153 bl_153 br_153 data_153 en vdd gnd sense_amp
Xsa_d154 bl_154 br_154 data_154 en vdd gnd sense_amp
Xsa_d155 bl_155 br_155 data_155 en vdd gnd sense_amp
Xsa_d156 bl_156 br_156 data_156 en vdd gnd sense_amp
Xsa_d157 bl_157 br_157 data_157 en vdd gnd sense_amp
Xsa_d158 bl_158 br_158 data_158 en vdd gnd sense_amp
Xsa_d159 bl_159 br_159 data_159 en vdd gnd sense_amp
Xsa_d160 bl_160 br_160 data_160 en vdd gnd sense_amp
Xsa_d161 bl_161 br_161 data_161 en vdd gnd sense_amp
Xsa_d162 bl_162 br_162 data_162 en vdd gnd sense_amp
Xsa_d163 bl_163 br_163 data_163 en vdd gnd sense_amp
Xsa_d164 bl_164 br_164 data_164 en vdd gnd sense_amp
Xsa_d165 bl_165 br_165 data_165 en vdd gnd sense_amp
Xsa_d166 bl_166 br_166 data_166 en vdd gnd sense_amp
Xsa_d167 bl_167 br_167 data_167 en vdd gnd sense_amp
Xsa_d168 bl_168 br_168 data_168 en vdd gnd sense_amp
Xsa_d169 bl_169 br_169 data_169 en vdd gnd sense_amp
Xsa_d170 bl_170 br_170 data_170 en vdd gnd sense_amp
Xsa_d171 bl_171 br_171 data_171 en vdd gnd sense_amp
Xsa_d172 bl_172 br_172 data_172 en vdd gnd sense_amp
Xsa_d173 bl_173 br_173 data_173 en vdd gnd sense_amp
Xsa_d174 bl_174 br_174 data_174 en vdd gnd sense_amp
Xsa_d175 bl_175 br_175 data_175 en vdd gnd sense_amp
Xsa_d176 bl_176 br_176 data_176 en vdd gnd sense_amp
Xsa_d177 bl_177 br_177 data_177 en vdd gnd sense_amp
Xsa_d178 bl_178 br_178 data_178 en vdd gnd sense_amp
Xsa_d179 bl_179 br_179 data_179 en vdd gnd sense_amp
Xsa_d180 bl_180 br_180 data_180 en vdd gnd sense_amp
Xsa_d181 bl_181 br_181 data_181 en vdd gnd sense_amp
Xsa_d182 bl_182 br_182 data_182 en vdd gnd sense_amp
Xsa_d183 bl_183 br_183 data_183 en vdd gnd sense_amp
Xsa_d184 bl_184 br_184 data_184 en vdd gnd sense_amp
Xsa_d185 bl_185 br_185 data_185 en vdd gnd sense_amp
Xsa_d186 bl_186 br_186 data_186 en vdd gnd sense_amp
Xsa_d187 bl_187 br_187 data_187 en vdd gnd sense_amp
Xsa_d188 bl_188 br_188 data_188 en vdd gnd sense_amp
Xsa_d189 bl_189 br_189 data_189 en vdd gnd sense_amp
Xsa_d190 bl_190 br_190 data_190 en vdd gnd sense_amp
Xsa_d191 bl_191 br_191 data_191 en vdd gnd sense_amp
Xsa_d192 bl_192 br_192 data_192 en vdd gnd sense_amp
Xsa_d193 bl_193 br_193 data_193 en vdd gnd sense_amp
Xsa_d194 bl_194 br_194 data_194 en vdd gnd sense_amp
Xsa_d195 bl_195 br_195 data_195 en vdd gnd sense_amp
Xsa_d196 bl_196 br_196 data_196 en vdd gnd sense_amp
Xsa_d197 bl_197 br_197 data_197 en vdd gnd sense_amp
Xsa_d198 bl_198 br_198 data_198 en vdd gnd sense_amp
Xsa_d199 bl_199 br_199 data_199 en vdd gnd sense_amp
Xsa_d200 bl_200 br_200 data_200 en vdd gnd sense_amp
Xsa_d201 bl_201 br_201 data_201 en vdd gnd sense_amp
Xsa_d202 bl_202 br_202 data_202 en vdd gnd sense_amp
Xsa_d203 bl_203 br_203 data_203 en vdd gnd sense_amp
Xsa_d204 bl_204 br_204 data_204 en vdd gnd sense_amp
Xsa_d205 bl_205 br_205 data_205 en vdd gnd sense_amp
Xsa_d206 bl_206 br_206 data_206 en vdd gnd sense_amp
Xsa_d207 bl_207 br_207 data_207 en vdd gnd sense_amp
Xsa_d208 bl_208 br_208 data_208 en vdd gnd sense_amp
Xsa_d209 bl_209 br_209 data_209 en vdd gnd sense_amp
Xsa_d210 bl_210 br_210 data_210 en vdd gnd sense_amp
Xsa_d211 bl_211 br_211 data_211 en vdd gnd sense_amp
Xsa_d212 bl_212 br_212 data_212 en vdd gnd sense_amp
Xsa_d213 bl_213 br_213 data_213 en vdd gnd sense_amp
Xsa_d214 bl_214 br_214 data_214 en vdd gnd sense_amp
Xsa_d215 bl_215 br_215 data_215 en vdd gnd sense_amp
Xsa_d216 bl_216 br_216 data_216 en vdd gnd sense_amp
Xsa_d217 bl_217 br_217 data_217 en vdd gnd sense_amp
Xsa_d218 bl_218 br_218 data_218 en vdd gnd sense_amp
Xsa_d219 bl_219 br_219 data_219 en vdd gnd sense_amp
Xsa_d220 bl_220 br_220 data_220 en vdd gnd sense_amp
Xsa_d221 bl_221 br_221 data_221 en vdd gnd sense_amp
Xsa_d222 bl_222 br_222 data_222 en vdd gnd sense_amp
Xsa_d223 bl_223 br_223 data_223 en vdd gnd sense_amp
Xsa_d224 bl_224 br_224 data_224 en vdd gnd sense_amp
Xsa_d225 bl_225 br_225 data_225 en vdd gnd sense_amp
Xsa_d226 bl_226 br_226 data_226 en vdd gnd sense_amp
Xsa_d227 bl_227 br_227 data_227 en vdd gnd sense_amp
Xsa_d228 bl_228 br_228 data_228 en vdd gnd sense_amp
Xsa_d229 bl_229 br_229 data_229 en vdd gnd sense_amp
Xsa_d230 bl_230 br_230 data_230 en vdd gnd sense_amp
Xsa_d231 bl_231 br_231 data_231 en vdd gnd sense_amp
Xsa_d232 bl_232 br_232 data_232 en vdd gnd sense_amp
Xsa_d233 bl_233 br_233 data_233 en vdd gnd sense_amp
Xsa_d234 bl_234 br_234 data_234 en vdd gnd sense_amp
Xsa_d235 bl_235 br_235 data_235 en vdd gnd sense_amp
Xsa_d236 bl_236 br_236 data_236 en vdd gnd sense_amp
Xsa_d237 bl_237 br_237 data_237 en vdd gnd sense_amp
Xsa_d238 bl_238 br_238 data_238 en vdd gnd sense_amp
Xsa_d239 bl_239 br_239 data_239 en vdd gnd sense_amp
Xsa_d240 bl_240 br_240 data_240 en vdd gnd sense_amp
Xsa_d241 bl_241 br_241 data_241 en vdd gnd sense_amp
Xsa_d242 bl_242 br_242 data_242 en vdd gnd sense_amp
Xsa_d243 bl_243 br_243 data_243 en vdd gnd sense_amp
Xsa_d244 bl_244 br_244 data_244 en vdd gnd sense_amp
Xsa_d245 bl_245 br_245 data_245 en vdd gnd sense_amp
Xsa_d246 bl_246 br_246 data_246 en vdd gnd sense_amp
Xsa_d247 bl_247 br_247 data_247 en vdd gnd sense_amp
Xsa_d248 bl_248 br_248 data_248 en vdd gnd sense_amp
Xsa_d249 bl_249 br_249 data_249 en vdd gnd sense_amp
Xsa_d250 bl_250 br_250 data_250 en vdd gnd sense_amp
Xsa_d251 bl_251 br_251 data_251 en vdd gnd sense_amp
Xsa_d252 bl_252 br_252 data_252 en vdd gnd sense_amp
Xsa_d253 bl_253 br_253 data_253 en vdd gnd sense_amp
Xsa_d254 bl_254 br_254 data_254 en vdd gnd sense_amp
Xsa_d255 bl_255 br_255 data_255 en vdd gnd sense_amp
.ENDS sense_amp_array_0

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT write_driver_array_0 data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9 data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17 data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25 data_26 data_27 data_28 data_29 data_30 data_31 data_32 data_33 data_34 data_35 data_36 data_37 data_38 data_39 data_40 data_41 data_42 data_43 data_44 data_45 data_46 data_47 data_48 data_49 data_50 data_51 data_52 data_53 data_54 data_55 data_56 data_57 data_58 data_59 data_60 data_61 data_62 data_63 data_64 data_65 data_66 data_67 data_68 data_69 data_70 data_71 data_72 data_73 data_74 data_75 data_76 data_77 data_78 data_79 data_80 data_81 data_82 data_83 data_84 data_85 data_86 data_87 data_88 data_89 data_90 data_91 data_92 data_93 data_94 data_95 data_96 data_97 data_98 data_99 data_100 data_101 data_102 data_103 data_104 data_105 data_106 data_107 data_108 data_109 data_110 data_111 data_112 data_113 data_114 data_115 data_116 data_117 data_118 data_119 data_120 data_121 data_122 data_123 data_124 data_125 data_126 data_127 data_128 data_129 data_130 data_131 data_132 data_133 data_134 data_135 data_136 data_137 data_138 data_139 data_140 data_141 data_142 data_143 data_144 data_145 data_146 data_147 data_148 data_149 data_150 data_151 data_152 data_153 data_154 data_155 data_156 data_157 data_158 data_159 data_160 data_161 data_162 data_163 data_164 data_165 data_166 data_167 data_168 data_169 data_170 data_171 data_172 data_173 data_174 data_175 data_176 data_177 data_178 data_179 data_180 data_181 data_182 data_183 data_184 data_185 data_186 data_187 data_188 data_189 data_190 data_191 data_192 data_193 data_194 data_195 data_196 data_197 data_198 data_199 data_200 data_201 data_202 data_203 data_204 data_205 data_206 data_207 data_208 data_209 data_210 data_211 data_212 data_213 data_214 data_215 data_216 data_217 data_218 data_219 data_220 data_221 data_222 data_223 data_224 data_225 data_226 data_227 data_228 data_229 data_230 data_231 data_232 data_233 data_234 data_235 data_236 data_237 data_238 data_239 data_240 data_241 data_242 data_243 data_244 data_245 data_246 data_247 data_248 data_249 data_250 data_251 data_252 data_253 data_254 data_255 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 en vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* INPUT : data_32 
* INPUT : data_33 
* INPUT : data_34 
* INPUT : data_35 
* INPUT : data_36 
* INPUT : data_37 
* INPUT : data_38 
* INPUT : data_39 
* INPUT : data_40 
* INPUT : data_41 
* INPUT : data_42 
* INPUT : data_43 
* INPUT : data_44 
* INPUT : data_45 
* INPUT : data_46 
* INPUT : data_47 
* INPUT : data_48 
* INPUT : data_49 
* INPUT : data_50 
* INPUT : data_51 
* INPUT : data_52 
* INPUT : data_53 
* INPUT : data_54 
* INPUT : data_55 
* INPUT : data_56 
* INPUT : data_57 
* INPUT : data_58 
* INPUT : data_59 
* INPUT : data_60 
* INPUT : data_61 
* INPUT : data_62 
* INPUT : data_63 
* INPUT : data_64 
* INPUT : data_65 
* INPUT : data_66 
* INPUT : data_67 
* INPUT : data_68 
* INPUT : data_69 
* INPUT : data_70 
* INPUT : data_71 
* INPUT : data_72 
* INPUT : data_73 
* INPUT : data_74 
* INPUT : data_75 
* INPUT : data_76 
* INPUT : data_77 
* INPUT : data_78 
* INPUT : data_79 
* INPUT : data_80 
* INPUT : data_81 
* INPUT : data_82 
* INPUT : data_83 
* INPUT : data_84 
* INPUT : data_85 
* INPUT : data_86 
* INPUT : data_87 
* INPUT : data_88 
* INPUT : data_89 
* INPUT : data_90 
* INPUT : data_91 
* INPUT : data_92 
* INPUT : data_93 
* INPUT : data_94 
* INPUT : data_95 
* INPUT : data_96 
* INPUT : data_97 
* INPUT : data_98 
* INPUT : data_99 
* INPUT : data_100 
* INPUT : data_101 
* INPUT : data_102 
* INPUT : data_103 
* INPUT : data_104 
* INPUT : data_105 
* INPUT : data_106 
* INPUT : data_107 
* INPUT : data_108 
* INPUT : data_109 
* INPUT : data_110 
* INPUT : data_111 
* INPUT : data_112 
* INPUT : data_113 
* INPUT : data_114 
* INPUT : data_115 
* INPUT : data_116 
* INPUT : data_117 
* INPUT : data_118 
* INPUT : data_119 
* INPUT : data_120 
* INPUT : data_121 
* INPUT : data_122 
* INPUT : data_123 
* INPUT : data_124 
* INPUT : data_125 
* INPUT : data_126 
* INPUT : data_127 
* INPUT : data_128 
* INPUT : data_129 
* INPUT : data_130 
* INPUT : data_131 
* INPUT : data_132 
* INPUT : data_133 
* INPUT : data_134 
* INPUT : data_135 
* INPUT : data_136 
* INPUT : data_137 
* INPUT : data_138 
* INPUT : data_139 
* INPUT : data_140 
* INPUT : data_141 
* INPUT : data_142 
* INPUT : data_143 
* INPUT : data_144 
* INPUT : data_145 
* INPUT : data_146 
* INPUT : data_147 
* INPUT : data_148 
* INPUT : data_149 
* INPUT : data_150 
* INPUT : data_151 
* INPUT : data_152 
* INPUT : data_153 
* INPUT : data_154 
* INPUT : data_155 
* INPUT : data_156 
* INPUT : data_157 
* INPUT : data_158 
* INPUT : data_159 
* INPUT : data_160 
* INPUT : data_161 
* INPUT : data_162 
* INPUT : data_163 
* INPUT : data_164 
* INPUT : data_165 
* INPUT : data_166 
* INPUT : data_167 
* INPUT : data_168 
* INPUT : data_169 
* INPUT : data_170 
* INPUT : data_171 
* INPUT : data_172 
* INPUT : data_173 
* INPUT : data_174 
* INPUT : data_175 
* INPUT : data_176 
* INPUT : data_177 
* INPUT : data_178 
* INPUT : data_179 
* INPUT : data_180 
* INPUT : data_181 
* INPUT : data_182 
* INPUT : data_183 
* INPUT : data_184 
* INPUT : data_185 
* INPUT : data_186 
* INPUT : data_187 
* INPUT : data_188 
* INPUT : data_189 
* INPUT : data_190 
* INPUT : data_191 
* INPUT : data_192 
* INPUT : data_193 
* INPUT : data_194 
* INPUT : data_195 
* INPUT : data_196 
* INPUT : data_197 
* INPUT : data_198 
* INPUT : data_199 
* INPUT : data_200 
* INPUT : data_201 
* INPUT : data_202 
* INPUT : data_203 
* INPUT : data_204 
* INPUT : data_205 
* INPUT : data_206 
* INPUT : data_207 
* INPUT : data_208 
* INPUT : data_209 
* INPUT : data_210 
* INPUT : data_211 
* INPUT : data_212 
* INPUT : data_213 
* INPUT : data_214 
* INPUT : data_215 
* INPUT : data_216 
* INPUT : data_217 
* INPUT : data_218 
* INPUT : data_219 
* INPUT : data_220 
* INPUT : data_221 
* INPUT : data_222 
* INPUT : data_223 
* INPUT : data_224 
* INPUT : data_225 
* INPUT : data_226 
* INPUT : data_227 
* INPUT : data_228 
* INPUT : data_229 
* INPUT : data_230 
* INPUT : data_231 
* INPUT : data_232 
* INPUT : data_233 
* INPUT : data_234 
* INPUT : data_235 
* INPUT : data_236 
* INPUT : data_237 
* INPUT : data_238 
* INPUT : data_239 
* INPUT : data_240 
* INPUT : data_241 
* INPUT : data_242 
* INPUT : data_243 
* INPUT : data_244 
* INPUT : data_245 
* INPUT : data_246 
* INPUT : data_247 
* INPUT : data_248 
* INPUT : data_249 
* INPUT : data_250 
* INPUT : data_251 
* INPUT : data_252 
* INPUT : data_253 
* INPUT : data_254 
* INPUT : data_255 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 256
Xwrite_driver0 data_0 bl_0 br_0 en vdd gnd write_driver
Xwrite_driver1 data_1 bl_1 br_1 en vdd gnd write_driver
Xwrite_driver2 data_2 bl_2 br_2 en vdd gnd write_driver
Xwrite_driver3 data_3 bl_3 br_3 en vdd gnd write_driver
Xwrite_driver4 data_4 bl_4 br_4 en vdd gnd write_driver
Xwrite_driver5 data_5 bl_5 br_5 en vdd gnd write_driver
Xwrite_driver6 data_6 bl_6 br_6 en vdd gnd write_driver
Xwrite_driver7 data_7 bl_7 br_7 en vdd gnd write_driver
Xwrite_driver8 data_8 bl_8 br_8 en vdd gnd write_driver
Xwrite_driver9 data_9 bl_9 br_9 en vdd gnd write_driver
Xwrite_driver10 data_10 bl_10 br_10 en vdd gnd write_driver
Xwrite_driver11 data_11 bl_11 br_11 en vdd gnd write_driver
Xwrite_driver12 data_12 bl_12 br_12 en vdd gnd write_driver
Xwrite_driver13 data_13 bl_13 br_13 en vdd gnd write_driver
Xwrite_driver14 data_14 bl_14 br_14 en vdd gnd write_driver
Xwrite_driver15 data_15 bl_15 br_15 en vdd gnd write_driver
Xwrite_driver16 data_16 bl_16 br_16 en vdd gnd write_driver
Xwrite_driver17 data_17 bl_17 br_17 en vdd gnd write_driver
Xwrite_driver18 data_18 bl_18 br_18 en vdd gnd write_driver
Xwrite_driver19 data_19 bl_19 br_19 en vdd gnd write_driver
Xwrite_driver20 data_20 bl_20 br_20 en vdd gnd write_driver
Xwrite_driver21 data_21 bl_21 br_21 en vdd gnd write_driver
Xwrite_driver22 data_22 bl_22 br_22 en vdd gnd write_driver
Xwrite_driver23 data_23 bl_23 br_23 en vdd gnd write_driver
Xwrite_driver24 data_24 bl_24 br_24 en vdd gnd write_driver
Xwrite_driver25 data_25 bl_25 br_25 en vdd gnd write_driver
Xwrite_driver26 data_26 bl_26 br_26 en vdd gnd write_driver
Xwrite_driver27 data_27 bl_27 br_27 en vdd gnd write_driver
Xwrite_driver28 data_28 bl_28 br_28 en vdd gnd write_driver
Xwrite_driver29 data_29 bl_29 br_29 en vdd gnd write_driver
Xwrite_driver30 data_30 bl_30 br_30 en vdd gnd write_driver
Xwrite_driver31 data_31 bl_31 br_31 en vdd gnd write_driver
Xwrite_driver32 data_32 bl_32 br_32 en vdd gnd write_driver
Xwrite_driver33 data_33 bl_33 br_33 en vdd gnd write_driver
Xwrite_driver34 data_34 bl_34 br_34 en vdd gnd write_driver
Xwrite_driver35 data_35 bl_35 br_35 en vdd gnd write_driver
Xwrite_driver36 data_36 bl_36 br_36 en vdd gnd write_driver
Xwrite_driver37 data_37 bl_37 br_37 en vdd gnd write_driver
Xwrite_driver38 data_38 bl_38 br_38 en vdd gnd write_driver
Xwrite_driver39 data_39 bl_39 br_39 en vdd gnd write_driver
Xwrite_driver40 data_40 bl_40 br_40 en vdd gnd write_driver
Xwrite_driver41 data_41 bl_41 br_41 en vdd gnd write_driver
Xwrite_driver42 data_42 bl_42 br_42 en vdd gnd write_driver
Xwrite_driver43 data_43 bl_43 br_43 en vdd gnd write_driver
Xwrite_driver44 data_44 bl_44 br_44 en vdd gnd write_driver
Xwrite_driver45 data_45 bl_45 br_45 en vdd gnd write_driver
Xwrite_driver46 data_46 bl_46 br_46 en vdd gnd write_driver
Xwrite_driver47 data_47 bl_47 br_47 en vdd gnd write_driver
Xwrite_driver48 data_48 bl_48 br_48 en vdd gnd write_driver
Xwrite_driver49 data_49 bl_49 br_49 en vdd gnd write_driver
Xwrite_driver50 data_50 bl_50 br_50 en vdd gnd write_driver
Xwrite_driver51 data_51 bl_51 br_51 en vdd gnd write_driver
Xwrite_driver52 data_52 bl_52 br_52 en vdd gnd write_driver
Xwrite_driver53 data_53 bl_53 br_53 en vdd gnd write_driver
Xwrite_driver54 data_54 bl_54 br_54 en vdd gnd write_driver
Xwrite_driver55 data_55 bl_55 br_55 en vdd gnd write_driver
Xwrite_driver56 data_56 bl_56 br_56 en vdd gnd write_driver
Xwrite_driver57 data_57 bl_57 br_57 en vdd gnd write_driver
Xwrite_driver58 data_58 bl_58 br_58 en vdd gnd write_driver
Xwrite_driver59 data_59 bl_59 br_59 en vdd gnd write_driver
Xwrite_driver60 data_60 bl_60 br_60 en vdd gnd write_driver
Xwrite_driver61 data_61 bl_61 br_61 en vdd gnd write_driver
Xwrite_driver62 data_62 bl_62 br_62 en vdd gnd write_driver
Xwrite_driver63 data_63 bl_63 br_63 en vdd gnd write_driver
Xwrite_driver64 data_64 bl_64 br_64 en vdd gnd write_driver
Xwrite_driver65 data_65 bl_65 br_65 en vdd gnd write_driver
Xwrite_driver66 data_66 bl_66 br_66 en vdd gnd write_driver
Xwrite_driver67 data_67 bl_67 br_67 en vdd gnd write_driver
Xwrite_driver68 data_68 bl_68 br_68 en vdd gnd write_driver
Xwrite_driver69 data_69 bl_69 br_69 en vdd gnd write_driver
Xwrite_driver70 data_70 bl_70 br_70 en vdd gnd write_driver
Xwrite_driver71 data_71 bl_71 br_71 en vdd gnd write_driver
Xwrite_driver72 data_72 bl_72 br_72 en vdd gnd write_driver
Xwrite_driver73 data_73 bl_73 br_73 en vdd gnd write_driver
Xwrite_driver74 data_74 bl_74 br_74 en vdd gnd write_driver
Xwrite_driver75 data_75 bl_75 br_75 en vdd gnd write_driver
Xwrite_driver76 data_76 bl_76 br_76 en vdd gnd write_driver
Xwrite_driver77 data_77 bl_77 br_77 en vdd gnd write_driver
Xwrite_driver78 data_78 bl_78 br_78 en vdd gnd write_driver
Xwrite_driver79 data_79 bl_79 br_79 en vdd gnd write_driver
Xwrite_driver80 data_80 bl_80 br_80 en vdd gnd write_driver
Xwrite_driver81 data_81 bl_81 br_81 en vdd gnd write_driver
Xwrite_driver82 data_82 bl_82 br_82 en vdd gnd write_driver
Xwrite_driver83 data_83 bl_83 br_83 en vdd gnd write_driver
Xwrite_driver84 data_84 bl_84 br_84 en vdd gnd write_driver
Xwrite_driver85 data_85 bl_85 br_85 en vdd gnd write_driver
Xwrite_driver86 data_86 bl_86 br_86 en vdd gnd write_driver
Xwrite_driver87 data_87 bl_87 br_87 en vdd gnd write_driver
Xwrite_driver88 data_88 bl_88 br_88 en vdd gnd write_driver
Xwrite_driver89 data_89 bl_89 br_89 en vdd gnd write_driver
Xwrite_driver90 data_90 bl_90 br_90 en vdd gnd write_driver
Xwrite_driver91 data_91 bl_91 br_91 en vdd gnd write_driver
Xwrite_driver92 data_92 bl_92 br_92 en vdd gnd write_driver
Xwrite_driver93 data_93 bl_93 br_93 en vdd gnd write_driver
Xwrite_driver94 data_94 bl_94 br_94 en vdd gnd write_driver
Xwrite_driver95 data_95 bl_95 br_95 en vdd gnd write_driver
Xwrite_driver96 data_96 bl_96 br_96 en vdd gnd write_driver
Xwrite_driver97 data_97 bl_97 br_97 en vdd gnd write_driver
Xwrite_driver98 data_98 bl_98 br_98 en vdd gnd write_driver
Xwrite_driver99 data_99 bl_99 br_99 en vdd gnd write_driver
Xwrite_driver100 data_100 bl_100 br_100 en vdd gnd write_driver
Xwrite_driver101 data_101 bl_101 br_101 en vdd gnd write_driver
Xwrite_driver102 data_102 bl_102 br_102 en vdd gnd write_driver
Xwrite_driver103 data_103 bl_103 br_103 en vdd gnd write_driver
Xwrite_driver104 data_104 bl_104 br_104 en vdd gnd write_driver
Xwrite_driver105 data_105 bl_105 br_105 en vdd gnd write_driver
Xwrite_driver106 data_106 bl_106 br_106 en vdd gnd write_driver
Xwrite_driver107 data_107 bl_107 br_107 en vdd gnd write_driver
Xwrite_driver108 data_108 bl_108 br_108 en vdd gnd write_driver
Xwrite_driver109 data_109 bl_109 br_109 en vdd gnd write_driver
Xwrite_driver110 data_110 bl_110 br_110 en vdd gnd write_driver
Xwrite_driver111 data_111 bl_111 br_111 en vdd gnd write_driver
Xwrite_driver112 data_112 bl_112 br_112 en vdd gnd write_driver
Xwrite_driver113 data_113 bl_113 br_113 en vdd gnd write_driver
Xwrite_driver114 data_114 bl_114 br_114 en vdd gnd write_driver
Xwrite_driver115 data_115 bl_115 br_115 en vdd gnd write_driver
Xwrite_driver116 data_116 bl_116 br_116 en vdd gnd write_driver
Xwrite_driver117 data_117 bl_117 br_117 en vdd gnd write_driver
Xwrite_driver118 data_118 bl_118 br_118 en vdd gnd write_driver
Xwrite_driver119 data_119 bl_119 br_119 en vdd gnd write_driver
Xwrite_driver120 data_120 bl_120 br_120 en vdd gnd write_driver
Xwrite_driver121 data_121 bl_121 br_121 en vdd gnd write_driver
Xwrite_driver122 data_122 bl_122 br_122 en vdd gnd write_driver
Xwrite_driver123 data_123 bl_123 br_123 en vdd gnd write_driver
Xwrite_driver124 data_124 bl_124 br_124 en vdd gnd write_driver
Xwrite_driver125 data_125 bl_125 br_125 en vdd gnd write_driver
Xwrite_driver126 data_126 bl_126 br_126 en vdd gnd write_driver
Xwrite_driver127 data_127 bl_127 br_127 en vdd gnd write_driver
Xwrite_driver128 data_128 bl_128 br_128 en vdd gnd write_driver
Xwrite_driver129 data_129 bl_129 br_129 en vdd gnd write_driver
Xwrite_driver130 data_130 bl_130 br_130 en vdd gnd write_driver
Xwrite_driver131 data_131 bl_131 br_131 en vdd gnd write_driver
Xwrite_driver132 data_132 bl_132 br_132 en vdd gnd write_driver
Xwrite_driver133 data_133 bl_133 br_133 en vdd gnd write_driver
Xwrite_driver134 data_134 bl_134 br_134 en vdd gnd write_driver
Xwrite_driver135 data_135 bl_135 br_135 en vdd gnd write_driver
Xwrite_driver136 data_136 bl_136 br_136 en vdd gnd write_driver
Xwrite_driver137 data_137 bl_137 br_137 en vdd gnd write_driver
Xwrite_driver138 data_138 bl_138 br_138 en vdd gnd write_driver
Xwrite_driver139 data_139 bl_139 br_139 en vdd gnd write_driver
Xwrite_driver140 data_140 bl_140 br_140 en vdd gnd write_driver
Xwrite_driver141 data_141 bl_141 br_141 en vdd gnd write_driver
Xwrite_driver142 data_142 bl_142 br_142 en vdd gnd write_driver
Xwrite_driver143 data_143 bl_143 br_143 en vdd gnd write_driver
Xwrite_driver144 data_144 bl_144 br_144 en vdd gnd write_driver
Xwrite_driver145 data_145 bl_145 br_145 en vdd gnd write_driver
Xwrite_driver146 data_146 bl_146 br_146 en vdd gnd write_driver
Xwrite_driver147 data_147 bl_147 br_147 en vdd gnd write_driver
Xwrite_driver148 data_148 bl_148 br_148 en vdd gnd write_driver
Xwrite_driver149 data_149 bl_149 br_149 en vdd gnd write_driver
Xwrite_driver150 data_150 bl_150 br_150 en vdd gnd write_driver
Xwrite_driver151 data_151 bl_151 br_151 en vdd gnd write_driver
Xwrite_driver152 data_152 bl_152 br_152 en vdd gnd write_driver
Xwrite_driver153 data_153 bl_153 br_153 en vdd gnd write_driver
Xwrite_driver154 data_154 bl_154 br_154 en vdd gnd write_driver
Xwrite_driver155 data_155 bl_155 br_155 en vdd gnd write_driver
Xwrite_driver156 data_156 bl_156 br_156 en vdd gnd write_driver
Xwrite_driver157 data_157 bl_157 br_157 en vdd gnd write_driver
Xwrite_driver158 data_158 bl_158 br_158 en vdd gnd write_driver
Xwrite_driver159 data_159 bl_159 br_159 en vdd gnd write_driver
Xwrite_driver160 data_160 bl_160 br_160 en vdd gnd write_driver
Xwrite_driver161 data_161 bl_161 br_161 en vdd gnd write_driver
Xwrite_driver162 data_162 bl_162 br_162 en vdd gnd write_driver
Xwrite_driver163 data_163 bl_163 br_163 en vdd gnd write_driver
Xwrite_driver164 data_164 bl_164 br_164 en vdd gnd write_driver
Xwrite_driver165 data_165 bl_165 br_165 en vdd gnd write_driver
Xwrite_driver166 data_166 bl_166 br_166 en vdd gnd write_driver
Xwrite_driver167 data_167 bl_167 br_167 en vdd gnd write_driver
Xwrite_driver168 data_168 bl_168 br_168 en vdd gnd write_driver
Xwrite_driver169 data_169 bl_169 br_169 en vdd gnd write_driver
Xwrite_driver170 data_170 bl_170 br_170 en vdd gnd write_driver
Xwrite_driver171 data_171 bl_171 br_171 en vdd gnd write_driver
Xwrite_driver172 data_172 bl_172 br_172 en vdd gnd write_driver
Xwrite_driver173 data_173 bl_173 br_173 en vdd gnd write_driver
Xwrite_driver174 data_174 bl_174 br_174 en vdd gnd write_driver
Xwrite_driver175 data_175 bl_175 br_175 en vdd gnd write_driver
Xwrite_driver176 data_176 bl_176 br_176 en vdd gnd write_driver
Xwrite_driver177 data_177 bl_177 br_177 en vdd gnd write_driver
Xwrite_driver178 data_178 bl_178 br_178 en vdd gnd write_driver
Xwrite_driver179 data_179 bl_179 br_179 en vdd gnd write_driver
Xwrite_driver180 data_180 bl_180 br_180 en vdd gnd write_driver
Xwrite_driver181 data_181 bl_181 br_181 en vdd gnd write_driver
Xwrite_driver182 data_182 bl_182 br_182 en vdd gnd write_driver
Xwrite_driver183 data_183 bl_183 br_183 en vdd gnd write_driver
Xwrite_driver184 data_184 bl_184 br_184 en vdd gnd write_driver
Xwrite_driver185 data_185 bl_185 br_185 en vdd gnd write_driver
Xwrite_driver186 data_186 bl_186 br_186 en vdd gnd write_driver
Xwrite_driver187 data_187 bl_187 br_187 en vdd gnd write_driver
Xwrite_driver188 data_188 bl_188 br_188 en vdd gnd write_driver
Xwrite_driver189 data_189 bl_189 br_189 en vdd gnd write_driver
Xwrite_driver190 data_190 bl_190 br_190 en vdd gnd write_driver
Xwrite_driver191 data_191 bl_191 br_191 en vdd gnd write_driver
Xwrite_driver192 data_192 bl_192 br_192 en vdd gnd write_driver
Xwrite_driver193 data_193 bl_193 br_193 en vdd gnd write_driver
Xwrite_driver194 data_194 bl_194 br_194 en vdd gnd write_driver
Xwrite_driver195 data_195 bl_195 br_195 en vdd gnd write_driver
Xwrite_driver196 data_196 bl_196 br_196 en vdd gnd write_driver
Xwrite_driver197 data_197 bl_197 br_197 en vdd gnd write_driver
Xwrite_driver198 data_198 bl_198 br_198 en vdd gnd write_driver
Xwrite_driver199 data_199 bl_199 br_199 en vdd gnd write_driver
Xwrite_driver200 data_200 bl_200 br_200 en vdd gnd write_driver
Xwrite_driver201 data_201 bl_201 br_201 en vdd gnd write_driver
Xwrite_driver202 data_202 bl_202 br_202 en vdd gnd write_driver
Xwrite_driver203 data_203 bl_203 br_203 en vdd gnd write_driver
Xwrite_driver204 data_204 bl_204 br_204 en vdd gnd write_driver
Xwrite_driver205 data_205 bl_205 br_205 en vdd gnd write_driver
Xwrite_driver206 data_206 bl_206 br_206 en vdd gnd write_driver
Xwrite_driver207 data_207 bl_207 br_207 en vdd gnd write_driver
Xwrite_driver208 data_208 bl_208 br_208 en vdd gnd write_driver
Xwrite_driver209 data_209 bl_209 br_209 en vdd gnd write_driver
Xwrite_driver210 data_210 bl_210 br_210 en vdd gnd write_driver
Xwrite_driver211 data_211 bl_211 br_211 en vdd gnd write_driver
Xwrite_driver212 data_212 bl_212 br_212 en vdd gnd write_driver
Xwrite_driver213 data_213 bl_213 br_213 en vdd gnd write_driver
Xwrite_driver214 data_214 bl_214 br_214 en vdd gnd write_driver
Xwrite_driver215 data_215 bl_215 br_215 en vdd gnd write_driver
Xwrite_driver216 data_216 bl_216 br_216 en vdd gnd write_driver
Xwrite_driver217 data_217 bl_217 br_217 en vdd gnd write_driver
Xwrite_driver218 data_218 bl_218 br_218 en vdd gnd write_driver
Xwrite_driver219 data_219 bl_219 br_219 en vdd gnd write_driver
Xwrite_driver220 data_220 bl_220 br_220 en vdd gnd write_driver
Xwrite_driver221 data_221 bl_221 br_221 en vdd gnd write_driver
Xwrite_driver222 data_222 bl_222 br_222 en vdd gnd write_driver
Xwrite_driver223 data_223 bl_223 br_223 en vdd gnd write_driver
Xwrite_driver224 data_224 bl_224 br_224 en vdd gnd write_driver
Xwrite_driver225 data_225 bl_225 br_225 en vdd gnd write_driver
Xwrite_driver226 data_226 bl_226 br_226 en vdd gnd write_driver
Xwrite_driver227 data_227 bl_227 br_227 en vdd gnd write_driver
Xwrite_driver228 data_228 bl_228 br_228 en vdd gnd write_driver
Xwrite_driver229 data_229 bl_229 br_229 en vdd gnd write_driver
Xwrite_driver230 data_230 bl_230 br_230 en vdd gnd write_driver
Xwrite_driver231 data_231 bl_231 br_231 en vdd gnd write_driver
Xwrite_driver232 data_232 bl_232 br_232 en vdd gnd write_driver
Xwrite_driver233 data_233 bl_233 br_233 en vdd gnd write_driver
Xwrite_driver234 data_234 bl_234 br_234 en vdd gnd write_driver
Xwrite_driver235 data_235 bl_235 br_235 en vdd gnd write_driver
Xwrite_driver236 data_236 bl_236 br_236 en vdd gnd write_driver
Xwrite_driver237 data_237 bl_237 br_237 en vdd gnd write_driver
Xwrite_driver238 data_238 bl_238 br_238 en vdd gnd write_driver
Xwrite_driver239 data_239 bl_239 br_239 en vdd gnd write_driver
Xwrite_driver240 data_240 bl_240 br_240 en vdd gnd write_driver
Xwrite_driver241 data_241 bl_241 br_241 en vdd gnd write_driver
Xwrite_driver242 data_242 bl_242 br_242 en vdd gnd write_driver
Xwrite_driver243 data_243 bl_243 br_243 en vdd gnd write_driver
Xwrite_driver244 data_244 bl_244 br_244 en vdd gnd write_driver
Xwrite_driver245 data_245 bl_245 br_245 en vdd gnd write_driver
Xwrite_driver246 data_246 bl_246 br_246 en vdd gnd write_driver
Xwrite_driver247 data_247 bl_247 br_247 en vdd gnd write_driver
Xwrite_driver248 data_248 bl_248 br_248 en vdd gnd write_driver
Xwrite_driver249 data_249 bl_249 br_249 en vdd gnd write_driver
Xwrite_driver250 data_250 bl_250 br_250 en vdd gnd write_driver
Xwrite_driver251 data_251 bl_251 br_251 en vdd gnd write_driver
Xwrite_driver252 data_252 bl_252 br_252 en vdd gnd write_driver
Xwrite_driver253 data_253 bl_253 br_253 en vdd gnd write_driver
Xwrite_driver254 data_254 bl_254 br_254 en vdd gnd write_driver
Xwrite_driver255 data_255 bl_255 br_255 en vdd gnd write_driver
.ENDS write_driver_array_0

.SUBCKT port_data_0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38 dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46 dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54 dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62 dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70 dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78 dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86 dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94 dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102 dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109 dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116 dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123 dout_124 dout_125 dout_126 dout_127 dout_128 dout_129 dout_130 dout_131 dout_132 dout_133 dout_134 dout_135 dout_136 dout_137 dout_138 dout_139 dout_140 dout_141 dout_142 dout_143 dout_144 dout_145 dout_146 dout_147 dout_148 dout_149 dout_150 dout_151 dout_152 dout_153 dout_154 dout_155 dout_156 dout_157 dout_158 dout_159 dout_160 dout_161 dout_162 dout_163 dout_164 dout_165 dout_166 dout_167 dout_168 dout_169 dout_170 dout_171 dout_172 dout_173 dout_174 dout_175 dout_176 dout_177 dout_178 dout_179 dout_180 dout_181 dout_182 dout_183 dout_184 dout_185 dout_186 dout_187 dout_188 dout_189 dout_190 dout_191 dout_192 dout_193 dout_194 dout_195 dout_196 dout_197 dout_198 dout_199 dout_200 dout_201 dout_202 dout_203 dout_204 dout_205 dout_206 dout_207 dout_208 dout_209 dout_210 dout_211 dout_212 dout_213 dout_214 dout_215 dout_216 dout_217 dout_218 dout_219 dout_220 dout_221 dout_222 dout_223 dout_224 dout_225 dout_226 dout_227 dout_228 dout_229 dout_230 dout_231 dout_232 dout_233 dout_234 dout_235 dout_236 dout_237 dout_238 dout_239 dout_240 dout_241 dout_242 dout_243 dout_244 dout_245 dout_246 dout_247 dout_248 dout_249 dout_250 dout_251 dout_252 dout_253 dout_254 dout_255 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 din_128 din_129 din_130 din_131 din_132 din_133 din_134 din_135 din_136 din_137 din_138 din_139 din_140 din_141 din_142 din_143 din_144 din_145 din_146 din_147 din_148 din_149 din_150 din_151 din_152 din_153 din_154 din_155 din_156 din_157 din_158 din_159 din_160 din_161 din_162 din_163 din_164 din_165 din_166 din_167 din_168 din_169 din_170 din_171 din_172 din_173 din_174 din_175 din_176 din_177 din_178 din_179 din_180 din_181 din_182 din_183 din_184 din_185 din_186 din_187 din_188 din_189 din_190 din_191 din_192 din_193 din_194 din_195 din_196 din_197 din_198 din_199 din_200 din_201 din_202 din_203 din_204 din_205 din_206 din_207 din_208 din_209 din_210 din_211 din_212 din_213 din_214 din_215 din_216 din_217 din_218 din_219 din_220 din_221 din_222 din_223 din_224 din_225 din_226 din_227 din_228 din_229 din_230 din_231 din_232 din_233 din_234 din_235 din_236 din_237 din_238 din_239 din_240 din_241 din_242 din_243 din_244 din_245 din_246 din_247 din_248 din_249 din_250 din_251 din_252 din_253 din_254 din_255 s_en p_en_bar w_en vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* OUTPUT: dout_128 
* OUTPUT: dout_129 
* OUTPUT: dout_130 
* OUTPUT: dout_131 
* OUTPUT: dout_132 
* OUTPUT: dout_133 
* OUTPUT: dout_134 
* OUTPUT: dout_135 
* OUTPUT: dout_136 
* OUTPUT: dout_137 
* OUTPUT: dout_138 
* OUTPUT: dout_139 
* OUTPUT: dout_140 
* OUTPUT: dout_141 
* OUTPUT: dout_142 
* OUTPUT: dout_143 
* OUTPUT: dout_144 
* OUTPUT: dout_145 
* OUTPUT: dout_146 
* OUTPUT: dout_147 
* OUTPUT: dout_148 
* OUTPUT: dout_149 
* OUTPUT: dout_150 
* OUTPUT: dout_151 
* OUTPUT: dout_152 
* OUTPUT: dout_153 
* OUTPUT: dout_154 
* OUTPUT: dout_155 
* OUTPUT: dout_156 
* OUTPUT: dout_157 
* OUTPUT: dout_158 
* OUTPUT: dout_159 
* OUTPUT: dout_160 
* OUTPUT: dout_161 
* OUTPUT: dout_162 
* OUTPUT: dout_163 
* OUTPUT: dout_164 
* OUTPUT: dout_165 
* OUTPUT: dout_166 
* OUTPUT: dout_167 
* OUTPUT: dout_168 
* OUTPUT: dout_169 
* OUTPUT: dout_170 
* OUTPUT: dout_171 
* OUTPUT: dout_172 
* OUTPUT: dout_173 
* OUTPUT: dout_174 
* OUTPUT: dout_175 
* OUTPUT: dout_176 
* OUTPUT: dout_177 
* OUTPUT: dout_178 
* OUTPUT: dout_179 
* OUTPUT: dout_180 
* OUTPUT: dout_181 
* OUTPUT: dout_182 
* OUTPUT: dout_183 
* OUTPUT: dout_184 
* OUTPUT: dout_185 
* OUTPUT: dout_186 
* OUTPUT: dout_187 
* OUTPUT: dout_188 
* OUTPUT: dout_189 
* OUTPUT: dout_190 
* OUTPUT: dout_191 
* OUTPUT: dout_192 
* OUTPUT: dout_193 
* OUTPUT: dout_194 
* OUTPUT: dout_195 
* OUTPUT: dout_196 
* OUTPUT: dout_197 
* OUTPUT: dout_198 
* OUTPUT: dout_199 
* OUTPUT: dout_200 
* OUTPUT: dout_201 
* OUTPUT: dout_202 
* OUTPUT: dout_203 
* OUTPUT: dout_204 
* OUTPUT: dout_205 
* OUTPUT: dout_206 
* OUTPUT: dout_207 
* OUTPUT: dout_208 
* OUTPUT: dout_209 
* OUTPUT: dout_210 
* OUTPUT: dout_211 
* OUTPUT: dout_212 
* OUTPUT: dout_213 
* OUTPUT: dout_214 
* OUTPUT: dout_215 
* OUTPUT: dout_216 
* OUTPUT: dout_217 
* OUTPUT: dout_218 
* OUTPUT: dout_219 
* OUTPUT: dout_220 
* OUTPUT: dout_221 
* OUTPUT: dout_222 
* OUTPUT: dout_223 
* OUTPUT: dout_224 
* OUTPUT: dout_225 
* OUTPUT: dout_226 
* OUTPUT: dout_227 
* OUTPUT: dout_228 
* OUTPUT: dout_229 
* OUTPUT: dout_230 
* OUTPUT: dout_231 
* OUTPUT: dout_232 
* OUTPUT: dout_233 
* OUTPUT: dout_234 
* OUTPUT: dout_235 
* OUTPUT: dout_236 
* OUTPUT: dout_237 
* OUTPUT: dout_238 
* OUTPUT: dout_239 
* OUTPUT: dout_240 
* OUTPUT: dout_241 
* OUTPUT: dout_242 
* OUTPUT: dout_243 
* OUTPUT: dout_244 
* OUTPUT: dout_245 
* OUTPUT: dout_246 
* OUTPUT: dout_247 
* OUTPUT: dout_248 
* OUTPUT: dout_249 
* OUTPUT: dout_250 
* OUTPUT: dout_251 
* OUTPUT: dout_252 
* OUTPUT: dout_253 
* OUTPUT: dout_254 
* OUTPUT: dout_255 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* INPUT : din_128 
* INPUT : din_129 
* INPUT : din_130 
* INPUT : din_131 
* INPUT : din_132 
* INPUT : din_133 
* INPUT : din_134 
* INPUT : din_135 
* INPUT : din_136 
* INPUT : din_137 
* INPUT : din_138 
* INPUT : din_139 
* INPUT : din_140 
* INPUT : din_141 
* INPUT : din_142 
* INPUT : din_143 
* INPUT : din_144 
* INPUT : din_145 
* INPUT : din_146 
* INPUT : din_147 
* INPUT : din_148 
* INPUT : din_149 
* INPUT : din_150 
* INPUT : din_151 
* INPUT : din_152 
* INPUT : din_153 
* INPUT : din_154 
* INPUT : din_155 
* INPUT : din_156 
* INPUT : din_157 
* INPUT : din_158 
* INPUT : din_159 
* INPUT : din_160 
* INPUT : din_161 
* INPUT : din_162 
* INPUT : din_163 
* INPUT : din_164 
* INPUT : din_165 
* INPUT : din_166 
* INPUT : din_167 
* INPUT : din_168 
* INPUT : din_169 
* INPUT : din_170 
* INPUT : din_171 
* INPUT : din_172 
* INPUT : din_173 
* INPUT : din_174 
* INPUT : din_175 
* INPUT : din_176 
* INPUT : din_177 
* INPUT : din_178 
* INPUT : din_179 
* INPUT : din_180 
* INPUT : din_181 
* INPUT : din_182 
* INPUT : din_183 
* INPUT : din_184 
* INPUT : din_185 
* INPUT : din_186 
* INPUT : din_187 
* INPUT : din_188 
* INPUT : din_189 
* INPUT : din_190 
* INPUT : din_191 
* INPUT : din_192 
* INPUT : din_193 
* INPUT : din_194 
* INPUT : din_195 
* INPUT : din_196 
* INPUT : din_197 
* INPUT : din_198 
* INPUT : din_199 
* INPUT : din_200 
* INPUT : din_201 
* INPUT : din_202 
* INPUT : din_203 
* INPUT : din_204 
* INPUT : din_205 
* INPUT : din_206 
* INPUT : din_207 
* INPUT : din_208 
* INPUT : din_209 
* INPUT : din_210 
* INPUT : din_211 
* INPUT : din_212 
* INPUT : din_213 
* INPUT : din_214 
* INPUT : din_215 
* INPUT : din_216 
* INPUT : din_217 
* INPUT : din_218 
* INPUT : din_219 
* INPUT : din_220 
* INPUT : din_221 
* INPUT : din_222 
* INPUT : din_223 
* INPUT : din_224 
* INPUT : din_225 
* INPUT : din_226 
* INPUT : din_227 
* INPUT : din_228 
* INPUT : din_229 
* INPUT : din_230 
* INPUT : din_231 
* INPUT : din_232 
* INPUT : din_233 
* INPUT : din_234 
* INPUT : din_235 
* INPUT : din_236 
* INPUT : din_237 
* INPUT : din_238 
* INPUT : din_239 
* INPUT : din_240 
* INPUT : din_241 
* INPUT : din_242 
* INPUT : din_243 
* INPUT : din_244 
* INPUT : din_245 
* INPUT : din_246 
* INPUT : din_247 
* INPUT : din_248 
* INPUT : din_249 
* INPUT : din_250 
* INPUT : din_251 
* INPUT : din_252 
* INPUT : din_253 
* INPUT : din_254 
* INPUT : din_255 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 p_en_bar vdd precharge_array_0
Xsense_amp_array0 dout_0 bl_0 br_0 dout_1 bl_1 br_1 dout_2 bl_2 br_2 dout_3 bl_3 br_3 dout_4 bl_4 br_4 dout_5 bl_5 br_5 dout_6 bl_6 br_6 dout_7 bl_7 br_7 dout_8 bl_8 br_8 dout_9 bl_9 br_9 dout_10 bl_10 br_10 dout_11 bl_11 br_11 dout_12 bl_12 br_12 dout_13 bl_13 br_13 dout_14 bl_14 br_14 dout_15 bl_15 br_15 dout_16 bl_16 br_16 dout_17 bl_17 br_17 dout_18 bl_18 br_18 dout_19 bl_19 br_19 dout_20 bl_20 br_20 dout_21 bl_21 br_21 dout_22 bl_22 br_22 dout_23 bl_23 br_23 dout_24 bl_24 br_24 dout_25 bl_25 br_25 dout_26 bl_26 br_26 dout_27 bl_27 br_27 dout_28 bl_28 br_28 dout_29 bl_29 br_29 dout_30 bl_30 br_30 dout_31 bl_31 br_31 dout_32 bl_32 br_32 dout_33 bl_33 br_33 dout_34 bl_34 br_34 dout_35 bl_35 br_35 dout_36 bl_36 br_36 dout_37 bl_37 br_37 dout_38 bl_38 br_38 dout_39 bl_39 br_39 dout_40 bl_40 br_40 dout_41 bl_41 br_41 dout_42 bl_42 br_42 dout_43 bl_43 br_43 dout_44 bl_44 br_44 dout_45 bl_45 br_45 dout_46 bl_46 br_46 dout_47 bl_47 br_47 dout_48 bl_48 br_48 dout_49 bl_49 br_49 dout_50 bl_50 br_50 dout_51 bl_51 br_51 dout_52 bl_52 br_52 dout_53 bl_53 br_53 dout_54 bl_54 br_54 dout_55 bl_55 br_55 dout_56 bl_56 br_56 dout_57 bl_57 br_57 dout_58 bl_58 br_58 dout_59 bl_59 br_59 dout_60 bl_60 br_60 dout_61 bl_61 br_61 dout_62 bl_62 br_62 dout_63 bl_63 br_63 dout_64 bl_64 br_64 dout_65 bl_65 br_65 dout_66 bl_66 br_66 dout_67 bl_67 br_67 dout_68 bl_68 br_68 dout_69 bl_69 br_69 dout_70 bl_70 br_70 dout_71 bl_71 br_71 dout_72 bl_72 br_72 dout_73 bl_73 br_73 dout_74 bl_74 br_74 dout_75 bl_75 br_75 dout_76 bl_76 br_76 dout_77 bl_77 br_77 dout_78 bl_78 br_78 dout_79 bl_79 br_79 dout_80 bl_80 br_80 dout_81 bl_81 br_81 dout_82 bl_82 br_82 dout_83 bl_83 br_83 dout_84 bl_84 br_84 dout_85 bl_85 br_85 dout_86 bl_86 br_86 dout_87 bl_87 br_87 dout_88 bl_88 br_88 dout_89 bl_89 br_89 dout_90 bl_90 br_90 dout_91 bl_91 br_91 dout_92 bl_92 br_92 dout_93 bl_93 br_93 dout_94 bl_94 br_94 dout_95 bl_95 br_95 dout_96 bl_96 br_96 dout_97 bl_97 br_97 dout_98 bl_98 br_98 dout_99 bl_99 br_99 dout_100 bl_100 br_100 dout_101 bl_101 br_101 dout_102 bl_102 br_102 dout_103 bl_103 br_103 dout_104 bl_104 br_104 dout_105 bl_105 br_105 dout_106 bl_106 br_106 dout_107 bl_107 br_107 dout_108 bl_108 br_108 dout_109 bl_109 br_109 dout_110 bl_110 br_110 dout_111 bl_111 br_111 dout_112 bl_112 br_112 dout_113 bl_113 br_113 dout_114 bl_114 br_114 dout_115 bl_115 br_115 dout_116 bl_116 br_116 dout_117 bl_117 br_117 dout_118 bl_118 br_118 dout_119 bl_119 br_119 dout_120 bl_120 br_120 dout_121 bl_121 br_121 dout_122 bl_122 br_122 dout_123 bl_123 br_123 dout_124 bl_124 br_124 dout_125 bl_125 br_125 dout_126 bl_126 br_126 dout_127 bl_127 br_127 dout_128 bl_128 br_128 dout_129 bl_129 br_129 dout_130 bl_130 br_130 dout_131 bl_131 br_131 dout_132 bl_132 br_132 dout_133 bl_133 br_133 dout_134 bl_134 br_134 dout_135 bl_135 br_135 dout_136 bl_136 br_136 dout_137 bl_137 br_137 dout_138 bl_138 br_138 dout_139 bl_139 br_139 dout_140 bl_140 br_140 dout_141 bl_141 br_141 dout_142 bl_142 br_142 dout_143 bl_143 br_143 dout_144 bl_144 br_144 dout_145 bl_145 br_145 dout_146 bl_146 br_146 dout_147 bl_147 br_147 dout_148 bl_148 br_148 dout_149 bl_149 br_149 dout_150 bl_150 br_150 dout_151 bl_151 br_151 dout_152 bl_152 br_152 dout_153 bl_153 br_153 dout_154 bl_154 br_154 dout_155 bl_155 br_155 dout_156 bl_156 br_156 dout_157 bl_157 br_157 dout_158 bl_158 br_158 dout_159 bl_159 br_159 dout_160 bl_160 br_160 dout_161 bl_161 br_161 dout_162 bl_162 br_162 dout_163 bl_163 br_163 dout_164 bl_164 br_164 dout_165 bl_165 br_165 dout_166 bl_166 br_166 dout_167 bl_167 br_167 dout_168 bl_168 br_168 dout_169 bl_169 br_169 dout_170 bl_170 br_170 dout_171 bl_171 br_171 dout_172 bl_172 br_172 dout_173 bl_173 br_173 dout_174 bl_174 br_174 dout_175 bl_175 br_175 dout_176 bl_176 br_176 dout_177 bl_177 br_177 dout_178 bl_178 br_178 dout_179 bl_179 br_179 dout_180 bl_180 br_180 dout_181 bl_181 br_181 dout_182 bl_182 br_182 dout_183 bl_183 br_183 dout_184 bl_184 br_184 dout_185 bl_185 br_185 dout_186 bl_186 br_186 dout_187 bl_187 br_187 dout_188 bl_188 br_188 dout_189 bl_189 br_189 dout_190 bl_190 br_190 dout_191 bl_191 br_191 dout_192 bl_192 br_192 dout_193 bl_193 br_193 dout_194 bl_194 br_194 dout_195 bl_195 br_195 dout_196 bl_196 br_196 dout_197 bl_197 br_197 dout_198 bl_198 br_198 dout_199 bl_199 br_199 dout_200 bl_200 br_200 dout_201 bl_201 br_201 dout_202 bl_202 br_202 dout_203 bl_203 br_203 dout_204 bl_204 br_204 dout_205 bl_205 br_205 dout_206 bl_206 br_206 dout_207 bl_207 br_207 dout_208 bl_208 br_208 dout_209 bl_209 br_209 dout_210 bl_210 br_210 dout_211 bl_211 br_211 dout_212 bl_212 br_212 dout_213 bl_213 br_213 dout_214 bl_214 br_214 dout_215 bl_215 br_215 dout_216 bl_216 br_216 dout_217 bl_217 br_217 dout_218 bl_218 br_218 dout_219 bl_219 br_219 dout_220 bl_220 br_220 dout_221 bl_221 br_221 dout_222 bl_222 br_222 dout_223 bl_223 br_223 dout_224 bl_224 br_224 dout_225 bl_225 br_225 dout_226 bl_226 br_226 dout_227 bl_227 br_227 dout_228 bl_228 br_228 dout_229 bl_229 br_229 dout_230 bl_230 br_230 dout_231 bl_231 br_231 dout_232 bl_232 br_232 dout_233 bl_233 br_233 dout_234 bl_234 br_234 dout_235 bl_235 br_235 dout_236 bl_236 br_236 dout_237 bl_237 br_237 dout_238 bl_238 br_238 dout_239 bl_239 br_239 dout_240 bl_240 br_240 dout_241 bl_241 br_241 dout_242 bl_242 br_242 dout_243 bl_243 br_243 dout_244 bl_244 br_244 dout_245 bl_245 br_245 dout_246 bl_246 br_246 dout_247 bl_247 br_247 dout_248 bl_248 br_248 dout_249 bl_249 br_249 dout_250 bl_250 br_250 dout_251 bl_251 br_251 dout_252 bl_252 br_252 dout_253 bl_253 br_253 dout_254 bl_254 br_254 dout_255 bl_255 br_255 s_en vdd gnd sense_amp_array_0
Xwrite_driver_array0 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 din_128 din_129 din_130 din_131 din_132 din_133 din_134 din_135 din_136 din_137 din_138 din_139 din_140 din_141 din_142 din_143 din_144 din_145 din_146 din_147 din_148 din_149 din_150 din_151 din_152 din_153 din_154 din_155 din_156 din_157 din_158 din_159 din_160 din_161 din_162 din_163 din_164 din_165 din_166 din_167 din_168 din_169 din_170 din_171 din_172 din_173 din_174 din_175 din_176 din_177 din_178 din_179 din_180 din_181 din_182 din_183 din_184 din_185 din_186 din_187 din_188 din_189 din_190 din_191 din_192 din_193 din_194 din_195 din_196 din_197 din_198 din_199 din_200 din_201 din_202 din_203 din_204 din_205 din_206 din_207 din_208 din_209 din_210 din_211 din_212 din_213 din_214 din_215 din_216 din_217 din_218 din_219 din_220 din_221 din_222 din_223 din_224 din_225 din_226 din_227 din_228 din_229 din_230 din_231 din_232 din_233 din_234 din_235 din_236 din_237 din_238 din_239 din_240 din_241 din_242 din_243 din_244 din_245 din_246 din_247 din_248 din_249 din_250 din_251 din_252 din_253 din_254 din_255 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 w_en vdd gnd write_driver_array_0
.ENDS port_data_0

* ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_0

* ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT pnand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_0

.SUBCKT pnand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_0

.SUBCKT hierarchical_predecode2x4_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
XXpre2x4_nand_0 inbar_0 inbar_1 Z_0 vdd gnd pnand2_0
XXpre2x4_nand_1 in_0 inbar_1 Z_1 vdd gnd pnand2_0
XXpre2x4_nand_2 inbar_0 in_1 Z_2 vdd gnd pnand2_0
XXpre2x4_nand_3 in_0 in_1 Z_3 vdd gnd pnand2_0
.ENDS hierarchical_predecode2x4_0

.SUBCKT hierarchical_predecode3x8_0 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
Xpre_nand_inv_4 Z_4 out_4 vdd gnd pinv_0
Xpre_nand_inv_5 Z_5 out_5 vdd gnd pinv_0
Xpre_nand_inv_6 Z_6 out_6 vdd gnd pinv_0
Xpre_nand_inv_7 Z_7 out_7 vdd gnd pinv_0
XXpre3x8_nand_0 inbar_0 inbar_1 inbar_2 Z_0 vdd gnd pnand3_0
XXpre3x8_nand_1 in_0 inbar_1 inbar_2 Z_1 vdd gnd pnand3_0
XXpre3x8_nand_2 inbar_0 in_1 inbar_2 Z_2 vdd gnd pnand3_0
XXpre3x8_nand_3 in_0 in_1 inbar_2 Z_3 vdd gnd pnand3_0
XXpre3x8_nand_4 inbar_0 inbar_1 in_2 Z_4 vdd gnd pnand3_0
XXpre3x8_nand_5 in_0 inbar_1 in_2 Z_5 vdd gnd pnand3_0
XXpre3x8_nand_6 inbar_0 in_1 in_2 Z_6 vdd gnd pnand3_0
XXpre3x8_nand_7 in_0 in_1 in_2 Z_7 vdd gnd pnand3_0
.ENDS hierarchical_predecode3x8_0

.SUBCKT hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 decode_0 decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* POWER : vdd 
* GROUND: gnd 
Xpre_0 addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd hierarchical_predecode2x4_0
Xpre_1 addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd hierarchical_predecode2x4_0
Xpre_2 addr_4 addr_5 out_8 out_9 out_10 out_11 vdd gnd hierarchical_predecode2x4_0
XDEC_NAND_0 out_0 out_4 out_8 Z_0 vdd gnd pnand3_0
XDEC_NAND_16 out_0 out_4 out_9 Z_16 vdd gnd pnand3_0
XDEC_NAND_32 out_0 out_4 out_10 Z_32 vdd gnd pnand3_0
XDEC_NAND_48 out_0 out_4 out_11 Z_48 vdd gnd pnand3_0
XDEC_NAND_4 out_0 out_5 out_8 Z_4 vdd gnd pnand3_0
XDEC_NAND_20 out_0 out_5 out_9 Z_20 vdd gnd pnand3_0
XDEC_NAND_36 out_0 out_5 out_10 Z_36 vdd gnd pnand3_0
XDEC_NAND_52 out_0 out_5 out_11 Z_52 vdd gnd pnand3_0
XDEC_NAND_8 out_0 out_6 out_8 Z_8 vdd gnd pnand3_0
XDEC_NAND_24 out_0 out_6 out_9 Z_24 vdd gnd pnand3_0
XDEC_NAND_40 out_0 out_6 out_10 Z_40 vdd gnd pnand3_0
XDEC_NAND_56 out_0 out_6 out_11 Z_56 vdd gnd pnand3_0
XDEC_NAND_12 out_0 out_7 out_8 Z_12 vdd gnd pnand3_0
XDEC_NAND_28 out_0 out_7 out_9 Z_28 vdd gnd pnand3_0
XDEC_NAND_44 out_0 out_7 out_10 Z_44 vdd gnd pnand3_0
XDEC_NAND_60 out_0 out_7 out_11 Z_60 vdd gnd pnand3_0
XDEC_NAND_1 out_1 out_4 out_8 Z_1 vdd gnd pnand3_0
XDEC_NAND_17 out_1 out_4 out_9 Z_17 vdd gnd pnand3_0
XDEC_NAND_33 out_1 out_4 out_10 Z_33 vdd gnd pnand3_0
XDEC_NAND_49 out_1 out_4 out_11 Z_49 vdd gnd pnand3_0
XDEC_NAND_5 out_1 out_5 out_8 Z_5 vdd gnd pnand3_0
XDEC_NAND_21 out_1 out_5 out_9 Z_21 vdd gnd pnand3_0
XDEC_NAND_37 out_1 out_5 out_10 Z_37 vdd gnd pnand3_0
XDEC_NAND_53 out_1 out_5 out_11 Z_53 vdd gnd pnand3_0
XDEC_NAND_9 out_1 out_6 out_8 Z_9 vdd gnd pnand3_0
XDEC_NAND_25 out_1 out_6 out_9 Z_25 vdd gnd pnand3_0
XDEC_NAND_41 out_1 out_6 out_10 Z_41 vdd gnd pnand3_0
XDEC_NAND_57 out_1 out_6 out_11 Z_57 vdd gnd pnand3_0
XDEC_NAND_13 out_1 out_7 out_8 Z_13 vdd gnd pnand3_0
XDEC_NAND_29 out_1 out_7 out_9 Z_29 vdd gnd pnand3_0
XDEC_NAND_45 out_1 out_7 out_10 Z_45 vdd gnd pnand3_0
XDEC_NAND_61 out_1 out_7 out_11 Z_61 vdd gnd pnand3_0
XDEC_NAND_2 out_2 out_4 out_8 Z_2 vdd gnd pnand3_0
XDEC_NAND_18 out_2 out_4 out_9 Z_18 vdd gnd pnand3_0
XDEC_NAND_34 out_2 out_4 out_10 Z_34 vdd gnd pnand3_0
XDEC_NAND_50 out_2 out_4 out_11 Z_50 vdd gnd pnand3_0
XDEC_NAND_6 out_2 out_5 out_8 Z_6 vdd gnd pnand3_0
XDEC_NAND_22 out_2 out_5 out_9 Z_22 vdd gnd pnand3_0
XDEC_NAND_38 out_2 out_5 out_10 Z_38 vdd gnd pnand3_0
XDEC_NAND_54 out_2 out_5 out_11 Z_54 vdd gnd pnand3_0
XDEC_NAND_10 out_2 out_6 out_8 Z_10 vdd gnd pnand3_0
XDEC_NAND_26 out_2 out_6 out_9 Z_26 vdd gnd pnand3_0
XDEC_NAND_42 out_2 out_6 out_10 Z_42 vdd gnd pnand3_0
XDEC_NAND_58 out_2 out_6 out_11 Z_58 vdd gnd pnand3_0
XDEC_NAND_14 out_2 out_7 out_8 Z_14 vdd gnd pnand3_0
XDEC_NAND_30 out_2 out_7 out_9 Z_30 vdd gnd pnand3_0
XDEC_NAND_46 out_2 out_7 out_10 Z_46 vdd gnd pnand3_0
XDEC_NAND_62 out_2 out_7 out_11 Z_62 vdd gnd pnand3_0
XDEC_NAND_3 out_3 out_4 out_8 Z_3 vdd gnd pnand3_0
XDEC_NAND_19 out_3 out_4 out_9 Z_19 vdd gnd pnand3_0
XDEC_NAND_35 out_3 out_4 out_10 Z_35 vdd gnd pnand3_0
XDEC_NAND_51 out_3 out_4 out_11 Z_51 vdd gnd pnand3_0
XDEC_NAND_7 out_3 out_5 out_8 Z_7 vdd gnd pnand3_0
XDEC_NAND_23 out_3 out_5 out_9 Z_23 vdd gnd pnand3_0
XDEC_NAND_39 out_3 out_5 out_10 Z_39 vdd gnd pnand3_0
XDEC_NAND_55 out_3 out_5 out_11 Z_55 vdd gnd pnand3_0
XDEC_NAND_11 out_3 out_6 out_8 Z_11 vdd gnd pnand3_0
XDEC_NAND_27 out_3 out_6 out_9 Z_27 vdd gnd pnand3_0
XDEC_NAND_43 out_3 out_6 out_10 Z_43 vdd gnd pnand3_0
XDEC_NAND_59 out_3 out_6 out_11 Z_59 vdd gnd pnand3_0
XDEC_NAND_15 out_3 out_7 out_8 Z_15 vdd gnd pnand3_0
XDEC_NAND_31 out_3 out_7 out_9 Z_31 vdd gnd pnand3_0
XDEC_NAND_47 out_3 out_7 out_10 Z_47 vdd gnd pnand3_0
XDEC_NAND_63 out_3 out_7 out_11 Z_63 vdd gnd pnand3_0
XDEC_INV_0 Z_0 decode_0 vdd gnd pinv_0
XDEC_INV_1 Z_1 decode_1 vdd gnd pinv_0
XDEC_INV_2 Z_2 decode_2 vdd gnd pinv_0
XDEC_INV_3 Z_3 decode_3 vdd gnd pinv_0
XDEC_INV_4 Z_4 decode_4 vdd gnd pinv_0
XDEC_INV_5 Z_5 decode_5 vdd gnd pinv_0
XDEC_INV_6 Z_6 decode_6 vdd gnd pinv_0
XDEC_INV_7 Z_7 decode_7 vdd gnd pinv_0
XDEC_INV_8 Z_8 decode_8 vdd gnd pinv_0
XDEC_INV_9 Z_9 decode_9 vdd gnd pinv_0
XDEC_INV_10 Z_10 decode_10 vdd gnd pinv_0
XDEC_INV_11 Z_11 decode_11 vdd gnd pinv_0
XDEC_INV_12 Z_12 decode_12 vdd gnd pinv_0
XDEC_INV_13 Z_13 decode_13 vdd gnd pinv_0
XDEC_INV_14 Z_14 decode_14 vdd gnd pinv_0
XDEC_INV_15 Z_15 decode_15 vdd gnd pinv_0
XDEC_INV_16 Z_16 decode_16 vdd gnd pinv_0
XDEC_INV_17 Z_17 decode_17 vdd gnd pinv_0
XDEC_INV_18 Z_18 decode_18 vdd gnd pinv_0
XDEC_INV_19 Z_19 decode_19 vdd gnd pinv_0
XDEC_INV_20 Z_20 decode_20 vdd gnd pinv_0
XDEC_INV_21 Z_21 decode_21 vdd gnd pinv_0
XDEC_INV_22 Z_22 decode_22 vdd gnd pinv_0
XDEC_INV_23 Z_23 decode_23 vdd gnd pinv_0
XDEC_INV_24 Z_24 decode_24 vdd gnd pinv_0
XDEC_INV_25 Z_25 decode_25 vdd gnd pinv_0
XDEC_INV_26 Z_26 decode_26 vdd gnd pinv_0
XDEC_INV_27 Z_27 decode_27 vdd gnd pinv_0
XDEC_INV_28 Z_28 decode_28 vdd gnd pinv_0
XDEC_INV_29 Z_29 decode_29 vdd gnd pinv_0
XDEC_INV_30 Z_30 decode_30 vdd gnd pinv_0
XDEC_INV_31 Z_31 decode_31 vdd gnd pinv_0
XDEC_INV_32 Z_32 decode_32 vdd gnd pinv_0
XDEC_INV_33 Z_33 decode_33 vdd gnd pinv_0
XDEC_INV_34 Z_34 decode_34 vdd gnd pinv_0
XDEC_INV_35 Z_35 decode_35 vdd gnd pinv_0
XDEC_INV_36 Z_36 decode_36 vdd gnd pinv_0
XDEC_INV_37 Z_37 decode_37 vdd gnd pinv_0
XDEC_INV_38 Z_38 decode_38 vdd gnd pinv_0
XDEC_INV_39 Z_39 decode_39 vdd gnd pinv_0
XDEC_INV_40 Z_40 decode_40 vdd gnd pinv_0
XDEC_INV_41 Z_41 decode_41 vdd gnd pinv_0
XDEC_INV_42 Z_42 decode_42 vdd gnd pinv_0
XDEC_INV_43 Z_43 decode_43 vdd gnd pinv_0
XDEC_INV_44 Z_44 decode_44 vdd gnd pinv_0
XDEC_INV_45 Z_45 decode_45 vdd gnd pinv_0
XDEC_INV_46 Z_46 decode_46 vdd gnd pinv_0
XDEC_INV_47 Z_47 decode_47 vdd gnd pinv_0
XDEC_INV_48 Z_48 decode_48 vdd gnd pinv_0
XDEC_INV_49 Z_49 decode_49 vdd gnd pinv_0
XDEC_INV_50 Z_50 decode_50 vdd gnd pinv_0
XDEC_INV_51 Z_51 decode_51 vdd gnd pinv_0
XDEC_INV_52 Z_52 decode_52 vdd gnd pinv_0
XDEC_INV_53 Z_53 decode_53 vdd gnd pinv_0
XDEC_INV_54 Z_54 decode_54 vdd gnd pinv_0
XDEC_INV_55 Z_55 decode_55 vdd gnd pinv_0
XDEC_INV_56 Z_56 decode_56 vdd gnd pinv_0
XDEC_INV_57 Z_57 decode_57 vdd gnd pinv_0
XDEC_INV_58 Z_58 decode_58 vdd gnd pinv_0
XDEC_INV_59 Z_59 decode_59 vdd gnd pinv_0
XDEC_INV_60 Z_60 decode_60 vdd gnd pinv_0
XDEC_INV_61 Z_61 decode_61 vdd gnd pinv_0
XDEC_INV_62 Z_62 decode_62 vdd gnd pinv_0
XDEC_INV_63 Z_63 decode_63 vdd gnd pinv_0
.ENDS hierarchical_decoder_0

.SUBCKT pinv_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_1

* ptx M{0} {1} nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_2

* ptx M{0} {1} nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_3

* ptx M{0} {1} nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

.SUBCKT pinv_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_4

* ptx M{0} {1} nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

.SUBCKT pinv_5 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_5

.SUBCKT pdriver_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_1
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_1
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_1
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_2
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_3
Xbuf_inv6 Zb5_int Zb6_int vdd gnd pinv_4
Xbuf_inv7 Zb6_int Z vdd gnd pinv_5
.ENDS pdriver_0

.SUBCKT wordline_driver_0 in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 64 cols: 256
Xwl_driver_nand0 en in_0 wl_bar_0 vdd gnd pnand2_0
Xwl_driver_inv0 wl_bar_0 wl_0 vdd gnd pdriver_0
Xwl_driver_nand1 en in_1 wl_bar_1 vdd gnd pnand2_0
Xwl_driver_inv1 wl_bar_1 wl_1 vdd gnd pdriver_0
Xwl_driver_nand2 en in_2 wl_bar_2 vdd gnd pnand2_0
Xwl_driver_inv2 wl_bar_2 wl_2 vdd gnd pdriver_0
Xwl_driver_nand3 en in_3 wl_bar_3 vdd gnd pnand2_0
Xwl_driver_inv3 wl_bar_3 wl_3 vdd gnd pdriver_0
Xwl_driver_nand4 en in_4 wl_bar_4 vdd gnd pnand2_0
Xwl_driver_inv4 wl_bar_4 wl_4 vdd gnd pdriver_0
Xwl_driver_nand5 en in_5 wl_bar_5 vdd gnd pnand2_0
Xwl_driver_inv5 wl_bar_5 wl_5 vdd gnd pdriver_0
Xwl_driver_nand6 en in_6 wl_bar_6 vdd gnd pnand2_0
Xwl_driver_inv6 wl_bar_6 wl_6 vdd gnd pdriver_0
Xwl_driver_nand7 en in_7 wl_bar_7 vdd gnd pnand2_0
Xwl_driver_inv7 wl_bar_7 wl_7 vdd gnd pdriver_0
Xwl_driver_nand8 en in_8 wl_bar_8 vdd gnd pnand2_0
Xwl_driver_inv8 wl_bar_8 wl_8 vdd gnd pdriver_0
Xwl_driver_nand9 en in_9 wl_bar_9 vdd gnd pnand2_0
Xwl_driver_inv9 wl_bar_9 wl_9 vdd gnd pdriver_0
Xwl_driver_nand10 en in_10 wl_bar_10 vdd gnd pnand2_0
Xwl_driver_inv10 wl_bar_10 wl_10 vdd gnd pdriver_0
Xwl_driver_nand11 en in_11 wl_bar_11 vdd gnd pnand2_0
Xwl_driver_inv11 wl_bar_11 wl_11 vdd gnd pdriver_0
Xwl_driver_nand12 en in_12 wl_bar_12 vdd gnd pnand2_0
Xwl_driver_inv12 wl_bar_12 wl_12 vdd gnd pdriver_0
Xwl_driver_nand13 en in_13 wl_bar_13 vdd gnd pnand2_0
Xwl_driver_inv13 wl_bar_13 wl_13 vdd gnd pdriver_0
Xwl_driver_nand14 en in_14 wl_bar_14 vdd gnd pnand2_0
Xwl_driver_inv14 wl_bar_14 wl_14 vdd gnd pdriver_0
Xwl_driver_nand15 en in_15 wl_bar_15 vdd gnd pnand2_0
Xwl_driver_inv15 wl_bar_15 wl_15 vdd gnd pdriver_0
Xwl_driver_nand16 en in_16 wl_bar_16 vdd gnd pnand2_0
Xwl_driver_inv16 wl_bar_16 wl_16 vdd gnd pdriver_0
Xwl_driver_nand17 en in_17 wl_bar_17 vdd gnd pnand2_0
Xwl_driver_inv17 wl_bar_17 wl_17 vdd gnd pdriver_0
Xwl_driver_nand18 en in_18 wl_bar_18 vdd gnd pnand2_0
Xwl_driver_inv18 wl_bar_18 wl_18 vdd gnd pdriver_0
Xwl_driver_nand19 en in_19 wl_bar_19 vdd gnd pnand2_0
Xwl_driver_inv19 wl_bar_19 wl_19 vdd gnd pdriver_0
Xwl_driver_nand20 en in_20 wl_bar_20 vdd gnd pnand2_0
Xwl_driver_inv20 wl_bar_20 wl_20 vdd gnd pdriver_0
Xwl_driver_nand21 en in_21 wl_bar_21 vdd gnd pnand2_0
Xwl_driver_inv21 wl_bar_21 wl_21 vdd gnd pdriver_0
Xwl_driver_nand22 en in_22 wl_bar_22 vdd gnd pnand2_0
Xwl_driver_inv22 wl_bar_22 wl_22 vdd gnd pdriver_0
Xwl_driver_nand23 en in_23 wl_bar_23 vdd gnd pnand2_0
Xwl_driver_inv23 wl_bar_23 wl_23 vdd gnd pdriver_0
Xwl_driver_nand24 en in_24 wl_bar_24 vdd gnd pnand2_0
Xwl_driver_inv24 wl_bar_24 wl_24 vdd gnd pdriver_0
Xwl_driver_nand25 en in_25 wl_bar_25 vdd gnd pnand2_0
Xwl_driver_inv25 wl_bar_25 wl_25 vdd gnd pdriver_0
Xwl_driver_nand26 en in_26 wl_bar_26 vdd gnd pnand2_0
Xwl_driver_inv26 wl_bar_26 wl_26 vdd gnd pdriver_0
Xwl_driver_nand27 en in_27 wl_bar_27 vdd gnd pnand2_0
Xwl_driver_inv27 wl_bar_27 wl_27 vdd gnd pdriver_0
Xwl_driver_nand28 en in_28 wl_bar_28 vdd gnd pnand2_0
Xwl_driver_inv28 wl_bar_28 wl_28 vdd gnd pdriver_0
Xwl_driver_nand29 en in_29 wl_bar_29 vdd gnd pnand2_0
Xwl_driver_inv29 wl_bar_29 wl_29 vdd gnd pdriver_0
Xwl_driver_nand30 en in_30 wl_bar_30 vdd gnd pnand2_0
Xwl_driver_inv30 wl_bar_30 wl_30 vdd gnd pdriver_0
Xwl_driver_nand31 en in_31 wl_bar_31 vdd gnd pnand2_0
Xwl_driver_inv31 wl_bar_31 wl_31 vdd gnd pdriver_0
Xwl_driver_nand32 en in_32 wl_bar_32 vdd gnd pnand2_0
Xwl_driver_inv32 wl_bar_32 wl_32 vdd gnd pdriver_0
Xwl_driver_nand33 en in_33 wl_bar_33 vdd gnd pnand2_0
Xwl_driver_inv33 wl_bar_33 wl_33 vdd gnd pdriver_0
Xwl_driver_nand34 en in_34 wl_bar_34 vdd gnd pnand2_0
Xwl_driver_inv34 wl_bar_34 wl_34 vdd gnd pdriver_0
Xwl_driver_nand35 en in_35 wl_bar_35 vdd gnd pnand2_0
Xwl_driver_inv35 wl_bar_35 wl_35 vdd gnd pdriver_0
Xwl_driver_nand36 en in_36 wl_bar_36 vdd gnd pnand2_0
Xwl_driver_inv36 wl_bar_36 wl_36 vdd gnd pdriver_0
Xwl_driver_nand37 en in_37 wl_bar_37 vdd gnd pnand2_0
Xwl_driver_inv37 wl_bar_37 wl_37 vdd gnd pdriver_0
Xwl_driver_nand38 en in_38 wl_bar_38 vdd gnd pnand2_0
Xwl_driver_inv38 wl_bar_38 wl_38 vdd gnd pdriver_0
Xwl_driver_nand39 en in_39 wl_bar_39 vdd gnd pnand2_0
Xwl_driver_inv39 wl_bar_39 wl_39 vdd gnd pdriver_0
Xwl_driver_nand40 en in_40 wl_bar_40 vdd gnd pnand2_0
Xwl_driver_inv40 wl_bar_40 wl_40 vdd gnd pdriver_0
Xwl_driver_nand41 en in_41 wl_bar_41 vdd gnd pnand2_0
Xwl_driver_inv41 wl_bar_41 wl_41 vdd gnd pdriver_0
Xwl_driver_nand42 en in_42 wl_bar_42 vdd gnd pnand2_0
Xwl_driver_inv42 wl_bar_42 wl_42 vdd gnd pdriver_0
Xwl_driver_nand43 en in_43 wl_bar_43 vdd gnd pnand2_0
Xwl_driver_inv43 wl_bar_43 wl_43 vdd gnd pdriver_0
Xwl_driver_nand44 en in_44 wl_bar_44 vdd gnd pnand2_0
Xwl_driver_inv44 wl_bar_44 wl_44 vdd gnd pdriver_0
Xwl_driver_nand45 en in_45 wl_bar_45 vdd gnd pnand2_0
Xwl_driver_inv45 wl_bar_45 wl_45 vdd gnd pdriver_0
Xwl_driver_nand46 en in_46 wl_bar_46 vdd gnd pnand2_0
Xwl_driver_inv46 wl_bar_46 wl_46 vdd gnd pdriver_0
Xwl_driver_nand47 en in_47 wl_bar_47 vdd gnd pnand2_0
Xwl_driver_inv47 wl_bar_47 wl_47 vdd gnd pdriver_0
Xwl_driver_nand48 en in_48 wl_bar_48 vdd gnd pnand2_0
Xwl_driver_inv48 wl_bar_48 wl_48 vdd gnd pdriver_0
Xwl_driver_nand49 en in_49 wl_bar_49 vdd gnd pnand2_0
Xwl_driver_inv49 wl_bar_49 wl_49 vdd gnd pdriver_0
Xwl_driver_nand50 en in_50 wl_bar_50 vdd gnd pnand2_0
Xwl_driver_inv50 wl_bar_50 wl_50 vdd gnd pdriver_0
Xwl_driver_nand51 en in_51 wl_bar_51 vdd gnd pnand2_0
Xwl_driver_inv51 wl_bar_51 wl_51 vdd gnd pdriver_0
Xwl_driver_nand52 en in_52 wl_bar_52 vdd gnd pnand2_0
Xwl_driver_inv52 wl_bar_52 wl_52 vdd gnd pdriver_0
Xwl_driver_nand53 en in_53 wl_bar_53 vdd gnd pnand2_0
Xwl_driver_inv53 wl_bar_53 wl_53 vdd gnd pdriver_0
Xwl_driver_nand54 en in_54 wl_bar_54 vdd gnd pnand2_0
Xwl_driver_inv54 wl_bar_54 wl_54 vdd gnd pdriver_0
Xwl_driver_nand55 en in_55 wl_bar_55 vdd gnd pnand2_0
Xwl_driver_inv55 wl_bar_55 wl_55 vdd gnd pdriver_0
Xwl_driver_nand56 en in_56 wl_bar_56 vdd gnd pnand2_0
Xwl_driver_inv56 wl_bar_56 wl_56 vdd gnd pdriver_0
Xwl_driver_nand57 en in_57 wl_bar_57 vdd gnd pnand2_0
Xwl_driver_inv57 wl_bar_57 wl_57 vdd gnd pdriver_0
Xwl_driver_nand58 en in_58 wl_bar_58 vdd gnd pnand2_0
Xwl_driver_inv58 wl_bar_58 wl_58 vdd gnd pdriver_0
Xwl_driver_nand59 en in_59 wl_bar_59 vdd gnd pnand2_0
Xwl_driver_inv59 wl_bar_59 wl_59 vdd gnd pdriver_0
Xwl_driver_nand60 en in_60 wl_bar_60 vdd gnd pnand2_0
Xwl_driver_inv60 wl_bar_60 wl_60 vdd gnd pdriver_0
Xwl_driver_nand61 en in_61 wl_bar_61 vdd gnd pnand2_0
Xwl_driver_inv61 wl_bar_61 wl_61 vdd gnd pdriver_0
Xwl_driver_nand62 en in_62 wl_bar_62 vdd gnd pnand2_0
Xwl_driver_inv62 wl_bar_62 wl_62 vdd gnd pdriver_0
Xwl_driver_nand63 en in_63 wl_bar_63 vdd gnd pnand2_0
Xwl_driver_inv63 wl_bar_63 wl_63 vdd gnd pdriver_0
.ENDS wordline_driver_0

.SUBCKT port_address_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 vdd gnd hierarchical_decoder_0
Xwordline_driver dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_en vdd gnd wordline_driver_0
.ENDS port_address_0

.SUBCKT cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* POWER : vdd 
* GROUND: gnd 
* rows: 64 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd cell_6t
Xbit_r1_c1 bl_1 br_1 wl_1 vdd gnd cell_6t
Xbit_r2_c1 bl_1 br_1 wl_2 vdd gnd cell_6t
Xbit_r3_c1 bl_1 br_1 wl_3 vdd gnd cell_6t
Xbit_r4_c1 bl_1 br_1 wl_4 vdd gnd cell_6t
Xbit_r5_c1 bl_1 br_1 wl_5 vdd gnd cell_6t
Xbit_r6_c1 bl_1 br_1 wl_6 vdd gnd cell_6t
Xbit_r7_c1 bl_1 br_1 wl_7 vdd gnd cell_6t
Xbit_r8_c1 bl_1 br_1 wl_8 vdd gnd cell_6t
Xbit_r9_c1 bl_1 br_1 wl_9 vdd gnd cell_6t
Xbit_r10_c1 bl_1 br_1 wl_10 vdd gnd cell_6t
Xbit_r11_c1 bl_1 br_1 wl_11 vdd gnd cell_6t
Xbit_r12_c1 bl_1 br_1 wl_12 vdd gnd cell_6t
Xbit_r13_c1 bl_1 br_1 wl_13 vdd gnd cell_6t
Xbit_r14_c1 bl_1 br_1 wl_14 vdd gnd cell_6t
Xbit_r15_c1 bl_1 br_1 wl_15 vdd gnd cell_6t
Xbit_r16_c1 bl_1 br_1 wl_16 vdd gnd cell_6t
Xbit_r17_c1 bl_1 br_1 wl_17 vdd gnd cell_6t
Xbit_r18_c1 bl_1 br_1 wl_18 vdd gnd cell_6t
Xbit_r19_c1 bl_1 br_1 wl_19 vdd gnd cell_6t
Xbit_r20_c1 bl_1 br_1 wl_20 vdd gnd cell_6t
Xbit_r21_c1 bl_1 br_1 wl_21 vdd gnd cell_6t
Xbit_r22_c1 bl_1 br_1 wl_22 vdd gnd cell_6t
Xbit_r23_c1 bl_1 br_1 wl_23 vdd gnd cell_6t
Xbit_r24_c1 bl_1 br_1 wl_24 vdd gnd cell_6t
Xbit_r25_c1 bl_1 br_1 wl_25 vdd gnd cell_6t
Xbit_r26_c1 bl_1 br_1 wl_26 vdd gnd cell_6t
Xbit_r27_c1 bl_1 br_1 wl_27 vdd gnd cell_6t
Xbit_r28_c1 bl_1 br_1 wl_28 vdd gnd cell_6t
Xbit_r29_c1 bl_1 br_1 wl_29 vdd gnd cell_6t
Xbit_r30_c1 bl_1 br_1 wl_30 vdd gnd cell_6t
Xbit_r31_c1 bl_1 br_1 wl_31 vdd gnd cell_6t
Xbit_r32_c1 bl_1 br_1 wl_32 vdd gnd cell_6t
Xbit_r33_c1 bl_1 br_1 wl_33 vdd gnd cell_6t
Xbit_r34_c1 bl_1 br_1 wl_34 vdd gnd cell_6t
Xbit_r35_c1 bl_1 br_1 wl_35 vdd gnd cell_6t
Xbit_r36_c1 bl_1 br_1 wl_36 vdd gnd cell_6t
Xbit_r37_c1 bl_1 br_1 wl_37 vdd gnd cell_6t
Xbit_r38_c1 bl_1 br_1 wl_38 vdd gnd cell_6t
Xbit_r39_c1 bl_1 br_1 wl_39 vdd gnd cell_6t
Xbit_r40_c1 bl_1 br_1 wl_40 vdd gnd cell_6t
Xbit_r41_c1 bl_1 br_1 wl_41 vdd gnd cell_6t
Xbit_r42_c1 bl_1 br_1 wl_42 vdd gnd cell_6t
Xbit_r43_c1 bl_1 br_1 wl_43 vdd gnd cell_6t
Xbit_r44_c1 bl_1 br_1 wl_44 vdd gnd cell_6t
Xbit_r45_c1 bl_1 br_1 wl_45 vdd gnd cell_6t
Xbit_r46_c1 bl_1 br_1 wl_46 vdd gnd cell_6t
Xbit_r47_c1 bl_1 br_1 wl_47 vdd gnd cell_6t
Xbit_r48_c1 bl_1 br_1 wl_48 vdd gnd cell_6t
Xbit_r49_c1 bl_1 br_1 wl_49 vdd gnd cell_6t
Xbit_r50_c1 bl_1 br_1 wl_50 vdd gnd cell_6t
Xbit_r51_c1 bl_1 br_1 wl_51 vdd gnd cell_6t
Xbit_r52_c1 bl_1 br_1 wl_52 vdd gnd cell_6t
Xbit_r53_c1 bl_1 br_1 wl_53 vdd gnd cell_6t
Xbit_r54_c1 bl_1 br_1 wl_54 vdd gnd cell_6t
Xbit_r55_c1 bl_1 br_1 wl_55 vdd gnd cell_6t
Xbit_r56_c1 bl_1 br_1 wl_56 vdd gnd cell_6t
Xbit_r57_c1 bl_1 br_1 wl_57 vdd gnd cell_6t
Xbit_r58_c1 bl_1 br_1 wl_58 vdd gnd cell_6t
Xbit_r59_c1 bl_1 br_1 wl_59 vdd gnd cell_6t
Xbit_r60_c1 bl_1 br_1 wl_60 vdd gnd cell_6t
Xbit_r61_c1 bl_1 br_1 wl_61 vdd gnd cell_6t
Xbit_r62_c1 bl_1 br_1 wl_62 vdd gnd cell_6t
Xbit_r63_c1 bl_1 br_1 wl_63 vdd gnd cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd cell_6t
Xbit_r1_c2 bl_2 br_2 wl_1 vdd gnd cell_6t
Xbit_r2_c2 bl_2 br_2 wl_2 vdd gnd cell_6t
Xbit_r3_c2 bl_2 br_2 wl_3 vdd gnd cell_6t
Xbit_r4_c2 bl_2 br_2 wl_4 vdd gnd cell_6t
Xbit_r5_c2 bl_2 br_2 wl_5 vdd gnd cell_6t
Xbit_r6_c2 bl_2 br_2 wl_6 vdd gnd cell_6t
Xbit_r7_c2 bl_2 br_2 wl_7 vdd gnd cell_6t
Xbit_r8_c2 bl_2 br_2 wl_8 vdd gnd cell_6t
Xbit_r9_c2 bl_2 br_2 wl_9 vdd gnd cell_6t
Xbit_r10_c2 bl_2 br_2 wl_10 vdd gnd cell_6t
Xbit_r11_c2 bl_2 br_2 wl_11 vdd gnd cell_6t
Xbit_r12_c2 bl_2 br_2 wl_12 vdd gnd cell_6t
Xbit_r13_c2 bl_2 br_2 wl_13 vdd gnd cell_6t
Xbit_r14_c2 bl_2 br_2 wl_14 vdd gnd cell_6t
Xbit_r15_c2 bl_2 br_2 wl_15 vdd gnd cell_6t
Xbit_r16_c2 bl_2 br_2 wl_16 vdd gnd cell_6t
Xbit_r17_c2 bl_2 br_2 wl_17 vdd gnd cell_6t
Xbit_r18_c2 bl_2 br_2 wl_18 vdd gnd cell_6t
Xbit_r19_c2 bl_2 br_2 wl_19 vdd gnd cell_6t
Xbit_r20_c2 bl_2 br_2 wl_20 vdd gnd cell_6t
Xbit_r21_c2 bl_2 br_2 wl_21 vdd gnd cell_6t
Xbit_r22_c2 bl_2 br_2 wl_22 vdd gnd cell_6t
Xbit_r23_c2 bl_2 br_2 wl_23 vdd gnd cell_6t
Xbit_r24_c2 bl_2 br_2 wl_24 vdd gnd cell_6t
Xbit_r25_c2 bl_2 br_2 wl_25 vdd gnd cell_6t
Xbit_r26_c2 bl_2 br_2 wl_26 vdd gnd cell_6t
Xbit_r27_c2 bl_2 br_2 wl_27 vdd gnd cell_6t
Xbit_r28_c2 bl_2 br_2 wl_28 vdd gnd cell_6t
Xbit_r29_c2 bl_2 br_2 wl_29 vdd gnd cell_6t
Xbit_r30_c2 bl_2 br_2 wl_30 vdd gnd cell_6t
Xbit_r31_c2 bl_2 br_2 wl_31 vdd gnd cell_6t
Xbit_r32_c2 bl_2 br_2 wl_32 vdd gnd cell_6t
Xbit_r33_c2 bl_2 br_2 wl_33 vdd gnd cell_6t
Xbit_r34_c2 bl_2 br_2 wl_34 vdd gnd cell_6t
Xbit_r35_c2 bl_2 br_2 wl_35 vdd gnd cell_6t
Xbit_r36_c2 bl_2 br_2 wl_36 vdd gnd cell_6t
Xbit_r37_c2 bl_2 br_2 wl_37 vdd gnd cell_6t
Xbit_r38_c2 bl_2 br_2 wl_38 vdd gnd cell_6t
Xbit_r39_c2 bl_2 br_2 wl_39 vdd gnd cell_6t
Xbit_r40_c2 bl_2 br_2 wl_40 vdd gnd cell_6t
Xbit_r41_c2 bl_2 br_2 wl_41 vdd gnd cell_6t
Xbit_r42_c2 bl_2 br_2 wl_42 vdd gnd cell_6t
Xbit_r43_c2 bl_2 br_2 wl_43 vdd gnd cell_6t
Xbit_r44_c2 bl_2 br_2 wl_44 vdd gnd cell_6t
Xbit_r45_c2 bl_2 br_2 wl_45 vdd gnd cell_6t
Xbit_r46_c2 bl_2 br_2 wl_46 vdd gnd cell_6t
Xbit_r47_c2 bl_2 br_2 wl_47 vdd gnd cell_6t
Xbit_r48_c2 bl_2 br_2 wl_48 vdd gnd cell_6t
Xbit_r49_c2 bl_2 br_2 wl_49 vdd gnd cell_6t
Xbit_r50_c2 bl_2 br_2 wl_50 vdd gnd cell_6t
Xbit_r51_c2 bl_2 br_2 wl_51 vdd gnd cell_6t
Xbit_r52_c2 bl_2 br_2 wl_52 vdd gnd cell_6t
Xbit_r53_c2 bl_2 br_2 wl_53 vdd gnd cell_6t
Xbit_r54_c2 bl_2 br_2 wl_54 vdd gnd cell_6t
Xbit_r55_c2 bl_2 br_2 wl_55 vdd gnd cell_6t
Xbit_r56_c2 bl_2 br_2 wl_56 vdd gnd cell_6t
Xbit_r57_c2 bl_2 br_2 wl_57 vdd gnd cell_6t
Xbit_r58_c2 bl_2 br_2 wl_58 vdd gnd cell_6t
Xbit_r59_c2 bl_2 br_2 wl_59 vdd gnd cell_6t
Xbit_r60_c2 bl_2 br_2 wl_60 vdd gnd cell_6t
Xbit_r61_c2 bl_2 br_2 wl_61 vdd gnd cell_6t
Xbit_r62_c2 bl_2 br_2 wl_62 vdd gnd cell_6t
Xbit_r63_c2 bl_2 br_2 wl_63 vdd gnd cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd cell_6t
Xbit_r1_c3 bl_3 br_3 wl_1 vdd gnd cell_6t
Xbit_r2_c3 bl_3 br_3 wl_2 vdd gnd cell_6t
Xbit_r3_c3 bl_3 br_3 wl_3 vdd gnd cell_6t
Xbit_r4_c3 bl_3 br_3 wl_4 vdd gnd cell_6t
Xbit_r5_c3 bl_3 br_3 wl_5 vdd gnd cell_6t
Xbit_r6_c3 bl_3 br_3 wl_6 vdd gnd cell_6t
Xbit_r7_c3 bl_3 br_3 wl_7 vdd gnd cell_6t
Xbit_r8_c3 bl_3 br_3 wl_8 vdd gnd cell_6t
Xbit_r9_c3 bl_3 br_3 wl_9 vdd gnd cell_6t
Xbit_r10_c3 bl_3 br_3 wl_10 vdd gnd cell_6t
Xbit_r11_c3 bl_3 br_3 wl_11 vdd gnd cell_6t
Xbit_r12_c3 bl_3 br_3 wl_12 vdd gnd cell_6t
Xbit_r13_c3 bl_3 br_3 wl_13 vdd gnd cell_6t
Xbit_r14_c3 bl_3 br_3 wl_14 vdd gnd cell_6t
Xbit_r15_c3 bl_3 br_3 wl_15 vdd gnd cell_6t
Xbit_r16_c3 bl_3 br_3 wl_16 vdd gnd cell_6t
Xbit_r17_c3 bl_3 br_3 wl_17 vdd gnd cell_6t
Xbit_r18_c3 bl_3 br_3 wl_18 vdd gnd cell_6t
Xbit_r19_c3 bl_3 br_3 wl_19 vdd gnd cell_6t
Xbit_r20_c3 bl_3 br_3 wl_20 vdd gnd cell_6t
Xbit_r21_c3 bl_3 br_3 wl_21 vdd gnd cell_6t
Xbit_r22_c3 bl_3 br_3 wl_22 vdd gnd cell_6t
Xbit_r23_c3 bl_3 br_3 wl_23 vdd gnd cell_6t
Xbit_r24_c3 bl_3 br_3 wl_24 vdd gnd cell_6t
Xbit_r25_c3 bl_3 br_3 wl_25 vdd gnd cell_6t
Xbit_r26_c3 bl_3 br_3 wl_26 vdd gnd cell_6t
Xbit_r27_c3 bl_3 br_3 wl_27 vdd gnd cell_6t
Xbit_r28_c3 bl_3 br_3 wl_28 vdd gnd cell_6t
Xbit_r29_c3 bl_3 br_3 wl_29 vdd gnd cell_6t
Xbit_r30_c3 bl_3 br_3 wl_30 vdd gnd cell_6t
Xbit_r31_c3 bl_3 br_3 wl_31 vdd gnd cell_6t
Xbit_r32_c3 bl_3 br_3 wl_32 vdd gnd cell_6t
Xbit_r33_c3 bl_3 br_3 wl_33 vdd gnd cell_6t
Xbit_r34_c3 bl_3 br_3 wl_34 vdd gnd cell_6t
Xbit_r35_c3 bl_3 br_3 wl_35 vdd gnd cell_6t
Xbit_r36_c3 bl_3 br_3 wl_36 vdd gnd cell_6t
Xbit_r37_c3 bl_3 br_3 wl_37 vdd gnd cell_6t
Xbit_r38_c3 bl_3 br_3 wl_38 vdd gnd cell_6t
Xbit_r39_c3 bl_3 br_3 wl_39 vdd gnd cell_6t
Xbit_r40_c3 bl_3 br_3 wl_40 vdd gnd cell_6t
Xbit_r41_c3 bl_3 br_3 wl_41 vdd gnd cell_6t
Xbit_r42_c3 bl_3 br_3 wl_42 vdd gnd cell_6t
Xbit_r43_c3 bl_3 br_3 wl_43 vdd gnd cell_6t
Xbit_r44_c3 bl_3 br_3 wl_44 vdd gnd cell_6t
Xbit_r45_c3 bl_3 br_3 wl_45 vdd gnd cell_6t
Xbit_r46_c3 bl_3 br_3 wl_46 vdd gnd cell_6t
Xbit_r47_c3 bl_3 br_3 wl_47 vdd gnd cell_6t
Xbit_r48_c3 bl_3 br_3 wl_48 vdd gnd cell_6t
Xbit_r49_c3 bl_3 br_3 wl_49 vdd gnd cell_6t
Xbit_r50_c3 bl_3 br_3 wl_50 vdd gnd cell_6t
Xbit_r51_c3 bl_3 br_3 wl_51 vdd gnd cell_6t
Xbit_r52_c3 bl_3 br_3 wl_52 vdd gnd cell_6t
Xbit_r53_c3 bl_3 br_3 wl_53 vdd gnd cell_6t
Xbit_r54_c3 bl_3 br_3 wl_54 vdd gnd cell_6t
Xbit_r55_c3 bl_3 br_3 wl_55 vdd gnd cell_6t
Xbit_r56_c3 bl_3 br_3 wl_56 vdd gnd cell_6t
Xbit_r57_c3 bl_3 br_3 wl_57 vdd gnd cell_6t
Xbit_r58_c3 bl_3 br_3 wl_58 vdd gnd cell_6t
Xbit_r59_c3 bl_3 br_3 wl_59 vdd gnd cell_6t
Xbit_r60_c3 bl_3 br_3 wl_60 vdd gnd cell_6t
Xbit_r61_c3 bl_3 br_3 wl_61 vdd gnd cell_6t
Xbit_r62_c3 bl_3 br_3 wl_62 vdd gnd cell_6t
Xbit_r63_c3 bl_3 br_3 wl_63 vdd gnd cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd cell_6t
Xbit_r1_c4 bl_4 br_4 wl_1 vdd gnd cell_6t
Xbit_r2_c4 bl_4 br_4 wl_2 vdd gnd cell_6t
Xbit_r3_c4 bl_4 br_4 wl_3 vdd gnd cell_6t
Xbit_r4_c4 bl_4 br_4 wl_4 vdd gnd cell_6t
Xbit_r5_c4 bl_4 br_4 wl_5 vdd gnd cell_6t
Xbit_r6_c4 bl_4 br_4 wl_6 vdd gnd cell_6t
Xbit_r7_c4 bl_4 br_4 wl_7 vdd gnd cell_6t
Xbit_r8_c4 bl_4 br_4 wl_8 vdd gnd cell_6t
Xbit_r9_c4 bl_4 br_4 wl_9 vdd gnd cell_6t
Xbit_r10_c4 bl_4 br_4 wl_10 vdd gnd cell_6t
Xbit_r11_c4 bl_4 br_4 wl_11 vdd gnd cell_6t
Xbit_r12_c4 bl_4 br_4 wl_12 vdd gnd cell_6t
Xbit_r13_c4 bl_4 br_4 wl_13 vdd gnd cell_6t
Xbit_r14_c4 bl_4 br_4 wl_14 vdd gnd cell_6t
Xbit_r15_c4 bl_4 br_4 wl_15 vdd gnd cell_6t
Xbit_r16_c4 bl_4 br_4 wl_16 vdd gnd cell_6t
Xbit_r17_c4 bl_4 br_4 wl_17 vdd gnd cell_6t
Xbit_r18_c4 bl_4 br_4 wl_18 vdd gnd cell_6t
Xbit_r19_c4 bl_4 br_4 wl_19 vdd gnd cell_6t
Xbit_r20_c4 bl_4 br_4 wl_20 vdd gnd cell_6t
Xbit_r21_c4 bl_4 br_4 wl_21 vdd gnd cell_6t
Xbit_r22_c4 bl_4 br_4 wl_22 vdd gnd cell_6t
Xbit_r23_c4 bl_4 br_4 wl_23 vdd gnd cell_6t
Xbit_r24_c4 bl_4 br_4 wl_24 vdd gnd cell_6t
Xbit_r25_c4 bl_4 br_4 wl_25 vdd gnd cell_6t
Xbit_r26_c4 bl_4 br_4 wl_26 vdd gnd cell_6t
Xbit_r27_c4 bl_4 br_4 wl_27 vdd gnd cell_6t
Xbit_r28_c4 bl_4 br_4 wl_28 vdd gnd cell_6t
Xbit_r29_c4 bl_4 br_4 wl_29 vdd gnd cell_6t
Xbit_r30_c4 bl_4 br_4 wl_30 vdd gnd cell_6t
Xbit_r31_c4 bl_4 br_4 wl_31 vdd gnd cell_6t
Xbit_r32_c4 bl_4 br_4 wl_32 vdd gnd cell_6t
Xbit_r33_c4 bl_4 br_4 wl_33 vdd gnd cell_6t
Xbit_r34_c4 bl_4 br_4 wl_34 vdd gnd cell_6t
Xbit_r35_c4 bl_4 br_4 wl_35 vdd gnd cell_6t
Xbit_r36_c4 bl_4 br_4 wl_36 vdd gnd cell_6t
Xbit_r37_c4 bl_4 br_4 wl_37 vdd gnd cell_6t
Xbit_r38_c4 bl_4 br_4 wl_38 vdd gnd cell_6t
Xbit_r39_c4 bl_4 br_4 wl_39 vdd gnd cell_6t
Xbit_r40_c4 bl_4 br_4 wl_40 vdd gnd cell_6t
Xbit_r41_c4 bl_4 br_4 wl_41 vdd gnd cell_6t
Xbit_r42_c4 bl_4 br_4 wl_42 vdd gnd cell_6t
Xbit_r43_c4 bl_4 br_4 wl_43 vdd gnd cell_6t
Xbit_r44_c4 bl_4 br_4 wl_44 vdd gnd cell_6t
Xbit_r45_c4 bl_4 br_4 wl_45 vdd gnd cell_6t
Xbit_r46_c4 bl_4 br_4 wl_46 vdd gnd cell_6t
Xbit_r47_c4 bl_4 br_4 wl_47 vdd gnd cell_6t
Xbit_r48_c4 bl_4 br_4 wl_48 vdd gnd cell_6t
Xbit_r49_c4 bl_4 br_4 wl_49 vdd gnd cell_6t
Xbit_r50_c4 bl_4 br_4 wl_50 vdd gnd cell_6t
Xbit_r51_c4 bl_4 br_4 wl_51 vdd gnd cell_6t
Xbit_r52_c4 bl_4 br_4 wl_52 vdd gnd cell_6t
Xbit_r53_c4 bl_4 br_4 wl_53 vdd gnd cell_6t
Xbit_r54_c4 bl_4 br_4 wl_54 vdd gnd cell_6t
Xbit_r55_c4 bl_4 br_4 wl_55 vdd gnd cell_6t
Xbit_r56_c4 bl_4 br_4 wl_56 vdd gnd cell_6t
Xbit_r57_c4 bl_4 br_4 wl_57 vdd gnd cell_6t
Xbit_r58_c4 bl_4 br_4 wl_58 vdd gnd cell_6t
Xbit_r59_c4 bl_4 br_4 wl_59 vdd gnd cell_6t
Xbit_r60_c4 bl_4 br_4 wl_60 vdd gnd cell_6t
Xbit_r61_c4 bl_4 br_4 wl_61 vdd gnd cell_6t
Xbit_r62_c4 bl_4 br_4 wl_62 vdd gnd cell_6t
Xbit_r63_c4 bl_4 br_4 wl_63 vdd gnd cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd cell_6t
Xbit_r1_c5 bl_5 br_5 wl_1 vdd gnd cell_6t
Xbit_r2_c5 bl_5 br_5 wl_2 vdd gnd cell_6t
Xbit_r3_c5 bl_5 br_5 wl_3 vdd gnd cell_6t
Xbit_r4_c5 bl_5 br_5 wl_4 vdd gnd cell_6t
Xbit_r5_c5 bl_5 br_5 wl_5 vdd gnd cell_6t
Xbit_r6_c5 bl_5 br_5 wl_6 vdd gnd cell_6t
Xbit_r7_c5 bl_5 br_5 wl_7 vdd gnd cell_6t
Xbit_r8_c5 bl_5 br_5 wl_8 vdd gnd cell_6t
Xbit_r9_c5 bl_5 br_5 wl_9 vdd gnd cell_6t
Xbit_r10_c5 bl_5 br_5 wl_10 vdd gnd cell_6t
Xbit_r11_c5 bl_5 br_5 wl_11 vdd gnd cell_6t
Xbit_r12_c5 bl_5 br_5 wl_12 vdd gnd cell_6t
Xbit_r13_c5 bl_5 br_5 wl_13 vdd gnd cell_6t
Xbit_r14_c5 bl_5 br_5 wl_14 vdd gnd cell_6t
Xbit_r15_c5 bl_5 br_5 wl_15 vdd gnd cell_6t
Xbit_r16_c5 bl_5 br_5 wl_16 vdd gnd cell_6t
Xbit_r17_c5 bl_5 br_5 wl_17 vdd gnd cell_6t
Xbit_r18_c5 bl_5 br_5 wl_18 vdd gnd cell_6t
Xbit_r19_c5 bl_5 br_5 wl_19 vdd gnd cell_6t
Xbit_r20_c5 bl_5 br_5 wl_20 vdd gnd cell_6t
Xbit_r21_c5 bl_5 br_5 wl_21 vdd gnd cell_6t
Xbit_r22_c5 bl_5 br_5 wl_22 vdd gnd cell_6t
Xbit_r23_c5 bl_5 br_5 wl_23 vdd gnd cell_6t
Xbit_r24_c5 bl_5 br_5 wl_24 vdd gnd cell_6t
Xbit_r25_c5 bl_5 br_5 wl_25 vdd gnd cell_6t
Xbit_r26_c5 bl_5 br_5 wl_26 vdd gnd cell_6t
Xbit_r27_c5 bl_5 br_5 wl_27 vdd gnd cell_6t
Xbit_r28_c5 bl_5 br_5 wl_28 vdd gnd cell_6t
Xbit_r29_c5 bl_5 br_5 wl_29 vdd gnd cell_6t
Xbit_r30_c5 bl_5 br_5 wl_30 vdd gnd cell_6t
Xbit_r31_c5 bl_5 br_5 wl_31 vdd gnd cell_6t
Xbit_r32_c5 bl_5 br_5 wl_32 vdd gnd cell_6t
Xbit_r33_c5 bl_5 br_5 wl_33 vdd gnd cell_6t
Xbit_r34_c5 bl_5 br_5 wl_34 vdd gnd cell_6t
Xbit_r35_c5 bl_5 br_5 wl_35 vdd gnd cell_6t
Xbit_r36_c5 bl_5 br_5 wl_36 vdd gnd cell_6t
Xbit_r37_c5 bl_5 br_5 wl_37 vdd gnd cell_6t
Xbit_r38_c5 bl_5 br_5 wl_38 vdd gnd cell_6t
Xbit_r39_c5 bl_5 br_5 wl_39 vdd gnd cell_6t
Xbit_r40_c5 bl_5 br_5 wl_40 vdd gnd cell_6t
Xbit_r41_c5 bl_5 br_5 wl_41 vdd gnd cell_6t
Xbit_r42_c5 bl_5 br_5 wl_42 vdd gnd cell_6t
Xbit_r43_c5 bl_5 br_5 wl_43 vdd gnd cell_6t
Xbit_r44_c5 bl_5 br_5 wl_44 vdd gnd cell_6t
Xbit_r45_c5 bl_5 br_5 wl_45 vdd gnd cell_6t
Xbit_r46_c5 bl_5 br_5 wl_46 vdd gnd cell_6t
Xbit_r47_c5 bl_5 br_5 wl_47 vdd gnd cell_6t
Xbit_r48_c5 bl_5 br_5 wl_48 vdd gnd cell_6t
Xbit_r49_c5 bl_5 br_5 wl_49 vdd gnd cell_6t
Xbit_r50_c5 bl_5 br_5 wl_50 vdd gnd cell_6t
Xbit_r51_c5 bl_5 br_5 wl_51 vdd gnd cell_6t
Xbit_r52_c5 bl_5 br_5 wl_52 vdd gnd cell_6t
Xbit_r53_c5 bl_5 br_5 wl_53 vdd gnd cell_6t
Xbit_r54_c5 bl_5 br_5 wl_54 vdd gnd cell_6t
Xbit_r55_c5 bl_5 br_5 wl_55 vdd gnd cell_6t
Xbit_r56_c5 bl_5 br_5 wl_56 vdd gnd cell_6t
Xbit_r57_c5 bl_5 br_5 wl_57 vdd gnd cell_6t
Xbit_r58_c5 bl_5 br_5 wl_58 vdd gnd cell_6t
Xbit_r59_c5 bl_5 br_5 wl_59 vdd gnd cell_6t
Xbit_r60_c5 bl_5 br_5 wl_60 vdd gnd cell_6t
Xbit_r61_c5 bl_5 br_5 wl_61 vdd gnd cell_6t
Xbit_r62_c5 bl_5 br_5 wl_62 vdd gnd cell_6t
Xbit_r63_c5 bl_5 br_5 wl_63 vdd gnd cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd cell_6t
Xbit_r1_c6 bl_6 br_6 wl_1 vdd gnd cell_6t
Xbit_r2_c6 bl_6 br_6 wl_2 vdd gnd cell_6t
Xbit_r3_c6 bl_6 br_6 wl_3 vdd gnd cell_6t
Xbit_r4_c6 bl_6 br_6 wl_4 vdd gnd cell_6t
Xbit_r5_c6 bl_6 br_6 wl_5 vdd gnd cell_6t
Xbit_r6_c6 bl_6 br_6 wl_6 vdd gnd cell_6t
Xbit_r7_c6 bl_6 br_6 wl_7 vdd gnd cell_6t
Xbit_r8_c6 bl_6 br_6 wl_8 vdd gnd cell_6t
Xbit_r9_c6 bl_6 br_6 wl_9 vdd gnd cell_6t
Xbit_r10_c6 bl_6 br_6 wl_10 vdd gnd cell_6t
Xbit_r11_c6 bl_6 br_6 wl_11 vdd gnd cell_6t
Xbit_r12_c6 bl_6 br_6 wl_12 vdd gnd cell_6t
Xbit_r13_c6 bl_6 br_6 wl_13 vdd gnd cell_6t
Xbit_r14_c6 bl_6 br_6 wl_14 vdd gnd cell_6t
Xbit_r15_c6 bl_6 br_6 wl_15 vdd gnd cell_6t
Xbit_r16_c6 bl_6 br_6 wl_16 vdd gnd cell_6t
Xbit_r17_c6 bl_6 br_6 wl_17 vdd gnd cell_6t
Xbit_r18_c6 bl_6 br_6 wl_18 vdd gnd cell_6t
Xbit_r19_c6 bl_6 br_6 wl_19 vdd gnd cell_6t
Xbit_r20_c6 bl_6 br_6 wl_20 vdd gnd cell_6t
Xbit_r21_c6 bl_6 br_6 wl_21 vdd gnd cell_6t
Xbit_r22_c6 bl_6 br_6 wl_22 vdd gnd cell_6t
Xbit_r23_c6 bl_6 br_6 wl_23 vdd gnd cell_6t
Xbit_r24_c6 bl_6 br_6 wl_24 vdd gnd cell_6t
Xbit_r25_c6 bl_6 br_6 wl_25 vdd gnd cell_6t
Xbit_r26_c6 bl_6 br_6 wl_26 vdd gnd cell_6t
Xbit_r27_c6 bl_6 br_6 wl_27 vdd gnd cell_6t
Xbit_r28_c6 bl_6 br_6 wl_28 vdd gnd cell_6t
Xbit_r29_c6 bl_6 br_6 wl_29 vdd gnd cell_6t
Xbit_r30_c6 bl_6 br_6 wl_30 vdd gnd cell_6t
Xbit_r31_c6 bl_6 br_6 wl_31 vdd gnd cell_6t
Xbit_r32_c6 bl_6 br_6 wl_32 vdd gnd cell_6t
Xbit_r33_c6 bl_6 br_6 wl_33 vdd gnd cell_6t
Xbit_r34_c6 bl_6 br_6 wl_34 vdd gnd cell_6t
Xbit_r35_c6 bl_6 br_6 wl_35 vdd gnd cell_6t
Xbit_r36_c6 bl_6 br_6 wl_36 vdd gnd cell_6t
Xbit_r37_c6 bl_6 br_6 wl_37 vdd gnd cell_6t
Xbit_r38_c6 bl_6 br_6 wl_38 vdd gnd cell_6t
Xbit_r39_c6 bl_6 br_6 wl_39 vdd gnd cell_6t
Xbit_r40_c6 bl_6 br_6 wl_40 vdd gnd cell_6t
Xbit_r41_c6 bl_6 br_6 wl_41 vdd gnd cell_6t
Xbit_r42_c6 bl_6 br_6 wl_42 vdd gnd cell_6t
Xbit_r43_c6 bl_6 br_6 wl_43 vdd gnd cell_6t
Xbit_r44_c6 bl_6 br_6 wl_44 vdd gnd cell_6t
Xbit_r45_c6 bl_6 br_6 wl_45 vdd gnd cell_6t
Xbit_r46_c6 bl_6 br_6 wl_46 vdd gnd cell_6t
Xbit_r47_c6 bl_6 br_6 wl_47 vdd gnd cell_6t
Xbit_r48_c6 bl_6 br_6 wl_48 vdd gnd cell_6t
Xbit_r49_c6 bl_6 br_6 wl_49 vdd gnd cell_6t
Xbit_r50_c6 bl_6 br_6 wl_50 vdd gnd cell_6t
Xbit_r51_c6 bl_6 br_6 wl_51 vdd gnd cell_6t
Xbit_r52_c6 bl_6 br_6 wl_52 vdd gnd cell_6t
Xbit_r53_c6 bl_6 br_6 wl_53 vdd gnd cell_6t
Xbit_r54_c6 bl_6 br_6 wl_54 vdd gnd cell_6t
Xbit_r55_c6 bl_6 br_6 wl_55 vdd gnd cell_6t
Xbit_r56_c6 bl_6 br_6 wl_56 vdd gnd cell_6t
Xbit_r57_c6 bl_6 br_6 wl_57 vdd gnd cell_6t
Xbit_r58_c6 bl_6 br_6 wl_58 vdd gnd cell_6t
Xbit_r59_c6 bl_6 br_6 wl_59 vdd gnd cell_6t
Xbit_r60_c6 bl_6 br_6 wl_60 vdd gnd cell_6t
Xbit_r61_c6 bl_6 br_6 wl_61 vdd gnd cell_6t
Xbit_r62_c6 bl_6 br_6 wl_62 vdd gnd cell_6t
Xbit_r63_c6 bl_6 br_6 wl_63 vdd gnd cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd cell_6t
Xbit_r1_c7 bl_7 br_7 wl_1 vdd gnd cell_6t
Xbit_r2_c7 bl_7 br_7 wl_2 vdd gnd cell_6t
Xbit_r3_c7 bl_7 br_7 wl_3 vdd gnd cell_6t
Xbit_r4_c7 bl_7 br_7 wl_4 vdd gnd cell_6t
Xbit_r5_c7 bl_7 br_7 wl_5 vdd gnd cell_6t
Xbit_r6_c7 bl_7 br_7 wl_6 vdd gnd cell_6t
Xbit_r7_c7 bl_7 br_7 wl_7 vdd gnd cell_6t
Xbit_r8_c7 bl_7 br_7 wl_8 vdd gnd cell_6t
Xbit_r9_c7 bl_7 br_7 wl_9 vdd gnd cell_6t
Xbit_r10_c7 bl_7 br_7 wl_10 vdd gnd cell_6t
Xbit_r11_c7 bl_7 br_7 wl_11 vdd gnd cell_6t
Xbit_r12_c7 bl_7 br_7 wl_12 vdd gnd cell_6t
Xbit_r13_c7 bl_7 br_7 wl_13 vdd gnd cell_6t
Xbit_r14_c7 bl_7 br_7 wl_14 vdd gnd cell_6t
Xbit_r15_c7 bl_7 br_7 wl_15 vdd gnd cell_6t
Xbit_r16_c7 bl_7 br_7 wl_16 vdd gnd cell_6t
Xbit_r17_c7 bl_7 br_7 wl_17 vdd gnd cell_6t
Xbit_r18_c7 bl_7 br_7 wl_18 vdd gnd cell_6t
Xbit_r19_c7 bl_7 br_7 wl_19 vdd gnd cell_6t
Xbit_r20_c7 bl_7 br_7 wl_20 vdd gnd cell_6t
Xbit_r21_c7 bl_7 br_7 wl_21 vdd gnd cell_6t
Xbit_r22_c7 bl_7 br_7 wl_22 vdd gnd cell_6t
Xbit_r23_c7 bl_7 br_7 wl_23 vdd gnd cell_6t
Xbit_r24_c7 bl_7 br_7 wl_24 vdd gnd cell_6t
Xbit_r25_c7 bl_7 br_7 wl_25 vdd gnd cell_6t
Xbit_r26_c7 bl_7 br_7 wl_26 vdd gnd cell_6t
Xbit_r27_c7 bl_7 br_7 wl_27 vdd gnd cell_6t
Xbit_r28_c7 bl_7 br_7 wl_28 vdd gnd cell_6t
Xbit_r29_c7 bl_7 br_7 wl_29 vdd gnd cell_6t
Xbit_r30_c7 bl_7 br_7 wl_30 vdd gnd cell_6t
Xbit_r31_c7 bl_7 br_7 wl_31 vdd gnd cell_6t
Xbit_r32_c7 bl_7 br_7 wl_32 vdd gnd cell_6t
Xbit_r33_c7 bl_7 br_7 wl_33 vdd gnd cell_6t
Xbit_r34_c7 bl_7 br_7 wl_34 vdd gnd cell_6t
Xbit_r35_c7 bl_7 br_7 wl_35 vdd gnd cell_6t
Xbit_r36_c7 bl_7 br_7 wl_36 vdd gnd cell_6t
Xbit_r37_c7 bl_7 br_7 wl_37 vdd gnd cell_6t
Xbit_r38_c7 bl_7 br_7 wl_38 vdd gnd cell_6t
Xbit_r39_c7 bl_7 br_7 wl_39 vdd gnd cell_6t
Xbit_r40_c7 bl_7 br_7 wl_40 vdd gnd cell_6t
Xbit_r41_c7 bl_7 br_7 wl_41 vdd gnd cell_6t
Xbit_r42_c7 bl_7 br_7 wl_42 vdd gnd cell_6t
Xbit_r43_c7 bl_7 br_7 wl_43 vdd gnd cell_6t
Xbit_r44_c7 bl_7 br_7 wl_44 vdd gnd cell_6t
Xbit_r45_c7 bl_7 br_7 wl_45 vdd gnd cell_6t
Xbit_r46_c7 bl_7 br_7 wl_46 vdd gnd cell_6t
Xbit_r47_c7 bl_7 br_7 wl_47 vdd gnd cell_6t
Xbit_r48_c7 bl_7 br_7 wl_48 vdd gnd cell_6t
Xbit_r49_c7 bl_7 br_7 wl_49 vdd gnd cell_6t
Xbit_r50_c7 bl_7 br_7 wl_50 vdd gnd cell_6t
Xbit_r51_c7 bl_7 br_7 wl_51 vdd gnd cell_6t
Xbit_r52_c7 bl_7 br_7 wl_52 vdd gnd cell_6t
Xbit_r53_c7 bl_7 br_7 wl_53 vdd gnd cell_6t
Xbit_r54_c7 bl_7 br_7 wl_54 vdd gnd cell_6t
Xbit_r55_c7 bl_7 br_7 wl_55 vdd gnd cell_6t
Xbit_r56_c7 bl_7 br_7 wl_56 vdd gnd cell_6t
Xbit_r57_c7 bl_7 br_7 wl_57 vdd gnd cell_6t
Xbit_r58_c7 bl_7 br_7 wl_58 vdd gnd cell_6t
Xbit_r59_c7 bl_7 br_7 wl_59 vdd gnd cell_6t
Xbit_r60_c7 bl_7 br_7 wl_60 vdd gnd cell_6t
Xbit_r61_c7 bl_7 br_7 wl_61 vdd gnd cell_6t
Xbit_r62_c7 bl_7 br_7 wl_62 vdd gnd cell_6t
Xbit_r63_c7 bl_7 br_7 wl_63 vdd gnd cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd cell_6t
Xbit_r1_c8 bl_8 br_8 wl_1 vdd gnd cell_6t
Xbit_r2_c8 bl_8 br_8 wl_2 vdd gnd cell_6t
Xbit_r3_c8 bl_8 br_8 wl_3 vdd gnd cell_6t
Xbit_r4_c8 bl_8 br_8 wl_4 vdd gnd cell_6t
Xbit_r5_c8 bl_8 br_8 wl_5 vdd gnd cell_6t
Xbit_r6_c8 bl_8 br_8 wl_6 vdd gnd cell_6t
Xbit_r7_c8 bl_8 br_8 wl_7 vdd gnd cell_6t
Xbit_r8_c8 bl_8 br_8 wl_8 vdd gnd cell_6t
Xbit_r9_c8 bl_8 br_8 wl_9 vdd gnd cell_6t
Xbit_r10_c8 bl_8 br_8 wl_10 vdd gnd cell_6t
Xbit_r11_c8 bl_8 br_8 wl_11 vdd gnd cell_6t
Xbit_r12_c8 bl_8 br_8 wl_12 vdd gnd cell_6t
Xbit_r13_c8 bl_8 br_8 wl_13 vdd gnd cell_6t
Xbit_r14_c8 bl_8 br_8 wl_14 vdd gnd cell_6t
Xbit_r15_c8 bl_8 br_8 wl_15 vdd gnd cell_6t
Xbit_r16_c8 bl_8 br_8 wl_16 vdd gnd cell_6t
Xbit_r17_c8 bl_8 br_8 wl_17 vdd gnd cell_6t
Xbit_r18_c8 bl_8 br_8 wl_18 vdd gnd cell_6t
Xbit_r19_c8 bl_8 br_8 wl_19 vdd gnd cell_6t
Xbit_r20_c8 bl_8 br_8 wl_20 vdd gnd cell_6t
Xbit_r21_c8 bl_8 br_8 wl_21 vdd gnd cell_6t
Xbit_r22_c8 bl_8 br_8 wl_22 vdd gnd cell_6t
Xbit_r23_c8 bl_8 br_8 wl_23 vdd gnd cell_6t
Xbit_r24_c8 bl_8 br_8 wl_24 vdd gnd cell_6t
Xbit_r25_c8 bl_8 br_8 wl_25 vdd gnd cell_6t
Xbit_r26_c8 bl_8 br_8 wl_26 vdd gnd cell_6t
Xbit_r27_c8 bl_8 br_8 wl_27 vdd gnd cell_6t
Xbit_r28_c8 bl_8 br_8 wl_28 vdd gnd cell_6t
Xbit_r29_c8 bl_8 br_8 wl_29 vdd gnd cell_6t
Xbit_r30_c8 bl_8 br_8 wl_30 vdd gnd cell_6t
Xbit_r31_c8 bl_8 br_8 wl_31 vdd gnd cell_6t
Xbit_r32_c8 bl_8 br_8 wl_32 vdd gnd cell_6t
Xbit_r33_c8 bl_8 br_8 wl_33 vdd gnd cell_6t
Xbit_r34_c8 bl_8 br_8 wl_34 vdd gnd cell_6t
Xbit_r35_c8 bl_8 br_8 wl_35 vdd gnd cell_6t
Xbit_r36_c8 bl_8 br_8 wl_36 vdd gnd cell_6t
Xbit_r37_c8 bl_8 br_8 wl_37 vdd gnd cell_6t
Xbit_r38_c8 bl_8 br_8 wl_38 vdd gnd cell_6t
Xbit_r39_c8 bl_8 br_8 wl_39 vdd gnd cell_6t
Xbit_r40_c8 bl_8 br_8 wl_40 vdd gnd cell_6t
Xbit_r41_c8 bl_8 br_8 wl_41 vdd gnd cell_6t
Xbit_r42_c8 bl_8 br_8 wl_42 vdd gnd cell_6t
Xbit_r43_c8 bl_8 br_8 wl_43 vdd gnd cell_6t
Xbit_r44_c8 bl_8 br_8 wl_44 vdd gnd cell_6t
Xbit_r45_c8 bl_8 br_8 wl_45 vdd gnd cell_6t
Xbit_r46_c8 bl_8 br_8 wl_46 vdd gnd cell_6t
Xbit_r47_c8 bl_8 br_8 wl_47 vdd gnd cell_6t
Xbit_r48_c8 bl_8 br_8 wl_48 vdd gnd cell_6t
Xbit_r49_c8 bl_8 br_8 wl_49 vdd gnd cell_6t
Xbit_r50_c8 bl_8 br_8 wl_50 vdd gnd cell_6t
Xbit_r51_c8 bl_8 br_8 wl_51 vdd gnd cell_6t
Xbit_r52_c8 bl_8 br_8 wl_52 vdd gnd cell_6t
Xbit_r53_c8 bl_8 br_8 wl_53 vdd gnd cell_6t
Xbit_r54_c8 bl_8 br_8 wl_54 vdd gnd cell_6t
Xbit_r55_c8 bl_8 br_8 wl_55 vdd gnd cell_6t
Xbit_r56_c8 bl_8 br_8 wl_56 vdd gnd cell_6t
Xbit_r57_c8 bl_8 br_8 wl_57 vdd gnd cell_6t
Xbit_r58_c8 bl_8 br_8 wl_58 vdd gnd cell_6t
Xbit_r59_c8 bl_8 br_8 wl_59 vdd gnd cell_6t
Xbit_r60_c8 bl_8 br_8 wl_60 vdd gnd cell_6t
Xbit_r61_c8 bl_8 br_8 wl_61 vdd gnd cell_6t
Xbit_r62_c8 bl_8 br_8 wl_62 vdd gnd cell_6t
Xbit_r63_c8 bl_8 br_8 wl_63 vdd gnd cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd cell_6t
Xbit_r1_c9 bl_9 br_9 wl_1 vdd gnd cell_6t
Xbit_r2_c9 bl_9 br_9 wl_2 vdd gnd cell_6t
Xbit_r3_c9 bl_9 br_9 wl_3 vdd gnd cell_6t
Xbit_r4_c9 bl_9 br_9 wl_4 vdd gnd cell_6t
Xbit_r5_c9 bl_9 br_9 wl_5 vdd gnd cell_6t
Xbit_r6_c9 bl_9 br_9 wl_6 vdd gnd cell_6t
Xbit_r7_c9 bl_9 br_9 wl_7 vdd gnd cell_6t
Xbit_r8_c9 bl_9 br_9 wl_8 vdd gnd cell_6t
Xbit_r9_c9 bl_9 br_9 wl_9 vdd gnd cell_6t
Xbit_r10_c9 bl_9 br_9 wl_10 vdd gnd cell_6t
Xbit_r11_c9 bl_9 br_9 wl_11 vdd gnd cell_6t
Xbit_r12_c9 bl_9 br_9 wl_12 vdd gnd cell_6t
Xbit_r13_c9 bl_9 br_9 wl_13 vdd gnd cell_6t
Xbit_r14_c9 bl_9 br_9 wl_14 vdd gnd cell_6t
Xbit_r15_c9 bl_9 br_9 wl_15 vdd gnd cell_6t
Xbit_r16_c9 bl_9 br_9 wl_16 vdd gnd cell_6t
Xbit_r17_c9 bl_9 br_9 wl_17 vdd gnd cell_6t
Xbit_r18_c9 bl_9 br_9 wl_18 vdd gnd cell_6t
Xbit_r19_c9 bl_9 br_9 wl_19 vdd gnd cell_6t
Xbit_r20_c9 bl_9 br_9 wl_20 vdd gnd cell_6t
Xbit_r21_c9 bl_9 br_9 wl_21 vdd gnd cell_6t
Xbit_r22_c9 bl_9 br_9 wl_22 vdd gnd cell_6t
Xbit_r23_c9 bl_9 br_9 wl_23 vdd gnd cell_6t
Xbit_r24_c9 bl_9 br_9 wl_24 vdd gnd cell_6t
Xbit_r25_c9 bl_9 br_9 wl_25 vdd gnd cell_6t
Xbit_r26_c9 bl_9 br_9 wl_26 vdd gnd cell_6t
Xbit_r27_c9 bl_9 br_9 wl_27 vdd gnd cell_6t
Xbit_r28_c9 bl_9 br_9 wl_28 vdd gnd cell_6t
Xbit_r29_c9 bl_9 br_9 wl_29 vdd gnd cell_6t
Xbit_r30_c9 bl_9 br_9 wl_30 vdd gnd cell_6t
Xbit_r31_c9 bl_9 br_9 wl_31 vdd gnd cell_6t
Xbit_r32_c9 bl_9 br_9 wl_32 vdd gnd cell_6t
Xbit_r33_c9 bl_9 br_9 wl_33 vdd gnd cell_6t
Xbit_r34_c9 bl_9 br_9 wl_34 vdd gnd cell_6t
Xbit_r35_c9 bl_9 br_9 wl_35 vdd gnd cell_6t
Xbit_r36_c9 bl_9 br_9 wl_36 vdd gnd cell_6t
Xbit_r37_c9 bl_9 br_9 wl_37 vdd gnd cell_6t
Xbit_r38_c9 bl_9 br_9 wl_38 vdd gnd cell_6t
Xbit_r39_c9 bl_9 br_9 wl_39 vdd gnd cell_6t
Xbit_r40_c9 bl_9 br_9 wl_40 vdd gnd cell_6t
Xbit_r41_c9 bl_9 br_9 wl_41 vdd gnd cell_6t
Xbit_r42_c9 bl_9 br_9 wl_42 vdd gnd cell_6t
Xbit_r43_c9 bl_9 br_9 wl_43 vdd gnd cell_6t
Xbit_r44_c9 bl_9 br_9 wl_44 vdd gnd cell_6t
Xbit_r45_c9 bl_9 br_9 wl_45 vdd gnd cell_6t
Xbit_r46_c9 bl_9 br_9 wl_46 vdd gnd cell_6t
Xbit_r47_c9 bl_9 br_9 wl_47 vdd gnd cell_6t
Xbit_r48_c9 bl_9 br_9 wl_48 vdd gnd cell_6t
Xbit_r49_c9 bl_9 br_9 wl_49 vdd gnd cell_6t
Xbit_r50_c9 bl_9 br_9 wl_50 vdd gnd cell_6t
Xbit_r51_c9 bl_9 br_9 wl_51 vdd gnd cell_6t
Xbit_r52_c9 bl_9 br_9 wl_52 vdd gnd cell_6t
Xbit_r53_c9 bl_9 br_9 wl_53 vdd gnd cell_6t
Xbit_r54_c9 bl_9 br_9 wl_54 vdd gnd cell_6t
Xbit_r55_c9 bl_9 br_9 wl_55 vdd gnd cell_6t
Xbit_r56_c9 bl_9 br_9 wl_56 vdd gnd cell_6t
Xbit_r57_c9 bl_9 br_9 wl_57 vdd gnd cell_6t
Xbit_r58_c9 bl_9 br_9 wl_58 vdd gnd cell_6t
Xbit_r59_c9 bl_9 br_9 wl_59 vdd gnd cell_6t
Xbit_r60_c9 bl_9 br_9 wl_60 vdd gnd cell_6t
Xbit_r61_c9 bl_9 br_9 wl_61 vdd gnd cell_6t
Xbit_r62_c9 bl_9 br_9 wl_62 vdd gnd cell_6t
Xbit_r63_c9 bl_9 br_9 wl_63 vdd gnd cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd cell_6t
Xbit_r1_c10 bl_10 br_10 wl_1 vdd gnd cell_6t
Xbit_r2_c10 bl_10 br_10 wl_2 vdd gnd cell_6t
Xbit_r3_c10 bl_10 br_10 wl_3 vdd gnd cell_6t
Xbit_r4_c10 bl_10 br_10 wl_4 vdd gnd cell_6t
Xbit_r5_c10 bl_10 br_10 wl_5 vdd gnd cell_6t
Xbit_r6_c10 bl_10 br_10 wl_6 vdd gnd cell_6t
Xbit_r7_c10 bl_10 br_10 wl_7 vdd gnd cell_6t
Xbit_r8_c10 bl_10 br_10 wl_8 vdd gnd cell_6t
Xbit_r9_c10 bl_10 br_10 wl_9 vdd gnd cell_6t
Xbit_r10_c10 bl_10 br_10 wl_10 vdd gnd cell_6t
Xbit_r11_c10 bl_10 br_10 wl_11 vdd gnd cell_6t
Xbit_r12_c10 bl_10 br_10 wl_12 vdd gnd cell_6t
Xbit_r13_c10 bl_10 br_10 wl_13 vdd gnd cell_6t
Xbit_r14_c10 bl_10 br_10 wl_14 vdd gnd cell_6t
Xbit_r15_c10 bl_10 br_10 wl_15 vdd gnd cell_6t
Xbit_r16_c10 bl_10 br_10 wl_16 vdd gnd cell_6t
Xbit_r17_c10 bl_10 br_10 wl_17 vdd gnd cell_6t
Xbit_r18_c10 bl_10 br_10 wl_18 vdd gnd cell_6t
Xbit_r19_c10 bl_10 br_10 wl_19 vdd gnd cell_6t
Xbit_r20_c10 bl_10 br_10 wl_20 vdd gnd cell_6t
Xbit_r21_c10 bl_10 br_10 wl_21 vdd gnd cell_6t
Xbit_r22_c10 bl_10 br_10 wl_22 vdd gnd cell_6t
Xbit_r23_c10 bl_10 br_10 wl_23 vdd gnd cell_6t
Xbit_r24_c10 bl_10 br_10 wl_24 vdd gnd cell_6t
Xbit_r25_c10 bl_10 br_10 wl_25 vdd gnd cell_6t
Xbit_r26_c10 bl_10 br_10 wl_26 vdd gnd cell_6t
Xbit_r27_c10 bl_10 br_10 wl_27 vdd gnd cell_6t
Xbit_r28_c10 bl_10 br_10 wl_28 vdd gnd cell_6t
Xbit_r29_c10 bl_10 br_10 wl_29 vdd gnd cell_6t
Xbit_r30_c10 bl_10 br_10 wl_30 vdd gnd cell_6t
Xbit_r31_c10 bl_10 br_10 wl_31 vdd gnd cell_6t
Xbit_r32_c10 bl_10 br_10 wl_32 vdd gnd cell_6t
Xbit_r33_c10 bl_10 br_10 wl_33 vdd gnd cell_6t
Xbit_r34_c10 bl_10 br_10 wl_34 vdd gnd cell_6t
Xbit_r35_c10 bl_10 br_10 wl_35 vdd gnd cell_6t
Xbit_r36_c10 bl_10 br_10 wl_36 vdd gnd cell_6t
Xbit_r37_c10 bl_10 br_10 wl_37 vdd gnd cell_6t
Xbit_r38_c10 bl_10 br_10 wl_38 vdd gnd cell_6t
Xbit_r39_c10 bl_10 br_10 wl_39 vdd gnd cell_6t
Xbit_r40_c10 bl_10 br_10 wl_40 vdd gnd cell_6t
Xbit_r41_c10 bl_10 br_10 wl_41 vdd gnd cell_6t
Xbit_r42_c10 bl_10 br_10 wl_42 vdd gnd cell_6t
Xbit_r43_c10 bl_10 br_10 wl_43 vdd gnd cell_6t
Xbit_r44_c10 bl_10 br_10 wl_44 vdd gnd cell_6t
Xbit_r45_c10 bl_10 br_10 wl_45 vdd gnd cell_6t
Xbit_r46_c10 bl_10 br_10 wl_46 vdd gnd cell_6t
Xbit_r47_c10 bl_10 br_10 wl_47 vdd gnd cell_6t
Xbit_r48_c10 bl_10 br_10 wl_48 vdd gnd cell_6t
Xbit_r49_c10 bl_10 br_10 wl_49 vdd gnd cell_6t
Xbit_r50_c10 bl_10 br_10 wl_50 vdd gnd cell_6t
Xbit_r51_c10 bl_10 br_10 wl_51 vdd gnd cell_6t
Xbit_r52_c10 bl_10 br_10 wl_52 vdd gnd cell_6t
Xbit_r53_c10 bl_10 br_10 wl_53 vdd gnd cell_6t
Xbit_r54_c10 bl_10 br_10 wl_54 vdd gnd cell_6t
Xbit_r55_c10 bl_10 br_10 wl_55 vdd gnd cell_6t
Xbit_r56_c10 bl_10 br_10 wl_56 vdd gnd cell_6t
Xbit_r57_c10 bl_10 br_10 wl_57 vdd gnd cell_6t
Xbit_r58_c10 bl_10 br_10 wl_58 vdd gnd cell_6t
Xbit_r59_c10 bl_10 br_10 wl_59 vdd gnd cell_6t
Xbit_r60_c10 bl_10 br_10 wl_60 vdd gnd cell_6t
Xbit_r61_c10 bl_10 br_10 wl_61 vdd gnd cell_6t
Xbit_r62_c10 bl_10 br_10 wl_62 vdd gnd cell_6t
Xbit_r63_c10 bl_10 br_10 wl_63 vdd gnd cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd cell_6t
Xbit_r1_c11 bl_11 br_11 wl_1 vdd gnd cell_6t
Xbit_r2_c11 bl_11 br_11 wl_2 vdd gnd cell_6t
Xbit_r3_c11 bl_11 br_11 wl_3 vdd gnd cell_6t
Xbit_r4_c11 bl_11 br_11 wl_4 vdd gnd cell_6t
Xbit_r5_c11 bl_11 br_11 wl_5 vdd gnd cell_6t
Xbit_r6_c11 bl_11 br_11 wl_6 vdd gnd cell_6t
Xbit_r7_c11 bl_11 br_11 wl_7 vdd gnd cell_6t
Xbit_r8_c11 bl_11 br_11 wl_8 vdd gnd cell_6t
Xbit_r9_c11 bl_11 br_11 wl_9 vdd gnd cell_6t
Xbit_r10_c11 bl_11 br_11 wl_10 vdd gnd cell_6t
Xbit_r11_c11 bl_11 br_11 wl_11 vdd gnd cell_6t
Xbit_r12_c11 bl_11 br_11 wl_12 vdd gnd cell_6t
Xbit_r13_c11 bl_11 br_11 wl_13 vdd gnd cell_6t
Xbit_r14_c11 bl_11 br_11 wl_14 vdd gnd cell_6t
Xbit_r15_c11 bl_11 br_11 wl_15 vdd gnd cell_6t
Xbit_r16_c11 bl_11 br_11 wl_16 vdd gnd cell_6t
Xbit_r17_c11 bl_11 br_11 wl_17 vdd gnd cell_6t
Xbit_r18_c11 bl_11 br_11 wl_18 vdd gnd cell_6t
Xbit_r19_c11 bl_11 br_11 wl_19 vdd gnd cell_6t
Xbit_r20_c11 bl_11 br_11 wl_20 vdd gnd cell_6t
Xbit_r21_c11 bl_11 br_11 wl_21 vdd gnd cell_6t
Xbit_r22_c11 bl_11 br_11 wl_22 vdd gnd cell_6t
Xbit_r23_c11 bl_11 br_11 wl_23 vdd gnd cell_6t
Xbit_r24_c11 bl_11 br_11 wl_24 vdd gnd cell_6t
Xbit_r25_c11 bl_11 br_11 wl_25 vdd gnd cell_6t
Xbit_r26_c11 bl_11 br_11 wl_26 vdd gnd cell_6t
Xbit_r27_c11 bl_11 br_11 wl_27 vdd gnd cell_6t
Xbit_r28_c11 bl_11 br_11 wl_28 vdd gnd cell_6t
Xbit_r29_c11 bl_11 br_11 wl_29 vdd gnd cell_6t
Xbit_r30_c11 bl_11 br_11 wl_30 vdd gnd cell_6t
Xbit_r31_c11 bl_11 br_11 wl_31 vdd gnd cell_6t
Xbit_r32_c11 bl_11 br_11 wl_32 vdd gnd cell_6t
Xbit_r33_c11 bl_11 br_11 wl_33 vdd gnd cell_6t
Xbit_r34_c11 bl_11 br_11 wl_34 vdd gnd cell_6t
Xbit_r35_c11 bl_11 br_11 wl_35 vdd gnd cell_6t
Xbit_r36_c11 bl_11 br_11 wl_36 vdd gnd cell_6t
Xbit_r37_c11 bl_11 br_11 wl_37 vdd gnd cell_6t
Xbit_r38_c11 bl_11 br_11 wl_38 vdd gnd cell_6t
Xbit_r39_c11 bl_11 br_11 wl_39 vdd gnd cell_6t
Xbit_r40_c11 bl_11 br_11 wl_40 vdd gnd cell_6t
Xbit_r41_c11 bl_11 br_11 wl_41 vdd gnd cell_6t
Xbit_r42_c11 bl_11 br_11 wl_42 vdd gnd cell_6t
Xbit_r43_c11 bl_11 br_11 wl_43 vdd gnd cell_6t
Xbit_r44_c11 bl_11 br_11 wl_44 vdd gnd cell_6t
Xbit_r45_c11 bl_11 br_11 wl_45 vdd gnd cell_6t
Xbit_r46_c11 bl_11 br_11 wl_46 vdd gnd cell_6t
Xbit_r47_c11 bl_11 br_11 wl_47 vdd gnd cell_6t
Xbit_r48_c11 bl_11 br_11 wl_48 vdd gnd cell_6t
Xbit_r49_c11 bl_11 br_11 wl_49 vdd gnd cell_6t
Xbit_r50_c11 bl_11 br_11 wl_50 vdd gnd cell_6t
Xbit_r51_c11 bl_11 br_11 wl_51 vdd gnd cell_6t
Xbit_r52_c11 bl_11 br_11 wl_52 vdd gnd cell_6t
Xbit_r53_c11 bl_11 br_11 wl_53 vdd gnd cell_6t
Xbit_r54_c11 bl_11 br_11 wl_54 vdd gnd cell_6t
Xbit_r55_c11 bl_11 br_11 wl_55 vdd gnd cell_6t
Xbit_r56_c11 bl_11 br_11 wl_56 vdd gnd cell_6t
Xbit_r57_c11 bl_11 br_11 wl_57 vdd gnd cell_6t
Xbit_r58_c11 bl_11 br_11 wl_58 vdd gnd cell_6t
Xbit_r59_c11 bl_11 br_11 wl_59 vdd gnd cell_6t
Xbit_r60_c11 bl_11 br_11 wl_60 vdd gnd cell_6t
Xbit_r61_c11 bl_11 br_11 wl_61 vdd gnd cell_6t
Xbit_r62_c11 bl_11 br_11 wl_62 vdd gnd cell_6t
Xbit_r63_c11 bl_11 br_11 wl_63 vdd gnd cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd cell_6t
Xbit_r1_c12 bl_12 br_12 wl_1 vdd gnd cell_6t
Xbit_r2_c12 bl_12 br_12 wl_2 vdd gnd cell_6t
Xbit_r3_c12 bl_12 br_12 wl_3 vdd gnd cell_6t
Xbit_r4_c12 bl_12 br_12 wl_4 vdd gnd cell_6t
Xbit_r5_c12 bl_12 br_12 wl_5 vdd gnd cell_6t
Xbit_r6_c12 bl_12 br_12 wl_6 vdd gnd cell_6t
Xbit_r7_c12 bl_12 br_12 wl_7 vdd gnd cell_6t
Xbit_r8_c12 bl_12 br_12 wl_8 vdd gnd cell_6t
Xbit_r9_c12 bl_12 br_12 wl_9 vdd gnd cell_6t
Xbit_r10_c12 bl_12 br_12 wl_10 vdd gnd cell_6t
Xbit_r11_c12 bl_12 br_12 wl_11 vdd gnd cell_6t
Xbit_r12_c12 bl_12 br_12 wl_12 vdd gnd cell_6t
Xbit_r13_c12 bl_12 br_12 wl_13 vdd gnd cell_6t
Xbit_r14_c12 bl_12 br_12 wl_14 vdd gnd cell_6t
Xbit_r15_c12 bl_12 br_12 wl_15 vdd gnd cell_6t
Xbit_r16_c12 bl_12 br_12 wl_16 vdd gnd cell_6t
Xbit_r17_c12 bl_12 br_12 wl_17 vdd gnd cell_6t
Xbit_r18_c12 bl_12 br_12 wl_18 vdd gnd cell_6t
Xbit_r19_c12 bl_12 br_12 wl_19 vdd gnd cell_6t
Xbit_r20_c12 bl_12 br_12 wl_20 vdd gnd cell_6t
Xbit_r21_c12 bl_12 br_12 wl_21 vdd gnd cell_6t
Xbit_r22_c12 bl_12 br_12 wl_22 vdd gnd cell_6t
Xbit_r23_c12 bl_12 br_12 wl_23 vdd gnd cell_6t
Xbit_r24_c12 bl_12 br_12 wl_24 vdd gnd cell_6t
Xbit_r25_c12 bl_12 br_12 wl_25 vdd gnd cell_6t
Xbit_r26_c12 bl_12 br_12 wl_26 vdd gnd cell_6t
Xbit_r27_c12 bl_12 br_12 wl_27 vdd gnd cell_6t
Xbit_r28_c12 bl_12 br_12 wl_28 vdd gnd cell_6t
Xbit_r29_c12 bl_12 br_12 wl_29 vdd gnd cell_6t
Xbit_r30_c12 bl_12 br_12 wl_30 vdd gnd cell_6t
Xbit_r31_c12 bl_12 br_12 wl_31 vdd gnd cell_6t
Xbit_r32_c12 bl_12 br_12 wl_32 vdd gnd cell_6t
Xbit_r33_c12 bl_12 br_12 wl_33 vdd gnd cell_6t
Xbit_r34_c12 bl_12 br_12 wl_34 vdd gnd cell_6t
Xbit_r35_c12 bl_12 br_12 wl_35 vdd gnd cell_6t
Xbit_r36_c12 bl_12 br_12 wl_36 vdd gnd cell_6t
Xbit_r37_c12 bl_12 br_12 wl_37 vdd gnd cell_6t
Xbit_r38_c12 bl_12 br_12 wl_38 vdd gnd cell_6t
Xbit_r39_c12 bl_12 br_12 wl_39 vdd gnd cell_6t
Xbit_r40_c12 bl_12 br_12 wl_40 vdd gnd cell_6t
Xbit_r41_c12 bl_12 br_12 wl_41 vdd gnd cell_6t
Xbit_r42_c12 bl_12 br_12 wl_42 vdd gnd cell_6t
Xbit_r43_c12 bl_12 br_12 wl_43 vdd gnd cell_6t
Xbit_r44_c12 bl_12 br_12 wl_44 vdd gnd cell_6t
Xbit_r45_c12 bl_12 br_12 wl_45 vdd gnd cell_6t
Xbit_r46_c12 bl_12 br_12 wl_46 vdd gnd cell_6t
Xbit_r47_c12 bl_12 br_12 wl_47 vdd gnd cell_6t
Xbit_r48_c12 bl_12 br_12 wl_48 vdd gnd cell_6t
Xbit_r49_c12 bl_12 br_12 wl_49 vdd gnd cell_6t
Xbit_r50_c12 bl_12 br_12 wl_50 vdd gnd cell_6t
Xbit_r51_c12 bl_12 br_12 wl_51 vdd gnd cell_6t
Xbit_r52_c12 bl_12 br_12 wl_52 vdd gnd cell_6t
Xbit_r53_c12 bl_12 br_12 wl_53 vdd gnd cell_6t
Xbit_r54_c12 bl_12 br_12 wl_54 vdd gnd cell_6t
Xbit_r55_c12 bl_12 br_12 wl_55 vdd gnd cell_6t
Xbit_r56_c12 bl_12 br_12 wl_56 vdd gnd cell_6t
Xbit_r57_c12 bl_12 br_12 wl_57 vdd gnd cell_6t
Xbit_r58_c12 bl_12 br_12 wl_58 vdd gnd cell_6t
Xbit_r59_c12 bl_12 br_12 wl_59 vdd gnd cell_6t
Xbit_r60_c12 bl_12 br_12 wl_60 vdd gnd cell_6t
Xbit_r61_c12 bl_12 br_12 wl_61 vdd gnd cell_6t
Xbit_r62_c12 bl_12 br_12 wl_62 vdd gnd cell_6t
Xbit_r63_c12 bl_12 br_12 wl_63 vdd gnd cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd cell_6t
Xbit_r1_c13 bl_13 br_13 wl_1 vdd gnd cell_6t
Xbit_r2_c13 bl_13 br_13 wl_2 vdd gnd cell_6t
Xbit_r3_c13 bl_13 br_13 wl_3 vdd gnd cell_6t
Xbit_r4_c13 bl_13 br_13 wl_4 vdd gnd cell_6t
Xbit_r5_c13 bl_13 br_13 wl_5 vdd gnd cell_6t
Xbit_r6_c13 bl_13 br_13 wl_6 vdd gnd cell_6t
Xbit_r7_c13 bl_13 br_13 wl_7 vdd gnd cell_6t
Xbit_r8_c13 bl_13 br_13 wl_8 vdd gnd cell_6t
Xbit_r9_c13 bl_13 br_13 wl_9 vdd gnd cell_6t
Xbit_r10_c13 bl_13 br_13 wl_10 vdd gnd cell_6t
Xbit_r11_c13 bl_13 br_13 wl_11 vdd gnd cell_6t
Xbit_r12_c13 bl_13 br_13 wl_12 vdd gnd cell_6t
Xbit_r13_c13 bl_13 br_13 wl_13 vdd gnd cell_6t
Xbit_r14_c13 bl_13 br_13 wl_14 vdd gnd cell_6t
Xbit_r15_c13 bl_13 br_13 wl_15 vdd gnd cell_6t
Xbit_r16_c13 bl_13 br_13 wl_16 vdd gnd cell_6t
Xbit_r17_c13 bl_13 br_13 wl_17 vdd gnd cell_6t
Xbit_r18_c13 bl_13 br_13 wl_18 vdd gnd cell_6t
Xbit_r19_c13 bl_13 br_13 wl_19 vdd gnd cell_6t
Xbit_r20_c13 bl_13 br_13 wl_20 vdd gnd cell_6t
Xbit_r21_c13 bl_13 br_13 wl_21 vdd gnd cell_6t
Xbit_r22_c13 bl_13 br_13 wl_22 vdd gnd cell_6t
Xbit_r23_c13 bl_13 br_13 wl_23 vdd gnd cell_6t
Xbit_r24_c13 bl_13 br_13 wl_24 vdd gnd cell_6t
Xbit_r25_c13 bl_13 br_13 wl_25 vdd gnd cell_6t
Xbit_r26_c13 bl_13 br_13 wl_26 vdd gnd cell_6t
Xbit_r27_c13 bl_13 br_13 wl_27 vdd gnd cell_6t
Xbit_r28_c13 bl_13 br_13 wl_28 vdd gnd cell_6t
Xbit_r29_c13 bl_13 br_13 wl_29 vdd gnd cell_6t
Xbit_r30_c13 bl_13 br_13 wl_30 vdd gnd cell_6t
Xbit_r31_c13 bl_13 br_13 wl_31 vdd gnd cell_6t
Xbit_r32_c13 bl_13 br_13 wl_32 vdd gnd cell_6t
Xbit_r33_c13 bl_13 br_13 wl_33 vdd gnd cell_6t
Xbit_r34_c13 bl_13 br_13 wl_34 vdd gnd cell_6t
Xbit_r35_c13 bl_13 br_13 wl_35 vdd gnd cell_6t
Xbit_r36_c13 bl_13 br_13 wl_36 vdd gnd cell_6t
Xbit_r37_c13 bl_13 br_13 wl_37 vdd gnd cell_6t
Xbit_r38_c13 bl_13 br_13 wl_38 vdd gnd cell_6t
Xbit_r39_c13 bl_13 br_13 wl_39 vdd gnd cell_6t
Xbit_r40_c13 bl_13 br_13 wl_40 vdd gnd cell_6t
Xbit_r41_c13 bl_13 br_13 wl_41 vdd gnd cell_6t
Xbit_r42_c13 bl_13 br_13 wl_42 vdd gnd cell_6t
Xbit_r43_c13 bl_13 br_13 wl_43 vdd gnd cell_6t
Xbit_r44_c13 bl_13 br_13 wl_44 vdd gnd cell_6t
Xbit_r45_c13 bl_13 br_13 wl_45 vdd gnd cell_6t
Xbit_r46_c13 bl_13 br_13 wl_46 vdd gnd cell_6t
Xbit_r47_c13 bl_13 br_13 wl_47 vdd gnd cell_6t
Xbit_r48_c13 bl_13 br_13 wl_48 vdd gnd cell_6t
Xbit_r49_c13 bl_13 br_13 wl_49 vdd gnd cell_6t
Xbit_r50_c13 bl_13 br_13 wl_50 vdd gnd cell_6t
Xbit_r51_c13 bl_13 br_13 wl_51 vdd gnd cell_6t
Xbit_r52_c13 bl_13 br_13 wl_52 vdd gnd cell_6t
Xbit_r53_c13 bl_13 br_13 wl_53 vdd gnd cell_6t
Xbit_r54_c13 bl_13 br_13 wl_54 vdd gnd cell_6t
Xbit_r55_c13 bl_13 br_13 wl_55 vdd gnd cell_6t
Xbit_r56_c13 bl_13 br_13 wl_56 vdd gnd cell_6t
Xbit_r57_c13 bl_13 br_13 wl_57 vdd gnd cell_6t
Xbit_r58_c13 bl_13 br_13 wl_58 vdd gnd cell_6t
Xbit_r59_c13 bl_13 br_13 wl_59 vdd gnd cell_6t
Xbit_r60_c13 bl_13 br_13 wl_60 vdd gnd cell_6t
Xbit_r61_c13 bl_13 br_13 wl_61 vdd gnd cell_6t
Xbit_r62_c13 bl_13 br_13 wl_62 vdd gnd cell_6t
Xbit_r63_c13 bl_13 br_13 wl_63 vdd gnd cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd cell_6t
Xbit_r1_c14 bl_14 br_14 wl_1 vdd gnd cell_6t
Xbit_r2_c14 bl_14 br_14 wl_2 vdd gnd cell_6t
Xbit_r3_c14 bl_14 br_14 wl_3 vdd gnd cell_6t
Xbit_r4_c14 bl_14 br_14 wl_4 vdd gnd cell_6t
Xbit_r5_c14 bl_14 br_14 wl_5 vdd gnd cell_6t
Xbit_r6_c14 bl_14 br_14 wl_6 vdd gnd cell_6t
Xbit_r7_c14 bl_14 br_14 wl_7 vdd gnd cell_6t
Xbit_r8_c14 bl_14 br_14 wl_8 vdd gnd cell_6t
Xbit_r9_c14 bl_14 br_14 wl_9 vdd gnd cell_6t
Xbit_r10_c14 bl_14 br_14 wl_10 vdd gnd cell_6t
Xbit_r11_c14 bl_14 br_14 wl_11 vdd gnd cell_6t
Xbit_r12_c14 bl_14 br_14 wl_12 vdd gnd cell_6t
Xbit_r13_c14 bl_14 br_14 wl_13 vdd gnd cell_6t
Xbit_r14_c14 bl_14 br_14 wl_14 vdd gnd cell_6t
Xbit_r15_c14 bl_14 br_14 wl_15 vdd gnd cell_6t
Xbit_r16_c14 bl_14 br_14 wl_16 vdd gnd cell_6t
Xbit_r17_c14 bl_14 br_14 wl_17 vdd gnd cell_6t
Xbit_r18_c14 bl_14 br_14 wl_18 vdd gnd cell_6t
Xbit_r19_c14 bl_14 br_14 wl_19 vdd gnd cell_6t
Xbit_r20_c14 bl_14 br_14 wl_20 vdd gnd cell_6t
Xbit_r21_c14 bl_14 br_14 wl_21 vdd gnd cell_6t
Xbit_r22_c14 bl_14 br_14 wl_22 vdd gnd cell_6t
Xbit_r23_c14 bl_14 br_14 wl_23 vdd gnd cell_6t
Xbit_r24_c14 bl_14 br_14 wl_24 vdd gnd cell_6t
Xbit_r25_c14 bl_14 br_14 wl_25 vdd gnd cell_6t
Xbit_r26_c14 bl_14 br_14 wl_26 vdd gnd cell_6t
Xbit_r27_c14 bl_14 br_14 wl_27 vdd gnd cell_6t
Xbit_r28_c14 bl_14 br_14 wl_28 vdd gnd cell_6t
Xbit_r29_c14 bl_14 br_14 wl_29 vdd gnd cell_6t
Xbit_r30_c14 bl_14 br_14 wl_30 vdd gnd cell_6t
Xbit_r31_c14 bl_14 br_14 wl_31 vdd gnd cell_6t
Xbit_r32_c14 bl_14 br_14 wl_32 vdd gnd cell_6t
Xbit_r33_c14 bl_14 br_14 wl_33 vdd gnd cell_6t
Xbit_r34_c14 bl_14 br_14 wl_34 vdd gnd cell_6t
Xbit_r35_c14 bl_14 br_14 wl_35 vdd gnd cell_6t
Xbit_r36_c14 bl_14 br_14 wl_36 vdd gnd cell_6t
Xbit_r37_c14 bl_14 br_14 wl_37 vdd gnd cell_6t
Xbit_r38_c14 bl_14 br_14 wl_38 vdd gnd cell_6t
Xbit_r39_c14 bl_14 br_14 wl_39 vdd gnd cell_6t
Xbit_r40_c14 bl_14 br_14 wl_40 vdd gnd cell_6t
Xbit_r41_c14 bl_14 br_14 wl_41 vdd gnd cell_6t
Xbit_r42_c14 bl_14 br_14 wl_42 vdd gnd cell_6t
Xbit_r43_c14 bl_14 br_14 wl_43 vdd gnd cell_6t
Xbit_r44_c14 bl_14 br_14 wl_44 vdd gnd cell_6t
Xbit_r45_c14 bl_14 br_14 wl_45 vdd gnd cell_6t
Xbit_r46_c14 bl_14 br_14 wl_46 vdd gnd cell_6t
Xbit_r47_c14 bl_14 br_14 wl_47 vdd gnd cell_6t
Xbit_r48_c14 bl_14 br_14 wl_48 vdd gnd cell_6t
Xbit_r49_c14 bl_14 br_14 wl_49 vdd gnd cell_6t
Xbit_r50_c14 bl_14 br_14 wl_50 vdd gnd cell_6t
Xbit_r51_c14 bl_14 br_14 wl_51 vdd gnd cell_6t
Xbit_r52_c14 bl_14 br_14 wl_52 vdd gnd cell_6t
Xbit_r53_c14 bl_14 br_14 wl_53 vdd gnd cell_6t
Xbit_r54_c14 bl_14 br_14 wl_54 vdd gnd cell_6t
Xbit_r55_c14 bl_14 br_14 wl_55 vdd gnd cell_6t
Xbit_r56_c14 bl_14 br_14 wl_56 vdd gnd cell_6t
Xbit_r57_c14 bl_14 br_14 wl_57 vdd gnd cell_6t
Xbit_r58_c14 bl_14 br_14 wl_58 vdd gnd cell_6t
Xbit_r59_c14 bl_14 br_14 wl_59 vdd gnd cell_6t
Xbit_r60_c14 bl_14 br_14 wl_60 vdd gnd cell_6t
Xbit_r61_c14 bl_14 br_14 wl_61 vdd gnd cell_6t
Xbit_r62_c14 bl_14 br_14 wl_62 vdd gnd cell_6t
Xbit_r63_c14 bl_14 br_14 wl_63 vdd gnd cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd cell_6t
Xbit_r1_c15 bl_15 br_15 wl_1 vdd gnd cell_6t
Xbit_r2_c15 bl_15 br_15 wl_2 vdd gnd cell_6t
Xbit_r3_c15 bl_15 br_15 wl_3 vdd gnd cell_6t
Xbit_r4_c15 bl_15 br_15 wl_4 vdd gnd cell_6t
Xbit_r5_c15 bl_15 br_15 wl_5 vdd gnd cell_6t
Xbit_r6_c15 bl_15 br_15 wl_6 vdd gnd cell_6t
Xbit_r7_c15 bl_15 br_15 wl_7 vdd gnd cell_6t
Xbit_r8_c15 bl_15 br_15 wl_8 vdd gnd cell_6t
Xbit_r9_c15 bl_15 br_15 wl_9 vdd gnd cell_6t
Xbit_r10_c15 bl_15 br_15 wl_10 vdd gnd cell_6t
Xbit_r11_c15 bl_15 br_15 wl_11 vdd gnd cell_6t
Xbit_r12_c15 bl_15 br_15 wl_12 vdd gnd cell_6t
Xbit_r13_c15 bl_15 br_15 wl_13 vdd gnd cell_6t
Xbit_r14_c15 bl_15 br_15 wl_14 vdd gnd cell_6t
Xbit_r15_c15 bl_15 br_15 wl_15 vdd gnd cell_6t
Xbit_r16_c15 bl_15 br_15 wl_16 vdd gnd cell_6t
Xbit_r17_c15 bl_15 br_15 wl_17 vdd gnd cell_6t
Xbit_r18_c15 bl_15 br_15 wl_18 vdd gnd cell_6t
Xbit_r19_c15 bl_15 br_15 wl_19 vdd gnd cell_6t
Xbit_r20_c15 bl_15 br_15 wl_20 vdd gnd cell_6t
Xbit_r21_c15 bl_15 br_15 wl_21 vdd gnd cell_6t
Xbit_r22_c15 bl_15 br_15 wl_22 vdd gnd cell_6t
Xbit_r23_c15 bl_15 br_15 wl_23 vdd gnd cell_6t
Xbit_r24_c15 bl_15 br_15 wl_24 vdd gnd cell_6t
Xbit_r25_c15 bl_15 br_15 wl_25 vdd gnd cell_6t
Xbit_r26_c15 bl_15 br_15 wl_26 vdd gnd cell_6t
Xbit_r27_c15 bl_15 br_15 wl_27 vdd gnd cell_6t
Xbit_r28_c15 bl_15 br_15 wl_28 vdd gnd cell_6t
Xbit_r29_c15 bl_15 br_15 wl_29 vdd gnd cell_6t
Xbit_r30_c15 bl_15 br_15 wl_30 vdd gnd cell_6t
Xbit_r31_c15 bl_15 br_15 wl_31 vdd gnd cell_6t
Xbit_r32_c15 bl_15 br_15 wl_32 vdd gnd cell_6t
Xbit_r33_c15 bl_15 br_15 wl_33 vdd gnd cell_6t
Xbit_r34_c15 bl_15 br_15 wl_34 vdd gnd cell_6t
Xbit_r35_c15 bl_15 br_15 wl_35 vdd gnd cell_6t
Xbit_r36_c15 bl_15 br_15 wl_36 vdd gnd cell_6t
Xbit_r37_c15 bl_15 br_15 wl_37 vdd gnd cell_6t
Xbit_r38_c15 bl_15 br_15 wl_38 vdd gnd cell_6t
Xbit_r39_c15 bl_15 br_15 wl_39 vdd gnd cell_6t
Xbit_r40_c15 bl_15 br_15 wl_40 vdd gnd cell_6t
Xbit_r41_c15 bl_15 br_15 wl_41 vdd gnd cell_6t
Xbit_r42_c15 bl_15 br_15 wl_42 vdd gnd cell_6t
Xbit_r43_c15 bl_15 br_15 wl_43 vdd gnd cell_6t
Xbit_r44_c15 bl_15 br_15 wl_44 vdd gnd cell_6t
Xbit_r45_c15 bl_15 br_15 wl_45 vdd gnd cell_6t
Xbit_r46_c15 bl_15 br_15 wl_46 vdd gnd cell_6t
Xbit_r47_c15 bl_15 br_15 wl_47 vdd gnd cell_6t
Xbit_r48_c15 bl_15 br_15 wl_48 vdd gnd cell_6t
Xbit_r49_c15 bl_15 br_15 wl_49 vdd gnd cell_6t
Xbit_r50_c15 bl_15 br_15 wl_50 vdd gnd cell_6t
Xbit_r51_c15 bl_15 br_15 wl_51 vdd gnd cell_6t
Xbit_r52_c15 bl_15 br_15 wl_52 vdd gnd cell_6t
Xbit_r53_c15 bl_15 br_15 wl_53 vdd gnd cell_6t
Xbit_r54_c15 bl_15 br_15 wl_54 vdd gnd cell_6t
Xbit_r55_c15 bl_15 br_15 wl_55 vdd gnd cell_6t
Xbit_r56_c15 bl_15 br_15 wl_56 vdd gnd cell_6t
Xbit_r57_c15 bl_15 br_15 wl_57 vdd gnd cell_6t
Xbit_r58_c15 bl_15 br_15 wl_58 vdd gnd cell_6t
Xbit_r59_c15 bl_15 br_15 wl_59 vdd gnd cell_6t
Xbit_r60_c15 bl_15 br_15 wl_60 vdd gnd cell_6t
Xbit_r61_c15 bl_15 br_15 wl_61 vdd gnd cell_6t
Xbit_r62_c15 bl_15 br_15 wl_62 vdd gnd cell_6t
Xbit_r63_c15 bl_15 br_15 wl_63 vdd gnd cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd cell_6t
Xbit_r1_c16 bl_16 br_16 wl_1 vdd gnd cell_6t
Xbit_r2_c16 bl_16 br_16 wl_2 vdd gnd cell_6t
Xbit_r3_c16 bl_16 br_16 wl_3 vdd gnd cell_6t
Xbit_r4_c16 bl_16 br_16 wl_4 vdd gnd cell_6t
Xbit_r5_c16 bl_16 br_16 wl_5 vdd gnd cell_6t
Xbit_r6_c16 bl_16 br_16 wl_6 vdd gnd cell_6t
Xbit_r7_c16 bl_16 br_16 wl_7 vdd gnd cell_6t
Xbit_r8_c16 bl_16 br_16 wl_8 vdd gnd cell_6t
Xbit_r9_c16 bl_16 br_16 wl_9 vdd gnd cell_6t
Xbit_r10_c16 bl_16 br_16 wl_10 vdd gnd cell_6t
Xbit_r11_c16 bl_16 br_16 wl_11 vdd gnd cell_6t
Xbit_r12_c16 bl_16 br_16 wl_12 vdd gnd cell_6t
Xbit_r13_c16 bl_16 br_16 wl_13 vdd gnd cell_6t
Xbit_r14_c16 bl_16 br_16 wl_14 vdd gnd cell_6t
Xbit_r15_c16 bl_16 br_16 wl_15 vdd gnd cell_6t
Xbit_r16_c16 bl_16 br_16 wl_16 vdd gnd cell_6t
Xbit_r17_c16 bl_16 br_16 wl_17 vdd gnd cell_6t
Xbit_r18_c16 bl_16 br_16 wl_18 vdd gnd cell_6t
Xbit_r19_c16 bl_16 br_16 wl_19 vdd gnd cell_6t
Xbit_r20_c16 bl_16 br_16 wl_20 vdd gnd cell_6t
Xbit_r21_c16 bl_16 br_16 wl_21 vdd gnd cell_6t
Xbit_r22_c16 bl_16 br_16 wl_22 vdd gnd cell_6t
Xbit_r23_c16 bl_16 br_16 wl_23 vdd gnd cell_6t
Xbit_r24_c16 bl_16 br_16 wl_24 vdd gnd cell_6t
Xbit_r25_c16 bl_16 br_16 wl_25 vdd gnd cell_6t
Xbit_r26_c16 bl_16 br_16 wl_26 vdd gnd cell_6t
Xbit_r27_c16 bl_16 br_16 wl_27 vdd gnd cell_6t
Xbit_r28_c16 bl_16 br_16 wl_28 vdd gnd cell_6t
Xbit_r29_c16 bl_16 br_16 wl_29 vdd gnd cell_6t
Xbit_r30_c16 bl_16 br_16 wl_30 vdd gnd cell_6t
Xbit_r31_c16 bl_16 br_16 wl_31 vdd gnd cell_6t
Xbit_r32_c16 bl_16 br_16 wl_32 vdd gnd cell_6t
Xbit_r33_c16 bl_16 br_16 wl_33 vdd gnd cell_6t
Xbit_r34_c16 bl_16 br_16 wl_34 vdd gnd cell_6t
Xbit_r35_c16 bl_16 br_16 wl_35 vdd gnd cell_6t
Xbit_r36_c16 bl_16 br_16 wl_36 vdd gnd cell_6t
Xbit_r37_c16 bl_16 br_16 wl_37 vdd gnd cell_6t
Xbit_r38_c16 bl_16 br_16 wl_38 vdd gnd cell_6t
Xbit_r39_c16 bl_16 br_16 wl_39 vdd gnd cell_6t
Xbit_r40_c16 bl_16 br_16 wl_40 vdd gnd cell_6t
Xbit_r41_c16 bl_16 br_16 wl_41 vdd gnd cell_6t
Xbit_r42_c16 bl_16 br_16 wl_42 vdd gnd cell_6t
Xbit_r43_c16 bl_16 br_16 wl_43 vdd gnd cell_6t
Xbit_r44_c16 bl_16 br_16 wl_44 vdd gnd cell_6t
Xbit_r45_c16 bl_16 br_16 wl_45 vdd gnd cell_6t
Xbit_r46_c16 bl_16 br_16 wl_46 vdd gnd cell_6t
Xbit_r47_c16 bl_16 br_16 wl_47 vdd gnd cell_6t
Xbit_r48_c16 bl_16 br_16 wl_48 vdd gnd cell_6t
Xbit_r49_c16 bl_16 br_16 wl_49 vdd gnd cell_6t
Xbit_r50_c16 bl_16 br_16 wl_50 vdd gnd cell_6t
Xbit_r51_c16 bl_16 br_16 wl_51 vdd gnd cell_6t
Xbit_r52_c16 bl_16 br_16 wl_52 vdd gnd cell_6t
Xbit_r53_c16 bl_16 br_16 wl_53 vdd gnd cell_6t
Xbit_r54_c16 bl_16 br_16 wl_54 vdd gnd cell_6t
Xbit_r55_c16 bl_16 br_16 wl_55 vdd gnd cell_6t
Xbit_r56_c16 bl_16 br_16 wl_56 vdd gnd cell_6t
Xbit_r57_c16 bl_16 br_16 wl_57 vdd gnd cell_6t
Xbit_r58_c16 bl_16 br_16 wl_58 vdd gnd cell_6t
Xbit_r59_c16 bl_16 br_16 wl_59 vdd gnd cell_6t
Xbit_r60_c16 bl_16 br_16 wl_60 vdd gnd cell_6t
Xbit_r61_c16 bl_16 br_16 wl_61 vdd gnd cell_6t
Xbit_r62_c16 bl_16 br_16 wl_62 vdd gnd cell_6t
Xbit_r63_c16 bl_16 br_16 wl_63 vdd gnd cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd cell_6t
Xbit_r1_c17 bl_17 br_17 wl_1 vdd gnd cell_6t
Xbit_r2_c17 bl_17 br_17 wl_2 vdd gnd cell_6t
Xbit_r3_c17 bl_17 br_17 wl_3 vdd gnd cell_6t
Xbit_r4_c17 bl_17 br_17 wl_4 vdd gnd cell_6t
Xbit_r5_c17 bl_17 br_17 wl_5 vdd gnd cell_6t
Xbit_r6_c17 bl_17 br_17 wl_6 vdd gnd cell_6t
Xbit_r7_c17 bl_17 br_17 wl_7 vdd gnd cell_6t
Xbit_r8_c17 bl_17 br_17 wl_8 vdd gnd cell_6t
Xbit_r9_c17 bl_17 br_17 wl_9 vdd gnd cell_6t
Xbit_r10_c17 bl_17 br_17 wl_10 vdd gnd cell_6t
Xbit_r11_c17 bl_17 br_17 wl_11 vdd gnd cell_6t
Xbit_r12_c17 bl_17 br_17 wl_12 vdd gnd cell_6t
Xbit_r13_c17 bl_17 br_17 wl_13 vdd gnd cell_6t
Xbit_r14_c17 bl_17 br_17 wl_14 vdd gnd cell_6t
Xbit_r15_c17 bl_17 br_17 wl_15 vdd gnd cell_6t
Xbit_r16_c17 bl_17 br_17 wl_16 vdd gnd cell_6t
Xbit_r17_c17 bl_17 br_17 wl_17 vdd gnd cell_6t
Xbit_r18_c17 bl_17 br_17 wl_18 vdd gnd cell_6t
Xbit_r19_c17 bl_17 br_17 wl_19 vdd gnd cell_6t
Xbit_r20_c17 bl_17 br_17 wl_20 vdd gnd cell_6t
Xbit_r21_c17 bl_17 br_17 wl_21 vdd gnd cell_6t
Xbit_r22_c17 bl_17 br_17 wl_22 vdd gnd cell_6t
Xbit_r23_c17 bl_17 br_17 wl_23 vdd gnd cell_6t
Xbit_r24_c17 bl_17 br_17 wl_24 vdd gnd cell_6t
Xbit_r25_c17 bl_17 br_17 wl_25 vdd gnd cell_6t
Xbit_r26_c17 bl_17 br_17 wl_26 vdd gnd cell_6t
Xbit_r27_c17 bl_17 br_17 wl_27 vdd gnd cell_6t
Xbit_r28_c17 bl_17 br_17 wl_28 vdd gnd cell_6t
Xbit_r29_c17 bl_17 br_17 wl_29 vdd gnd cell_6t
Xbit_r30_c17 bl_17 br_17 wl_30 vdd gnd cell_6t
Xbit_r31_c17 bl_17 br_17 wl_31 vdd gnd cell_6t
Xbit_r32_c17 bl_17 br_17 wl_32 vdd gnd cell_6t
Xbit_r33_c17 bl_17 br_17 wl_33 vdd gnd cell_6t
Xbit_r34_c17 bl_17 br_17 wl_34 vdd gnd cell_6t
Xbit_r35_c17 bl_17 br_17 wl_35 vdd gnd cell_6t
Xbit_r36_c17 bl_17 br_17 wl_36 vdd gnd cell_6t
Xbit_r37_c17 bl_17 br_17 wl_37 vdd gnd cell_6t
Xbit_r38_c17 bl_17 br_17 wl_38 vdd gnd cell_6t
Xbit_r39_c17 bl_17 br_17 wl_39 vdd gnd cell_6t
Xbit_r40_c17 bl_17 br_17 wl_40 vdd gnd cell_6t
Xbit_r41_c17 bl_17 br_17 wl_41 vdd gnd cell_6t
Xbit_r42_c17 bl_17 br_17 wl_42 vdd gnd cell_6t
Xbit_r43_c17 bl_17 br_17 wl_43 vdd gnd cell_6t
Xbit_r44_c17 bl_17 br_17 wl_44 vdd gnd cell_6t
Xbit_r45_c17 bl_17 br_17 wl_45 vdd gnd cell_6t
Xbit_r46_c17 bl_17 br_17 wl_46 vdd gnd cell_6t
Xbit_r47_c17 bl_17 br_17 wl_47 vdd gnd cell_6t
Xbit_r48_c17 bl_17 br_17 wl_48 vdd gnd cell_6t
Xbit_r49_c17 bl_17 br_17 wl_49 vdd gnd cell_6t
Xbit_r50_c17 bl_17 br_17 wl_50 vdd gnd cell_6t
Xbit_r51_c17 bl_17 br_17 wl_51 vdd gnd cell_6t
Xbit_r52_c17 bl_17 br_17 wl_52 vdd gnd cell_6t
Xbit_r53_c17 bl_17 br_17 wl_53 vdd gnd cell_6t
Xbit_r54_c17 bl_17 br_17 wl_54 vdd gnd cell_6t
Xbit_r55_c17 bl_17 br_17 wl_55 vdd gnd cell_6t
Xbit_r56_c17 bl_17 br_17 wl_56 vdd gnd cell_6t
Xbit_r57_c17 bl_17 br_17 wl_57 vdd gnd cell_6t
Xbit_r58_c17 bl_17 br_17 wl_58 vdd gnd cell_6t
Xbit_r59_c17 bl_17 br_17 wl_59 vdd gnd cell_6t
Xbit_r60_c17 bl_17 br_17 wl_60 vdd gnd cell_6t
Xbit_r61_c17 bl_17 br_17 wl_61 vdd gnd cell_6t
Xbit_r62_c17 bl_17 br_17 wl_62 vdd gnd cell_6t
Xbit_r63_c17 bl_17 br_17 wl_63 vdd gnd cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd cell_6t
Xbit_r1_c18 bl_18 br_18 wl_1 vdd gnd cell_6t
Xbit_r2_c18 bl_18 br_18 wl_2 vdd gnd cell_6t
Xbit_r3_c18 bl_18 br_18 wl_3 vdd gnd cell_6t
Xbit_r4_c18 bl_18 br_18 wl_4 vdd gnd cell_6t
Xbit_r5_c18 bl_18 br_18 wl_5 vdd gnd cell_6t
Xbit_r6_c18 bl_18 br_18 wl_6 vdd gnd cell_6t
Xbit_r7_c18 bl_18 br_18 wl_7 vdd gnd cell_6t
Xbit_r8_c18 bl_18 br_18 wl_8 vdd gnd cell_6t
Xbit_r9_c18 bl_18 br_18 wl_9 vdd gnd cell_6t
Xbit_r10_c18 bl_18 br_18 wl_10 vdd gnd cell_6t
Xbit_r11_c18 bl_18 br_18 wl_11 vdd gnd cell_6t
Xbit_r12_c18 bl_18 br_18 wl_12 vdd gnd cell_6t
Xbit_r13_c18 bl_18 br_18 wl_13 vdd gnd cell_6t
Xbit_r14_c18 bl_18 br_18 wl_14 vdd gnd cell_6t
Xbit_r15_c18 bl_18 br_18 wl_15 vdd gnd cell_6t
Xbit_r16_c18 bl_18 br_18 wl_16 vdd gnd cell_6t
Xbit_r17_c18 bl_18 br_18 wl_17 vdd gnd cell_6t
Xbit_r18_c18 bl_18 br_18 wl_18 vdd gnd cell_6t
Xbit_r19_c18 bl_18 br_18 wl_19 vdd gnd cell_6t
Xbit_r20_c18 bl_18 br_18 wl_20 vdd gnd cell_6t
Xbit_r21_c18 bl_18 br_18 wl_21 vdd gnd cell_6t
Xbit_r22_c18 bl_18 br_18 wl_22 vdd gnd cell_6t
Xbit_r23_c18 bl_18 br_18 wl_23 vdd gnd cell_6t
Xbit_r24_c18 bl_18 br_18 wl_24 vdd gnd cell_6t
Xbit_r25_c18 bl_18 br_18 wl_25 vdd gnd cell_6t
Xbit_r26_c18 bl_18 br_18 wl_26 vdd gnd cell_6t
Xbit_r27_c18 bl_18 br_18 wl_27 vdd gnd cell_6t
Xbit_r28_c18 bl_18 br_18 wl_28 vdd gnd cell_6t
Xbit_r29_c18 bl_18 br_18 wl_29 vdd gnd cell_6t
Xbit_r30_c18 bl_18 br_18 wl_30 vdd gnd cell_6t
Xbit_r31_c18 bl_18 br_18 wl_31 vdd gnd cell_6t
Xbit_r32_c18 bl_18 br_18 wl_32 vdd gnd cell_6t
Xbit_r33_c18 bl_18 br_18 wl_33 vdd gnd cell_6t
Xbit_r34_c18 bl_18 br_18 wl_34 vdd gnd cell_6t
Xbit_r35_c18 bl_18 br_18 wl_35 vdd gnd cell_6t
Xbit_r36_c18 bl_18 br_18 wl_36 vdd gnd cell_6t
Xbit_r37_c18 bl_18 br_18 wl_37 vdd gnd cell_6t
Xbit_r38_c18 bl_18 br_18 wl_38 vdd gnd cell_6t
Xbit_r39_c18 bl_18 br_18 wl_39 vdd gnd cell_6t
Xbit_r40_c18 bl_18 br_18 wl_40 vdd gnd cell_6t
Xbit_r41_c18 bl_18 br_18 wl_41 vdd gnd cell_6t
Xbit_r42_c18 bl_18 br_18 wl_42 vdd gnd cell_6t
Xbit_r43_c18 bl_18 br_18 wl_43 vdd gnd cell_6t
Xbit_r44_c18 bl_18 br_18 wl_44 vdd gnd cell_6t
Xbit_r45_c18 bl_18 br_18 wl_45 vdd gnd cell_6t
Xbit_r46_c18 bl_18 br_18 wl_46 vdd gnd cell_6t
Xbit_r47_c18 bl_18 br_18 wl_47 vdd gnd cell_6t
Xbit_r48_c18 bl_18 br_18 wl_48 vdd gnd cell_6t
Xbit_r49_c18 bl_18 br_18 wl_49 vdd gnd cell_6t
Xbit_r50_c18 bl_18 br_18 wl_50 vdd gnd cell_6t
Xbit_r51_c18 bl_18 br_18 wl_51 vdd gnd cell_6t
Xbit_r52_c18 bl_18 br_18 wl_52 vdd gnd cell_6t
Xbit_r53_c18 bl_18 br_18 wl_53 vdd gnd cell_6t
Xbit_r54_c18 bl_18 br_18 wl_54 vdd gnd cell_6t
Xbit_r55_c18 bl_18 br_18 wl_55 vdd gnd cell_6t
Xbit_r56_c18 bl_18 br_18 wl_56 vdd gnd cell_6t
Xbit_r57_c18 bl_18 br_18 wl_57 vdd gnd cell_6t
Xbit_r58_c18 bl_18 br_18 wl_58 vdd gnd cell_6t
Xbit_r59_c18 bl_18 br_18 wl_59 vdd gnd cell_6t
Xbit_r60_c18 bl_18 br_18 wl_60 vdd gnd cell_6t
Xbit_r61_c18 bl_18 br_18 wl_61 vdd gnd cell_6t
Xbit_r62_c18 bl_18 br_18 wl_62 vdd gnd cell_6t
Xbit_r63_c18 bl_18 br_18 wl_63 vdd gnd cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd cell_6t
Xbit_r1_c19 bl_19 br_19 wl_1 vdd gnd cell_6t
Xbit_r2_c19 bl_19 br_19 wl_2 vdd gnd cell_6t
Xbit_r3_c19 bl_19 br_19 wl_3 vdd gnd cell_6t
Xbit_r4_c19 bl_19 br_19 wl_4 vdd gnd cell_6t
Xbit_r5_c19 bl_19 br_19 wl_5 vdd gnd cell_6t
Xbit_r6_c19 bl_19 br_19 wl_6 vdd gnd cell_6t
Xbit_r7_c19 bl_19 br_19 wl_7 vdd gnd cell_6t
Xbit_r8_c19 bl_19 br_19 wl_8 vdd gnd cell_6t
Xbit_r9_c19 bl_19 br_19 wl_9 vdd gnd cell_6t
Xbit_r10_c19 bl_19 br_19 wl_10 vdd gnd cell_6t
Xbit_r11_c19 bl_19 br_19 wl_11 vdd gnd cell_6t
Xbit_r12_c19 bl_19 br_19 wl_12 vdd gnd cell_6t
Xbit_r13_c19 bl_19 br_19 wl_13 vdd gnd cell_6t
Xbit_r14_c19 bl_19 br_19 wl_14 vdd gnd cell_6t
Xbit_r15_c19 bl_19 br_19 wl_15 vdd gnd cell_6t
Xbit_r16_c19 bl_19 br_19 wl_16 vdd gnd cell_6t
Xbit_r17_c19 bl_19 br_19 wl_17 vdd gnd cell_6t
Xbit_r18_c19 bl_19 br_19 wl_18 vdd gnd cell_6t
Xbit_r19_c19 bl_19 br_19 wl_19 vdd gnd cell_6t
Xbit_r20_c19 bl_19 br_19 wl_20 vdd gnd cell_6t
Xbit_r21_c19 bl_19 br_19 wl_21 vdd gnd cell_6t
Xbit_r22_c19 bl_19 br_19 wl_22 vdd gnd cell_6t
Xbit_r23_c19 bl_19 br_19 wl_23 vdd gnd cell_6t
Xbit_r24_c19 bl_19 br_19 wl_24 vdd gnd cell_6t
Xbit_r25_c19 bl_19 br_19 wl_25 vdd gnd cell_6t
Xbit_r26_c19 bl_19 br_19 wl_26 vdd gnd cell_6t
Xbit_r27_c19 bl_19 br_19 wl_27 vdd gnd cell_6t
Xbit_r28_c19 bl_19 br_19 wl_28 vdd gnd cell_6t
Xbit_r29_c19 bl_19 br_19 wl_29 vdd gnd cell_6t
Xbit_r30_c19 bl_19 br_19 wl_30 vdd gnd cell_6t
Xbit_r31_c19 bl_19 br_19 wl_31 vdd gnd cell_6t
Xbit_r32_c19 bl_19 br_19 wl_32 vdd gnd cell_6t
Xbit_r33_c19 bl_19 br_19 wl_33 vdd gnd cell_6t
Xbit_r34_c19 bl_19 br_19 wl_34 vdd gnd cell_6t
Xbit_r35_c19 bl_19 br_19 wl_35 vdd gnd cell_6t
Xbit_r36_c19 bl_19 br_19 wl_36 vdd gnd cell_6t
Xbit_r37_c19 bl_19 br_19 wl_37 vdd gnd cell_6t
Xbit_r38_c19 bl_19 br_19 wl_38 vdd gnd cell_6t
Xbit_r39_c19 bl_19 br_19 wl_39 vdd gnd cell_6t
Xbit_r40_c19 bl_19 br_19 wl_40 vdd gnd cell_6t
Xbit_r41_c19 bl_19 br_19 wl_41 vdd gnd cell_6t
Xbit_r42_c19 bl_19 br_19 wl_42 vdd gnd cell_6t
Xbit_r43_c19 bl_19 br_19 wl_43 vdd gnd cell_6t
Xbit_r44_c19 bl_19 br_19 wl_44 vdd gnd cell_6t
Xbit_r45_c19 bl_19 br_19 wl_45 vdd gnd cell_6t
Xbit_r46_c19 bl_19 br_19 wl_46 vdd gnd cell_6t
Xbit_r47_c19 bl_19 br_19 wl_47 vdd gnd cell_6t
Xbit_r48_c19 bl_19 br_19 wl_48 vdd gnd cell_6t
Xbit_r49_c19 bl_19 br_19 wl_49 vdd gnd cell_6t
Xbit_r50_c19 bl_19 br_19 wl_50 vdd gnd cell_6t
Xbit_r51_c19 bl_19 br_19 wl_51 vdd gnd cell_6t
Xbit_r52_c19 bl_19 br_19 wl_52 vdd gnd cell_6t
Xbit_r53_c19 bl_19 br_19 wl_53 vdd gnd cell_6t
Xbit_r54_c19 bl_19 br_19 wl_54 vdd gnd cell_6t
Xbit_r55_c19 bl_19 br_19 wl_55 vdd gnd cell_6t
Xbit_r56_c19 bl_19 br_19 wl_56 vdd gnd cell_6t
Xbit_r57_c19 bl_19 br_19 wl_57 vdd gnd cell_6t
Xbit_r58_c19 bl_19 br_19 wl_58 vdd gnd cell_6t
Xbit_r59_c19 bl_19 br_19 wl_59 vdd gnd cell_6t
Xbit_r60_c19 bl_19 br_19 wl_60 vdd gnd cell_6t
Xbit_r61_c19 bl_19 br_19 wl_61 vdd gnd cell_6t
Xbit_r62_c19 bl_19 br_19 wl_62 vdd gnd cell_6t
Xbit_r63_c19 bl_19 br_19 wl_63 vdd gnd cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd cell_6t
Xbit_r1_c20 bl_20 br_20 wl_1 vdd gnd cell_6t
Xbit_r2_c20 bl_20 br_20 wl_2 vdd gnd cell_6t
Xbit_r3_c20 bl_20 br_20 wl_3 vdd gnd cell_6t
Xbit_r4_c20 bl_20 br_20 wl_4 vdd gnd cell_6t
Xbit_r5_c20 bl_20 br_20 wl_5 vdd gnd cell_6t
Xbit_r6_c20 bl_20 br_20 wl_6 vdd gnd cell_6t
Xbit_r7_c20 bl_20 br_20 wl_7 vdd gnd cell_6t
Xbit_r8_c20 bl_20 br_20 wl_8 vdd gnd cell_6t
Xbit_r9_c20 bl_20 br_20 wl_9 vdd gnd cell_6t
Xbit_r10_c20 bl_20 br_20 wl_10 vdd gnd cell_6t
Xbit_r11_c20 bl_20 br_20 wl_11 vdd gnd cell_6t
Xbit_r12_c20 bl_20 br_20 wl_12 vdd gnd cell_6t
Xbit_r13_c20 bl_20 br_20 wl_13 vdd gnd cell_6t
Xbit_r14_c20 bl_20 br_20 wl_14 vdd gnd cell_6t
Xbit_r15_c20 bl_20 br_20 wl_15 vdd gnd cell_6t
Xbit_r16_c20 bl_20 br_20 wl_16 vdd gnd cell_6t
Xbit_r17_c20 bl_20 br_20 wl_17 vdd gnd cell_6t
Xbit_r18_c20 bl_20 br_20 wl_18 vdd gnd cell_6t
Xbit_r19_c20 bl_20 br_20 wl_19 vdd gnd cell_6t
Xbit_r20_c20 bl_20 br_20 wl_20 vdd gnd cell_6t
Xbit_r21_c20 bl_20 br_20 wl_21 vdd gnd cell_6t
Xbit_r22_c20 bl_20 br_20 wl_22 vdd gnd cell_6t
Xbit_r23_c20 bl_20 br_20 wl_23 vdd gnd cell_6t
Xbit_r24_c20 bl_20 br_20 wl_24 vdd gnd cell_6t
Xbit_r25_c20 bl_20 br_20 wl_25 vdd gnd cell_6t
Xbit_r26_c20 bl_20 br_20 wl_26 vdd gnd cell_6t
Xbit_r27_c20 bl_20 br_20 wl_27 vdd gnd cell_6t
Xbit_r28_c20 bl_20 br_20 wl_28 vdd gnd cell_6t
Xbit_r29_c20 bl_20 br_20 wl_29 vdd gnd cell_6t
Xbit_r30_c20 bl_20 br_20 wl_30 vdd gnd cell_6t
Xbit_r31_c20 bl_20 br_20 wl_31 vdd gnd cell_6t
Xbit_r32_c20 bl_20 br_20 wl_32 vdd gnd cell_6t
Xbit_r33_c20 bl_20 br_20 wl_33 vdd gnd cell_6t
Xbit_r34_c20 bl_20 br_20 wl_34 vdd gnd cell_6t
Xbit_r35_c20 bl_20 br_20 wl_35 vdd gnd cell_6t
Xbit_r36_c20 bl_20 br_20 wl_36 vdd gnd cell_6t
Xbit_r37_c20 bl_20 br_20 wl_37 vdd gnd cell_6t
Xbit_r38_c20 bl_20 br_20 wl_38 vdd gnd cell_6t
Xbit_r39_c20 bl_20 br_20 wl_39 vdd gnd cell_6t
Xbit_r40_c20 bl_20 br_20 wl_40 vdd gnd cell_6t
Xbit_r41_c20 bl_20 br_20 wl_41 vdd gnd cell_6t
Xbit_r42_c20 bl_20 br_20 wl_42 vdd gnd cell_6t
Xbit_r43_c20 bl_20 br_20 wl_43 vdd gnd cell_6t
Xbit_r44_c20 bl_20 br_20 wl_44 vdd gnd cell_6t
Xbit_r45_c20 bl_20 br_20 wl_45 vdd gnd cell_6t
Xbit_r46_c20 bl_20 br_20 wl_46 vdd gnd cell_6t
Xbit_r47_c20 bl_20 br_20 wl_47 vdd gnd cell_6t
Xbit_r48_c20 bl_20 br_20 wl_48 vdd gnd cell_6t
Xbit_r49_c20 bl_20 br_20 wl_49 vdd gnd cell_6t
Xbit_r50_c20 bl_20 br_20 wl_50 vdd gnd cell_6t
Xbit_r51_c20 bl_20 br_20 wl_51 vdd gnd cell_6t
Xbit_r52_c20 bl_20 br_20 wl_52 vdd gnd cell_6t
Xbit_r53_c20 bl_20 br_20 wl_53 vdd gnd cell_6t
Xbit_r54_c20 bl_20 br_20 wl_54 vdd gnd cell_6t
Xbit_r55_c20 bl_20 br_20 wl_55 vdd gnd cell_6t
Xbit_r56_c20 bl_20 br_20 wl_56 vdd gnd cell_6t
Xbit_r57_c20 bl_20 br_20 wl_57 vdd gnd cell_6t
Xbit_r58_c20 bl_20 br_20 wl_58 vdd gnd cell_6t
Xbit_r59_c20 bl_20 br_20 wl_59 vdd gnd cell_6t
Xbit_r60_c20 bl_20 br_20 wl_60 vdd gnd cell_6t
Xbit_r61_c20 bl_20 br_20 wl_61 vdd gnd cell_6t
Xbit_r62_c20 bl_20 br_20 wl_62 vdd gnd cell_6t
Xbit_r63_c20 bl_20 br_20 wl_63 vdd gnd cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd cell_6t
Xbit_r1_c21 bl_21 br_21 wl_1 vdd gnd cell_6t
Xbit_r2_c21 bl_21 br_21 wl_2 vdd gnd cell_6t
Xbit_r3_c21 bl_21 br_21 wl_3 vdd gnd cell_6t
Xbit_r4_c21 bl_21 br_21 wl_4 vdd gnd cell_6t
Xbit_r5_c21 bl_21 br_21 wl_5 vdd gnd cell_6t
Xbit_r6_c21 bl_21 br_21 wl_6 vdd gnd cell_6t
Xbit_r7_c21 bl_21 br_21 wl_7 vdd gnd cell_6t
Xbit_r8_c21 bl_21 br_21 wl_8 vdd gnd cell_6t
Xbit_r9_c21 bl_21 br_21 wl_9 vdd gnd cell_6t
Xbit_r10_c21 bl_21 br_21 wl_10 vdd gnd cell_6t
Xbit_r11_c21 bl_21 br_21 wl_11 vdd gnd cell_6t
Xbit_r12_c21 bl_21 br_21 wl_12 vdd gnd cell_6t
Xbit_r13_c21 bl_21 br_21 wl_13 vdd gnd cell_6t
Xbit_r14_c21 bl_21 br_21 wl_14 vdd gnd cell_6t
Xbit_r15_c21 bl_21 br_21 wl_15 vdd gnd cell_6t
Xbit_r16_c21 bl_21 br_21 wl_16 vdd gnd cell_6t
Xbit_r17_c21 bl_21 br_21 wl_17 vdd gnd cell_6t
Xbit_r18_c21 bl_21 br_21 wl_18 vdd gnd cell_6t
Xbit_r19_c21 bl_21 br_21 wl_19 vdd gnd cell_6t
Xbit_r20_c21 bl_21 br_21 wl_20 vdd gnd cell_6t
Xbit_r21_c21 bl_21 br_21 wl_21 vdd gnd cell_6t
Xbit_r22_c21 bl_21 br_21 wl_22 vdd gnd cell_6t
Xbit_r23_c21 bl_21 br_21 wl_23 vdd gnd cell_6t
Xbit_r24_c21 bl_21 br_21 wl_24 vdd gnd cell_6t
Xbit_r25_c21 bl_21 br_21 wl_25 vdd gnd cell_6t
Xbit_r26_c21 bl_21 br_21 wl_26 vdd gnd cell_6t
Xbit_r27_c21 bl_21 br_21 wl_27 vdd gnd cell_6t
Xbit_r28_c21 bl_21 br_21 wl_28 vdd gnd cell_6t
Xbit_r29_c21 bl_21 br_21 wl_29 vdd gnd cell_6t
Xbit_r30_c21 bl_21 br_21 wl_30 vdd gnd cell_6t
Xbit_r31_c21 bl_21 br_21 wl_31 vdd gnd cell_6t
Xbit_r32_c21 bl_21 br_21 wl_32 vdd gnd cell_6t
Xbit_r33_c21 bl_21 br_21 wl_33 vdd gnd cell_6t
Xbit_r34_c21 bl_21 br_21 wl_34 vdd gnd cell_6t
Xbit_r35_c21 bl_21 br_21 wl_35 vdd gnd cell_6t
Xbit_r36_c21 bl_21 br_21 wl_36 vdd gnd cell_6t
Xbit_r37_c21 bl_21 br_21 wl_37 vdd gnd cell_6t
Xbit_r38_c21 bl_21 br_21 wl_38 vdd gnd cell_6t
Xbit_r39_c21 bl_21 br_21 wl_39 vdd gnd cell_6t
Xbit_r40_c21 bl_21 br_21 wl_40 vdd gnd cell_6t
Xbit_r41_c21 bl_21 br_21 wl_41 vdd gnd cell_6t
Xbit_r42_c21 bl_21 br_21 wl_42 vdd gnd cell_6t
Xbit_r43_c21 bl_21 br_21 wl_43 vdd gnd cell_6t
Xbit_r44_c21 bl_21 br_21 wl_44 vdd gnd cell_6t
Xbit_r45_c21 bl_21 br_21 wl_45 vdd gnd cell_6t
Xbit_r46_c21 bl_21 br_21 wl_46 vdd gnd cell_6t
Xbit_r47_c21 bl_21 br_21 wl_47 vdd gnd cell_6t
Xbit_r48_c21 bl_21 br_21 wl_48 vdd gnd cell_6t
Xbit_r49_c21 bl_21 br_21 wl_49 vdd gnd cell_6t
Xbit_r50_c21 bl_21 br_21 wl_50 vdd gnd cell_6t
Xbit_r51_c21 bl_21 br_21 wl_51 vdd gnd cell_6t
Xbit_r52_c21 bl_21 br_21 wl_52 vdd gnd cell_6t
Xbit_r53_c21 bl_21 br_21 wl_53 vdd gnd cell_6t
Xbit_r54_c21 bl_21 br_21 wl_54 vdd gnd cell_6t
Xbit_r55_c21 bl_21 br_21 wl_55 vdd gnd cell_6t
Xbit_r56_c21 bl_21 br_21 wl_56 vdd gnd cell_6t
Xbit_r57_c21 bl_21 br_21 wl_57 vdd gnd cell_6t
Xbit_r58_c21 bl_21 br_21 wl_58 vdd gnd cell_6t
Xbit_r59_c21 bl_21 br_21 wl_59 vdd gnd cell_6t
Xbit_r60_c21 bl_21 br_21 wl_60 vdd gnd cell_6t
Xbit_r61_c21 bl_21 br_21 wl_61 vdd gnd cell_6t
Xbit_r62_c21 bl_21 br_21 wl_62 vdd gnd cell_6t
Xbit_r63_c21 bl_21 br_21 wl_63 vdd gnd cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd cell_6t
Xbit_r1_c22 bl_22 br_22 wl_1 vdd gnd cell_6t
Xbit_r2_c22 bl_22 br_22 wl_2 vdd gnd cell_6t
Xbit_r3_c22 bl_22 br_22 wl_3 vdd gnd cell_6t
Xbit_r4_c22 bl_22 br_22 wl_4 vdd gnd cell_6t
Xbit_r5_c22 bl_22 br_22 wl_5 vdd gnd cell_6t
Xbit_r6_c22 bl_22 br_22 wl_6 vdd gnd cell_6t
Xbit_r7_c22 bl_22 br_22 wl_7 vdd gnd cell_6t
Xbit_r8_c22 bl_22 br_22 wl_8 vdd gnd cell_6t
Xbit_r9_c22 bl_22 br_22 wl_9 vdd gnd cell_6t
Xbit_r10_c22 bl_22 br_22 wl_10 vdd gnd cell_6t
Xbit_r11_c22 bl_22 br_22 wl_11 vdd gnd cell_6t
Xbit_r12_c22 bl_22 br_22 wl_12 vdd gnd cell_6t
Xbit_r13_c22 bl_22 br_22 wl_13 vdd gnd cell_6t
Xbit_r14_c22 bl_22 br_22 wl_14 vdd gnd cell_6t
Xbit_r15_c22 bl_22 br_22 wl_15 vdd gnd cell_6t
Xbit_r16_c22 bl_22 br_22 wl_16 vdd gnd cell_6t
Xbit_r17_c22 bl_22 br_22 wl_17 vdd gnd cell_6t
Xbit_r18_c22 bl_22 br_22 wl_18 vdd gnd cell_6t
Xbit_r19_c22 bl_22 br_22 wl_19 vdd gnd cell_6t
Xbit_r20_c22 bl_22 br_22 wl_20 vdd gnd cell_6t
Xbit_r21_c22 bl_22 br_22 wl_21 vdd gnd cell_6t
Xbit_r22_c22 bl_22 br_22 wl_22 vdd gnd cell_6t
Xbit_r23_c22 bl_22 br_22 wl_23 vdd gnd cell_6t
Xbit_r24_c22 bl_22 br_22 wl_24 vdd gnd cell_6t
Xbit_r25_c22 bl_22 br_22 wl_25 vdd gnd cell_6t
Xbit_r26_c22 bl_22 br_22 wl_26 vdd gnd cell_6t
Xbit_r27_c22 bl_22 br_22 wl_27 vdd gnd cell_6t
Xbit_r28_c22 bl_22 br_22 wl_28 vdd gnd cell_6t
Xbit_r29_c22 bl_22 br_22 wl_29 vdd gnd cell_6t
Xbit_r30_c22 bl_22 br_22 wl_30 vdd gnd cell_6t
Xbit_r31_c22 bl_22 br_22 wl_31 vdd gnd cell_6t
Xbit_r32_c22 bl_22 br_22 wl_32 vdd gnd cell_6t
Xbit_r33_c22 bl_22 br_22 wl_33 vdd gnd cell_6t
Xbit_r34_c22 bl_22 br_22 wl_34 vdd gnd cell_6t
Xbit_r35_c22 bl_22 br_22 wl_35 vdd gnd cell_6t
Xbit_r36_c22 bl_22 br_22 wl_36 vdd gnd cell_6t
Xbit_r37_c22 bl_22 br_22 wl_37 vdd gnd cell_6t
Xbit_r38_c22 bl_22 br_22 wl_38 vdd gnd cell_6t
Xbit_r39_c22 bl_22 br_22 wl_39 vdd gnd cell_6t
Xbit_r40_c22 bl_22 br_22 wl_40 vdd gnd cell_6t
Xbit_r41_c22 bl_22 br_22 wl_41 vdd gnd cell_6t
Xbit_r42_c22 bl_22 br_22 wl_42 vdd gnd cell_6t
Xbit_r43_c22 bl_22 br_22 wl_43 vdd gnd cell_6t
Xbit_r44_c22 bl_22 br_22 wl_44 vdd gnd cell_6t
Xbit_r45_c22 bl_22 br_22 wl_45 vdd gnd cell_6t
Xbit_r46_c22 bl_22 br_22 wl_46 vdd gnd cell_6t
Xbit_r47_c22 bl_22 br_22 wl_47 vdd gnd cell_6t
Xbit_r48_c22 bl_22 br_22 wl_48 vdd gnd cell_6t
Xbit_r49_c22 bl_22 br_22 wl_49 vdd gnd cell_6t
Xbit_r50_c22 bl_22 br_22 wl_50 vdd gnd cell_6t
Xbit_r51_c22 bl_22 br_22 wl_51 vdd gnd cell_6t
Xbit_r52_c22 bl_22 br_22 wl_52 vdd gnd cell_6t
Xbit_r53_c22 bl_22 br_22 wl_53 vdd gnd cell_6t
Xbit_r54_c22 bl_22 br_22 wl_54 vdd gnd cell_6t
Xbit_r55_c22 bl_22 br_22 wl_55 vdd gnd cell_6t
Xbit_r56_c22 bl_22 br_22 wl_56 vdd gnd cell_6t
Xbit_r57_c22 bl_22 br_22 wl_57 vdd gnd cell_6t
Xbit_r58_c22 bl_22 br_22 wl_58 vdd gnd cell_6t
Xbit_r59_c22 bl_22 br_22 wl_59 vdd gnd cell_6t
Xbit_r60_c22 bl_22 br_22 wl_60 vdd gnd cell_6t
Xbit_r61_c22 bl_22 br_22 wl_61 vdd gnd cell_6t
Xbit_r62_c22 bl_22 br_22 wl_62 vdd gnd cell_6t
Xbit_r63_c22 bl_22 br_22 wl_63 vdd gnd cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd cell_6t
Xbit_r1_c23 bl_23 br_23 wl_1 vdd gnd cell_6t
Xbit_r2_c23 bl_23 br_23 wl_2 vdd gnd cell_6t
Xbit_r3_c23 bl_23 br_23 wl_3 vdd gnd cell_6t
Xbit_r4_c23 bl_23 br_23 wl_4 vdd gnd cell_6t
Xbit_r5_c23 bl_23 br_23 wl_5 vdd gnd cell_6t
Xbit_r6_c23 bl_23 br_23 wl_6 vdd gnd cell_6t
Xbit_r7_c23 bl_23 br_23 wl_7 vdd gnd cell_6t
Xbit_r8_c23 bl_23 br_23 wl_8 vdd gnd cell_6t
Xbit_r9_c23 bl_23 br_23 wl_9 vdd gnd cell_6t
Xbit_r10_c23 bl_23 br_23 wl_10 vdd gnd cell_6t
Xbit_r11_c23 bl_23 br_23 wl_11 vdd gnd cell_6t
Xbit_r12_c23 bl_23 br_23 wl_12 vdd gnd cell_6t
Xbit_r13_c23 bl_23 br_23 wl_13 vdd gnd cell_6t
Xbit_r14_c23 bl_23 br_23 wl_14 vdd gnd cell_6t
Xbit_r15_c23 bl_23 br_23 wl_15 vdd gnd cell_6t
Xbit_r16_c23 bl_23 br_23 wl_16 vdd gnd cell_6t
Xbit_r17_c23 bl_23 br_23 wl_17 vdd gnd cell_6t
Xbit_r18_c23 bl_23 br_23 wl_18 vdd gnd cell_6t
Xbit_r19_c23 bl_23 br_23 wl_19 vdd gnd cell_6t
Xbit_r20_c23 bl_23 br_23 wl_20 vdd gnd cell_6t
Xbit_r21_c23 bl_23 br_23 wl_21 vdd gnd cell_6t
Xbit_r22_c23 bl_23 br_23 wl_22 vdd gnd cell_6t
Xbit_r23_c23 bl_23 br_23 wl_23 vdd gnd cell_6t
Xbit_r24_c23 bl_23 br_23 wl_24 vdd gnd cell_6t
Xbit_r25_c23 bl_23 br_23 wl_25 vdd gnd cell_6t
Xbit_r26_c23 bl_23 br_23 wl_26 vdd gnd cell_6t
Xbit_r27_c23 bl_23 br_23 wl_27 vdd gnd cell_6t
Xbit_r28_c23 bl_23 br_23 wl_28 vdd gnd cell_6t
Xbit_r29_c23 bl_23 br_23 wl_29 vdd gnd cell_6t
Xbit_r30_c23 bl_23 br_23 wl_30 vdd gnd cell_6t
Xbit_r31_c23 bl_23 br_23 wl_31 vdd gnd cell_6t
Xbit_r32_c23 bl_23 br_23 wl_32 vdd gnd cell_6t
Xbit_r33_c23 bl_23 br_23 wl_33 vdd gnd cell_6t
Xbit_r34_c23 bl_23 br_23 wl_34 vdd gnd cell_6t
Xbit_r35_c23 bl_23 br_23 wl_35 vdd gnd cell_6t
Xbit_r36_c23 bl_23 br_23 wl_36 vdd gnd cell_6t
Xbit_r37_c23 bl_23 br_23 wl_37 vdd gnd cell_6t
Xbit_r38_c23 bl_23 br_23 wl_38 vdd gnd cell_6t
Xbit_r39_c23 bl_23 br_23 wl_39 vdd gnd cell_6t
Xbit_r40_c23 bl_23 br_23 wl_40 vdd gnd cell_6t
Xbit_r41_c23 bl_23 br_23 wl_41 vdd gnd cell_6t
Xbit_r42_c23 bl_23 br_23 wl_42 vdd gnd cell_6t
Xbit_r43_c23 bl_23 br_23 wl_43 vdd gnd cell_6t
Xbit_r44_c23 bl_23 br_23 wl_44 vdd gnd cell_6t
Xbit_r45_c23 bl_23 br_23 wl_45 vdd gnd cell_6t
Xbit_r46_c23 bl_23 br_23 wl_46 vdd gnd cell_6t
Xbit_r47_c23 bl_23 br_23 wl_47 vdd gnd cell_6t
Xbit_r48_c23 bl_23 br_23 wl_48 vdd gnd cell_6t
Xbit_r49_c23 bl_23 br_23 wl_49 vdd gnd cell_6t
Xbit_r50_c23 bl_23 br_23 wl_50 vdd gnd cell_6t
Xbit_r51_c23 bl_23 br_23 wl_51 vdd gnd cell_6t
Xbit_r52_c23 bl_23 br_23 wl_52 vdd gnd cell_6t
Xbit_r53_c23 bl_23 br_23 wl_53 vdd gnd cell_6t
Xbit_r54_c23 bl_23 br_23 wl_54 vdd gnd cell_6t
Xbit_r55_c23 bl_23 br_23 wl_55 vdd gnd cell_6t
Xbit_r56_c23 bl_23 br_23 wl_56 vdd gnd cell_6t
Xbit_r57_c23 bl_23 br_23 wl_57 vdd gnd cell_6t
Xbit_r58_c23 bl_23 br_23 wl_58 vdd gnd cell_6t
Xbit_r59_c23 bl_23 br_23 wl_59 vdd gnd cell_6t
Xbit_r60_c23 bl_23 br_23 wl_60 vdd gnd cell_6t
Xbit_r61_c23 bl_23 br_23 wl_61 vdd gnd cell_6t
Xbit_r62_c23 bl_23 br_23 wl_62 vdd gnd cell_6t
Xbit_r63_c23 bl_23 br_23 wl_63 vdd gnd cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd cell_6t
Xbit_r1_c24 bl_24 br_24 wl_1 vdd gnd cell_6t
Xbit_r2_c24 bl_24 br_24 wl_2 vdd gnd cell_6t
Xbit_r3_c24 bl_24 br_24 wl_3 vdd gnd cell_6t
Xbit_r4_c24 bl_24 br_24 wl_4 vdd gnd cell_6t
Xbit_r5_c24 bl_24 br_24 wl_5 vdd gnd cell_6t
Xbit_r6_c24 bl_24 br_24 wl_6 vdd gnd cell_6t
Xbit_r7_c24 bl_24 br_24 wl_7 vdd gnd cell_6t
Xbit_r8_c24 bl_24 br_24 wl_8 vdd gnd cell_6t
Xbit_r9_c24 bl_24 br_24 wl_9 vdd gnd cell_6t
Xbit_r10_c24 bl_24 br_24 wl_10 vdd gnd cell_6t
Xbit_r11_c24 bl_24 br_24 wl_11 vdd gnd cell_6t
Xbit_r12_c24 bl_24 br_24 wl_12 vdd gnd cell_6t
Xbit_r13_c24 bl_24 br_24 wl_13 vdd gnd cell_6t
Xbit_r14_c24 bl_24 br_24 wl_14 vdd gnd cell_6t
Xbit_r15_c24 bl_24 br_24 wl_15 vdd gnd cell_6t
Xbit_r16_c24 bl_24 br_24 wl_16 vdd gnd cell_6t
Xbit_r17_c24 bl_24 br_24 wl_17 vdd gnd cell_6t
Xbit_r18_c24 bl_24 br_24 wl_18 vdd gnd cell_6t
Xbit_r19_c24 bl_24 br_24 wl_19 vdd gnd cell_6t
Xbit_r20_c24 bl_24 br_24 wl_20 vdd gnd cell_6t
Xbit_r21_c24 bl_24 br_24 wl_21 vdd gnd cell_6t
Xbit_r22_c24 bl_24 br_24 wl_22 vdd gnd cell_6t
Xbit_r23_c24 bl_24 br_24 wl_23 vdd gnd cell_6t
Xbit_r24_c24 bl_24 br_24 wl_24 vdd gnd cell_6t
Xbit_r25_c24 bl_24 br_24 wl_25 vdd gnd cell_6t
Xbit_r26_c24 bl_24 br_24 wl_26 vdd gnd cell_6t
Xbit_r27_c24 bl_24 br_24 wl_27 vdd gnd cell_6t
Xbit_r28_c24 bl_24 br_24 wl_28 vdd gnd cell_6t
Xbit_r29_c24 bl_24 br_24 wl_29 vdd gnd cell_6t
Xbit_r30_c24 bl_24 br_24 wl_30 vdd gnd cell_6t
Xbit_r31_c24 bl_24 br_24 wl_31 vdd gnd cell_6t
Xbit_r32_c24 bl_24 br_24 wl_32 vdd gnd cell_6t
Xbit_r33_c24 bl_24 br_24 wl_33 vdd gnd cell_6t
Xbit_r34_c24 bl_24 br_24 wl_34 vdd gnd cell_6t
Xbit_r35_c24 bl_24 br_24 wl_35 vdd gnd cell_6t
Xbit_r36_c24 bl_24 br_24 wl_36 vdd gnd cell_6t
Xbit_r37_c24 bl_24 br_24 wl_37 vdd gnd cell_6t
Xbit_r38_c24 bl_24 br_24 wl_38 vdd gnd cell_6t
Xbit_r39_c24 bl_24 br_24 wl_39 vdd gnd cell_6t
Xbit_r40_c24 bl_24 br_24 wl_40 vdd gnd cell_6t
Xbit_r41_c24 bl_24 br_24 wl_41 vdd gnd cell_6t
Xbit_r42_c24 bl_24 br_24 wl_42 vdd gnd cell_6t
Xbit_r43_c24 bl_24 br_24 wl_43 vdd gnd cell_6t
Xbit_r44_c24 bl_24 br_24 wl_44 vdd gnd cell_6t
Xbit_r45_c24 bl_24 br_24 wl_45 vdd gnd cell_6t
Xbit_r46_c24 bl_24 br_24 wl_46 vdd gnd cell_6t
Xbit_r47_c24 bl_24 br_24 wl_47 vdd gnd cell_6t
Xbit_r48_c24 bl_24 br_24 wl_48 vdd gnd cell_6t
Xbit_r49_c24 bl_24 br_24 wl_49 vdd gnd cell_6t
Xbit_r50_c24 bl_24 br_24 wl_50 vdd gnd cell_6t
Xbit_r51_c24 bl_24 br_24 wl_51 vdd gnd cell_6t
Xbit_r52_c24 bl_24 br_24 wl_52 vdd gnd cell_6t
Xbit_r53_c24 bl_24 br_24 wl_53 vdd gnd cell_6t
Xbit_r54_c24 bl_24 br_24 wl_54 vdd gnd cell_6t
Xbit_r55_c24 bl_24 br_24 wl_55 vdd gnd cell_6t
Xbit_r56_c24 bl_24 br_24 wl_56 vdd gnd cell_6t
Xbit_r57_c24 bl_24 br_24 wl_57 vdd gnd cell_6t
Xbit_r58_c24 bl_24 br_24 wl_58 vdd gnd cell_6t
Xbit_r59_c24 bl_24 br_24 wl_59 vdd gnd cell_6t
Xbit_r60_c24 bl_24 br_24 wl_60 vdd gnd cell_6t
Xbit_r61_c24 bl_24 br_24 wl_61 vdd gnd cell_6t
Xbit_r62_c24 bl_24 br_24 wl_62 vdd gnd cell_6t
Xbit_r63_c24 bl_24 br_24 wl_63 vdd gnd cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd cell_6t
Xbit_r1_c25 bl_25 br_25 wl_1 vdd gnd cell_6t
Xbit_r2_c25 bl_25 br_25 wl_2 vdd gnd cell_6t
Xbit_r3_c25 bl_25 br_25 wl_3 vdd gnd cell_6t
Xbit_r4_c25 bl_25 br_25 wl_4 vdd gnd cell_6t
Xbit_r5_c25 bl_25 br_25 wl_5 vdd gnd cell_6t
Xbit_r6_c25 bl_25 br_25 wl_6 vdd gnd cell_6t
Xbit_r7_c25 bl_25 br_25 wl_7 vdd gnd cell_6t
Xbit_r8_c25 bl_25 br_25 wl_8 vdd gnd cell_6t
Xbit_r9_c25 bl_25 br_25 wl_9 vdd gnd cell_6t
Xbit_r10_c25 bl_25 br_25 wl_10 vdd gnd cell_6t
Xbit_r11_c25 bl_25 br_25 wl_11 vdd gnd cell_6t
Xbit_r12_c25 bl_25 br_25 wl_12 vdd gnd cell_6t
Xbit_r13_c25 bl_25 br_25 wl_13 vdd gnd cell_6t
Xbit_r14_c25 bl_25 br_25 wl_14 vdd gnd cell_6t
Xbit_r15_c25 bl_25 br_25 wl_15 vdd gnd cell_6t
Xbit_r16_c25 bl_25 br_25 wl_16 vdd gnd cell_6t
Xbit_r17_c25 bl_25 br_25 wl_17 vdd gnd cell_6t
Xbit_r18_c25 bl_25 br_25 wl_18 vdd gnd cell_6t
Xbit_r19_c25 bl_25 br_25 wl_19 vdd gnd cell_6t
Xbit_r20_c25 bl_25 br_25 wl_20 vdd gnd cell_6t
Xbit_r21_c25 bl_25 br_25 wl_21 vdd gnd cell_6t
Xbit_r22_c25 bl_25 br_25 wl_22 vdd gnd cell_6t
Xbit_r23_c25 bl_25 br_25 wl_23 vdd gnd cell_6t
Xbit_r24_c25 bl_25 br_25 wl_24 vdd gnd cell_6t
Xbit_r25_c25 bl_25 br_25 wl_25 vdd gnd cell_6t
Xbit_r26_c25 bl_25 br_25 wl_26 vdd gnd cell_6t
Xbit_r27_c25 bl_25 br_25 wl_27 vdd gnd cell_6t
Xbit_r28_c25 bl_25 br_25 wl_28 vdd gnd cell_6t
Xbit_r29_c25 bl_25 br_25 wl_29 vdd gnd cell_6t
Xbit_r30_c25 bl_25 br_25 wl_30 vdd gnd cell_6t
Xbit_r31_c25 bl_25 br_25 wl_31 vdd gnd cell_6t
Xbit_r32_c25 bl_25 br_25 wl_32 vdd gnd cell_6t
Xbit_r33_c25 bl_25 br_25 wl_33 vdd gnd cell_6t
Xbit_r34_c25 bl_25 br_25 wl_34 vdd gnd cell_6t
Xbit_r35_c25 bl_25 br_25 wl_35 vdd gnd cell_6t
Xbit_r36_c25 bl_25 br_25 wl_36 vdd gnd cell_6t
Xbit_r37_c25 bl_25 br_25 wl_37 vdd gnd cell_6t
Xbit_r38_c25 bl_25 br_25 wl_38 vdd gnd cell_6t
Xbit_r39_c25 bl_25 br_25 wl_39 vdd gnd cell_6t
Xbit_r40_c25 bl_25 br_25 wl_40 vdd gnd cell_6t
Xbit_r41_c25 bl_25 br_25 wl_41 vdd gnd cell_6t
Xbit_r42_c25 bl_25 br_25 wl_42 vdd gnd cell_6t
Xbit_r43_c25 bl_25 br_25 wl_43 vdd gnd cell_6t
Xbit_r44_c25 bl_25 br_25 wl_44 vdd gnd cell_6t
Xbit_r45_c25 bl_25 br_25 wl_45 vdd gnd cell_6t
Xbit_r46_c25 bl_25 br_25 wl_46 vdd gnd cell_6t
Xbit_r47_c25 bl_25 br_25 wl_47 vdd gnd cell_6t
Xbit_r48_c25 bl_25 br_25 wl_48 vdd gnd cell_6t
Xbit_r49_c25 bl_25 br_25 wl_49 vdd gnd cell_6t
Xbit_r50_c25 bl_25 br_25 wl_50 vdd gnd cell_6t
Xbit_r51_c25 bl_25 br_25 wl_51 vdd gnd cell_6t
Xbit_r52_c25 bl_25 br_25 wl_52 vdd gnd cell_6t
Xbit_r53_c25 bl_25 br_25 wl_53 vdd gnd cell_6t
Xbit_r54_c25 bl_25 br_25 wl_54 vdd gnd cell_6t
Xbit_r55_c25 bl_25 br_25 wl_55 vdd gnd cell_6t
Xbit_r56_c25 bl_25 br_25 wl_56 vdd gnd cell_6t
Xbit_r57_c25 bl_25 br_25 wl_57 vdd gnd cell_6t
Xbit_r58_c25 bl_25 br_25 wl_58 vdd gnd cell_6t
Xbit_r59_c25 bl_25 br_25 wl_59 vdd gnd cell_6t
Xbit_r60_c25 bl_25 br_25 wl_60 vdd gnd cell_6t
Xbit_r61_c25 bl_25 br_25 wl_61 vdd gnd cell_6t
Xbit_r62_c25 bl_25 br_25 wl_62 vdd gnd cell_6t
Xbit_r63_c25 bl_25 br_25 wl_63 vdd gnd cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd cell_6t
Xbit_r1_c26 bl_26 br_26 wl_1 vdd gnd cell_6t
Xbit_r2_c26 bl_26 br_26 wl_2 vdd gnd cell_6t
Xbit_r3_c26 bl_26 br_26 wl_3 vdd gnd cell_6t
Xbit_r4_c26 bl_26 br_26 wl_4 vdd gnd cell_6t
Xbit_r5_c26 bl_26 br_26 wl_5 vdd gnd cell_6t
Xbit_r6_c26 bl_26 br_26 wl_6 vdd gnd cell_6t
Xbit_r7_c26 bl_26 br_26 wl_7 vdd gnd cell_6t
Xbit_r8_c26 bl_26 br_26 wl_8 vdd gnd cell_6t
Xbit_r9_c26 bl_26 br_26 wl_9 vdd gnd cell_6t
Xbit_r10_c26 bl_26 br_26 wl_10 vdd gnd cell_6t
Xbit_r11_c26 bl_26 br_26 wl_11 vdd gnd cell_6t
Xbit_r12_c26 bl_26 br_26 wl_12 vdd gnd cell_6t
Xbit_r13_c26 bl_26 br_26 wl_13 vdd gnd cell_6t
Xbit_r14_c26 bl_26 br_26 wl_14 vdd gnd cell_6t
Xbit_r15_c26 bl_26 br_26 wl_15 vdd gnd cell_6t
Xbit_r16_c26 bl_26 br_26 wl_16 vdd gnd cell_6t
Xbit_r17_c26 bl_26 br_26 wl_17 vdd gnd cell_6t
Xbit_r18_c26 bl_26 br_26 wl_18 vdd gnd cell_6t
Xbit_r19_c26 bl_26 br_26 wl_19 vdd gnd cell_6t
Xbit_r20_c26 bl_26 br_26 wl_20 vdd gnd cell_6t
Xbit_r21_c26 bl_26 br_26 wl_21 vdd gnd cell_6t
Xbit_r22_c26 bl_26 br_26 wl_22 vdd gnd cell_6t
Xbit_r23_c26 bl_26 br_26 wl_23 vdd gnd cell_6t
Xbit_r24_c26 bl_26 br_26 wl_24 vdd gnd cell_6t
Xbit_r25_c26 bl_26 br_26 wl_25 vdd gnd cell_6t
Xbit_r26_c26 bl_26 br_26 wl_26 vdd gnd cell_6t
Xbit_r27_c26 bl_26 br_26 wl_27 vdd gnd cell_6t
Xbit_r28_c26 bl_26 br_26 wl_28 vdd gnd cell_6t
Xbit_r29_c26 bl_26 br_26 wl_29 vdd gnd cell_6t
Xbit_r30_c26 bl_26 br_26 wl_30 vdd gnd cell_6t
Xbit_r31_c26 bl_26 br_26 wl_31 vdd gnd cell_6t
Xbit_r32_c26 bl_26 br_26 wl_32 vdd gnd cell_6t
Xbit_r33_c26 bl_26 br_26 wl_33 vdd gnd cell_6t
Xbit_r34_c26 bl_26 br_26 wl_34 vdd gnd cell_6t
Xbit_r35_c26 bl_26 br_26 wl_35 vdd gnd cell_6t
Xbit_r36_c26 bl_26 br_26 wl_36 vdd gnd cell_6t
Xbit_r37_c26 bl_26 br_26 wl_37 vdd gnd cell_6t
Xbit_r38_c26 bl_26 br_26 wl_38 vdd gnd cell_6t
Xbit_r39_c26 bl_26 br_26 wl_39 vdd gnd cell_6t
Xbit_r40_c26 bl_26 br_26 wl_40 vdd gnd cell_6t
Xbit_r41_c26 bl_26 br_26 wl_41 vdd gnd cell_6t
Xbit_r42_c26 bl_26 br_26 wl_42 vdd gnd cell_6t
Xbit_r43_c26 bl_26 br_26 wl_43 vdd gnd cell_6t
Xbit_r44_c26 bl_26 br_26 wl_44 vdd gnd cell_6t
Xbit_r45_c26 bl_26 br_26 wl_45 vdd gnd cell_6t
Xbit_r46_c26 bl_26 br_26 wl_46 vdd gnd cell_6t
Xbit_r47_c26 bl_26 br_26 wl_47 vdd gnd cell_6t
Xbit_r48_c26 bl_26 br_26 wl_48 vdd gnd cell_6t
Xbit_r49_c26 bl_26 br_26 wl_49 vdd gnd cell_6t
Xbit_r50_c26 bl_26 br_26 wl_50 vdd gnd cell_6t
Xbit_r51_c26 bl_26 br_26 wl_51 vdd gnd cell_6t
Xbit_r52_c26 bl_26 br_26 wl_52 vdd gnd cell_6t
Xbit_r53_c26 bl_26 br_26 wl_53 vdd gnd cell_6t
Xbit_r54_c26 bl_26 br_26 wl_54 vdd gnd cell_6t
Xbit_r55_c26 bl_26 br_26 wl_55 vdd gnd cell_6t
Xbit_r56_c26 bl_26 br_26 wl_56 vdd gnd cell_6t
Xbit_r57_c26 bl_26 br_26 wl_57 vdd gnd cell_6t
Xbit_r58_c26 bl_26 br_26 wl_58 vdd gnd cell_6t
Xbit_r59_c26 bl_26 br_26 wl_59 vdd gnd cell_6t
Xbit_r60_c26 bl_26 br_26 wl_60 vdd gnd cell_6t
Xbit_r61_c26 bl_26 br_26 wl_61 vdd gnd cell_6t
Xbit_r62_c26 bl_26 br_26 wl_62 vdd gnd cell_6t
Xbit_r63_c26 bl_26 br_26 wl_63 vdd gnd cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd cell_6t
Xbit_r1_c27 bl_27 br_27 wl_1 vdd gnd cell_6t
Xbit_r2_c27 bl_27 br_27 wl_2 vdd gnd cell_6t
Xbit_r3_c27 bl_27 br_27 wl_3 vdd gnd cell_6t
Xbit_r4_c27 bl_27 br_27 wl_4 vdd gnd cell_6t
Xbit_r5_c27 bl_27 br_27 wl_5 vdd gnd cell_6t
Xbit_r6_c27 bl_27 br_27 wl_6 vdd gnd cell_6t
Xbit_r7_c27 bl_27 br_27 wl_7 vdd gnd cell_6t
Xbit_r8_c27 bl_27 br_27 wl_8 vdd gnd cell_6t
Xbit_r9_c27 bl_27 br_27 wl_9 vdd gnd cell_6t
Xbit_r10_c27 bl_27 br_27 wl_10 vdd gnd cell_6t
Xbit_r11_c27 bl_27 br_27 wl_11 vdd gnd cell_6t
Xbit_r12_c27 bl_27 br_27 wl_12 vdd gnd cell_6t
Xbit_r13_c27 bl_27 br_27 wl_13 vdd gnd cell_6t
Xbit_r14_c27 bl_27 br_27 wl_14 vdd gnd cell_6t
Xbit_r15_c27 bl_27 br_27 wl_15 vdd gnd cell_6t
Xbit_r16_c27 bl_27 br_27 wl_16 vdd gnd cell_6t
Xbit_r17_c27 bl_27 br_27 wl_17 vdd gnd cell_6t
Xbit_r18_c27 bl_27 br_27 wl_18 vdd gnd cell_6t
Xbit_r19_c27 bl_27 br_27 wl_19 vdd gnd cell_6t
Xbit_r20_c27 bl_27 br_27 wl_20 vdd gnd cell_6t
Xbit_r21_c27 bl_27 br_27 wl_21 vdd gnd cell_6t
Xbit_r22_c27 bl_27 br_27 wl_22 vdd gnd cell_6t
Xbit_r23_c27 bl_27 br_27 wl_23 vdd gnd cell_6t
Xbit_r24_c27 bl_27 br_27 wl_24 vdd gnd cell_6t
Xbit_r25_c27 bl_27 br_27 wl_25 vdd gnd cell_6t
Xbit_r26_c27 bl_27 br_27 wl_26 vdd gnd cell_6t
Xbit_r27_c27 bl_27 br_27 wl_27 vdd gnd cell_6t
Xbit_r28_c27 bl_27 br_27 wl_28 vdd gnd cell_6t
Xbit_r29_c27 bl_27 br_27 wl_29 vdd gnd cell_6t
Xbit_r30_c27 bl_27 br_27 wl_30 vdd gnd cell_6t
Xbit_r31_c27 bl_27 br_27 wl_31 vdd gnd cell_6t
Xbit_r32_c27 bl_27 br_27 wl_32 vdd gnd cell_6t
Xbit_r33_c27 bl_27 br_27 wl_33 vdd gnd cell_6t
Xbit_r34_c27 bl_27 br_27 wl_34 vdd gnd cell_6t
Xbit_r35_c27 bl_27 br_27 wl_35 vdd gnd cell_6t
Xbit_r36_c27 bl_27 br_27 wl_36 vdd gnd cell_6t
Xbit_r37_c27 bl_27 br_27 wl_37 vdd gnd cell_6t
Xbit_r38_c27 bl_27 br_27 wl_38 vdd gnd cell_6t
Xbit_r39_c27 bl_27 br_27 wl_39 vdd gnd cell_6t
Xbit_r40_c27 bl_27 br_27 wl_40 vdd gnd cell_6t
Xbit_r41_c27 bl_27 br_27 wl_41 vdd gnd cell_6t
Xbit_r42_c27 bl_27 br_27 wl_42 vdd gnd cell_6t
Xbit_r43_c27 bl_27 br_27 wl_43 vdd gnd cell_6t
Xbit_r44_c27 bl_27 br_27 wl_44 vdd gnd cell_6t
Xbit_r45_c27 bl_27 br_27 wl_45 vdd gnd cell_6t
Xbit_r46_c27 bl_27 br_27 wl_46 vdd gnd cell_6t
Xbit_r47_c27 bl_27 br_27 wl_47 vdd gnd cell_6t
Xbit_r48_c27 bl_27 br_27 wl_48 vdd gnd cell_6t
Xbit_r49_c27 bl_27 br_27 wl_49 vdd gnd cell_6t
Xbit_r50_c27 bl_27 br_27 wl_50 vdd gnd cell_6t
Xbit_r51_c27 bl_27 br_27 wl_51 vdd gnd cell_6t
Xbit_r52_c27 bl_27 br_27 wl_52 vdd gnd cell_6t
Xbit_r53_c27 bl_27 br_27 wl_53 vdd gnd cell_6t
Xbit_r54_c27 bl_27 br_27 wl_54 vdd gnd cell_6t
Xbit_r55_c27 bl_27 br_27 wl_55 vdd gnd cell_6t
Xbit_r56_c27 bl_27 br_27 wl_56 vdd gnd cell_6t
Xbit_r57_c27 bl_27 br_27 wl_57 vdd gnd cell_6t
Xbit_r58_c27 bl_27 br_27 wl_58 vdd gnd cell_6t
Xbit_r59_c27 bl_27 br_27 wl_59 vdd gnd cell_6t
Xbit_r60_c27 bl_27 br_27 wl_60 vdd gnd cell_6t
Xbit_r61_c27 bl_27 br_27 wl_61 vdd gnd cell_6t
Xbit_r62_c27 bl_27 br_27 wl_62 vdd gnd cell_6t
Xbit_r63_c27 bl_27 br_27 wl_63 vdd gnd cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd cell_6t
Xbit_r1_c28 bl_28 br_28 wl_1 vdd gnd cell_6t
Xbit_r2_c28 bl_28 br_28 wl_2 vdd gnd cell_6t
Xbit_r3_c28 bl_28 br_28 wl_3 vdd gnd cell_6t
Xbit_r4_c28 bl_28 br_28 wl_4 vdd gnd cell_6t
Xbit_r5_c28 bl_28 br_28 wl_5 vdd gnd cell_6t
Xbit_r6_c28 bl_28 br_28 wl_6 vdd gnd cell_6t
Xbit_r7_c28 bl_28 br_28 wl_7 vdd gnd cell_6t
Xbit_r8_c28 bl_28 br_28 wl_8 vdd gnd cell_6t
Xbit_r9_c28 bl_28 br_28 wl_9 vdd gnd cell_6t
Xbit_r10_c28 bl_28 br_28 wl_10 vdd gnd cell_6t
Xbit_r11_c28 bl_28 br_28 wl_11 vdd gnd cell_6t
Xbit_r12_c28 bl_28 br_28 wl_12 vdd gnd cell_6t
Xbit_r13_c28 bl_28 br_28 wl_13 vdd gnd cell_6t
Xbit_r14_c28 bl_28 br_28 wl_14 vdd gnd cell_6t
Xbit_r15_c28 bl_28 br_28 wl_15 vdd gnd cell_6t
Xbit_r16_c28 bl_28 br_28 wl_16 vdd gnd cell_6t
Xbit_r17_c28 bl_28 br_28 wl_17 vdd gnd cell_6t
Xbit_r18_c28 bl_28 br_28 wl_18 vdd gnd cell_6t
Xbit_r19_c28 bl_28 br_28 wl_19 vdd gnd cell_6t
Xbit_r20_c28 bl_28 br_28 wl_20 vdd gnd cell_6t
Xbit_r21_c28 bl_28 br_28 wl_21 vdd gnd cell_6t
Xbit_r22_c28 bl_28 br_28 wl_22 vdd gnd cell_6t
Xbit_r23_c28 bl_28 br_28 wl_23 vdd gnd cell_6t
Xbit_r24_c28 bl_28 br_28 wl_24 vdd gnd cell_6t
Xbit_r25_c28 bl_28 br_28 wl_25 vdd gnd cell_6t
Xbit_r26_c28 bl_28 br_28 wl_26 vdd gnd cell_6t
Xbit_r27_c28 bl_28 br_28 wl_27 vdd gnd cell_6t
Xbit_r28_c28 bl_28 br_28 wl_28 vdd gnd cell_6t
Xbit_r29_c28 bl_28 br_28 wl_29 vdd gnd cell_6t
Xbit_r30_c28 bl_28 br_28 wl_30 vdd gnd cell_6t
Xbit_r31_c28 bl_28 br_28 wl_31 vdd gnd cell_6t
Xbit_r32_c28 bl_28 br_28 wl_32 vdd gnd cell_6t
Xbit_r33_c28 bl_28 br_28 wl_33 vdd gnd cell_6t
Xbit_r34_c28 bl_28 br_28 wl_34 vdd gnd cell_6t
Xbit_r35_c28 bl_28 br_28 wl_35 vdd gnd cell_6t
Xbit_r36_c28 bl_28 br_28 wl_36 vdd gnd cell_6t
Xbit_r37_c28 bl_28 br_28 wl_37 vdd gnd cell_6t
Xbit_r38_c28 bl_28 br_28 wl_38 vdd gnd cell_6t
Xbit_r39_c28 bl_28 br_28 wl_39 vdd gnd cell_6t
Xbit_r40_c28 bl_28 br_28 wl_40 vdd gnd cell_6t
Xbit_r41_c28 bl_28 br_28 wl_41 vdd gnd cell_6t
Xbit_r42_c28 bl_28 br_28 wl_42 vdd gnd cell_6t
Xbit_r43_c28 bl_28 br_28 wl_43 vdd gnd cell_6t
Xbit_r44_c28 bl_28 br_28 wl_44 vdd gnd cell_6t
Xbit_r45_c28 bl_28 br_28 wl_45 vdd gnd cell_6t
Xbit_r46_c28 bl_28 br_28 wl_46 vdd gnd cell_6t
Xbit_r47_c28 bl_28 br_28 wl_47 vdd gnd cell_6t
Xbit_r48_c28 bl_28 br_28 wl_48 vdd gnd cell_6t
Xbit_r49_c28 bl_28 br_28 wl_49 vdd gnd cell_6t
Xbit_r50_c28 bl_28 br_28 wl_50 vdd gnd cell_6t
Xbit_r51_c28 bl_28 br_28 wl_51 vdd gnd cell_6t
Xbit_r52_c28 bl_28 br_28 wl_52 vdd gnd cell_6t
Xbit_r53_c28 bl_28 br_28 wl_53 vdd gnd cell_6t
Xbit_r54_c28 bl_28 br_28 wl_54 vdd gnd cell_6t
Xbit_r55_c28 bl_28 br_28 wl_55 vdd gnd cell_6t
Xbit_r56_c28 bl_28 br_28 wl_56 vdd gnd cell_6t
Xbit_r57_c28 bl_28 br_28 wl_57 vdd gnd cell_6t
Xbit_r58_c28 bl_28 br_28 wl_58 vdd gnd cell_6t
Xbit_r59_c28 bl_28 br_28 wl_59 vdd gnd cell_6t
Xbit_r60_c28 bl_28 br_28 wl_60 vdd gnd cell_6t
Xbit_r61_c28 bl_28 br_28 wl_61 vdd gnd cell_6t
Xbit_r62_c28 bl_28 br_28 wl_62 vdd gnd cell_6t
Xbit_r63_c28 bl_28 br_28 wl_63 vdd gnd cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd cell_6t
Xbit_r1_c29 bl_29 br_29 wl_1 vdd gnd cell_6t
Xbit_r2_c29 bl_29 br_29 wl_2 vdd gnd cell_6t
Xbit_r3_c29 bl_29 br_29 wl_3 vdd gnd cell_6t
Xbit_r4_c29 bl_29 br_29 wl_4 vdd gnd cell_6t
Xbit_r5_c29 bl_29 br_29 wl_5 vdd gnd cell_6t
Xbit_r6_c29 bl_29 br_29 wl_6 vdd gnd cell_6t
Xbit_r7_c29 bl_29 br_29 wl_7 vdd gnd cell_6t
Xbit_r8_c29 bl_29 br_29 wl_8 vdd gnd cell_6t
Xbit_r9_c29 bl_29 br_29 wl_9 vdd gnd cell_6t
Xbit_r10_c29 bl_29 br_29 wl_10 vdd gnd cell_6t
Xbit_r11_c29 bl_29 br_29 wl_11 vdd gnd cell_6t
Xbit_r12_c29 bl_29 br_29 wl_12 vdd gnd cell_6t
Xbit_r13_c29 bl_29 br_29 wl_13 vdd gnd cell_6t
Xbit_r14_c29 bl_29 br_29 wl_14 vdd gnd cell_6t
Xbit_r15_c29 bl_29 br_29 wl_15 vdd gnd cell_6t
Xbit_r16_c29 bl_29 br_29 wl_16 vdd gnd cell_6t
Xbit_r17_c29 bl_29 br_29 wl_17 vdd gnd cell_6t
Xbit_r18_c29 bl_29 br_29 wl_18 vdd gnd cell_6t
Xbit_r19_c29 bl_29 br_29 wl_19 vdd gnd cell_6t
Xbit_r20_c29 bl_29 br_29 wl_20 vdd gnd cell_6t
Xbit_r21_c29 bl_29 br_29 wl_21 vdd gnd cell_6t
Xbit_r22_c29 bl_29 br_29 wl_22 vdd gnd cell_6t
Xbit_r23_c29 bl_29 br_29 wl_23 vdd gnd cell_6t
Xbit_r24_c29 bl_29 br_29 wl_24 vdd gnd cell_6t
Xbit_r25_c29 bl_29 br_29 wl_25 vdd gnd cell_6t
Xbit_r26_c29 bl_29 br_29 wl_26 vdd gnd cell_6t
Xbit_r27_c29 bl_29 br_29 wl_27 vdd gnd cell_6t
Xbit_r28_c29 bl_29 br_29 wl_28 vdd gnd cell_6t
Xbit_r29_c29 bl_29 br_29 wl_29 vdd gnd cell_6t
Xbit_r30_c29 bl_29 br_29 wl_30 vdd gnd cell_6t
Xbit_r31_c29 bl_29 br_29 wl_31 vdd gnd cell_6t
Xbit_r32_c29 bl_29 br_29 wl_32 vdd gnd cell_6t
Xbit_r33_c29 bl_29 br_29 wl_33 vdd gnd cell_6t
Xbit_r34_c29 bl_29 br_29 wl_34 vdd gnd cell_6t
Xbit_r35_c29 bl_29 br_29 wl_35 vdd gnd cell_6t
Xbit_r36_c29 bl_29 br_29 wl_36 vdd gnd cell_6t
Xbit_r37_c29 bl_29 br_29 wl_37 vdd gnd cell_6t
Xbit_r38_c29 bl_29 br_29 wl_38 vdd gnd cell_6t
Xbit_r39_c29 bl_29 br_29 wl_39 vdd gnd cell_6t
Xbit_r40_c29 bl_29 br_29 wl_40 vdd gnd cell_6t
Xbit_r41_c29 bl_29 br_29 wl_41 vdd gnd cell_6t
Xbit_r42_c29 bl_29 br_29 wl_42 vdd gnd cell_6t
Xbit_r43_c29 bl_29 br_29 wl_43 vdd gnd cell_6t
Xbit_r44_c29 bl_29 br_29 wl_44 vdd gnd cell_6t
Xbit_r45_c29 bl_29 br_29 wl_45 vdd gnd cell_6t
Xbit_r46_c29 bl_29 br_29 wl_46 vdd gnd cell_6t
Xbit_r47_c29 bl_29 br_29 wl_47 vdd gnd cell_6t
Xbit_r48_c29 bl_29 br_29 wl_48 vdd gnd cell_6t
Xbit_r49_c29 bl_29 br_29 wl_49 vdd gnd cell_6t
Xbit_r50_c29 bl_29 br_29 wl_50 vdd gnd cell_6t
Xbit_r51_c29 bl_29 br_29 wl_51 vdd gnd cell_6t
Xbit_r52_c29 bl_29 br_29 wl_52 vdd gnd cell_6t
Xbit_r53_c29 bl_29 br_29 wl_53 vdd gnd cell_6t
Xbit_r54_c29 bl_29 br_29 wl_54 vdd gnd cell_6t
Xbit_r55_c29 bl_29 br_29 wl_55 vdd gnd cell_6t
Xbit_r56_c29 bl_29 br_29 wl_56 vdd gnd cell_6t
Xbit_r57_c29 bl_29 br_29 wl_57 vdd gnd cell_6t
Xbit_r58_c29 bl_29 br_29 wl_58 vdd gnd cell_6t
Xbit_r59_c29 bl_29 br_29 wl_59 vdd gnd cell_6t
Xbit_r60_c29 bl_29 br_29 wl_60 vdd gnd cell_6t
Xbit_r61_c29 bl_29 br_29 wl_61 vdd gnd cell_6t
Xbit_r62_c29 bl_29 br_29 wl_62 vdd gnd cell_6t
Xbit_r63_c29 bl_29 br_29 wl_63 vdd gnd cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd cell_6t
Xbit_r1_c30 bl_30 br_30 wl_1 vdd gnd cell_6t
Xbit_r2_c30 bl_30 br_30 wl_2 vdd gnd cell_6t
Xbit_r3_c30 bl_30 br_30 wl_3 vdd gnd cell_6t
Xbit_r4_c30 bl_30 br_30 wl_4 vdd gnd cell_6t
Xbit_r5_c30 bl_30 br_30 wl_5 vdd gnd cell_6t
Xbit_r6_c30 bl_30 br_30 wl_6 vdd gnd cell_6t
Xbit_r7_c30 bl_30 br_30 wl_7 vdd gnd cell_6t
Xbit_r8_c30 bl_30 br_30 wl_8 vdd gnd cell_6t
Xbit_r9_c30 bl_30 br_30 wl_9 vdd gnd cell_6t
Xbit_r10_c30 bl_30 br_30 wl_10 vdd gnd cell_6t
Xbit_r11_c30 bl_30 br_30 wl_11 vdd gnd cell_6t
Xbit_r12_c30 bl_30 br_30 wl_12 vdd gnd cell_6t
Xbit_r13_c30 bl_30 br_30 wl_13 vdd gnd cell_6t
Xbit_r14_c30 bl_30 br_30 wl_14 vdd gnd cell_6t
Xbit_r15_c30 bl_30 br_30 wl_15 vdd gnd cell_6t
Xbit_r16_c30 bl_30 br_30 wl_16 vdd gnd cell_6t
Xbit_r17_c30 bl_30 br_30 wl_17 vdd gnd cell_6t
Xbit_r18_c30 bl_30 br_30 wl_18 vdd gnd cell_6t
Xbit_r19_c30 bl_30 br_30 wl_19 vdd gnd cell_6t
Xbit_r20_c30 bl_30 br_30 wl_20 vdd gnd cell_6t
Xbit_r21_c30 bl_30 br_30 wl_21 vdd gnd cell_6t
Xbit_r22_c30 bl_30 br_30 wl_22 vdd gnd cell_6t
Xbit_r23_c30 bl_30 br_30 wl_23 vdd gnd cell_6t
Xbit_r24_c30 bl_30 br_30 wl_24 vdd gnd cell_6t
Xbit_r25_c30 bl_30 br_30 wl_25 vdd gnd cell_6t
Xbit_r26_c30 bl_30 br_30 wl_26 vdd gnd cell_6t
Xbit_r27_c30 bl_30 br_30 wl_27 vdd gnd cell_6t
Xbit_r28_c30 bl_30 br_30 wl_28 vdd gnd cell_6t
Xbit_r29_c30 bl_30 br_30 wl_29 vdd gnd cell_6t
Xbit_r30_c30 bl_30 br_30 wl_30 vdd gnd cell_6t
Xbit_r31_c30 bl_30 br_30 wl_31 vdd gnd cell_6t
Xbit_r32_c30 bl_30 br_30 wl_32 vdd gnd cell_6t
Xbit_r33_c30 bl_30 br_30 wl_33 vdd gnd cell_6t
Xbit_r34_c30 bl_30 br_30 wl_34 vdd gnd cell_6t
Xbit_r35_c30 bl_30 br_30 wl_35 vdd gnd cell_6t
Xbit_r36_c30 bl_30 br_30 wl_36 vdd gnd cell_6t
Xbit_r37_c30 bl_30 br_30 wl_37 vdd gnd cell_6t
Xbit_r38_c30 bl_30 br_30 wl_38 vdd gnd cell_6t
Xbit_r39_c30 bl_30 br_30 wl_39 vdd gnd cell_6t
Xbit_r40_c30 bl_30 br_30 wl_40 vdd gnd cell_6t
Xbit_r41_c30 bl_30 br_30 wl_41 vdd gnd cell_6t
Xbit_r42_c30 bl_30 br_30 wl_42 vdd gnd cell_6t
Xbit_r43_c30 bl_30 br_30 wl_43 vdd gnd cell_6t
Xbit_r44_c30 bl_30 br_30 wl_44 vdd gnd cell_6t
Xbit_r45_c30 bl_30 br_30 wl_45 vdd gnd cell_6t
Xbit_r46_c30 bl_30 br_30 wl_46 vdd gnd cell_6t
Xbit_r47_c30 bl_30 br_30 wl_47 vdd gnd cell_6t
Xbit_r48_c30 bl_30 br_30 wl_48 vdd gnd cell_6t
Xbit_r49_c30 bl_30 br_30 wl_49 vdd gnd cell_6t
Xbit_r50_c30 bl_30 br_30 wl_50 vdd gnd cell_6t
Xbit_r51_c30 bl_30 br_30 wl_51 vdd gnd cell_6t
Xbit_r52_c30 bl_30 br_30 wl_52 vdd gnd cell_6t
Xbit_r53_c30 bl_30 br_30 wl_53 vdd gnd cell_6t
Xbit_r54_c30 bl_30 br_30 wl_54 vdd gnd cell_6t
Xbit_r55_c30 bl_30 br_30 wl_55 vdd gnd cell_6t
Xbit_r56_c30 bl_30 br_30 wl_56 vdd gnd cell_6t
Xbit_r57_c30 bl_30 br_30 wl_57 vdd gnd cell_6t
Xbit_r58_c30 bl_30 br_30 wl_58 vdd gnd cell_6t
Xbit_r59_c30 bl_30 br_30 wl_59 vdd gnd cell_6t
Xbit_r60_c30 bl_30 br_30 wl_60 vdd gnd cell_6t
Xbit_r61_c30 bl_30 br_30 wl_61 vdd gnd cell_6t
Xbit_r62_c30 bl_30 br_30 wl_62 vdd gnd cell_6t
Xbit_r63_c30 bl_30 br_30 wl_63 vdd gnd cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd cell_6t
Xbit_r1_c31 bl_31 br_31 wl_1 vdd gnd cell_6t
Xbit_r2_c31 bl_31 br_31 wl_2 vdd gnd cell_6t
Xbit_r3_c31 bl_31 br_31 wl_3 vdd gnd cell_6t
Xbit_r4_c31 bl_31 br_31 wl_4 vdd gnd cell_6t
Xbit_r5_c31 bl_31 br_31 wl_5 vdd gnd cell_6t
Xbit_r6_c31 bl_31 br_31 wl_6 vdd gnd cell_6t
Xbit_r7_c31 bl_31 br_31 wl_7 vdd gnd cell_6t
Xbit_r8_c31 bl_31 br_31 wl_8 vdd gnd cell_6t
Xbit_r9_c31 bl_31 br_31 wl_9 vdd gnd cell_6t
Xbit_r10_c31 bl_31 br_31 wl_10 vdd gnd cell_6t
Xbit_r11_c31 bl_31 br_31 wl_11 vdd gnd cell_6t
Xbit_r12_c31 bl_31 br_31 wl_12 vdd gnd cell_6t
Xbit_r13_c31 bl_31 br_31 wl_13 vdd gnd cell_6t
Xbit_r14_c31 bl_31 br_31 wl_14 vdd gnd cell_6t
Xbit_r15_c31 bl_31 br_31 wl_15 vdd gnd cell_6t
Xbit_r16_c31 bl_31 br_31 wl_16 vdd gnd cell_6t
Xbit_r17_c31 bl_31 br_31 wl_17 vdd gnd cell_6t
Xbit_r18_c31 bl_31 br_31 wl_18 vdd gnd cell_6t
Xbit_r19_c31 bl_31 br_31 wl_19 vdd gnd cell_6t
Xbit_r20_c31 bl_31 br_31 wl_20 vdd gnd cell_6t
Xbit_r21_c31 bl_31 br_31 wl_21 vdd gnd cell_6t
Xbit_r22_c31 bl_31 br_31 wl_22 vdd gnd cell_6t
Xbit_r23_c31 bl_31 br_31 wl_23 vdd gnd cell_6t
Xbit_r24_c31 bl_31 br_31 wl_24 vdd gnd cell_6t
Xbit_r25_c31 bl_31 br_31 wl_25 vdd gnd cell_6t
Xbit_r26_c31 bl_31 br_31 wl_26 vdd gnd cell_6t
Xbit_r27_c31 bl_31 br_31 wl_27 vdd gnd cell_6t
Xbit_r28_c31 bl_31 br_31 wl_28 vdd gnd cell_6t
Xbit_r29_c31 bl_31 br_31 wl_29 vdd gnd cell_6t
Xbit_r30_c31 bl_31 br_31 wl_30 vdd gnd cell_6t
Xbit_r31_c31 bl_31 br_31 wl_31 vdd gnd cell_6t
Xbit_r32_c31 bl_31 br_31 wl_32 vdd gnd cell_6t
Xbit_r33_c31 bl_31 br_31 wl_33 vdd gnd cell_6t
Xbit_r34_c31 bl_31 br_31 wl_34 vdd gnd cell_6t
Xbit_r35_c31 bl_31 br_31 wl_35 vdd gnd cell_6t
Xbit_r36_c31 bl_31 br_31 wl_36 vdd gnd cell_6t
Xbit_r37_c31 bl_31 br_31 wl_37 vdd gnd cell_6t
Xbit_r38_c31 bl_31 br_31 wl_38 vdd gnd cell_6t
Xbit_r39_c31 bl_31 br_31 wl_39 vdd gnd cell_6t
Xbit_r40_c31 bl_31 br_31 wl_40 vdd gnd cell_6t
Xbit_r41_c31 bl_31 br_31 wl_41 vdd gnd cell_6t
Xbit_r42_c31 bl_31 br_31 wl_42 vdd gnd cell_6t
Xbit_r43_c31 bl_31 br_31 wl_43 vdd gnd cell_6t
Xbit_r44_c31 bl_31 br_31 wl_44 vdd gnd cell_6t
Xbit_r45_c31 bl_31 br_31 wl_45 vdd gnd cell_6t
Xbit_r46_c31 bl_31 br_31 wl_46 vdd gnd cell_6t
Xbit_r47_c31 bl_31 br_31 wl_47 vdd gnd cell_6t
Xbit_r48_c31 bl_31 br_31 wl_48 vdd gnd cell_6t
Xbit_r49_c31 bl_31 br_31 wl_49 vdd gnd cell_6t
Xbit_r50_c31 bl_31 br_31 wl_50 vdd gnd cell_6t
Xbit_r51_c31 bl_31 br_31 wl_51 vdd gnd cell_6t
Xbit_r52_c31 bl_31 br_31 wl_52 vdd gnd cell_6t
Xbit_r53_c31 bl_31 br_31 wl_53 vdd gnd cell_6t
Xbit_r54_c31 bl_31 br_31 wl_54 vdd gnd cell_6t
Xbit_r55_c31 bl_31 br_31 wl_55 vdd gnd cell_6t
Xbit_r56_c31 bl_31 br_31 wl_56 vdd gnd cell_6t
Xbit_r57_c31 bl_31 br_31 wl_57 vdd gnd cell_6t
Xbit_r58_c31 bl_31 br_31 wl_58 vdd gnd cell_6t
Xbit_r59_c31 bl_31 br_31 wl_59 vdd gnd cell_6t
Xbit_r60_c31 bl_31 br_31 wl_60 vdd gnd cell_6t
Xbit_r61_c31 bl_31 br_31 wl_61 vdd gnd cell_6t
Xbit_r62_c31 bl_31 br_31 wl_62 vdd gnd cell_6t
Xbit_r63_c31 bl_31 br_31 wl_63 vdd gnd cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd cell_6t
Xbit_r1_c32 bl_32 br_32 wl_1 vdd gnd cell_6t
Xbit_r2_c32 bl_32 br_32 wl_2 vdd gnd cell_6t
Xbit_r3_c32 bl_32 br_32 wl_3 vdd gnd cell_6t
Xbit_r4_c32 bl_32 br_32 wl_4 vdd gnd cell_6t
Xbit_r5_c32 bl_32 br_32 wl_5 vdd gnd cell_6t
Xbit_r6_c32 bl_32 br_32 wl_6 vdd gnd cell_6t
Xbit_r7_c32 bl_32 br_32 wl_7 vdd gnd cell_6t
Xbit_r8_c32 bl_32 br_32 wl_8 vdd gnd cell_6t
Xbit_r9_c32 bl_32 br_32 wl_9 vdd gnd cell_6t
Xbit_r10_c32 bl_32 br_32 wl_10 vdd gnd cell_6t
Xbit_r11_c32 bl_32 br_32 wl_11 vdd gnd cell_6t
Xbit_r12_c32 bl_32 br_32 wl_12 vdd gnd cell_6t
Xbit_r13_c32 bl_32 br_32 wl_13 vdd gnd cell_6t
Xbit_r14_c32 bl_32 br_32 wl_14 vdd gnd cell_6t
Xbit_r15_c32 bl_32 br_32 wl_15 vdd gnd cell_6t
Xbit_r16_c32 bl_32 br_32 wl_16 vdd gnd cell_6t
Xbit_r17_c32 bl_32 br_32 wl_17 vdd gnd cell_6t
Xbit_r18_c32 bl_32 br_32 wl_18 vdd gnd cell_6t
Xbit_r19_c32 bl_32 br_32 wl_19 vdd gnd cell_6t
Xbit_r20_c32 bl_32 br_32 wl_20 vdd gnd cell_6t
Xbit_r21_c32 bl_32 br_32 wl_21 vdd gnd cell_6t
Xbit_r22_c32 bl_32 br_32 wl_22 vdd gnd cell_6t
Xbit_r23_c32 bl_32 br_32 wl_23 vdd gnd cell_6t
Xbit_r24_c32 bl_32 br_32 wl_24 vdd gnd cell_6t
Xbit_r25_c32 bl_32 br_32 wl_25 vdd gnd cell_6t
Xbit_r26_c32 bl_32 br_32 wl_26 vdd gnd cell_6t
Xbit_r27_c32 bl_32 br_32 wl_27 vdd gnd cell_6t
Xbit_r28_c32 bl_32 br_32 wl_28 vdd gnd cell_6t
Xbit_r29_c32 bl_32 br_32 wl_29 vdd gnd cell_6t
Xbit_r30_c32 bl_32 br_32 wl_30 vdd gnd cell_6t
Xbit_r31_c32 bl_32 br_32 wl_31 vdd gnd cell_6t
Xbit_r32_c32 bl_32 br_32 wl_32 vdd gnd cell_6t
Xbit_r33_c32 bl_32 br_32 wl_33 vdd gnd cell_6t
Xbit_r34_c32 bl_32 br_32 wl_34 vdd gnd cell_6t
Xbit_r35_c32 bl_32 br_32 wl_35 vdd gnd cell_6t
Xbit_r36_c32 bl_32 br_32 wl_36 vdd gnd cell_6t
Xbit_r37_c32 bl_32 br_32 wl_37 vdd gnd cell_6t
Xbit_r38_c32 bl_32 br_32 wl_38 vdd gnd cell_6t
Xbit_r39_c32 bl_32 br_32 wl_39 vdd gnd cell_6t
Xbit_r40_c32 bl_32 br_32 wl_40 vdd gnd cell_6t
Xbit_r41_c32 bl_32 br_32 wl_41 vdd gnd cell_6t
Xbit_r42_c32 bl_32 br_32 wl_42 vdd gnd cell_6t
Xbit_r43_c32 bl_32 br_32 wl_43 vdd gnd cell_6t
Xbit_r44_c32 bl_32 br_32 wl_44 vdd gnd cell_6t
Xbit_r45_c32 bl_32 br_32 wl_45 vdd gnd cell_6t
Xbit_r46_c32 bl_32 br_32 wl_46 vdd gnd cell_6t
Xbit_r47_c32 bl_32 br_32 wl_47 vdd gnd cell_6t
Xbit_r48_c32 bl_32 br_32 wl_48 vdd gnd cell_6t
Xbit_r49_c32 bl_32 br_32 wl_49 vdd gnd cell_6t
Xbit_r50_c32 bl_32 br_32 wl_50 vdd gnd cell_6t
Xbit_r51_c32 bl_32 br_32 wl_51 vdd gnd cell_6t
Xbit_r52_c32 bl_32 br_32 wl_52 vdd gnd cell_6t
Xbit_r53_c32 bl_32 br_32 wl_53 vdd gnd cell_6t
Xbit_r54_c32 bl_32 br_32 wl_54 vdd gnd cell_6t
Xbit_r55_c32 bl_32 br_32 wl_55 vdd gnd cell_6t
Xbit_r56_c32 bl_32 br_32 wl_56 vdd gnd cell_6t
Xbit_r57_c32 bl_32 br_32 wl_57 vdd gnd cell_6t
Xbit_r58_c32 bl_32 br_32 wl_58 vdd gnd cell_6t
Xbit_r59_c32 bl_32 br_32 wl_59 vdd gnd cell_6t
Xbit_r60_c32 bl_32 br_32 wl_60 vdd gnd cell_6t
Xbit_r61_c32 bl_32 br_32 wl_61 vdd gnd cell_6t
Xbit_r62_c32 bl_32 br_32 wl_62 vdd gnd cell_6t
Xbit_r63_c32 bl_32 br_32 wl_63 vdd gnd cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd cell_6t
Xbit_r1_c33 bl_33 br_33 wl_1 vdd gnd cell_6t
Xbit_r2_c33 bl_33 br_33 wl_2 vdd gnd cell_6t
Xbit_r3_c33 bl_33 br_33 wl_3 vdd gnd cell_6t
Xbit_r4_c33 bl_33 br_33 wl_4 vdd gnd cell_6t
Xbit_r5_c33 bl_33 br_33 wl_5 vdd gnd cell_6t
Xbit_r6_c33 bl_33 br_33 wl_6 vdd gnd cell_6t
Xbit_r7_c33 bl_33 br_33 wl_7 vdd gnd cell_6t
Xbit_r8_c33 bl_33 br_33 wl_8 vdd gnd cell_6t
Xbit_r9_c33 bl_33 br_33 wl_9 vdd gnd cell_6t
Xbit_r10_c33 bl_33 br_33 wl_10 vdd gnd cell_6t
Xbit_r11_c33 bl_33 br_33 wl_11 vdd gnd cell_6t
Xbit_r12_c33 bl_33 br_33 wl_12 vdd gnd cell_6t
Xbit_r13_c33 bl_33 br_33 wl_13 vdd gnd cell_6t
Xbit_r14_c33 bl_33 br_33 wl_14 vdd gnd cell_6t
Xbit_r15_c33 bl_33 br_33 wl_15 vdd gnd cell_6t
Xbit_r16_c33 bl_33 br_33 wl_16 vdd gnd cell_6t
Xbit_r17_c33 bl_33 br_33 wl_17 vdd gnd cell_6t
Xbit_r18_c33 bl_33 br_33 wl_18 vdd gnd cell_6t
Xbit_r19_c33 bl_33 br_33 wl_19 vdd gnd cell_6t
Xbit_r20_c33 bl_33 br_33 wl_20 vdd gnd cell_6t
Xbit_r21_c33 bl_33 br_33 wl_21 vdd gnd cell_6t
Xbit_r22_c33 bl_33 br_33 wl_22 vdd gnd cell_6t
Xbit_r23_c33 bl_33 br_33 wl_23 vdd gnd cell_6t
Xbit_r24_c33 bl_33 br_33 wl_24 vdd gnd cell_6t
Xbit_r25_c33 bl_33 br_33 wl_25 vdd gnd cell_6t
Xbit_r26_c33 bl_33 br_33 wl_26 vdd gnd cell_6t
Xbit_r27_c33 bl_33 br_33 wl_27 vdd gnd cell_6t
Xbit_r28_c33 bl_33 br_33 wl_28 vdd gnd cell_6t
Xbit_r29_c33 bl_33 br_33 wl_29 vdd gnd cell_6t
Xbit_r30_c33 bl_33 br_33 wl_30 vdd gnd cell_6t
Xbit_r31_c33 bl_33 br_33 wl_31 vdd gnd cell_6t
Xbit_r32_c33 bl_33 br_33 wl_32 vdd gnd cell_6t
Xbit_r33_c33 bl_33 br_33 wl_33 vdd gnd cell_6t
Xbit_r34_c33 bl_33 br_33 wl_34 vdd gnd cell_6t
Xbit_r35_c33 bl_33 br_33 wl_35 vdd gnd cell_6t
Xbit_r36_c33 bl_33 br_33 wl_36 vdd gnd cell_6t
Xbit_r37_c33 bl_33 br_33 wl_37 vdd gnd cell_6t
Xbit_r38_c33 bl_33 br_33 wl_38 vdd gnd cell_6t
Xbit_r39_c33 bl_33 br_33 wl_39 vdd gnd cell_6t
Xbit_r40_c33 bl_33 br_33 wl_40 vdd gnd cell_6t
Xbit_r41_c33 bl_33 br_33 wl_41 vdd gnd cell_6t
Xbit_r42_c33 bl_33 br_33 wl_42 vdd gnd cell_6t
Xbit_r43_c33 bl_33 br_33 wl_43 vdd gnd cell_6t
Xbit_r44_c33 bl_33 br_33 wl_44 vdd gnd cell_6t
Xbit_r45_c33 bl_33 br_33 wl_45 vdd gnd cell_6t
Xbit_r46_c33 bl_33 br_33 wl_46 vdd gnd cell_6t
Xbit_r47_c33 bl_33 br_33 wl_47 vdd gnd cell_6t
Xbit_r48_c33 bl_33 br_33 wl_48 vdd gnd cell_6t
Xbit_r49_c33 bl_33 br_33 wl_49 vdd gnd cell_6t
Xbit_r50_c33 bl_33 br_33 wl_50 vdd gnd cell_6t
Xbit_r51_c33 bl_33 br_33 wl_51 vdd gnd cell_6t
Xbit_r52_c33 bl_33 br_33 wl_52 vdd gnd cell_6t
Xbit_r53_c33 bl_33 br_33 wl_53 vdd gnd cell_6t
Xbit_r54_c33 bl_33 br_33 wl_54 vdd gnd cell_6t
Xbit_r55_c33 bl_33 br_33 wl_55 vdd gnd cell_6t
Xbit_r56_c33 bl_33 br_33 wl_56 vdd gnd cell_6t
Xbit_r57_c33 bl_33 br_33 wl_57 vdd gnd cell_6t
Xbit_r58_c33 bl_33 br_33 wl_58 vdd gnd cell_6t
Xbit_r59_c33 bl_33 br_33 wl_59 vdd gnd cell_6t
Xbit_r60_c33 bl_33 br_33 wl_60 vdd gnd cell_6t
Xbit_r61_c33 bl_33 br_33 wl_61 vdd gnd cell_6t
Xbit_r62_c33 bl_33 br_33 wl_62 vdd gnd cell_6t
Xbit_r63_c33 bl_33 br_33 wl_63 vdd gnd cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd cell_6t
Xbit_r1_c34 bl_34 br_34 wl_1 vdd gnd cell_6t
Xbit_r2_c34 bl_34 br_34 wl_2 vdd gnd cell_6t
Xbit_r3_c34 bl_34 br_34 wl_3 vdd gnd cell_6t
Xbit_r4_c34 bl_34 br_34 wl_4 vdd gnd cell_6t
Xbit_r5_c34 bl_34 br_34 wl_5 vdd gnd cell_6t
Xbit_r6_c34 bl_34 br_34 wl_6 vdd gnd cell_6t
Xbit_r7_c34 bl_34 br_34 wl_7 vdd gnd cell_6t
Xbit_r8_c34 bl_34 br_34 wl_8 vdd gnd cell_6t
Xbit_r9_c34 bl_34 br_34 wl_9 vdd gnd cell_6t
Xbit_r10_c34 bl_34 br_34 wl_10 vdd gnd cell_6t
Xbit_r11_c34 bl_34 br_34 wl_11 vdd gnd cell_6t
Xbit_r12_c34 bl_34 br_34 wl_12 vdd gnd cell_6t
Xbit_r13_c34 bl_34 br_34 wl_13 vdd gnd cell_6t
Xbit_r14_c34 bl_34 br_34 wl_14 vdd gnd cell_6t
Xbit_r15_c34 bl_34 br_34 wl_15 vdd gnd cell_6t
Xbit_r16_c34 bl_34 br_34 wl_16 vdd gnd cell_6t
Xbit_r17_c34 bl_34 br_34 wl_17 vdd gnd cell_6t
Xbit_r18_c34 bl_34 br_34 wl_18 vdd gnd cell_6t
Xbit_r19_c34 bl_34 br_34 wl_19 vdd gnd cell_6t
Xbit_r20_c34 bl_34 br_34 wl_20 vdd gnd cell_6t
Xbit_r21_c34 bl_34 br_34 wl_21 vdd gnd cell_6t
Xbit_r22_c34 bl_34 br_34 wl_22 vdd gnd cell_6t
Xbit_r23_c34 bl_34 br_34 wl_23 vdd gnd cell_6t
Xbit_r24_c34 bl_34 br_34 wl_24 vdd gnd cell_6t
Xbit_r25_c34 bl_34 br_34 wl_25 vdd gnd cell_6t
Xbit_r26_c34 bl_34 br_34 wl_26 vdd gnd cell_6t
Xbit_r27_c34 bl_34 br_34 wl_27 vdd gnd cell_6t
Xbit_r28_c34 bl_34 br_34 wl_28 vdd gnd cell_6t
Xbit_r29_c34 bl_34 br_34 wl_29 vdd gnd cell_6t
Xbit_r30_c34 bl_34 br_34 wl_30 vdd gnd cell_6t
Xbit_r31_c34 bl_34 br_34 wl_31 vdd gnd cell_6t
Xbit_r32_c34 bl_34 br_34 wl_32 vdd gnd cell_6t
Xbit_r33_c34 bl_34 br_34 wl_33 vdd gnd cell_6t
Xbit_r34_c34 bl_34 br_34 wl_34 vdd gnd cell_6t
Xbit_r35_c34 bl_34 br_34 wl_35 vdd gnd cell_6t
Xbit_r36_c34 bl_34 br_34 wl_36 vdd gnd cell_6t
Xbit_r37_c34 bl_34 br_34 wl_37 vdd gnd cell_6t
Xbit_r38_c34 bl_34 br_34 wl_38 vdd gnd cell_6t
Xbit_r39_c34 bl_34 br_34 wl_39 vdd gnd cell_6t
Xbit_r40_c34 bl_34 br_34 wl_40 vdd gnd cell_6t
Xbit_r41_c34 bl_34 br_34 wl_41 vdd gnd cell_6t
Xbit_r42_c34 bl_34 br_34 wl_42 vdd gnd cell_6t
Xbit_r43_c34 bl_34 br_34 wl_43 vdd gnd cell_6t
Xbit_r44_c34 bl_34 br_34 wl_44 vdd gnd cell_6t
Xbit_r45_c34 bl_34 br_34 wl_45 vdd gnd cell_6t
Xbit_r46_c34 bl_34 br_34 wl_46 vdd gnd cell_6t
Xbit_r47_c34 bl_34 br_34 wl_47 vdd gnd cell_6t
Xbit_r48_c34 bl_34 br_34 wl_48 vdd gnd cell_6t
Xbit_r49_c34 bl_34 br_34 wl_49 vdd gnd cell_6t
Xbit_r50_c34 bl_34 br_34 wl_50 vdd gnd cell_6t
Xbit_r51_c34 bl_34 br_34 wl_51 vdd gnd cell_6t
Xbit_r52_c34 bl_34 br_34 wl_52 vdd gnd cell_6t
Xbit_r53_c34 bl_34 br_34 wl_53 vdd gnd cell_6t
Xbit_r54_c34 bl_34 br_34 wl_54 vdd gnd cell_6t
Xbit_r55_c34 bl_34 br_34 wl_55 vdd gnd cell_6t
Xbit_r56_c34 bl_34 br_34 wl_56 vdd gnd cell_6t
Xbit_r57_c34 bl_34 br_34 wl_57 vdd gnd cell_6t
Xbit_r58_c34 bl_34 br_34 wl_58 vdd gnd cell_6t
Xbit_r59_c34 bl_34 br_34 wl_59 vdd gnd cell_6t
Xbit_r60_c34 bl_34 br_34 wl_60 vdd gnd cell_6t
Xbit_r61_c34 bl_34 br_34 wl_61 vdd gnd cell_6t
Xbit_r62_c34 bl_34 br_34 wl_62 vdd gnd cell_6t
Xbit_r63_c34 bl_34 br_34 wl_63 vdd gnd cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd cell_6t
Xbit_r1_c35 bl_35 br_35 wl_1 vdd gnd cell_6t
Xbit_r2_c35 bl_35 br_35 wl_2 vdd gnd cell_6t
Xbit_r3_c35 bl_35 br_35 wl_3 vdd gnd cell_6t
Xbit_r4_c35 bl_35 br_35 wl_4 vdd gnd cell_6t
Xbit_r5_c35 bl_35 br_35 wl_5 vdd gnd cell_6t
Xbit_r6_c35 bl_35 br_35 wl_6 vdd gnd cell_6t
Xbit_r7_c35 bl_35 br_35 wl_7 vdd gnd cell_6t
Xbit_r8_c35 bl_35 br_35 wl_8 vdd gnd cell_6t
Xbit_r9_c35 bl_35 br_35 wl_9 vdd gnd cell_6t
Xbit_r10_c35 bl_35 br_35 wl_10 vdd gnd cell_6t
Xbit_r11_c35 bl_35 br_35 wl_11 vdd gnd cell_6t
Xbit_r12_c35 bl_35 br_35 wl_12 vdd gnd cell_6t
Xbit_r13_c35 bl_35 br_35 wl_13 vdd gnd cell_6t
Xbit_r14_c35 bl_35 br_35 wl_14 vdd gnd cell_6t
Xbit_r15_c35 bl_35 br_35 wl_15 vdd gnd cell_6t
Xbit_r16_c35 bl_35 br_35 wl_16 vdd gnd cell_6t
Xbit_r17_c35 bl_35 br_35 wl_17 vdd gnd cell_6t
Xbit_r18_c35 bl_35 br_35 wl_18 vdd gnd cell_6t
Xbit_r19_c35 bl_35 br_35 wl_19 vdd gnd cell_6t
Xbit_r20_c35 bl_35 br_35 wl_20 vdd gnd cell_6t
Xbit_r21_c35 bl_35 br_35 wl_21 vdd gnd cell_6t
Xbit_r22_c35 bl_35 br_35 wl_22 vdd gnd cell_6t
Xbit_r23_c35 bl_35 br_35 wl_23 vdd gnd cell_6t
Xbit_r24_c35 bl_35 br_35 wl_24 vdd gnd cell_6t
Xbit_r25_c35 bl_35 br_35 wl_25 vdd gnd cell_6t
Xbit_r26_c35 bl_35 br_35 wl_26 vdd gnd cell_6t
Xbit_r27_c35 bl_35 br_35 wl_27 vdd gnd cell_6t
Xbit_r28_c35 bl_35 br_35 wl_28 vdd gnd cell_6t
Xbit_r29_c35 bl_35 br_35 wl_29 vdd gnd cell_6t
Xbit_r30_c35 bl_35 br_35 wl_30 vdd gnd cell_6t
Xbit_r31_c35 bl_35 br_35 wl_31 vdd gnd cell_6t
Xbit_r32_c35 bl_35 br_35 wl_32 vdd gnd cell_6t
Xbit_r33_c35 bl_35 br_35 wl_33 vdd gnd cell_6t
Xbit_r34_c35 bl_35 br_35 wl_34 vdd gnd cell_6t
Xbit_r35_c35 bl_35 br_35 wl_35 vdd gnd cell_6t
Xbit_r36_c35 bl_35 br_35 wl_36 vdd gnd cell_6t
Xbit_r37_c35 bl_35 br_35 wl_37 vdd gnd cell_6t
Xbit_r38_c35 bl_35 br_35 wl_38 vdd gnd cell_6t
Xbit_r39_c35 bl_35 br_35 wl_39 vdd gnd cell_6t
Xbit_r40_c35 bl_35 br_35 wl_40 vdd gnd cell_6t
Xbit_r41_c35 bl_35 br_35 wl_41 vdd gnd cell_6t
Xbit_r42_c35 bl_35 br_35 wl_42 vdd gnd cell_6t
Xbit_r43_c35 bl_35 br_35 wl_43 vdd gnd cell_6t
Xbit_r44_c35 bl_35 br_35 wl_44 vdd gnd cell_6t
Xbit_r45_c35 bl_35 br_35 wl_45 vdd gnd cell_6t
Xbit_r46_c35 bl_35 br_35 wl_46 vdd gnd cell_6t
Xbit_r47_c35 bl_35 br_35 wl_47 vdd gnd cell_6t
Xbit_r48_c35 bl_35 br_35 wl_48 vdd gnd cell_6t
Xbit_r49_c35 bl_35 br_35 wl_49 vdd gnd cell_6t
Xbit_r50_c35 bl_35 br_35 wl_50 vdd gnd cell_6t
Xbit_r51_c35 bl_35 br_35 wl_51 vdd gnd cell_6t
Xbit_r52_c35 bl_35 br_35 wl_52 vdd gnd cell_6t
Xbit_r53_c35 bl_35 br_35 wl_53 vdd gnd cell_6t
Xbit_r54_c35 bl_35 br_35 wl_54 vdd gnd cell_6t
Xbit_r55_c35 bl_35 br_35 wl_55 vdd gnd cell_6t
Xbit_r56_c35 bl_35 br_35 wl_56 vdd gnd cell_6t
Xbit_r57_c35 bl_35 br_35 wl_57 vdd gnd cell_6t
Xbit_r58_c35 bl_35 br_35 wl_58 vdd gnd cell_6t
Xbit_r59_c35 bl_35 br_35 wl_59 vdd gnd cell_6t
Xbit_r60_c35 bl_35 br_35 wl_60 vdd gnd cell_6t
Xbit_r61_c35 bl_35 br_35 wl_61 vdd gnd cell_6t
Xbit_r62_c35 bl_35 br_35 wl_62 vdd gnd cell_6t
Xbit_r63_c35 bl_35 br_35 wl_63 vdd gnd cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd cell_6t
Xbit_r1_c36 bl_36 br_36 wl_1 vdd gnd cell_6t
Xbit_r2_c36 bl_36 br_36 wl_2 vdd gnd cell_6t
Xbit_r3_c36 bl_36 br_36 wl_3 vdd gnd cell_6t
Xbit_r4_c36 bl_36 br_36 wl_4 vdd gnd cell_6t
Xbit_r5_c36 bl_36 br_36 wl_5 vdd gnd cell_6t
Xbit_r6_c36 bl_36 br_36 wl_6 vdd gnd cell_6t
Xbit_r7_c36 bl_36 br_36 wl_7 vdd gnd cell_6t
Xbit_r8_c36 bl_36 br_36 wl_8 vdd gnd cell_6t
Xbit_r9_c36 bl_36 br_36 wl_9 vdd gnd cell_6t
Xbit_r10_c36 bl_36 br_36 wl_10 vdd gnd cell_6t
Xbit_r11_c36 bl_36 br_36 wl_11 vdd gnd cell_6t
Xbit_r12_c36 bl_36 br_36 wl_12 vdd gnd cell_6t
Xbit_r13_c36 bl_36 br_36 wl_13 vdd gnd cell_6t
Xbit_r14_c36 bl_36 br_36 wl_14 vdd gnd cell_6t
Xbit_r15_c36 bl_36 br_36 wl_15 vdd gnd cell_6t
Xbit_r16_c36 bl_36 br_36 wl_16 vdd gnd cell_6t
Xbit_r17_c36 bl_36 br_36 wl_17 vdd gnd cell_6t
Xbit_r18_c36 bl_36 br_36 wl_18 vdd gnd cell_6t
Xbit_r19_c36 bl_36 br_36 wl_19 vdd gnd cell_6t
Xbit_r20_c36 bl_36 br_36 wl_20 vdd gnd cell_6t
Xbit_r21_c36 bl_36 br_36 wl_21 vdd gnd cell_6t
Xbit_r22_c36 bl_36 br_36 wl_22 vdd gnd cell_6t
Xbit_r23_c36 bl_36 br_36 wl_23 vdd gnd cell_6t
Xbit_r24_c36 bl_36 br_36 wl_24 vdd gnd cell_6t
Xbit_r25_c36 bl_36 br_36 wl_25 vdd gnd cell_6t
Xbit_r26_c36 bl_36 br_36 wl_26 vdd gnd cell_6t
Xbit_r27_c36 bl_36 br_36 wl_27 vdd gnd cell_6t
Xbit_r28_c36 bl_36 br_36 wl_28 vdd gnd cell_6t
Xbit_r29_c36 bl_36 br_36 wl_29 vdd gnd cell_6t
Xbit_r30_c36 bl_36 br_36 wl_30 vdd gnd cell_6t
Xbit_r31_c36 bl_36 br_36 wl_31 vdd gnd cell_6t
Xbit_r32_c36 bl_36 br_36 wl_32 vdd gnd cell_6t
Xbit_r33_c36 bl_36 br_36 wl_33 vdd gnd cell_6t
Xbit_r34_c36 bl_36 br_36 wl_34 vdd gnd cell_6t
Xbit_r35_c36 bl_36 br_36 wl_35 vdd gnd cell_6t
Xbit_r36_c36 bl_36 br_36 wl_36 vdd gnd cell_6t
Xbit_r37_c36 bl_36 br_36 wl_37 vdd gnd cell_6t
Xbit_r38_c36 bl_36 br_36 wl_38 vdd gnd cell_6t
Xbit_r39_c36 bl_36 br_36 wl_39 vdd gnd cell_6t
Xbit_r40_c36 bl_36 br_36 wl_40 vdd gnd cell_6t
Xbit_r41_c36 bl_36 br_36 wl_41 vdd gnd cell_6t
Xbit_r42_c36 bl_36 br_36 wl_42 vdd gnd cell_6t
Xbit_r43_c36 bl_36 br_36 wl_43 vdd gnd cell_6t
Xbit_r44_c36 bl_36 br_36 wl_44 vdd gnd cell_6t
Xbit_r45_c36 bl_36 br_36 wl_45 vdd gnd cell_6t
Xbit_r46_c36 bl_36 br_36 wl_46 vdd gnd cell_6t
Xbit_r47_c36 bl_36 br_36 wl_47 vdd gnd cell_6t
Xbit_r48_c36 bl_36 br_36 wl_48 vdd gnd cell_6t
Xbit_r49_c36 bl_36 br_36 wl_49 vdd gnd cell_6t
Xbit_r50_c36 bl_36 br_36 wl_50 vdd gnd cell_6t
Xbit_r51_c36 bl_36 br_36 wl_51 vdd gnd cell_6t
Xbit_r52_c36 bl_36 br_36 wl_52 vdd gnd cell_6t
Xbit_r53_c36 bl_36 br_36 wl_53 vdd gnd cell_6t
Xbit_r54_c36 bl_36 br_36 wl_54 vdd gnd cell_6t
Xbit_r55_c36 bl_36 br_36 wl_55 vdd gnd cell_6t
Xbit_r56_c36 bl_36 br_36 wl_56 vdd gnd cell_6t
Xbit_r57_c36 bl_36 br_36 wl_57 vdd gnd cell_6t
Xbit_r58_c36 bl_36 br_36 wl_58 vdd gnd cell_6t
Xbit_r59_c36 bl_36 br_36 wl_59 vdd gnd cell_6t
Xbit_r60_c36 bl_36 br_36 wl_60 vdd gnd cell_6t
Xbit_r61_c36 bl_36 br_36 wl_61 vdd gnd cell_6t
Xbit_r62_c36 bl_36 br_36 wl_62 vdd gnd cell_6t
Xbit_r63_c36 bl_36 br_36 wl_63 vdd gnd cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd cell_6t
Xbit_r1_c37 bl_37 br_37 wl_1 vdd gnd cell_6t
Xbit_r2_c37 bl_37 br_37 wl_2 vdd gnd cell_6t
Xbit_r3_c37 bl_37 br_37 wl_3 vdd gnd cell_6t
Xbit_r4_c37 bl_37 br_37 wl_4 vdd gnd cell_6t
Xbit_r5_c37 bl_37 br_37 wl_5 vdd gnd cell_6t
Xbit_r6_c37 bl_37 br_37 wl_6 vdd gnd cell_6t
Xbit_r7_c37 bl_37 br_37 wl_7 vdd gnd cell_6t
Xbit_r8_c37 bl_37 br_37 wl_8 vdd gnd cell_6t
Xbit_r9_c37 bl_37 br_37 wl_9 vdd gnd cell_6t
Xbit_r10_c37 bl_37 br_37 wl_10 vdd gnd cell_6t
Xbit_r11_c37 bl_37 br_37 wl_11 vdd gnd cell_6t
Xbit_r12_c37 bl_37 br_37 wl_12 vdd gnd cell_6t
Xbit_r13_c37 bl_37 br_37 wl_13 vdd gnd cell_6t
Xbit_r14_c37 bl_37 br_37 wl_14 vdd gnd cell_6t
Xbit_r15_c37 bl_37 br_37 wl_15 vdd gnd cell_6t
Xbit_r16_c37 bl_37 br_37 wl_16 vdd gnd cell_6t
Xbit_r17_c37 bl_37 br_37 wl_17 vdd gnd cell_6t
Xbit_r18_c37 bl_37 br_37 wl_18 vdd gnd cell_6t
Xbit_r19_c37 bl_37 br_37 wl_19 vdd gnd cell_6t
Xbit_r20_c37 bl_37 br_37 wl_20 vdd gnd cell_6t
Xbit_r21_c37 bl_37 br_37 wl_21 vdd gnd cell_6t
Xbit_r22_c37 bl_37 br_37 wl_22 vdd gnd cell_6t
Xbit_r23_c37 bl_37 br_37 wl_23 vdd gnd cell_6t
Xbit_r24_c37 bl_37 br_37 wl_24 vdd gnd cell_6t
Xbit_r25_c37 bl_37 br_37 wl_25 vdd gnd cell_6t
Xbit_r26_c37 bl_37 br_37 wl_26 vdd gnd cell_6t
Xbit_r27_c37 bl_37 br_37 wl_27 vdd gnd cell_6t
Xbit_r28_c37 bl_37 br_37 wl_28 vdd gnd cell_6t
Xbit_r29_c37 bl_37 br_37 wl_29 vdd gnd cell_6t
Xbit_r30_c37 bl_37 br_37 wl_30 vdd gnd cell_6t
Xbit_r31_c37 bl_37 br_37 wl_31 vdd gnd cell_6t
Xbit_r32_c37 bl_37 br_37 wl_32 vdd gnd cell_6t
Xbit_r33_c37 bl_37 br_37 wl_33 vdd gnd cell_6t
Xbit_r34_c37 bl_37 br_37 wl_34 vdd gnd cell_6t
Xbit_r35_c37 bl_37 br_37 wl_35 vdd gnd cell_6t
Xbit_r36_c37 bl_37 br_37 wl_36 vdd gnd cell_6t
Xbit_r37_c37 bl_37 br_37 wl_37 vdd gnd cell_6t
Xbit_r38_c37 bl_37 br_37 wl_38 vdd gnd cell_6t
Xbit_r39_c37 bl_37 br_37 wl_39 vdd gnd cell_6t
Xbit_r40_c37 bl_37 br_37 wl_40 vdd gnd cell_6t
Xbit_r41_c37 bl_37 br_37 wl_41 vdd gnd cell_6t
Xbit_r42_c37 bl_37 br_37 wl_42 vdd gnd cell_6t
Xbit_r43_c37 bl_37 br_37 wl_43 vdd gnd cell_6t
Xbit_r44_c37 bl_37 br_37 wl_44 vdd gnd cell_6t
Xbit_r45_c37 bl_37 br_37 wl_45 vdd gnd cell_6t
Xbit_r46_c37 bl_37 br_37 wl_46 vdd gnd cell_6t
Xbit_r47_c37 bl_37 br_37 wl_47 vdd gnd cell_6t
Xbit_r48_c37 bl_37 br_37 wl_48 vdd gnd cell_6t
Xbit_r49_c37 bl_37 br_37 wl_49 vdd gnd cell_6t
Xbit_r50_c37 bl_37 br_37 wl_50 vdd gnd cell_6t
Xbit_r51_c37 bl_37 br_37 wl_51 vdd gnd cell_6t
Xbit_r52_c37 bl_37 br_37 wl_52 vdd gnd cell_6t
Xbit_r53_c37 bl_37 br_37 wl_53 vdd gnd cell_6t
Xbit_r54_c37 bl_37 br_37 wl_54 vdd gnd cell_6t
Xbit_r55_c37 bl_37 br_37 wl_55 vdd gnd cell_6t
Xbit_r56_c37 bl_37 br_37 wl_56 vdd gnd cell_6t
Xbit_r57_c37 bl_37 br_37 wl_57 vdd gnd cell_6t
Xbit_r58_c37 bl_37 br_37 wl_58 vdd gnd cell_6t
Xbit_r59_c37 bl_37 br_37 wl_59 vdd gnd cell_6t
Xbit_r60_c37 bl_37 br_37 wl_60 vdd gnd cell_6t
Xbit_r61_c37 bl_37 br_37 wl_61 vdd gnd cell_6t
Xbit_r62_c37 bl_37 br_37 wl_62 vdd gnd cell_6t
Xbit_r63_c37 bl_37 br_37 wl_63 vdd gnd cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd cell_6t
Xbit_r1_c38 bl_38 br_38 wl_1 vdd gnd cell_6t
Xbit_r2_c38 bl_38 br_38 wl_2 vdd gnd cell_6t
Xbit_r3_c38 bl_38 br_38 wl_3 vdd gnd cell_6t
Xbit_r4_c38 bl_38 br_38 wl_4 vdd gnd cell_6t
Xbit_r5_c38 bl_38 br_38 wl_5 vdd gnd cell_6t
Xbit_r6_c38 bl_38 br_38 wl_6 vdd gnd cell_6t
Xbit_r7_c38 bl_38 br_38 wl_7 vdd gnd cell_6t
Xbit_r8_c38 bl_38 br_38 wl_8 vdd gnd cell_6t
Xbit_r9_c38 bl_38 br_38 wl_9 vdd gnd cell_6t
Xbit_r10_c38 bl_38 br_38 wl_10 vdd gnd cell_6t
Xbit_r11_c38 bl_38 br_38 wl_11 vdd gnd cell_6t
Xbit_r12_c38 bl_38 br_38 wl_12 vdd gnd cell_6t
Xbit_r13_c38 bl_38 br_38 wl_13 vdd gnd cell_6t
Xbit_r14_c38 bl_38 br_38 wl_14 vdd gnd cell_6t
Xbit_r15_c38 bl_38 br_38 wl_15 vdd gnd cell_6t
Xbit_r16_c38 bl_38 br_38 wl_16 vdd gnd cell_6t
Xbit_r17_c38 bl_38 br_38 wl_17 vdd gnd cell_6t
Xbit_r18_c38 bl_38 br_38 wl_18 vdd gnd cell_6t
Xbit_r19_c38 bl_38 br_38 wl_19 vdd gnd cell_6t
Xbit_r20_c38 bl_38 br_38 wl_20 vdd gnd cell_6t
Xbit_r21_c38 bl_38 br_38 wl_21 vdd gnd cell_6t
Xbit_r22_c38 bl_38 br_38 wl_22 vdd gnd cell_6t
Xbit_r23_c38 bl_38 br_38 wl_23 vdd gnd cell_6t
Xbit_r24_c38 bl_38 br_38 wl_24 vdd gnd cell_6t
Xbit_r25_c38 bl_38 br_38 wl_25 vdd gnd cell_6t
Xbit_r26_c38 bl_38 br_38 wl_26 vdd gnd cell_6t
Xbit_r27_c38 bl_38 br_38 wl_27 vdd gnd cell_6t
Xbit_r28_c38 bl_38 br_38 wl_28 vdd gnd cell_6t
Xbit_r29_c38 bl_38 br_38 wl_29 vdd gnd cell_6t
Xbit_r30_c38 bl_38 br_38 wl_30 vdd gnd cell_6t
Xbit_r31_c38 bl_38 br_38 wl_31 vdd gnd cell_6t
Xbit_r32_c38 bl_38 br_38 wl_32 vdd gnd cell_6t
Xbit_r33_c38 bl_38 br_38 wl_33 vdd gnd cell_6t
Xbit_r34_c38 bl_38 br_38 wl_34 vdd gnd cell_6t
Xbit_r35_c38 bl_38 br_38 wl_35 vdd gnd cell_6t
Xbit_r36_c38 bl_38 br_38 wl_36 vdd gnd cell_6t
Xbit_r37_c38 bl_38 br_38 wl_37 vdd gnd cell_6t
Xbit_r38_c38 bl_38 br_38 wl_38 vdd gnd cell_6t
Xbit_r39_c38 bl_38 br_38 wl_39 vdd gnd cell_6t
Xbit_r40_c38 bl_38 br_38 wl_40 vdd gnd cell_6t
Xbit_r41_c38 bl_38 br_38 wl_41 vdd gnd cell_6t
Xbit_r42_c38 bl_38 br_38 wl_42 vdd gnd cell_6t
Xbit_r43_c38 bl_38 br_38 wl_43 vdd gnd cell_6t
Xbit_r44_c38 bl_38 br_38 wl_44 vdd gnd cell_6t
Xbit_r45_c38 bl_38 br_38 wl_45 vdd gnd cell_6t
Xbit_r46_c38 bl_38 br_38 wl_46 vdd gnd cell_6t
Xbit_r47_c38 bl_38 br_38 wl_47 vdd gnd cell_6t
Xbit_r48_c38 bl_38 br_38 wl_48 vdd gnd cell_6t
Xbit_r49_c38 bl_38 br_38 wl_49 vdd gnd cell_6t
Xbit_r50_c38 bl_38 br_38 wl_50 vdd gnd cell_6t
Xbit_r51_c38 bl_38 br_38 wl_51 vdd gnd cell_6t
Xbit_r52_c38 bl_38 br_38 wl_52 vdd gnd cell_6t
Xbit_r53_c38 bl_38 br_38 wl_53 vdd gnd cell_6t
Xbit_r54_c38 bl_38 br_38 wl_54 vdd gnd cell_6t
Xbit_r55_c38 bl_38 br_38 wl_55 vdd gnd cell_6t
Xbit_r56_c38 bl_38 br_38 wl_56 vdd gnd cell_6t
Xbit_r57_c38 bl_38 br_38 wl_57 vdd gnd cell_6t
Xbit_r58_c38 bl_38 br_38 wl_58 vdd gnd cell_6t
Xbit_r59_c38 bl_38 br_38 wl_59 vdd gnd cell_6t
Xbit_r60_c38 bl_38 br_38 wl_60 vdd gnd cell_6t
Xbit_r61_c38 bl_38 br_38 wl_61 vdd gnd cell_6t
Xbit_r62_c38 bl_38 br_38 wl_62 vdd gnd cell_6t
Xbit_r63_c38 bl_38 br_38 wl_63 vdd gnd cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd cell_6t
Xbit_r1_c39 bl_39 br_39 wl_1 vdd gnd cell_6t
Xbit_r2_c39 bl_39 br_39 wl_2 vdd gnd cell_6t
Xbit_r3_c39 bl_39 br_39 wl_3 vdd gnd cell_6t
Xbit_r4_c39 bl_39 br_39 wl_4 vdd gnd cell_6t
Xbit_r5_c39 bl_39 br_39 wl_5 vdd gnd cell_6t
Xbit_r6_c39 bl_39 br_39 wl_6 vdd gnd cell_6t
Xbit_r7_c39 bl_39 br_39 wl_7 vdd gnd cell_6t
Xbit_r8_c39 bl_39 br_39 wl_8 vdd gnd cell_6t
Xbit_r9_c39 bl_39 br_39 wl_9 vdd gnd cell_6t
Xbit_r10_c39 bl_39 br_39 wl_10 vdd gnd cell_6t
Xbit_r11_c39 bl_39 br_39 wl_11 vdd gnd cell_6t
Xbit_r12_c39 bl_39 br_39 wl_12 vdd gnd cell_6t
Xbit_r13_c39 bl_39 br_39 wl_13 vdd gnd cell_6t
Xbit_r14_c39 bl_39 br_39 wl_14 vdd gnd cell_6t
Xbit_r15_c39 bl_39 br_39 wl_15 vdd gnd cell_6t
Xbit_r16_c39 bl_39 br_39 wl_16 vdd gnd cell_6t
Xbit_r17_c39 bl_39 br_39 wl_17 vdd gnd cell_6t
Xbit_r18_c39 bl_39 br_39 wl_18 vdd gnd cell_6t
Xbit_r19_c39 bl_39 br_39 wl_19 vdd gnd cell_6t
Xbit_r20_c39 bl_39 br_39 wl_20 vdd gnd cell_6t
Xbit_r21_c39 bl_39 br_39 wl_21 vdd gnd cell_6t
Xbit_r22_c39 bl_39 br_39 wl_22 vdd gnd cell_6t
Xbit_r23_c39 bl_39 br_39 wl_23 vdd gnd cell_6t
Xbit_r24_c39 bl_39 br_39 wl_24 vdd gnd cell_6t
Xbit_r25_c39 bl_39 br_39 wl_25 vdd gnd cell_6t
Xbit_r26_c39 bl_39 br_39 wl_26 vdd gnd cell_6t
Xbit_r27_c39 bl_39 br_39 wl_27 vdd gnd cell_6t
Xbit_r28_c39 bl_39 br_39 wl_28 vdd gnd cell_6t
Xbit_r29_c39 bl_39 br_39 wl_29 vdd gnd cell_6t
Xbit_r30_c39 bl_39 br_39 wl_30 vdd gnd cell_6t
Xbit_r31_c39 bl_39 br_39 wl_31 vdd gnd cell_6t
Xbit_r32_c39 bl_39 br_39 wl_32 vdd gnd cell_6t
Xbit_r33_c39 bl_39 br_39 wl_33 vdd gnd cell_6t
Xbit_r34_c39 bl_39 br_39 wl_34 vdd gnd cell_6t
Xbit_r35_c39 bl_39 br_39 wl_35 vdd gnd cell_6t
Xbit_r36_c39 bl_39 br_39 wl_36 vdd gnd cell_6t
Xbit_r37_c39 bl_39 br_39 wl_37 vdd gnd cell_6t
Xbit_r38_c39 bl_39 br_39 wl_38 vdd gnd cell_6t
Xbit_r39_c39 bl_39 br_39 wl_39 vdd gnd cell_6t
Xbit_r40_c39 bl_39 br_39 wl_40 vdd gnd cell_6t
Xbit_r41_c39 bl_39 br_39 wl_41 vdd gnd cell_6t
Xbit_r42_c39 bl_39 br_39 wl_42 vdd gnd cell_6t
Xbit_r43_c39 bl_39 br_39 wl_43 vdd gnd cell_6t
Xbit_r44_c39 bl_39 br_39 wl_44 vdd gnd cell_6t
Xbit_r45_c39 bl_39 br_39 wl_45 vdd gnd cell_6t
Xbit_r46_c39 bl_39 br_39 wl_46 vdd gnd cell_6t
Xbit_r47_c39 bl_39 br_39 wl_47 vdd gnd cell_6t
Xbit_r48_c39 bl_39 br_39 wl_48 vdd gnd cell_6t
Xbit_r49_c39 bl_39 br_39 wl_49 vdd gnd cell_6t
Xbit_r50_c39 bl_39 br_39 wl_50 vdd gnd cell_6t
Xbit_r51_c39 bl_39 br_39 wl_51 vdd gnd cell_6t
Xbit_r52_c39 bl_39 br_39 wl_52 vdd gnd cell_6t
Xbit_r53_c39 bl_39 br_39 wl_53 vdd gnd cell_6t
Xbit_r54_c39 bl_39 br_39 wl_54 vdd gnd cell_6t
Xbit_r55_c39 bl_39 br_39 wl_55 vdd gnd cell_6t
Xbit_r56_c39 bl_39 br_39 wl_56 vdd gnd cell_6t
Xbit_r57_c39 bl_39 br_39 wl_57 vdd gnd cell_6t
Xbit_r58_c39 bl_39 br_39 wl_58 vdd gnd cell_6t
Xbit_r59_c39 bl_39 br_39 wl_59 vdd gnd cell_6t
Xbit_r60_c39 bl_39 br_39 wl_60 vdd gnd cell_6t
Xbit_r61_c39 bl_39 br_39 wl_61 vdd gnd cell_6t
Xbit_r62_c39 bl_39 br_39 wl_62 vdd gnd cell_6t
Xbit_r63_c39 bl_39 br_39 wl_63 vdd gnd cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd cell_6t
Xbit_r1_c40 bl_40 br_40 wl_1 vdd gnd cell_6t
Xbit_r2_c40 bl_40 br_40 wl_2 vdd gnd cell_6t
Xbit_r3_c40 bl_40 br_40 wl_3 vdd gnd cell_6t
Xbit_r4_c40 bl_40 br_40 wl_4 vdd gnd cell_6t
Xbit_r5_c40 bl_40 br_40 wl_5 vdd gnd cell_6t
Xbit_r6_c40 bl_40 br_40 wl_6 vdd gnd cell_6t
Xbit_r7_c40 bl_40 br_40 wl_7 vdd gnd cell_6t
Xbit_r8_c40 bl_40 br_40 wl_8 vdd gnd cell_6t
Xbit_r9_c40 bl_40 br_40 wl_9 vdd gnd cell_6t
Xbit_r10_c40 bl_40 br_40 wl_10 vdd gnd cell_6t
Xbit_r11_c40 bl_40 br_40 wl_11 vdd gnd cell_6t
Xbit_r12_c40 bl_40 br_40 wl_12 vdd gnd cell_6t
Xbit_r13_c40 bl_40 br_40 wl_13 vdd gnd cell_6t
Xbit_r14_c40 bl_40 br_40 wl_14 vdd gnd cell_6t
Xbit_r15_c40 bl_40 br_40 wl_15 vdd gnd cell_6t
Xbit_r16_c40 bl_40 br_40 wl_16 vdd gnd cell_6t
Xbit_r17_c40 bl_40 br_40 wl_17 vdd gnd cell_6t
Xbit_r18_c40 bl_40 br_40 wl_18 vdd gnd cell_6t
Xbit_r19_c40 bl_40 br_40 wl_19 vdd gnd cell_6t
Xbit_r20_c40 bl_40 br_40 wl_20 vdd gnd cell_6t
Xbit_r21_c40 bl_40 br_40 wl_21 vdd gnd cell_6t
Xbit_r22_c40 bl_40 br_40 wl_22 vdd gnd cell_6t
Xbit_r23_c40 bl_40 br_40 wl_23 vdd gnd cell_6t
Xbit_r24_c40 bl_40 br_40 wl_24 vdd gnd cell_6t
Xbit_r25_c40 bl_40 br_40 wl_25 vdd gnd cell_6t
Xbit_r26_c40 bl_40 br_40 wl_26 vdd gnd cell_6t
Xbit_r27_c40 bl_40 br_40 wl_27 vdd gnd cell_6t
Xbit_r28_c40 bl_40 br_40 wl_28 vdd gnd cell_6t
Xbit_r29_c40 bl_40 br_40 wl_29 vdd gnd cell_6t
Xbit_r30_c40 bl_40 br_40 wl_30 vdd gnd cell_6t
Xbit_r31_c40 bl_40 br_40 wl_31 vdd gnd cell_6t
Xbit_r32_c40 bl_40 br_40 wl_32 vdd gnd cell_6t
Xbit_r33_c40 bl_40 br_40 wl_33 vdd gnd cell_6t
Xbit_r34_c40 bl_40 br_40 wl_34 vdd gnd cell_6t
Xbit_r35_c40 bl_40 br_40 wl_35 vdd gnd cell_6t
Xbit_r36_c40 bl_40 br_40 wl_36 vdd gnd cell_6t
Xbit_r37_c40 bl_40 br_40 wl_37 vdd gnd cell_6t
Xbit_r38_c40 bl_40 br_40 wl_38 vdd gnd cell_6t
Xbit_r39_c40 bl_40 br_40 wl_39 vdd gnd cell_6t
Xbit_r40_c40 bl_40 br_40 wl_40 vdd gnd cell_6t
Xbit_r41_c40 bl_40 br_40 wl_41 vdd gnd cell_6t
Xbit_r42_c40 bl_40 br_40 wl_42 vdd gnd cell_6t
Xbit_r43_c40 bl_40 br_40 wl_43 vdd gnd cell_6t
Xbit_r44_c40 bl_40 br_40 wl_44 vdd gnd cell_6t
Xbit_r45_c40 bl_40 br_40 wl_45 vdd gnd cell_6t
Xbit_r46_c40 bl_40 br_40 wl_46 vdd gnd cell_6t
Xbit_r47_c40 bl_40 br_40 wl_47 vdd gnd cell_6t
Xbit_r48_c40 bl_40 br_40 wl_48 vdd gnd cell_6t
Xbit_r49_c40 bl_40 br_40 wl_49 vdd gnd cell_6t
Xbit_r50_c40 bl_40 br_40 wl_50 vdd gnd cell_6t
Xbit_r51_c40 bl_40 br_40 wl_51 vdd gnd cell_6t
Xbit_r52_c40 bl_40 br_40 wl_52 vdd gnd cell_6t
Xbit_r53_c40 bl_40 br_40 wl_53 vdd gnd cell_6t
Xbit_r54_c40 bl_40 br_40 wl_54 vdd gnd cell_6t
Xbit_r55_c40 bl_40 br_40 wl_55 vdd gnd cell_6t
Xbit_r56_c40 bl_40 br_40 wl_56 vdd gnd cell_6t
Xbit_r57_c40 bl_40 br_40 wl_57 vdd gnd cell_6t
Xbit_r58_c40 bl_40 br_40 wl_58 vdd gnd cell_6t
Xbit_r59_c40 bl_40 br_40 wl_59 vdd gnd cell_6t
Xbit_r60_c40 bl_40 br_40 wl_60 vdd gnd cell_6t
Xbit_r61_c40 bl_40 br_40 wl_61 vdd gnd cell_6t
Xbit_r62_c40 bl_40 br_40 wl_62 vdd gnd cell_6t
Xbit_r63_c40 bl_40 br_40 wl_63 vdd gnd cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd cell_6t
Xbit_r1_c41 bl_41 br_41 wl_1 vdd gnd cell_6t
Xbit_r2_c41 bl_41 br_41 wl_2 vdd gnd cell_6t
Xbit_r3_c41 bl_41 br_41 wl_3 vdd gnd cell_6t
Xbit_r4_c41 bl_41 br_41 wl_4 vdd gnd cell_6t
Xbit_r5_c41 bl_41 br_41 wl_5 vdd gnd cell_6t
Xbit_r6_c41 bl_41 br_41 wl_6 vdd gnd cell_6t
Xbit_r7_c41 bl_41 br_41 wl_7 vdd gnd cell_6t
Xbit_r8_c41 bl_41 br_41 wl_8 vdd gnd cell_6t
Xbit_r9_c41 bl_41 br_41 wl_9 vdd gnd cell_6t
Xbit_r10_c41 bl_41 br_41 wl_10 vdd gnd cell_6t
Xbit_r11_c41 bl_41 br_41 wl_11 vdd gnd cell_6t
Xbit_r12_c41 bl_41 br_41 wl_12 vdd gnd cell_6t
Xbit_r13_c41 bl_41 br_41 wl_13 vdd gnd cell_6t
Xbit_r14_c41 bl_41 br_41 wl_14 vdd gnd cell_6t
Xbit_r15_c41 bl_41 br_41 wl_15 vdd gnd cell_6t
Xbit_r16_c41 bl_41 br_41 wl_16 vdd gnd cell_6t
Xbit_r17_c41 bl_41 br_41 wl_17 vdd gnd cell_6t
Xbit_r18_c41 bl_41 br_41 wl_18 vdd gnd cell_6t
Xbit_r19_c41 bl_41 br_41 wl_19 vdd gnd cell_6t
Xbit_r20_c41 bl_41 br_41 wl_20 vdd gnd cell_6t
Xbit_r21_c41 bl_41 br_41 wl_21 vdd gnd cell_6t
Xbit_r22_c41 bl_41 br_41 wl_22 vdd gnd cell_6t
Xbit_r23_c41 bl_41 br_41 wl_23 vdd gnd cell_6t
Xbit_r24_c41 bl_41 br_41 wl_24 vdd gnd cell_6t
Xbit_r25_c41 bl_41 br_41 wl_25 vdd gnd cell_6t
Xbit_r26_c41 bl_41 br_41 wl_26 vdd gnd cell_6t
Xbit_r27_c41 bl_41 br_41 wl_27 vdd gnd cell_6t
Xbit_r28_c41 bl_41 br_41 wl_28 vdd gnd cell_6t
Xbit_r29_c41 bl_41 br_41 wl_29 vdd gnd cell_6t
Xbit_r30_c41 bl_41 br_41 wl_30 vdd gnd cell_6t
Xbit_r31_c41 bl_41 br_41 wl_31 vdd gnd cell_6t
Xbit_r32_c41 bl_41 br_41 wl_32 vdd gnd cell_6t
Xbit_r33_c41 bl_41 br_41 wl_33 vdd gnd cell_6t
Xbit_r34_c41 bl_41 br_41 wl_34 vdd gnd cell_6t
Xbit_r35_c41 bl_41 br_41 wl_35 vdd gnd cell_6t
Xbit_r36_c41 bl_41 br_41 wl_36 vdd gnd cell_6t
Xbit_r37_c41 bl_41 br_41 wl_37 vdd gnd cell_6t
Xbit_r38_c41 bl_41 br_41 wl_38 vdd gnd cell_6t
Xbit_r39_c41 bl_41 br_41 wl_39 vdd gnd cell_6t
Xbit_r40_c41 bl_41 br_41 wl_40 vdd gnd cell_6t
Xbit_r41_c41 bl_41 br_41 wl_41 vdd gnd cell_6t
Xbit_r42_c41 bl_41 br_41 wl_42 vdd gnd cell_6t
Xbit_r43_c41 bl_41 br_41 wl_43 vdd gnd cell_6t
Xbit_r44_c41 bl_41 br_41 wl_44 vdd gnd cell_6t
Xbit_r45_c41 bl_41 br_41 wl_45 vdd gnd cell_6t
Xbit_r46_c41 bl_41 br_41 wl_46 vdd gnd cell_6t
Xbit_r47_c41 bl_41 br_41 wl_47 vdd gnd cell_6t
Xbit_r48_c41 bl_41 br_41 wl_48 vdd gnd cell_6t
Xbit_r49_c41 bl_41 br_41 wl_49 vdd gnd cell_6t
Xbit_r50_c41 bl_41 br_41 wl_50 vdd gnd cell_6t
Xbit_r51_c41 bl_41 br_41 wl_51 vdd gnd cell_6t
Xbit_r52_c41 bl_41 br_41 wl_52 vdd gnd cell_6t
Xbit_r53_c41 bl_41 br_41 wl_53 vdd gnd cell_6t
Xbit_r54_c41 bl_41 br_41 wl_54 vdd gnd cell_6t
Xbit_r55_c41 bl_41 br_41 wl_55 vdd gnd cell_6t
Xbit_r56_c41 bl_41 br_41 wl_56 vdd gnd cell_6t
Xbit_r57_c41 bl_41 br_41 wl_57 vdd gnd cell_6t
Xbit_r58_c41 bl_41 br_41 wl_58 vdd gnd cell_6t
Xbit_r59_c41 bl_41 br_41 wl_59 vdd gnd cell_6t
Xbit_r60_c41 bl_41 br_41 wl_60 vdd gnd cell_6t
Xbit_r61_c41 bl_41 br_41 wl_61 vdd gnd cell_6t
Xbit_r62_c41 bl_41 br_41 wl_62 vdd gnd cell_6t
Xbit_r63_c41 bl_41 br_41 wl_63 vdd gnd cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd cell_6t
Xbit_r1_c42 bl_42 br_42 wl_1 vdd gnd cell_6t
Xbit_r2_c42 bl_42 br_42 wl_2 vdd gnd cell_6t
Xbit_r3_c42 bl_42 br_42 wl_3 vdd gnd cell_6t
Xbit_r4_c42 bl_42 br_42 wl_4 vdd gnd cell_6t
Xbit_r5_c42 bl_42 br_42 wl_5 vdd gnd cell_6t
Xbit_r6_c42 bl_42 br_42 wl_6 vdd gnd cell_6t
Xbit_r7_c42 bl_42 br_42 wl_7 vdd gnd cell_6t
Xbit_r8_c42 bl_42 br_42 wl_8 vdd gnd cell_6t
Xbit_r9_c42 bl_42 br_42 wl_9 vdd gnd cell_6t
Xbit_r10_c42 bl_42 br_42 wl_10 vdd gnd cell_6t
Xbit_r11_c42 bl_42 br_42 wl_11 vdd gnd cell_6t
Xbit_r12_c42 bl_42 br_42 wl_12 vdd gnd cell_6t
Xbit_r13_c42 bl_42 br_42 wl_13 vdd gnd cell_6t
Xbit_r14_c42 bl_42 br_42 wl_14 vdd gnd cell_6t
Xbit_r15_c42 bl_42 br_42 wl_15 vdd gnd cell_6t
Xbit_r16_c42 bl_42 br_42 wl_16 vdd gnd cell_6t
Xbit_r17_c42 bl_42 br_42 wl_17 vdd gnd cell_6t
Xbit_r18_c42 bl_42 br_42 wl_18 vdd gnd cell_6t
Xbit_r19_c42 bl_42 br_42 wl_19 vdd gnd cell_6t
Xbit_r20_c42 bl_42 br_42 wl_20 vdd gnd cell_6t
Xbit_r21_c42 bl_42 br_42 wl_21 vdd gnd cell_6t
Xbit_r22_c42 bl_42 br_42 wl_22 vdd gnd cell_6t
Xbit_r23_c42 bl_42 br_42 wl_23 vdd gnd cell_6t
Xbit_r24_c42 bl_42 br_42 wl_24 vdd gnd cell_6t
Xbit_r25_c42 bl_42 br_42 wl_25 vdd gnd cell_6t
Xbit_r26_c42 bl_42 br_42 wl_26 vdd gnd cell_6t
Xbit_r27_c42 bl_42 br_42 wl_27 vdd gnd cell_6t
Xbit_r28_c42 bl_42 br_42 wl_28 vdd gnd cell_6t
Xbit_r29_c42 bl_42 br_42 wl_29 vdd gnd cell_6t
Xbit_r30_c42 bl_42 br_42 wl_30 vdd gnd cell_6t
Xbit_r31_c42 bl_42 br_42 wl_31 vdd gnd cell_6t
Xbit_r32_c42 bl_42 br_42 wl_32 vdd gnd cell_6t
Xbit_r33_c42 bl_42 br_42 wl_33 vdd gnd cell_6t
Xbit_r34_c42 bl_42 br_42 wl_34 vdd gnd cell_6t
Xbit_r35_c42 bl_42 br_42 wl_35 vdd gnd cell_6t
Xbit_r36_c42 bl_42 br_42 wl_36 vdd gnd cell_6t
Xbit_r37_c42 bl_42 br_42 wl_37 vdd gnd cell_6t
Xbit_r38_c42 bl_42 br_42 wl_38 vdd gnd cell_6t
Xbit_r39_c42 bl_42 br_42 wl_39 vdd gnd cell_6t
Xbit_r40_c42 bl_42 br_42 wl_40 vdd gnd cell_6t
Xbit_r41_c42 bl_42 br_42 wl_41 vdd gnd cell_6t
Xbit_r42_c42 bl_42 br_42 wl_42 vdd gnd cell_6t
Xbit_r43_c42 bl_42 br_42 wl_43 vdd gnd cell_6t
Xbit_r44_c42 bl_42 br_42 wl_44 vdd gnd cell_6t
Xbit_r45_c42 bl_42 br_42 wl_45 vdd gnd cell_6t
Xbit_r46_c42 bl_42 br_42 wl_46 vdd gnd cell_6t
Xbit_r47_c42 bl_42 br_42 wl_47 vdd gnd cell_6t
Xbit_r48_c42 bl_42 br_42 wl_48 vdd gnd cell_6t
Xbit_r49_c42 bl_42 br_42 wl_49 vdd gnd cell_6t
Xbit_r50_c42 bl_42 br_42 wl_50 vdd gnd cell_6t
Xbit_r51_c42 bl_42 br_42 wl_51 vdd gnd cell_6t
Xbit_r52_c42 bl_42 br_42 wl_52 vdd gnd cell_6t
Xbit_r53_c42 bl_42 br_42 wl_53 vdd gnd cell_6t
Xbit_r54_c42 bl_42 br_42 wl_54 vdd gnd cell_6t
Xbit_r55_c42 bl_42 br_42 wl_55 vdd gnd cell_6t
Xbit_r56_c42 bl_42 br_42 wl_56 vdd gnd cell_6t
Xbit_r57_c42 bl_42 br_42 wl_57 vdd gnd cell_6t
Xbit_r58_c42 bl_42 br_42 wl_58 vdd gnd cell_6t
Xbit_r59_c42 bl_42 br_42 wl_59 vdd gnd cell_6t
Xbit_r60_c42 bl_42 br_42 wl_60 vdd gnd cell_6t
Xbit_r61_c42 bl_42 br_42 wl_61 vdd gnd cell_6t
Xbit_r62_c42 bl_42 br_42 wl_62 vdd gnd cell_6t
Xbit_r63_c42 bl_42 br_42 wl_63 vdd gnd cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd cell_6t
Xbit_r1_c43 bl_43 br_43 wl_1 vdd gnd cell_6t
Xbit_r2_c43 bl_43 br_43 wl_2 vdd gnd cell_6t
Xbit_r3_c43 bl_43 br_43 wl_3 vdd gnd cell_6t
Xbit_r4_c43 bl_43 br_43 wl_4 vdd gnd cell_6t
Xbit_r5_c43 bl_43 br_43 wl_5 vdd gnd cell_6t
Xbit_r6_c43 bl_43 br_43 wl_6 vdd gnd cell_6t
Xbit_r7_c43 bl_43 br_43 wl_7 vdd gnd cell_6t
Xbit_r8_c43 bl_43 br_43 wl_8 vdd gnd cell_6t
Xbit_r9_c43 bl_43 br_43 wl_9 vdd gnd cell_6t
Xbit_r10_c43 bl_43 br_43 wl_10 vdd gnd cell_6t
Xbit_r11_c43 bl_43 br_43 wl_11 vdd gnd cell_6t
Xbit_r12_c43 bl_43 br_43 wl_12 vdd gnd cell_6t
Xbit_r13_c43 bl_43 br_43 wl_13 vdd gnd cell_6t
Xbit_r14_c43 bl_43 br_43 wl_14 vdd gnd cell_6t
Xbit_r15_c43 bl_43 br_43 wl_15 vdd gnd cell_6t
Xbit_r16_c43 bl_43 br_43 wl_16 vdd gnd cell_6t
Xbit_r17_c43 bl_43 br_43 wl_17 vdd gnd cell_6t
Xbit_r18_c43 bl_43 br_43 wl_18 vdd gnd cell_6t
Xbit_r19_c43 bl_43 br_43 wl_19 vdd gnd cell_6t
Xbit_r20_c43 bl_43 br_43 wl_20 vdd gnd cell_6t
Xbit_r21_c43 bl_43 br_43 wl_21 vdd gnd cell_6t
Xbit_r22_c43 bl_43 br_43 wl_22 vdd gnd cell_6t
Xbit_r23_c43 bl_43 br_43 wl_23 vdd gnd cell_6t
Xbit_r24_c43 bl_43 br_43 wl_24 vdd gnd cell_6t
Xbit_r25_c43 bl_43 br_43 wl_25 vdd gnd cell_6t
Xbit_r26_c43 bl_43 br_43 wl_26 vdd gnd cell_6t
Xbit_r27_c43 bl_43 br_43 wl_27 vdd gnd cell_6t
Xbit_r28_c43 bl_43 br_43 wl_28 vdd gnd cell_6t
Xbit_r29_c43 bl_43 br_43 wl_29 vdd gnd cell_6t
Xbit_r30_c43 bl_43 br_43 wl_30 vdd gnd cell_6t
Xbit_r31_c43 bl_43 br_43 wl_31 vdd gnd cell_6t
Xbit_r32_c43 bl_43 br_43 wl_32 vdd gnd cell_6t
Xbit_r33_c43 bl_43 br_43 wl_33 vdd gnd cell_6t
Xbit_r34_c43 bl_43 br_43 wl_34 vdd gnd cell_6t
Xbit_r35_c43 bl_43 br_43 wl_35 vdd gnd cell_6t
Xbit_r36_c43 bl_43 br_43 wl_36 vdd gnd cell_6t
Xbit_r37_c43 bl_43 br_43 wl_37 vdd gnd cell_6t
Xbit_r38_c43 bl_43 br_43 wl_38 vdd gnd cell_6t
Xbit_r39_c43 bl_43 br_43 wl_39 vdd gnd cell_6t
Xbit_r40_c43 bl_43 br_43 wl_40 vdd gnd cell_6t
Xbit_r41_c43 bl_43 br_43 wl_41 vdd gnd cell_6t
Xbit_r42_c43 bl_43 br_43 wl_42 vdd gnd cell_6t
Xbit_r43_c43 bl_43 br_43 wl_43 vdd gnd cell_6t
Xbit_r44_c43 bl_43 br_43 wl_44 vdd gnd cell_6t
Xbit_r45_c43 bl_43 br_43 wl_45 vdd gnd cell_6t
Xbit_r46_c43 bl_43 br_43 wl_46 vdd gnd cell_6t
Xbit_r47_c43 bl_43 br_43 wl_47 vdd gnd cell_6t
Xbit_r48_c43 bl_43 br_43 wl_48 vdd gnd cell_6t
Xbit_r49_c43 bl_43 br_43 wl_49 vdd gnd cell_6t
Xbit_r50_c43 bl_43 br_43 wl_50 vdd gnd cell_6t
Xbit_r51_c43 bl_43 br_43 wl_51 vdd gnd cell_6t
Xbit_r52_c43 bl_43 br_43 wl_52 vdd gnd cell_6t
Xbit_r53_c43 bl_43 br_43 wl_53 vdd gnd cell_6t
Xbit_r54_c43 bl_43 br_43 wl_54 vdd gnd cell_6t
Xbit_r55_c43 bl_43 br_43 wl_55 vdd gnd cell_6t
Xbit_r56_c43 bl_43 br_43 wl_56 vdd gnd cell_6t
Xbit_r57_c43 bl_43 br_43 wl_57 vdd gnd cell_6t
Xbit_r58_c43 bl_43 br_43 wl_58 vdd gnd cell_6t
Xbit_r59_c43 bl_43 br_43 wl_59 vdd gnd cell_6t
Xbit_r60_c43 bl_43 br_43 wl_60 vdd gnd cell_6t
Xbit_r61_c43 bl_43 br_43 wl_61 vdd gnd cell_6t
Xbit_r62_c43 bl_43 br_43 wl_62 vdd gnd cell_6t
Xbit_r63_c43 bl_43 br_43 wl_63 vdd gnd cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd cell_6t
Xbit_r1_c44 bl_44 br_44 wl_1 vdd gnd cell_6t
Xbit_r2_c44 bl_44 br_44 wl_2 vdd gnd cell_6t
Xbit_r3_c44 bl_44 br_44 wl_3 vdd gnd cell_6t
Xbit_r4_c44 bl_44 br_44 wl_4 vdd gnd cell_6t
Xbit_r5_c44 bl_44 br_44 wl_5 vdd gnd cell_6t
Xbit_r6_c44 bl_44 br_44 wl_6 vdd gnd cell_6t
Xbit_r7_c44 bl_44 br_44 wl_7 vdd gnd cell_6t
Xbit_r8_c44 bl_44 br_44 wl_8 vdd gnd cell_6t
Xbit_r9_c44 bl_44 br_44 wl_9 vdd gnd cell_6t
Xbit_r10_c44 bl_44 br_44 wl_10 vdd gnd cell_6t
Xbit_r11_c44 bl_44 br_44 wl_11 vdd gnd cell_6t
Xbit_r12_c44 bl_44 br_44 wl_12 vdd gnd cell_6t
Xbit_r13_c44 bl_44 br_44 wl_13 vdd gnd cell_6t
Xbit_r14_c44 bl_44 br_44 wl_14 vdd gnd cell_6t
Xbit_r15_c44 bl_44 br_44 wl_15 vdd gnd cell_6t
Xbit_r16_c44 bl_44 br_44 wl_16 vdd gnd cell_6t
Xbit_r17_c44 bl_44 br_44 wl_17 vdd gnd cell_6t
Xbit_r18_c44 bl_44 br_44 wl_18 vdd gnd cell_6t
Xbit_r19_c44 bl_44 br_44 wl_19 vdd gnd cell_6t
Xbit_r20_c44 bl_44 br_44 wl_20 vdd gnd cell_6t
Xbit_r21_c44 bl_44 br_44 wl_21 vdd gnd cell_6t
Xbit_r22_c44 bl_44 br_44 wl_22 vdd gnd cell_6t
Xbit_r23_c44 bl_44 br_44 wl_23 vdd gnd cell_6t
Xbit_r24_c44 bl_44 br_44 wl_24 vdd gnd cell_6t
Xbit_r25_c44 bl_44 br_44 wl_25 vdd gnd cell_6t
Xbit_r26_c44 bl_44 br_44 wl_26 vdd gnd cell_6t
Xbit_r27_c44 bl_44 br_44 wl_27 vdd gnd cell_6t
Xbit_r28_c44 bl_44 br_44 wl_28 vdd gnd cell_6t
Xbit_r29_c44 bl_44 br_44 wl_29 vdd gnd cell_6t
Xbit_r30_c44 bl_44 br_44 wl_30 vdd gnd cell_6t
Xbit_r31_c44 bl_44 br_44 wl_31 vdd gnd cell_6t
Xbit_r32_c44 bl_44 br_44 wl_32 vdd gnd cell_6t
Xbit_r33_c44 bl_44 br_44 wl_33 vdd gnd cell_6t
Xbit_r34_c44 bl_44 br_44 wl_34 vdd gnd cell_6t
Xbit_r35_c44 bl_44 br_44 wl_35 vdd gnd cell_6t
Xbit_r36_c44 bl_44 br_44 wl_36 vdd gnd cell_6t
Xbit_r37_c44 bl_44 br_44 wl_37 vdd gnd cell_6t
Xbit_r38_c44 bl_44 br_44 wl_38 vdd gnd cell_6t
Xbit_r39_c44 bl_44 br_44 wl_39 vdd gnd cell_6t
Xbit_r40_c44 bl_44 br_44 wl_40 vdd gnd cell_6t
Xbit_r41_c44 bl_44 br_44 wl_41 vdd gnd cell_6t
Xbit_r42_c44 bl_44 br_44 wl_42 vdd gnd cell_6t
Xbit_r43_c44 bl_44 br_44 wl_43 vdd gnd cell_6t
Xbit_r44_c44 bl_44 br_44 wl_44 vdd gnd cell_6t
Xbit_r45_c44 bl_44 br_44 wl_45 vdd gnd cell_6t
Xbit_r46_c44 bl_44 br_44 wl_46 vdd gnd cell_6t
Xbit_r47_c44 bl_44 br_44 wl_47 vdd gnd cell_6t
Xbit_r48_c44 bl_44 br_44 wl_48 vdd gnd cell_6t
Xbit_r49_c44 bl_44 br_44 wl_49 vdd gnd cell_6t
Xbit_r50_c44 bl_44 br_44 wl_50 vdd gnd cell_6t
Xbit_r51_c44 bl_44 br_44 wl_51 vdd gnd cell_6t
Xbit_r52_c44 bl_44 br_44 wl_52 vdd gnd cell_6t
Xbit_r53_c44 bl_44 br_44 wl_53 vdd gnd cell_6t
Xbit_r54_c44 bl_44 br_44 wl_54 vdd gnd cell_6t
Xbit_r55_c44 bl_44 br_44 wl_55 vdd gnd cell_6t
Xbit_r56_c44 bl_44 br_44 wl_56 vdd gnd cell_6t
Xbit_r57_c44 bl_44 br_44 wl_57 vdd gnd cell_6t
Xbit_r58_c44 bl_44 br_44 wl_58 vdd gnd cell_6t
Xbit_r59_c44 bl_44 br_44 wl_59 vdd gnd cell_6t
Xbit_r60_c44 bl_44 br_44 wl_60 vdd gnd cell_6t
Xbit_r61_c44 bl_44 br_44 wl_61 vdd gnd cell_6t
Xbit_r62_c44 bl_44 br_44 wl_62 vdd gnd cell_6t
Xbit_r63_c44 bl_44 br_44 wl_63 vdd gnd cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd cell_6t
Xbit_r1_c45 bl_45 br_45 wl_1 vdd gnd cell_6t
Xbit_r2_c45 bl_45 br_45 wl_2 vdd gnd cell_6t
Xbit_r3_c45 bl_45 br_45 wl_3 vdd gnd cell_6t
Xbit_r4_c45 bl_45 br_45 wl_4 vdd gnd cell_6t
Xbit_r5_c45 bl_45 br_45 wl_5 vdd gnd cell_6t
Xbit_r6_c45 bl_45 br_45 wl_6 vdd gnd cell_6t
Xbit_r7_c45 bl_45 br_45 wl_7 vdd gnd cell_6t
Xbit_r8_c45 bl_45 br_45 wl_8 vdd gnd cell_6t
Xbit_r9_c45 bl_45 br_45 wl_9 vdd gnd cell_6t
Xbit_r10_c45 bl_45 br_45 wl_10 vdd gnd cell_6t
Xbit_r11_c45 bl_45 br_45 wl_11 vdd gnd cell_6t
Xbit_r12_c45 bl_45 br_45 wl_12 vdd gnd cell_6t
Xbit_r13_c45 bl_45 br_45 wl_13 vdd gnd cell_6t
Xbit_r14_c45 bl_45 br_45 wl_14 vdd gnd cell_6t
Xbit_r15_c45 bl_45 br_45 wl_15 vdd gnd cell_6t
Xbit_r16_c45 bl_45 br_45 wl_16 vdd gnd cell_6t
Xbit_r17_c45 bl_45 br_45 wl_17 vdd gnd cell_6t
Xbit_r18_c45 bl_45 br_45 wl_18 vdd gnd cell_6t
Xbit_r19_c45 bl_45 br_45 wl_19 vdd gnd cell_6t
Xbit_r20_c45 bl_45 br_45 wl_20 vdd gnd cell_6t
Xbit_r21_c45 bl_45 br_45 wl_21 vdd gnd cell_6t
Xbit_r22_c45 bl_45 br_45 wl_22 vdd gnd cell_6t
Xbit_r23_c45 bl_45 br_45 wl_23 vdd gnd cell_6t
Xbit_r24_c45 bl_45 br_45 wl_24 vdd gnd cell_6t
Xbit_r25_c45 bl_45 br_45 wl_25 vdd gnd cell_6t
Xbit_r26_c45 bl_45 br_45 wl_26 vdd gnd cell_6t
Xbit_r27_c45 bl_45 br_45 wl_27 vdd gnd cell_6t
Xbit_r28_c45 bl_45 br_45 wl_28 vdd gnd cell_6t
Xbit_r29_c45 bl_45 br_45 wl_29 vdd gnd cell_6t
Xbit_r30_c45 bl_45 br_45 wl_30 vdd gnd cell_6t
Xbit_r31_c45 bl_45 br_45 wl_31 vdd gnd cell_6t
Xbit_r32_c45 bl_45 br_45 wl_32 vdd gnd cell_6t
Xbit_r33_c45 bl_45 br_45 wl_33 vdd gnd cell_6t
Xbit_r34_c45 bl_45 br_45 wl_34 vdd gnd cell_6t
Xbit_r35_c45 bl_45 br_45 wl_35 vdd gnd cell_6t
Xbit_r36_c45 bl_45 br_45 wl_36 vdd gnd cell_6t
Xbit_r37_c45 bl_45 br_45 wl_37 vdd gnd cell_6t
Xbit_r38_c45 bl_45 br_45 wl_38 vdd gnd cell_6t
Xbit_r39_c45 bl_45 br_45 wl_39 vdd gnd cell_6t
Xbit_r40_c45 bl_45 br_45 wl_40 vdd gnd cell_6t
Xbit_r41_c45 bl_45 br_45 wl_41 vdd gnd cell_6t
Xbit_r42_c45 bl_45 br_45 wl_42 vdd gnd cell_6t
Xbit_r43_c45 bl_45 br_45 wl_43 vdd gnd cell_6t
Xbit_r44_c45 bl_45 br_45 wl_44 vdd gnd cell_6t
Xbit_r45_c45 bl_45 br_45 wl_45 vdd gnd cell_6t
Xbit_r46_c45 bl_45 br_45 wl_46 vdd gnd cell_6t
Xbit_r47_c45 bl_45 br_45 wl_47 vdd gnd cell_6t
Xbit_r48_c45 bl_45 br_45 wl_48 vdd gnd cell_6t
Xbit_r49_c45 bl_45 br_45 wl_49 vdd gnd cell_6t
Xbit_r50_c45 bl_45 br_45 wl_50 vdd gnd cell_6t
Xbit_r51_c45 bl_45 br_45 wl_51 vdd gnd cell_6t
Xbit_r52_c45 bl_45 br_45 wl_52 vdd gnd cell_6t
Xbit_r53_c45 bl_45 br_45 wl_53 vdd gnd cell_6t
Xbit_r54_c45 bl_45 br_45 wl_54 vdd gnd cell_6t
Xbit_r55_c45 bl_45 br_45 wl_55 vdd gnd cell_6t
Xbit_r56_c45 bl_45 br_45 wl_56 vdd gnd cell_6t
Xbit_r57_c45 bl_45 br_45 wl_57 vdd gnd cell_6t
Xbit_r58_c45 bl_45 br_45 wl_58 vdd gnd cell_6t
Xbit_r59_c45 bl_45 br_45 wl_59 vdd gnd cell_6t
Xbit_r60_c45 bl_45 br_45 wl_60 vdd gnd cell_6t
Xbit_r61_c45 bl_45 br_45 wl_61 vdd gnd cell_6t
Xbit_r62_c45 bl_45 br_45 wl_62 vdd gnd cell_6t
Xbit_r63_c45 bl_45 br_45 wl_63 vdd gnd cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd cell_6t
Xbit_r1_c46 bl_46 br_46 wl_1 vdd gnd cell_6t
Xbit_r2_c46 bl_46 br_46 wl_2 vdd gnd cell_6t
Xbit_r3_c46 bl_46 br_46 wl_3 vdd gnd cell_6t
Xbit_r4_c46 bl_46 br_46 wl_4 vdd gnd cell_6t
Xbit_r5_c46 bl_46 br_46 wl_5 vdd gnd cell_6t
Xbit_r6_c46 bl_46 br_46 wl_6 vdd gnd cell_6t
Xbit_r7_c46 bl_46 br_46 wl_7 vdd gnd cell_6t
Xbit_r8_c46 bl_46 br_46 wl_8 vdd gnd cell_6t
Xbit_r9_c46 bl_46 br_46 wl_9 vdd gnd cell_6t
Xbit_r10_c46 bl_46 br_46 wl_10 vdd gnd cell_6t
Xbit_r11_c46 bl_46 br_46 wl_11 vdd gnd cell_6t
Xbit_r12_c46 bl_46 br_46 wl_12 vdd gnd cell_6t
Xbit_r13_c46 bl_46 br_46 wl_13 vdd gnd cell_6t
Xbit_r14_c46 bl_46 br_46 wl_14 vdd gnd cell_6t
Xbit_r15_c46 bl_46 br_46 wl_15 vdd gnd cell_6t
Xbit_r16_c46 bl_46 br_46 wl_16 vdd gnd cell_6t
Xbit_r17_c46 bl_46 br_46 wl_17 vdd gnd cell_6t
Xbit_r18_c46 bl_46 br_46 wl_18 vdd gnd cell_6t
Xbit_r19_c46 bl_46 br_46 wl_19 vdd gnd cell_6t
Xbit_r20_c46 bl_46 br_46 wl_20 vdd gnd cell_6t
Xbit_r21_c46 bl_46 br_46 wl_21 vdd gnd cell_6t
Xbit_r22_c46 bl_46 br_46 wl_22 vdd gnd cell_6t
Xbit_r23_c46 bl_46 br_46 wl_23 vdd gnd cell_6t
Xbit_r24_c46 bl_46 br_46 wl_24 vdd gnd cell_6t
Xbit_r25_c46 bl_46 br_46 wl_25 vdd gnd cell_6t
Xbit_r26_c46 bl_46 br_46 wl_26 vdd gnd cell_6t
Xbit_r27_c46 bl_46 br_46 wl_27 vdd gnd cell_6t
Xbit_r28_c46 bl_46 br_46 wl_28 vdd gnd cell_6t
Xbit_r29_c46 bl_46 br_46 wl_29 vdd gnd cell_6t
Xbit_r30_c46 bl_46 br_46 wl_30 vdd gnd cell_6t
Xbit_r31_c46 bl_46 br_46 wl_31 vdd gnd cell_6t
Xbit_r32_c46 bl_46 br_46 wl_32 vdd gnd cell_6t
Xbit_r33_c46 bl_46 br_46 wl_33 vdd gnd cell_6t
Xbit_r34_c46 bl_46 br_46 wl_34 vdd gnd cell_6t
Xbit_r35_c46 bl_46 br_46 wl_35 vdd gnd cell_6t
Xbit_r36_c46 bl_46 br_46 wl_36 vdd gnd cell_6t
Xbit_r37_c46 bl_46 br_46 wl_37 vdd gnd cell_6t
Xbit_r38_c46 bl_46 br_46 wl_38 vdd gnd cell_6t
Xbit_r39_c46 bl_46 br_46 wl_39 vdd gnd cell_6t
Xbit_r40_c46 bl_46 br_46 wl_40 vdd gnd cell_6t
Xbit_r41_c46 bl_46 br_46 wl_41 vdd gnd cell_6t
Xbit_r42_c46 bl_46 br_46 wl_42 vdd gnd cell_6t
Xbit_r43_c46 bl_46 br_46 wl_43 vdd gnd cell_6t
Xbit_r44_c46 bl_46 br_46 wl_44 vdd gnd cell_6t
Xbit_r45_c46 bl_46 br_46 wl_45 vdd gnd cell_6t
Xbit_r46_c46 bl_46 br_46 wl_46 vdd gnd cell_6t
Xbit_r47_c46 bl_46 br_46 wl_47 vdd gnd cell_6t
Xbit_r48_c46 bl_46 br_46 wl_48 vdd gnd cell_6t
Xbit_r49_c46 bl_46 br_46 wl_49 vdd gnd cell_6t
Xbit_r50_c46 bl_46 br_46 wl_50 vdd gnd cell_6t
Xbit_r51_c46 bl_46 br_46 wl_51 vdd gnd cell_6t
Xbit_r52_c46 bl_46 br_46 wl_52 vdd gnd cell_6t
Xbit_r53_c46 bl_46 br_46 wl_53 vdd gnd cell_6t
Xbit_r54_c46 bl_46 br_46 wl_54 vdd gnd cell_6t
Xbit_r55_c46 bl_46 br_46 wl_55 vdd gnd cell_6t
Xbit_r56_c46 bl_46 br_46 wl_56 vdd gnd cell_6t
Xbit_r57_c46 bl_46 br_46 wl_57 vdd gnd cell_6t
Xbit_r58_c46 bl_46 br_46 wl_58 vdd gnd cell_6t
Xbit_r59_c46 bl_46 br_46 wl_59 vdd gnd cell_6t
Xbit_r60_c46 bl_46 br_46 wl_60 vdd gnd cell_6t
Xbit_r61_c46 bl_46 br_46 wl_61 vdd gnd cell_6t
Xbit_r62_c46 bl_46 br_46 wl_62 vdd gnd cell_6t
Xbit_r63_c46 bl_46 br_46 wl_63 vdd gnd cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd cell_6t
Xbit_r1_c47 bl_47 br_47 wl_1 vdd gnd cell_6t
Xbit_r2_c47 bl_47 br_47 wl_2 vdd gnd cell_6t
Xbit_r3_c47 bl_47 br_47 wl_3 vdd gnd cell_6t
Xbit_r4_c47 bl_47 br_47 wl_4 vdd gnd cell_6t
Xbit_r5_c47 bl_47 br_47 wl_5 vdd gnd cell_6t
Xbit_r6_c47 bl_47 br_47 wl_6 vdd gnd cell_6t
Xbit_r7_c47 bl_47 br_47 wl_7 vdd gnd cell_6t
Xbit_r8_c47 bl_47 br_47 wl_8 vdd gnd cell_6t
Xbit_r9_c47 bl_47 br_47 wl_9 vdd gnd cell_6t
Xbit_r10_c47 bl_47 br_47 wl_10 vdd gnd cell_6t
Xbit_r11_c47 bl_47 br_47 wl_11 vdd gnd cell_6t
Xbit_r12_c47 bl_47 br_47 wl_12 vdd gnd cell_6t
Xbit_r13_c47 bl_47 br_47 wl_13 vdd gnd cell_6t
Xbit_r14_c47 bl_47 br_47 wl_14 vdd gnd cell_6t
Xbit_r15_c47 bl_47 br_47 wl_15 vdd gnd cell_6t
Xbit_r16_c47 bl_47 br_47 wl_16 vdd gnd cell_6t
Xbit_r17_c47 bl_47 br_47 wl_17 vdd gnd cell_6t
Xbit_r18_c47 bl_47 br_47 wl_18 vdd gnd cell_6t
Xbit_r19_c47 bl_47 br_47 wl_19 vdd gnd cell_6t
Xbit_r20_c47 bl_47 br_47 wl_20 vdd gnd cell_6t
Xbit_r21_c47 bl_47 br_47 wl_21 vdd gnd cell_6t
Xbit_r22_c47 bl_47 br_47 wl_22 vdd gnd cell_6t
Xbit_r23_c47 bl_47 br_47 wl_23 vdd gnd cell_6t
Xbit_r24_c47 bl_47 br_47 wl_24 vdd gnd cell_6t
Xbit_r25_c47 bl_47 br_47 wl_25 vdd gnd cell_6t
Xbit_r26_c47 bl_47 br_47 wl_26 vdd gnd cell_6t
Xbit_r27_c47 bl_47 br_47 wl_27 vdd gnd cell_6t
Xbit_r28_c47 bl_47 br_47 wl_28 vdd gnd cell_6t
Xbit_r29_c47 bl_47 br_47 wl_29 vdd gnd cell_6t
Xbit_r30_c47 bl_47 br_47 wl_30 vdd gnd cell_6t
Xbit_r31_c47 bl_47 br_47 wl_31 vdd gnd cell_6t
Xbit_r32_c47 bl_47 br_47 wl_32 vdd gnd cell_6t
Xbit_r33_c47 bl_47 br_47 wl_33 vdd gnd cell_6t
Xbit_r34_c47 bl_47 br_47 wl_34 vdd gnd cell_6t
Xbit_r35_c47 bl_47 br_47 wl_35 vdd gnd cell_6t
Xbit_r36_c47 bl_47 br_47 wl_36 vdd gnd cell_6t
Xbit_r37_c47 bl_47 br_47 wl_37 vdd gnd cell_6t
Xbit_r38_c47 bl_47 br_47 wl_38 vdd gnd cell_6t
Xbit_r39_c47 bl_47 br_47 wl_39 vdd gnd cell_6t
Xbit_r40_c47 bl_47 br_47 wl_40 vdd gnd cell_6t
Xbit_r41_c47 bl_47 br_47 wl_41 vdd gnd cell_6t
Xbit_r42_c47 bl_47 br_47 wl_42 vdd gnd cell_6t
Xbit_r43_c47 bl_47 br_47 wl_43 vdd gnd cell_6t
Xbit_r44_c47 bl_47 br_47 wl_44 vdd gnd cell_6t
Xbit_r45_c47 bl_47 br_47 wl_45 vdd gnd cell_6t
Xbit_r46_c47 bl_47 br_47 wl_46 vdd gnd cell_6t
Xbit_r47_c47 bl_47 br_47 wl_47 vdd gnd cell_6t
Xbit_r48_c47 bl_47 br_47 wl_48 vdd gnd cell_6t
Xbit_r49_c47 bl_47 br_47 wl_49 vdd gnd cell_6t
Xbit_r50_c47 bl_47 br_47 wl_50 vdd gnd cell_6t
Xbit_r51_c47 bl_47 br_47 wl_51 vdd gnd cell_6t
Xbit_r52_c47 bl_47 br_47 wl_52 vdd gnd cell_6t
Xbit_r53_c47 bl_47 br_47 wl_53 vdd gnd cell_6t
Xbit_r54_c47 bl_47 br_47 wl_54 vdd gnd cell_6t
Xbit_r55_c47 bl_47 br_47 wl_55 vdd gnd cell_6t
Xbit_r56_c47 bl_47 br_47 wl_56 vdd gnd cell_6t
Xbit_r57_c47 bl_47 br_47 wl_57 vdd gnd cell_6t
Xbit_r58_c47 bl_47 br_47 wl_58 vdd gnd cell_6t
Xbit_r59_c47 bl_47 br_47 wl_59 vdd gnd cell_6t
Xbit_r60_c47 bl_47 br_47 wl_60 vdd gnd cell_6t
Xbit_r61_c47 bl_47 br_47 wl_61 vdd gnd cell_6t
Xbit_r62_c47 bl_47 br_47 wl_62 vdd gnd cell_6t
Xbit_r63_c47 bl_47 br_47 wl_63 vdd gnd cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd cell_6t
Xbit_r1_c48 bl_48 br_48 wl_1 vdd gnd cell_6t
Xbit_r2_c48 bl_48 br_48 wl_2 vdd gnd cell_6t
Xbit_r3_c48 bl_48 br_48 wl_3 vdd gnd cell_6t
Xbit_r4_c48 bl_48 br_48 wl_4 vdd gnd cell_6t
Xbit_r5_c48 bl_48 br_48 wl_5 vdd gnd cell_6t
Xbit_r6_c48 bl_48 br_48 wl_6 vdd gnd cell_6t
Xbit_r7_c48 bl_48 br_48 wl_7 vdd gnd cell_6t
Xbit_r8_c48 bl_48 br_48 wl_8 vdd gnd cell_6t
Xbit_r9_c48 bl_48 br_48 wl_9 vdd gnd cell_6t
Xbit_r10_c48 bl_48 br_48 wl_10 vdd gnd cell_6t
Xbit_r11_c48 bl_48 br_48 wl_11 vdd gnd cell_6t
Xbit_r12_c48 bl_48 br_48 wl_12 vdd gnd cell_6t
Xbit_r13_c48 bl_48 br_48 wl_13 vdd gnd cell_6t
Xbit_r14_c48 bl_48 br_48 wl_14 vdd gnd cell_6t
Xbit_r15_c48 bl_48 br_48 wl_15 vdd gnd cell_6t
Xbit_r16_c48 bl_48 br_48 wl_16 vdd gnd cell_6t
Xbit_r17_c48 bl_48 br_48 wl_17 vdd gnd cell_6t
Xbit_r18_c48 bl_48 br_48 wl_18 vdd gnd cell_6t
Xbit_r19_c48 bl_48 br_48 wl_19 vdd gnd cell_6t
Xbit_r20_c48 bl_48 br_48 wl_20 vdd gnd cell_6t
Xbit_r21_c48 bl_48 br_48 wl_21 vdd gnd cell_6t
Xbit_r22_c48 bl_48 br_48 wl_22 vdd gnd cell_6t
Xbit_r23_c48 bl_48 br_48 wl_23 vdd gnd cell_6t
Xbit_r24_c48 bl_48 br_48 wl_24 vdd gnd cell_6t
Xbit_r25_c48 bl_48 br_48 wl_25 vdd gnd cell_6t
Xbit_r26_c48 bl_48 br_48 wl_26 vdd gnd cell_6t
Xbit_r27_c48 bl_48 br_48 wl_27 vdd gnd cell_6t
Xbit_r28_c48 bl_48 br_48 wl_28 vdd gnd cell_6t
Xbit_r29_c48 bl_48 br_48 wl_29 vdd gnd cell_6t
Xbit_r30_c48 bl_48 br_48 wl_30 vdd gnd cell_6t
Xbit_r31_c48 bl_48 br_48 wl_31 vdd gnd cell_6t
Xbit_r32_c48 bl_48 br_48 wl_32 vdd gnd cell_6t
Xbit_r33_c48 bl_48 br_48 wl_33 vdd gnd cell_6t
Xbit_r34_c48 bl_48 br_48 wl_34 vdd gnd cell_6t
Xbit_r35_c48 bl_48 br_48 wl_35 vdd gnd cell_6t
Xbit_r36_c48 bl_48 br_48 wl_36 vdd gnd cell_6t
Xbit_r37_c48 bl_48 br_48 wl_37 vdd gnd cell_6t
Xbit_r38_c48 bl_48 br_48 wl_38 vdd gnd cell_6t
Xbit_r39_c48 bl_48 br_48 wl_39 vdd gnd cell_6t
Xbit_r40_c48 bl_48 br_48 wl_40 vdd gnd cell_6t
Xbit_r41_c48 bl_48 br_48 wl_41 vdd gnd cell_6t
Xbit_r42_c48 bl_48 br_48 wl_42 vdd gnd cell_6t
Xbit_r43_c48 bl_48 br_48 wl_43 vdd gnd cell_6t
Xbit_r44_c48 bl_48 br_48 wl_44 vdd gnd cell_6t
Xbit_r45_c48 bl_48 br_48 wl_45 vdd gnd cell_6t
Xbit_r46_c48 bl_48 br_48 wl_46 vdd gnd cell_6t
Xbit_r47_c48 bl_48 br_48 wl_47 vdd gnd cell_6t
Xbit_r48_c48 bl_48 br_48 wl_48 vdd gnd cell_6t
Xbit_r49_c48 bl_48 br_48 wl_49 vdd gnd cell_6t
Xbit_r50_c48 bl_48 br_48 wl_50 vdd gnd cell_6t
Xbit_r51_c48 bl_48 br_48 wl_51 vdd gnd cell_6t
Xbit_r52_c48 bl_48 br_48 wl_52 vdd gnd cell_6t
Xbit_r53_c48 bl_48 br_48 wl_53 vdd gnd cell_6t
Xbit_r54_c48 bl_48 br_48 wl_54 vdd gnd cell_6t
Xbit_r55_c48 bl_48 br_48 wl_55 vdd gnd cell_6t
Xbit_r56_c48 bl_48 br_48 wl_56 vdd gnd cell_6t
Xbit_r57_c48 bl_48 br_48 wl_57 vdd gnd cell_6t
Xbit_r58_c48 bl_48 br_48 wl_58 vdd gnd cell_6t
Xbit_r59_c48 bl_48 br_48 wl_59 vdd gnd cell_6t
Xbit_r60_c48 bl_48 br_48 wl_60 vdd gnd cell_6t
Xbit_r61_c48 bl_48 br_48 wl_61 vdd gnd cell_6t
Xbit_r62_c48 bl_48 br_48 wl_62 vdd gnd cell_6t
Xbit_r63_c48 bl_48 br_48 wl_63 vdd gnd cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd cell_6t
Xbit_r1_c49 bl_49 br_49 wl_1 vdd gnd cell_6t
Xbit_r2_c49 bl_49 br_49 wl_2 vdd gnd cell_6t
Xbit_r3_c49 bl_49 br_49 wl_3 vdd gnd cell_6t
Xbit_r4_c49 bl_49 br_49 wl_4 vdd gnd cell_6t
Xbit_r5_c49 bl_49 br_49 wl_5 vdd gnd cell_6t
Xbit_r6_c49 bl_49 br_49 wl_6 vdd gnd cell_6t
Xbit_r7_c49 bl_49 br_49 wl_7 vdd gnd cell_6t
Xbit_r8_c49 bl_49 br_49 wl_8 vdd gnd cell_6t
Xbit_r9_c49 bl_49 br_49 wl_9 vdd gnd cell_6t
Xbit_r10_c49 bl_49 br_49 wl_10 vdd gnd cell_6t
Xbit_r11_c49 bl_49 br_49 wl_11 vdd gnd cell_6t
Xbit_r12_c49 bl_49 br_49 wl_12 vdd gnd cell_6t
Xbit_r13_c49 bl_49 br_49 wl_13 vdd gnd cell_6t
Xbit_r14_c49 bl_49 br_49 wl_14 vdd gnd cell_6t
Xbit_r15_c49 bl_49 br_49 wl_15 vdd gnd cell_6t
Xbit_r16_c49 bl_49 br_49 wl_16 vdd gnd cell_6t
Xbit_r17_c49 bl_49 br_49 wl_17 vdd gnd cell_6t
Xbit_r18_c49 bl_49 br_49 wl_18 vdd gnd cell_6t
Xbit_r19_c49 bl_49 br_49 wl_19 vdd gnd cell_6t
Xbit_r20_c49 bl_49 br_49 wl_20 vdd gnd cell_6t
Xbit_r21_c49 bl_49 br_49 wl_21 vdd gnd cell_6t
Xbit_r22_c49 bl_49 br_49 wl_22 vdd gnd cell_6t
Xbit_r23_c49 bl_49 br_49 wl_23 vdd gnd cell_6t
Xbit_r24_c49 bl_49 br_49 wl_24 vdd gnd cell_6t
Xbit_r25_c49 bl_49 br_49 wl_25 vdd gnd cell_6t
Xbit_r26_c49 bl_49 br_49 wl_26 vdd gnd cell_6t
Xbit_r27_c49 bl_49 br_49 wl_27 vdd gnd cell_6t
Xbit_r28_c49 bl_49 br_49 wl_28 vdd gnd cell_6t
Xbit_r29_c49 bl_49 br_49 wl_29 vdd gnd cell_6t
Xbit_r30_c49 bl_49 br_49 wl_30 vdd gnd cell_6t
Xbit_r31_c49 bl_49 br_49 wl_31 vdd gnd cell_6t
Xbit_r32_c49 bl_49 br_49 wl_32 vdd gnd cell_6t
Xbit_r33_c49 bl_49 br_49 wl_33 vdd gnd cell_6t
Xbit_r34_c49 bl_49 br_49 wl_34 vdd gnd cell_6t
Xbit_r35_c49 bl_49 br_49 wl_35 vdd gnd cell_6t
Xbit_r36_c49 bl_49 br_49 wl_36 vdd gnd cell_6t
Xbit_r37_c49 bl_49 br_49 wl_37 vdd gnd cell_6t
Xbit_r38_c49 bl_49 br_49 wl_38 vdd gnd cell_6t
Xbit_r39_c49 bl_49 br_49 wl_39 vdd gnd cell_6t
Xbit_r40_c49 bl_49 br_49 wl_40 vdd gnd cell_6t
Xbit_r41_c49 bl_49 br_49 wl_41 vdd gnd cell_6t
Xbit_r42_c49 bl_49 br_49 wl_42 vdd gnd cell_6t
Xbit_r43_c49 bl_49 br_49 wl_43 vdd gnd cell_6t
Xbit_r44_c49 bl_49 br_49 wl_44 vdd gnd cell_6t
Xbit_r45_c49 bl_49 br_49 wl_45 vdd gnd cell_6t
Xbit_r46_c49 bl_49 br_49 wl_46 vdd gnd cell_6t
Xbit_r47_c49 bl_49 br_49 wl_47 vdd gnd cell_6t
Xbit_r48_c49 bl_49 br_49 wl_48 vdd gnd cell_6t
Xbit_r49_c49 bl_49 br_49 wl_49 vdd gnd cell_6t
Xbit_r50_c49 bl_49 br_49 wl_50 vdd gnd cell_6t
Xbit_r51_c49 bl_49 br_49 wl_51 vdd gnd cell_6t
Xbit_r52_c49 bl_49 br_49 wl_52 vdd gnd cell_6t
Xbit_r53_c49 bl_49 br_49 wl_53 vdd gnd cell_6t
Xbit_r54_c49 bl_49 br_49 wl_54 vdd gnd cell_6t
Xbit_r55_c49 bl_49 br_49 wl_55 vdd gnd cell_6t
Xbit_r56_c49 bl_49 br_49 wl_56 vdd gnd cell_6t
Xbit_r57_c49 bl_49 br_49 wl_57 vdd gnd cell_6t
Xbit_r58_c49 bl_49 br_49 wl_58 vdd gnd cell_6t
Xbit_r59_c49 bl_49 br_49 wl_59 vdd gnd cell_6t
Xbit_r60_c49 bl_49 br_49 wl_60 vdd gnd cell_6t
Xbit_r61_c49 bl_49 br_49 wl_61 vdd gnd cell_6t
Xbit_r62_c49 bl_49 br_49 wl_62 vdd gnd cell_6t
Xbit_r63_c49 bl_49 br_49 wl_63 vdd gnd cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd cell_6t
Xbit_r1_c50 bl_50 br_50 wl_1 vdd gnd cell_6t
Xbit_r2_c50 bl_50 br_50 wl_2 vdd gnd cell_6t
Xbit_r3_c50 bl_50 br_50 wl_3 vdd gnd cell_6t
Xbit_r4_c50 bl_50 br_50 wl_4 vdd gnd cell_6t
Xbit_r5_c50 bl_50 br_50 wl_5 vdd gnd cell_6t
Xbit_r6_c50 bl_50 br_50 wl_6 vdd gnd cell_6t
Xbit_r7_c50 bl_50 br_50 wl_7 vdd gnd cell_6t
Xbit_r8_c50 bl_50 br_50 wl_8 vdd gnd cell_6t
Xbit_r9_c50 bl_50 br_50 wl_9 vdd gnd cell_6t
Xbit_r10_c50 bl_50 br_50 wl_10 vdd gnd cell_6t
Xbit_r11_c50 bl_50 br_50 wl_11 vdd gnd cell_6t
Xbit_r12_c50 bl_50 br_50 wl_12 vdd gnd cell_6t
Xbit_r13_c50 bl_50 br_50 wl_13 vdd gnd cell_6t
Xbit_r14_c50 bl_50 br_50 wl_14 vdd gnd cell_6t
Xbit_r15_c50 bl_50 br_50 wl_15 vdd gnd cell_6t
Xbit_r16_c50 bl_50 br_50 wl_16 vdd gnd cell_6t
Xbit_r17_c50 bl_50 br_50 wl_17 vdd gnd cell_6t
Xbit_r18_c50 bl_50 br_50 wl_18 vdd gnd cell_6t
Xbit_r19_c50 bl_50 br_50 wl_19 vdd gnd cell_6t
Xbit_r20_c50 bl_50 br_50 wl_20 vdd gnd cell_6t
Xbit_r21_c50 bl_50 br_50 wl_21 vdd gnd cell_6t
Xbit_r22_c50 bl_50 br_50 wl_22 vdd gnd cell_6t
Xbit_r23_c50 bl_50 br_50 wl_23 vdd gnd cell_6t
Xbit_r24_c50 bl_50 br_50 wl_24 vdd gnd cell_6t
Xbit_r25_c50 bl_50 br_50 wl_25 vdd gnd cell_6t
Xbit_r26_c50 bl_50 br_50 wl_26 vdd gnd cell_6t
Xbit_r27_c50 bl_50 br_50 wl_27 vdd gnd cell_6t
Xbit_r28_c50 bl_50 br_50 wl_28 vdd gnd cell_6t
Xbit_r29_c50 bl_50 br_50 wl_29 vdd gnd cell_6t
Xbit_r30_c50 bl_50 br_50 wl_30 vdd gnd cell_6t
Xbit_r31_c50 bl_50 br_50 wl_31 vdd gnd cell_6t
Xbit_r32_c50 bl_50 br_50 wl_32 vdd gnd cell_6t
Xbit_r33_c50 bl_50 br_50 wl_33 vdd gnd cell_6t
Xbit_r34_c50 bl_50 br_50 wl_34 vdd gnd cell_6t
Xbit_r35_c50 bl_50 br_50 wl_35 vdd gnd cell_6t
Xbit_r36_c50 bl_50 br_50 wl_36 vdd gnd cell_6t
Xbit_r37_c50 bl_50 br_50 wl_37 vdd gnd cell_6t
Xbit_r38_c50 bl_50 br_50 wl_38 vdd gnd cell_6t
Xbit_r39_c50 bl_50 br_50 wl_39 vdd gnd cell_6t
Xbit_r40_c50 bl_50 br_50 wl_40 vdd gnd cell_6t
Xbit_r41_c50 bl_50 br_50 wl_41 vdd gnd cell_6t
Xbit_r42_c50 bl_50 br_50 wl_42 vdd gnd cell_6t
Xbit_r43_c50 bl_50 br_50 wl_43 vdd gnd cell_6t
Xbit_r44_c50 bl_50 br_50 wl_44 vdd gnd cell_6t
Xbit_r45_c50 bl_50 br_50 wl_45 vdd gnd cell_6t
Xbit_r46_c50 bl_50 br_50 wl_46 vdd gnd cell_6t
Xbit_r47_c50 bl_50 br_50 wl_47 vdd gnd cell_6t
Xbit_r48_c50 bl_50 br_50 wl_48 vdd gnd cell_6t
Xbit_r49_c50 bl_50 br_50 wl_49 vdd gnd cell_6t
Xbit_r50_c50 bl_50 br_50 wl_50 vdd gnd cell_6t
Xbit_r51_c50 bl_50 br_50 wl_51 vdd gnd cell_6t
Xbit_r52_c50 bl_50 br_50 wl_52 vdd gnd cell_6t
Xbit_r53_c50 bl_50 br_50 wl_53 vdd gnd cell_6t
Xbit_r54_c50 bl_50 br_50 wl_54 vdd gnd cell_6t
Xbit_r55_c50 bl_50 br_50 wl_55 vdd gnd cell_6t
Xbit_r56_c50 bl_50 br_50 wl_56 vdd gnd cell_6t
Xbit_r57_c50 bl_50 br_50 wl_57 vdd gnd cell_6t
Xbit_r58_c50 bl_50 br_50 wl_58 vdd gnd cell_6t
Xbit_r59_c50 bl_50 br_50 wl_59 vdd gnd cell_6t
Xbit_r60_c50 bl_50 br_50 wl_60 vdd gnd cell_6t
Xbit_r61_c50 bl_50 br_50 wl_61 vdd gnd cell_6t
Xbit_r62_c50 bl_50 br_50 wl_62 vdd gnd cell_6t
Xbit_r63_c50 bl_50 br_50 wl_63 vdd gnd cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd cell_6t
Xbit_r1_c51 bl_51 br_51 wl_1 vdd gnd cell_6t
Xbit_r2_c51 bl_51 br_51 wl_2 vdd gnd cell_6t
Xbit_r3_c51 bl_51 br_51 wl_3 vdd gnd cell_6t
Xbit_r4_c51 bl_51 br_51 wl_4 vdd gnd cell_6t
Xbit_r5_c51 bl_51 br_51 wl_5 vdd gnd cell_6t
Xbit_r6_c51 bl_51 br_51 wl_6 vdd gnd cell_6t
Xbit_r7_c51 bl_51 br_51 wl_7 vdd gnd cell_6t
Xbit_r8_c51 bl_51 br_51 wl_8 vdd gnd cell_6t
Xbit_r9_c51 bl_51 br_51 wl_9 vdd gnd cell_6t
Xbit_r10_c51 bl_51 br_51 wl_10 vdd gnd cell_6t
Xbit_r11_c51 bl_51 br_51 wl_11 vdd gnd cell_6t
Xbit_r12_c51 bl_51 br_51 wl_12 vdd gnd cell_6t
Xbit_r13_c51 bl_51 br_51 wl_13 vdd gnd cell_6t
Xbit_r14_c51 bl_51 br_51 wl_14 vdd gnd cell_6t
Xbit_r15_c51 bl_51 br_51 wl_15 vdd gnd cell_6t
Xbit_r16_c51 bl_51 br_51 wl_16 vdd gnd cell_6t
Xbit_r17_c51 bl_51 br_51 wl_17 vdd gnd cell_6t
Xbit_r18_c51 bl_51 br_51 wl_18 vdd gnd cell_6t
Xbit_r19_c51 bl_51 br_51 wl_19 vdd gnd cell_6t
Xbit_r20_c51 bl_51 br_51 wl_20 vdd gnd cell_6t
Xbit_r21_c51 bl_51 br_51 wl_21 vdd gnd cell_6t
Xbit_r22_c51 bl_51 br_51 wl_22 vdd gnd cell_6t
Xbit_r23_c51 bl_51 br_51 wl_23 vdd gnd cell_6t
Xbit_r24_c51 bl_51 br_51 wl_24 vdd gnd cell_6t
Xbit_r25_c51 bl_51 br_51 wl_25 vdd gnd cell_6t
Xbit_r26_c51 bl_51 br_51 wl_26 vdd gnd cell_6t
Xbit_r27_c51 bl_51 br_51 wl_27 vdd gnd cell_6t
Xbit_r28_c51 bl_51 br_51 wl_28 vdd gnd cell_6t
Xbit_r29_c51 bl_51 br_51 wl_29 vdd gnd cell_6t
Xbit_r30_c51 bl_51 br_51 wl_30 vdd gnd cell_6t
Xbit_r31_c51 bl_51 br_51 wl_31 vdd gnd cell_6t
Xbit_r32_c51 bl_51 br_51 wl_32 vdd gnd cell_6t
Xbit_r33_c51 bl_51 br_51 wl_33 vdd gnd cell_6t
Xbit_r34_c51 bl_51 br_51 wl_34 vdd gnd cell_6t
Xbit_r35_c51 bl_51 br_51 wl_35 vdd gnd cell_6t
Xbit_r36_c51 bl_51 br_51 wl_36 vdd gnd cell_6t
Xbit_r37_c51 bl_51 br_51 wl_37 vdd gnd cell_6t
Xbit_r38_c51 bl_51 br_51 wl_38 vdd gnd cell_6t
Xbit_r39_c51 bl_51 br_51 wl_39 vdd gnd cell_6t
Xbit_r40_c51 bl_51 br_51 wl_40 vdd gnd cell_6t
Xbit_r41_c51 bl_51 br_51 wl_41 vdd gnd cell_6t
Xbit_r42_c51 bl_51 br_51 wl_42 vdd gnd cell_6t
Xbit_r43_c51 bl_51 br_51 wl_43 vdd gnd cell_6t
Xbit_r44_c51 bl_51 br_51 wl_44 vdd gnd cell_6t
Xbit_r45_c51 bl_51 br_51 wl_45 vdd gnd cell_6t
Xbit_r46_c51 bl_51 br_51 wl_46 vdd gnd cell_6t
Xbit_r47_c51 bl_51 br_51 wl_47 vdd gnd cell_6t
Xbit_r48_c51 bl_51 br_51 wl_48 vdd gnd cell_6t
Xbit_r49_c51 bl_51 br_51 wl_49 vdd gnd cell_6t
Xbit_r50_c51 bl_51 br_51 wl_50 vdd gnd cell_6t
Xbit_r51_c51 bl_51 br_51 wl_51 vdd gnd cell_6t
Xbit_r52_c51 bl_51 br_51 wl_52 vdd gnd cell_6t
Xbit_r53_c51 bl_51 br_51 wl_53 vdd gnd cell_6t
Xbit_r54_c51 bl_51 br_51 wl_54 vdd gnd cell_6t
Xbit_r55_c51 bl_51 br_51 wl_55 vdd gnd cell_6t
Xbit_r56_c51 bl_51 br_51 wl_56 vdd gnd cell_6t
Xbit_r57_c51 bl_51 br_51 wl_57 vdd gnd cell_6t
Xbit_r58_c51 bl_51 br_51 wl_58 vdd gnd cell_6t
Xbit_r59_c51 bl_51 br_51 wl_59 vdd gnd cell_6t
Xbit_r60_c51 bl_51 br_51 wl_60 vdd gnd cell_6t
Xbit_r61_c51 bl_51 br_51 wl_61 vdd gnd cell_6t
Xbit_r62_c51 bl_51 br_51 wl_62 vdd gnd cell_6t
Xbit_r63_c51 bl_51 br_51 wl_63 vdd gnd cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd cell_6t
Xbit_r1_c52 bl_52 br_52 wl_1 vdd gnd cell_6t
Xbit_r2_c52 bl_52 br_52 wl_2 vdd gnd cell_6t
Xbit_r3_c52 bl_52 br_52 wl_3 vdd gnd cell_6t
Xbit_r4_c52 bl_52 br_52 wl_4 vdd gnd cell_6t
Xbit_r5_c52 bl_52 br_52 wl_5 vdd gnd cell_6t
Xbit_r6_c52 bl_52 br_52 wl_6 vdd gnd cell_6t
Xbit_r7_c52 bl_52 br_52 wl_7 vdd gnd cell_6t
Xbit_r8_c52 bl_52 br_52 wl_8 vdd gnd cell_6t
Xbit_r9_c52 bl_52 br_52 wl_9 vdd gnd cell_6t
Xbit_r10_c52 bl_52 br_52 wl_10 vdd gnd cell_6t
Xbit_r11_c52 bl_52 br_52 wl_11 vdd gnd cell_6t
Xbit_r12_c52 bl_52 br_52 wl_12 vdd gnd cell_6t
Xbit_r13_c52 bl_52 br_52 wl_13 vdd gnd cell_6t
Xbit_r14_c52 bl_52 br_52 wl_14 vdd gnd cell_6t
Xbit_r15_c52 bl_52 br_52 wl_15 vdd gnd cell_6t
Xbit_r16_c52 bl_52 br_52 wl_16 vdd gnd cell_6t
Xbit_r17_c52 bl_52 br_52 wl_17 vdd gnd cell_6t
Xbit_r18_c52 bl_52 br_52 wl_18 vdd gnd cell_6t
Xbit_r19_c52 bl_52 br_52 wl_19 vdd gnd cell_6t
Xbit_r20_c52 bl_52 br_52 wl_20 vdd gnd cell_6t
Xbit_r21_c52 bl_52 br_52 wl_21 vdd gnd cell_6t
Xbit_r22_c52 bl_52 br_52 wl_22 vdd gnd cell_6t
Xbit_r23_c52 bl_52 br_52 wl_23 vdd gnd cell_6t
Xbit_r24_c52 bl_52 br_52 wl_24 vdd gnd cell_6t
Xbit_r25_c52 bl_52 br_52 wl_25 vdd gnd cell_6t
Xbit_r26_c52 bl_52 br_52 wl_26 vdd gnd cell_6t
Xbit_r27_c52 bl_52 br_52 wl_27 vdd gnd cell_6t
Xbit_r28_c52 bl_52 br_52 wl_28 vdd gnd cell_6t
Xbit_r29_c52 bl_52 br_52 wl_29 vdd gnd cell_6t
Xbit_r30_c52 bl_52 br_52 wl_30 vdd gnd cell_6t
Xbit_r31_c52 bl_52 br_52 wl_31 vdd gnd cell_6t
Xbit_r32_c52 bl_52 br_52 wl_32 vdd gnd cell_6t
Xbit_r33_c52 bl_52 br_52 wl_33 vdd gnd cell_6t
Xbit_r34_c52 bl_52 br_52 wl_34 vdd gnd cell_6t
Xbit_r35_c52 bl_52 br_52 wl_35 vdd gnd cell_6t
Xbit_r36_c52 bl_52 br_52 wl_36 vdd gnd cell_6t
Xbit_r37_c52 bl_52 br_52 wl_37 vdd gnd cell_6t
Xbit_r38_c52 bl_52 br_52 wl_38 vdd gnd cell_6t
Xbit_r39_c52 bl_52 br_52 wl_39 vdd gnd cell_6t
Xbit_r40_c52 bl_52 br_52 wl_40 vdd gnd cell_6t
Xbit_r41_c52 bl_52 br_52 wl_41 vdd gnd cell_6t
Xbit_r42_c52 bl_52 br_52 wl_42 vdd gnd cell_6t
Xbit_r43_c52 bl_52 br_52 wl_43 vdd gnd cell_6t
Xbit_r44_c52 bl_52 br_52 wl_44 vdd gnd cell_6t
Xbit_r45_c52 bl_52 br_52 wl_45 vdd gnd cell_6t
Xbit_r46_c52 bl_52 br_52 wl_46 vdd gnd cell_6t
Xbit_r47_c52 bl_52 br_52 wl_47 vdd gnd cell_6t
Xbit_r48_c52 bl_52 br_52 wl_48 vdd gnd cell_6t
Xbit_r49_c52 bl_52 br_52 wl_49 vdd gnd cell_6t
Xbit_r50_c52 bl_52 br_52 wl_50 vdd gnd cell_6t
Xbit_r51_c52 bl_52 br_52 wl_51 vdd gnd cell_6t
Xbit_r52_c52 bl_52 br_52 wl_52 vdd gnd cell_6t
Xbit_r53_c52 bl_52 br_52 wl_53 vdd gnd cell_6t
Xbit_r54_c52 bl_52 br_52 wl_54 vdd gnd cell_6t
Xbit_r55_c52 bl_52 br_52 wl_55 vdd gnd cell_6t
Xbit_r56_c52 bl_52 br_52 wl_56 vdd gnd cell_6t
Xbit_r57_c52 bl_52 br_52 wl_57 vdd gnd cell_6t
Xbit_r58_c52 bl_52 br_52 wl_58 vdd gnd cell_6t
Xbit_r59_c52 bl_52 br_52 wl_59 vdd gnd cell_6t
Xbit_r60_c52 bl_52 br_52 wl_60 vdd gnd cell_6t
Xbit_r61_c52 bl_52 br_52 wl_61 vdd gnd cell_6t
Xbit_r62_c52 bl_52 br_52 wl_62 vdd gnd cell_6t
Xbit_r63_c52 bl_52 br_52 wl_63 vdd gnd cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd cell_6t
Xbit_r1_c53 bl_53 br_53 wl_1 vdd gnd cell_6t
Xbit_r2_c53 bl_53 br_53 wl_2 vdd gnd cell_6t
Xbit_r3_c53 bl_53 br_53 wl_3 vdd gnd cell_6t
Xbit_r4_c53 bl_53 br_53 wl_4 vdd gnd cell_6t
Xbit_r5_c53 bl_53 br_53 wl_5 vdd gnd cell_6t
Xbit_r6_c53 bl_53 br_53 wl_6 vdd gnd cell_6t
Xbit_r7_c53 bl_53 br_53 wl_7 vdd gnd cell_6t
Xbit_r8_c53 bl_53 br_53 wl_8 vdd gnd cell_6t
Xbit_r9_c53 bl_53 br_53 wl_9 vdd gnd cell_6t
Xbit_r10_c53 bl_53 br_53 wl_10 vdd gnd cell_6t
Xbit_r11_c53 bl_53 br_53 wl_11 vdd gnd cell_6t
Xbit_r12_c53 bl_53 br_53 wl_12 vdd gnd cell_6t
Xbit_r13_c53 bl_53 br_53 wl_13 vdd gnd cell_6t
Xbit_r14_c53 bl_53 br_53 wl_14 vdd gnd cell_6t
Xbit_r15_c53 bl_53 br_53 wl_15 vdd gnd cell_6t
Xbit_r16_c53 bl_53 br_53 wl_16 vdd gnd cell_6t
Xbit_r17_c53 bl_53 br_53 wl_17 vdd gnd cell_6t
Xbit_r18_c53 bl_53 br_53 wl_18 vdd gnd cell_6t
Xbit_r19_c53 bl_53 br_53 wl_19 vdd gnd cell_6t
Xbit_r20_c53 bl_53 br_53 wl_20 vdd gnd cell_6t
Xbit_r21_c53 bl_53 br_53 wl_21 vdd gnd cell_6t
Xbit_r22_c53 bl_53 br_53 wl_22 vdd gnd cell_6t
Xbit_r23_c53 bl_53 br_53 wl_23 vdd gnd cell_6t
Xbit_r24_c53 bl_53 br_53 wl_24 vdd gnd cell_6t
Xbit_r25_c53 bl_53 br_53 wl_25 vdd gnd cell_6t
Xbit_r26_c53 bl_53 br_53 wl_26 vdd gnd cell_6t
Xbit_r27_c53 bl_53 br_53 wl_27 vdd gnd cell_6t
Xbit_r28_c53 bl_53 br_53 wl_28 vdd gnd cell_6t
Xbit_r29_c53 bl_53 br_53 wl_29 vdd gnd cell_6t
Xbit_r30_c53 bl_53 br_53 wl_30 vdd gnd cell_6t
Xbit_r31_c53 bl_53 br_53 wl_31 vdd gnd cell_6t
Xbit_r32_c53 bl_53 br_53 wl_32 vdd gnd cell_6t
Xbit_r33_c53 bl_53 br_53 wl_33 vdd gnd cell_6t
Xbit_r34_c53 bl_53 br_53 wl_34 vdd gnd cell_6t
Xbit_r35_c53 bl_53 br_53 wl_35 vdd gnd cell_6t
Xbit_r36_c53 bl_53 br_53 wl_36 vdd gnd cell_6t
Xbit_r37_c53 bl_53 br_53 wl_37 vdd gnd cell_6t
Xbit_r38_c53 bl_53 br_53 wl_38 vdd gnd cell_6t
Xbit_r39_c53 bl_53 br_53 wl_39 vdd gnd cell_6t
Xbit_r40_c53 bl_53 br_53 wl_40 vdd gnd cell_6t
Xbit_r41_c53 bl_53 br_53 wl_41 vdd gnd cell_6t
Xbit_r42_c53 bl_53 br_53 wl_42 vdd gnd cell_6t
Xbit_r43_c53 bl_53 br_53 wl_43 vdd gnd cell_6t
Xbit_r44_c53 bl_53 br_53 wl_44 vdd gnd cell_6t
Xbit_r45_c53 bl_53 br_53 wl_45 vdd gnd cell_6t
Xbit_r46_c53 bl_53 br_53 wl_46 vdd gnd cell_6t
Xbit_r47_c53 bl_53 br_53 wl_47 vdd gnd cell_6t
Xbit_r48_c53 bl_53 br_53 wl_48 vdd gnd cell_6t
Xbit_r49_c53 bl_53 br_53 wl_49 vdd gnd cell_6t
Xbit_r50_c53 bl_53 br_53 wl_50 vdd gnd cell_6t
Xbit_r51_c53 bl_53 br_53 wl_51 vdd gnd cell_6t
Xbit_r52_c53 bl_53 br_53 wl_52 vdd gnd cell_6t
Xbit_r53_c53 bl_53 br_53 wl_53 vdd gnd cell_6t
Xbit_r54_c53 bl_53 br_53 wl_54 vdd gnd cell_6t
Xbit_r55_c53 bl_53 br_53 wl_55 vdd gnd cell_6t
Xbit_r56_c53 bl_53 br_53 wl_56 vdd gnd cell_6t
Xbit_r57_c53 bl_53 br_53 wl_57 vdd gnd cell_6t
Xbit_r58_c53 bl_53 br_53 wl_58 vdd gnd cell_6t
Xbit_r59_c53 bl_53 br_53 wl_59 vdd gnd cell_6t
Xbit_r60_c53 bl_53 br_53 wl_60 vdd gnd cell_6t
Xbit_r61_c53 bl_53 br_53 wl_61 vdd gnd cell_6t
Xbit_r62_c53 bl_53 br_53 wl_62 vdd gnd cell_6t
Xbit_r63_c53 bl_53 br_53 wl_63 vdd gnd cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd cell_6t
Xbit_r1_c54 bl_54 br_54 wl_1 vdd gnd cell_6t
Xbit_r2_c54 bl_54 br_54 wl_2 vdd gnd cell_6t
Xbit_r3_c54 bl_54 br_54 wl_3 vdd gnd cell_6t
Xbit_r4_c54 bl_54 br_54 wl_4 vdd gnd cell_6t
Xbit_r5_c54 bl_54 br_54 wl_5 vdd gnd cell_6t
Xbit_r6_c54 bl_54 br_54 wl_6 vdd gnd cell_6t
Xbit_r7_c54 bl_54 br_54 wl_7 vdd gnd cell_6t
Xbit_r8_c54 bl_54 br_54 wl_8 vdd gnd cell_6t
Xbit_r9_c54 bl_54 br_54 wl_9 vdd gnd cell_6t
Xbit_r10_c54 bl_54 br_54 wl_10 vdd gnd cell_6t
Xbit_r11_c54 bl_54 br_54 wl_11 vdd gnd cell_6t
Xbit_r12_c54 bl_54 br_54 wl_12 vdd gnd cell_6t
Xbit_r13_c54 bl_54 br_54 wl_13 vdd gnd cell_6t
Xbit_r14_c54 bl_54 br_54 wl_14 vdd gnd cell_6t
Xbit_r15_c54 bl_54 br_54 wl_15 vdd gnd cell_6t
Xbit_r16_c54 bl_54 br_54 wl_16 vdd gnd cell_6t
Xbit_r17_c54 bl_54 br_54 wl_17 vdd gnd cell_6t
Xbit_r18_c54 bl_54 br_54 wl_18 vdd gnd cell_6t
Xbit_r19_c54 bl_54 br_54 wl_19 vdd gnd cell_6t
Xbit_r20_c54 bl_54 br_54 wl_20 vdd gnd cell_6t
Xbit_r21_c54 bl_54 br_54 wl_21 vdd gnd cell_6t
Xbit_r22_c54 bl_54 br_54 wl_22 vdd gnd cell_6t
Xbit_r23_c54 bl_54 br_54 wl_23 vdd gnd cell_6t
Xbit_r24_c54 bl_54 br_54 wl_24 vdd gnd cell_6t
Xbit_r25_c54 bl_54 br_54 wl_25 vdd gnd cell_6t
Xbit_r26_c54 bl_54 br_54 wl_26 vdd gnd cell_6t
Xbit_r27_c54 bl_54 br_54 wl_27 vdd gnd cell_6t
Xbit_r28_c54 bl_54 br_54 wl_28 vdd gnd cell_6t
Xbit_r29_c54 bl_54 br_54 wl_29 vdd gnd cell_6t
Xbit_r30_c54 bl_54 br_54 wl_30 vdd gnd cell_6t
Xbit_r31_c54 bl_54 br_54 wl_31 vdd gnd cell_6t
Xbit_r32_c54 bl_54 br_54 wl_32 vdd gnd cell_6t
Xbit_r33_c54 bl_54 br_54 wl_33 vdd gnd cell_6t
Xbit_r34_c54 bl_54 br_54 wl_34 vdd gnd cell_6t
Xbit_r35_c54 bl_54 br_54 wl_35 vdd gnd cell_6t
Xbit_r36_c54 bl_54 br_54 wl_36 vdd gnd cell_6t
Xbit_r37_c54 bl_54 br_54 wl_37 vdd gnd cell_6t
Xbit_r38_c54 bl_54 br_54 wl_38 vdd gnd cell_6t
Xbit_r39_c54 bl_54 br_54 wl_39 vdd gnd cell_6t
Xbit_r40_c54 bl_54 br_54 wl_40 vdd gnd cell_6t
Xbit_r41_c54 bl_54 br_54 wl_41 vdd gnd cell_6t
Xbit_r42_c54 bl_54 br_54 wl_42 vdd gnd cell_6t
Xbit_r43_c54 bl_54 br_54 wl_43 vdd gnd cell_6t
Xbit_r44_c54 bl_54 br_54 wl_44 vdd gnd cell_6t
Xbit_r45_c54 bl_54 br_54 wl_45 vdd gnd cell_6t
Xbit_r46_c54 bl_54 br_54 wl_46 vdd gnd cell_6t
Xbit_r47_c54 bl_54 br_54 wl_47 vdd gnd cell_6t
Xbit_r48_c54 bl_54 br_54 wl_48 vdd gnd cell_6t
Xbit_r49_c54 bl_54 br_54 wl_49 vdd gnd cell_6t
Xbit_r50_c54 bl_54 br_54 wl_50 vdd gnd cell_6t
Xbit_r51_c54 bl_54 br_54 wl_51 vdd gnd cell_6t
Xbit_r52_c54 bl_54 br_54 wl_52 vdd gnd cell_6t
Xbit_r53_c54 bl_54 br_54 wl_53 vdd gnd cell_6t
Xbit_r54_c54 bl_54 br_54 wl_54 vdd gnd cell_6t
Xbit_r55_c54 bl_54 br_54 wl_55 vdd gnd cell_6t
Xbit_r56_c54 bl_54 br_54 wl_56 vdd gnd cell_6t
Xbit_r57_c54 bl_54 br_54 wl_57 vdd gnd cell_6t
Xbit_r58_c54 bl_54 br_54 wl_58 vdd gnd cell_6t
Xbit_r59_c54 bl_54 br_54 wl_59 vdd gnd cell_6t
Xbit_r60_c54 bl_54 br_54 wl_60 vdd gnd cell_6t
Xbit_r61_c54 bl_54 br_54 wl_61 vdd gnd cell_6t
Xbit_r62_c54 bl_54 br_54 wl_62 vdd gnd cell_6t
Xbit_r63_c54 bl_54 br_54 wl_63 vdd gnd cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd cell_6t
Xbit_r1_c55 bl_55 br_55 wl_1 vdd gnd cell_6t
Xbit_r2_c55 bl_55 br_55 wl_2 vdd gnd cell_6t
Xbit_r3_c55 bl_55 br_55 wl_3 vdd gnd cell_6t
Xbit_r4_c55 bl_55 br_55 wl_4 vdd gnd cell_6t
Xbit_r5_c55 bl_55 br_55 wl_5 vdd gnd cell_6t
Xbit_r6_c55 bl_55 br_55 wl_6 vdd gnd cell_6t
Xbit_r7_c55 bl_55 br_55 wl_7 vdd gnd cell_6t
Xbit_r8_c55 bl_55 br_55 wl_8 vdd gnd cell_6t
Xbit_r9_c55 bl_55 br_55 wl_9 vdd gnd cell_6t
Xbit_r10_c55 bl_55 br_55 wl_10 vdd gnd cell_6t
Xbit_r11_c55 bl_55 br_55 wl_11 vdd gnd cell_6t
Xbit_r12_c55 bl_55 br_55 wl_12 vdd gnd cell_6t
Xbit_r13_c55 bl_55 br_55 wl_13 vdd gnd cell_6t
Xbit_r14_c55 bl_55 br_55 wl_14 vdd gnd cell_6t
Xbit_r15_c55 bl_55 br_55 wl_15 vdd gnd cell_6t
Xbit_r16_c55 bl_55 br_55 wl_16 vdd gnd cell_6t
Xbit_r17_c55 bl_55 br_55 wl_17 vdd gnd cell_6t
Xbit_r18_c55 bl_55 br_55 wl_18 vdd gnd cell_6t
Xbit_r19_c55 bl_55 br_55 wl_19 vdd gnd cell_6t
Xbit_r20_c55 bl_55 br_55 wl_20 vdd gnd cell_6t
Xbit_r21_c55 bl_55 br_55 wl_21 vdd gnd cell_6t
Xbit_r22_c55 bl_55 br_55 wl_22 vdd gnd cell_6t
Xbit_r23_c55 bl_55 br_55 wl_23 vdd gnd cell_6t
Xbit_r24_c55 bl_55 br_55 wl_24 vdd gnd cell_6t
Xbit_r25_c55 bl_55 br_55 wl_25 vdd gnd cell_6t
Xbit_r26_c55 bl_55 br_55 wl_26 vdd gnd cell_6t
Xbit_r27_c55 bl_55 br_55 wl_27 vdd gnd cell_6t
Xbit_r28_c55 bl_55 br_55 wl_28 vdd gnd cell_6t
Xbit_r29_c55 bl_55 br_55 wl_29 vdd gnd cell_6t
Xbit_r30_c55 bl_55 br_55 wl_30 vdd gnd cell_6t
Xbit_r31_c55 bl_55 br_55 wl_31 vdd gnd cell_6t
Xbit_r32_c55 bl_55 br_55 wl_32 vdd gnd cell_6t
Xbit_r33_c55 bl_55 br_55 wl_33 vdd gnd cell_6t
Xbit_r34_c55 bl_55 br_55 wl_34 vdd gnd cell_6t
Xbit_r35_c55 bl_55 br_55 wl_35 vdd gnd cell_6t
Xbit_r36_c55 bl_55 br_55 wl_36 vdd gnd cell_6t
Xbit_r37_c55 bl_55 br_55 wl_37 vdd gnd cell_6t
Xbit_r38_c55 bl_55 br_55 wl_38 vdd gnd cell_6t
Xbit_r39_c55 bl_55 br_55 wl_39 vdd gnd cell_6t
Xbit_r40_c55 bl_55 br_55 wl_40 vdd gnd cell_6t
Xbit_r41_c55 bl_55 br_55 wl_41 vdd gnd cell_6t
Xbit_r42_c55 bl_55 br_55 wl_42 vdd gnd cell_6t
Xbit_r43_c55 bl_55 br_55 wl_43 vdd gnd cell_6t
Xbit_r44_c55 bl_55 br_55 wl_44 vdd gnd cell_6t
Xbit_r45_c55 bl_55 br_55 wl_45 vdd gnd cell_6t
Xbit_r46_c55 bl_55 br_55 wl_46 vdd gnd cell_6t
Xbit_r47_c55 bl_55 br_55 wl_47 vdd gnd cell_6t
Xbit_r48_c55 bl_55 br_55 wl_48 vdd gnd cell_6t
Xbit_r49_c55 bl_55 br_55 wl_49 vdd gnd cell_6t
Xbit_r50_c55 bl_55 br_55 wl_50 vdd gnd cell_6t
Xbit_r51_c55 bl_55 br_55 wl_51 vdd gnd cell_6t
Xbit_r52_c55 bl_55 br_55 wl_52 vdd gnd cell_6t
Xbit_r53_c55 bl_55 br_55 wl_53 vdd gnd cell_6t
Xbit_r54_c55 bl_55 br_55 wl_54 vdd gnd cell_6t
Xbit_r55_c55 bl_55 br_55 wl_55 vdd gnd cell_6t
Xbit_r56_c55 bl_55 br_55 wl_56 vdd gnd cell_6t
Xbit_r57_c55 bl_55 br_55 wl_57 vdd gnd cell_6t
Xbit_r58_c55 bl_55 br_55 wl_58 vdd gnd cell_6t
Xbit_r59_c55 bl_55 br_55 wl_59 vdd gnd cell_6t
Xbit_r60_c55 bl_55 br_55 wl_60 vdd gnd cell_6t
Xbit_r61_c55 bl_55 br_55 wl_61 vdd gnd cell_6t
Xbit_r62_c55 bl_55 br_55 wl_62 vdd gnd cell_6t
Xbit_r63_c55 bl_55 br_55 wl_63 vdd gnd cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd cell_6t
Xbit_r1_c56 bl_56 br_56 wl_1 vdd gnd cell_6t
Xbit_r2_c56 bl_56 br_56 wl_2 vdd gnd cell_6t
Xbit_r3_c56 bl_56 br_56 wl_3 vdd gnd cell_6t
Xbit_r4_c56 bl_56 br_56 wl_4 vdd gnd cell_6t
Xbit_r5_c56 bl_56 br_56 wl_5 vdd gnd cell_6t
Xbit_r6_c56 bl_56 br_56 wl_6 vdd gnd cell_6t
Xbit_r7_c56 bl_56 br_56 wl_7 vdd gnd cell_6t
Xbit_r8_c56 bl_56 br_56 wl_8 vdd gnd cell_6t
Xbit_r9_c56 bl_56 br_56 wl_9 vdd gnd cell_6t
Xbit_r10_c56 bl_56 br_56 wl_10 vdd gnd cell_6t
Xbit_r11_c56 bl_56 br_56 wl_11 vdd gnd cell_6t
Xbit_r12_c56 bl_56 br_56 wl_12 vdd gnd cell_6t
Xbit_r13_c56 bl_56 br_56 wl_13 vdd gnd cell_6t
Xbit_r14_c56 bl_56 br_56 wl_14 vdd gnd cell_6t
Xbit_r15_c56 bl_56 br_56 wl_15 vdd gnd cell_6t
Xbit_r16_c56 bl_56 br_56 wl_16 vdd gnd cell_6t
Xbit_r17_c56 bl_56 br_56 wl_17 vdd gnd cell_6t
Xbit_r18_c56 bl_56 br_56 wl_18 vdd gnd cell_6t
Xbit_r19_c56 bl_56 br_56 wl_19 vdd gnd cell_6t
Xbit_r20_c56 bl_56 br_56 wl_20 vdd gnd cell_6t
Xbit_r21_c56 bl_56 br_56 wl_21 vdd gnd cell_6t
Xbit_r22_c56 bl_56 br_56 wl_22 vdd gnd cell_6t
Xbit_r23_c56 bl_56 br_56 wl_23 vdd gnd cell_6t
Xbit_r24_c56 bl_56 br_56 wl_24 vdd gnd cell_6t
Xbit_r25_c56 bl_56 br_56 wl_25 vdd gnd cell_6t
Xbit_r26_c56 bl_56 br_56 wl_26 vdd gnd cell_6t
Xbit_r27_c56 bl_56 br_56 wl_27 vdd gnd cell_6t
Xbit_r28_c56 bl_56 br_56 wl_28 vdd gnd cell_6t
Xbit_r29_c56 bl_56 br_56 wl_29 vdd gnd cell_6t
Xbit_r30_c56 bl_56 br_56 wl_30 vdd gnd cell_6t
Xbit_r31_c56 bl_56 br_56 wl_31 vdd gnd cell_6t
Xbit_r32_c56 bl_56 br_56 wl_32 vdd gnd cell_6t
Xbit_r33_c56 bl_56 br_56 wl_33 vdd gnd cell_6t
Xbit_r34_c56 bl_56 br_56 wl_34 vdd gnd cell_6t
Xbit_r35_c56 bl_56 br_56 wl_35 vdd gnd cell_6t
Xbit_r36_c56 bl_56 br_56 wl_36 vdd gnd cell_6t
Xbit_r37_c56 bl_56 br_56 wl_37 vdd gnd cell_6t
Xbit_r38_c56 bl_56 br_56 wl_38 vdd gnd cell_6t
Xbit_r39_c56 bl_56 br_56 wl_39 vdd gnd cell_6t
Xbit_r40_c56 bl_56 br_56 wl_40 vdd gnd cell_6t
Xbit_r41_c56 bl_56 br_56 wl_41 vdd gnd cell_6t
Xbit_r42_c56 bl_56 br_56 wl_42 vdd gnd cell_6t
Xbit_r43_c56 bl_56 br_56 wl_43 vdd gnd cell_6t
Xbit_r44_c56 bl_56 br_56 wl_44 vdd gnd cell_6t
Xbit_r45_c56 bl_56 br_56 wl_45 vdd gnd cell_6t
Xbit_r46_c56 bl_56 br_56 wl_46 vdd gnd cell_6t
Xbit_r47_c56 bl_56 br_56 wl_47 vdd gnd cell_6t
Xbit_r48_c56 bl_56 br_56 wl_48 vdd gnd cell_6t
Xbit_r49_c56 bl_56 br_56 wl_49 vdd gnd cell_6t
Xbit_r50_c56 bl_56 br_56 wl_50 vdd gnd cell_6t
Xbit_r51_c56 bl_56 br_56 wl_51 vdd gnd cell_6t
Xbit_r52_c56 bl_56 br_56 wl_52 vdd gnd cell_6t
Xbit_r53_c56 bl_56 br_56 wl_53 vdd gnd cell_6t
Xbit_r54_c56 bl_56 br_56 wl_54 vdd gnd cell_6t
Xbit_r55_c56 bl_56 br_56 wl_55 vdd gnd cell_6t
Xbit_r56_c56 bl_56 br_56 wl_56 vdd gnd cell_6t
Xbit_r57_c56 bl_56 br_56 wl_57 vdd gnd cell_6t
Xbit_r58_c56 bl_56 br_56 wl_58 vdd gnd cell_6t
Xbit_r59_c56 bl_56 br_56 wl_59 vdd gnd cell_6t
Xbit_r60_c56 bl_56 br_56 wl_60 vdd gnd cell_6t
Xbit_r61_c56 bl_56 br_56 wl_61 vdd gnd cell_6t
Xbit_r62_c56 bl_56 br_56 wl_62 vdd gnd cell_6t
Xbit_r63_c56 bl_56 br_56 wl_63 vdd gnd cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd cell_6t
Xbit_r1_c57 bl_57 br_57 wl_1 vdd gnd cell_6t
Xbit_r2_c57 bl_57 br_57 wl_2 vdd gnd cell_6t
Xbit_r3_c57 bl_57 br_57 wl_3 vdd gnd cell_6t
Xbit_r4_c57 bl_57 br_57 wl_4 vdd gnd cell_6t
Xbit_r5_c57 bl_57 br_57 wl_5 vdd gnd cell_6t
Xbit_r6_c57 bl_57 br_57 wl_6 vdd gnd cell_6t
Xbit_r7_c57 bl_57 br_57 wl_7 vdd gnd cell_6t
Xbit_r8_c57 bl_57 br_57 wl_8 vdd gnd cell_6t
Xbit_r9_c57 bl_57 br_57 wl_9 vdd gnd cell_6t
Xbit_r10_c57 bl_57 br_57 wl_10 vdd gnd cell_6t
Xbit_r11_c57 bl_57 br_57 wl_11 vdd gnd cell_6t
Xbit_r12_c57 bl_57 br_57 wl_12 vdd gnd cell_6t
Xbit_r13_c57 bl_57 br_57 wl_13 vdd gnd cell_6t
Xbit_r14_c57 bl_57 br_57 wl_14 vdd gnd cell_6t
Xbit_r15_c57 bl_57 br_57 wl_15 vdd gnd cell_6t
Xbit_r16_c57 bl_57 br_57 wl_16 vdd gnd cell_6t
Xbit_r17_c57 bl_57 br_57 wl_17 vdd gnd cell_6t
Xbit_r18_c57 bl_57 br_57 wl_18 vdd gnd cell_6t
Xbit_r19_c57 bl_57 br_57 wl_19 vdd gnd cell_6t
Xbit_r20_c57 bl_57 br_57 wl_20 vdd gnd cell_6t
Xbit_r21_c57 bl_57 br_57 wl_21 vdd gnd cell_6t
Xbit_r22_c57 bl_57 br_57 wl_22 vdd gnd cell_6t
Xbit_r23_c57 bl_57 br_57 wl_23 vdd gnd cell_6t
Xbit_r24_c57 bl_57 br_57 wl_24 vdd gnd cell_6t
Xbit_r25_c57 bl_57 br_57 wl_25 vdd gnd cell_6t
Xbit_r26_c57 bl_57 br_57 wl_26 vdd gnd cell_6t
Xbit_r27_c57 bl_57 br_57 wl_27 vdd gnd cell_6t
Xbit_r28_c57 bl_57 br_57 wl_28 vdd gnd cell_6t
Xbit_r29_c57 bl_57 br_57 wl_29 vdd gnd cell_6t
Xbit_r30_c57 bl_57 br_57 wl_30 vdd gnd cell_6t
Xbit_r31_c57 bl_57 br_57 wl_31 vdd gnd cell_6t
Xbit_r32_c57 bl_57 br_57 wl_32 vdd gnd cell_6t
Xbit_r33_c57 bl_57 br_57 wl_33 vdd gnd cell_6t
Xbit_r34_c57 bl_57 br_57 wl_34 vdd gnd cell_6t
Xbit_r35_c57 bl_57 br_57 wl_35 vdd gnd cell_6t
Xbit_r36_c57 bl_57 br_57 wl_36 vdd gnd cell_6t
Xbit_r37_c57 bl_57 br_57 wl_37 vdd gnd cell_6t
Xbit_r38_c57 bl_57 br_57 wl_38 vdd gnd cell_6t
Xbit_r39_c57 bl_57 br_57 wl_39 vdd gnd cell_6t
Xbit_r40_c57 bl_57 br_57 wl_40 vdd gnd cell_6t
Xbit_r41_c57 bl_57 br_57 wl_41 vdd gnd cell_6t
Xbit_r42_c57 bl_57 br_57 wl_42 vdd gnd cell_6t
Xbit_r43_c57 bl_57 br_57 wl_43 vdd gnd cell_6t
Xbit_r44_c57 bl_57 br_57 wl_44 vdd gnd cell_6t
Xbit_r45_c57 bl_57 br_57 wl_45 vdd gnd cell_6t
Xbit_r46_c57 bl_57 br_57 wl_46 vdd gnd cell_6t
Xbit_r47_c57 bl_57 br_57 wl_47 vdd gnd cell_6t
Xbit_r48_c57 bl_57 br_57 wl_48 vdd gnd cell_6t
Xbit_r49_c57 bl_57 br_57 wl_49 vdd gnd cell_6t
Xbit_r50_c57 bl_57 br_57 wl_50 vdd gnd cell_6t
Xbit_r51_c57 bl_57 br_57 wl_51 vdd gnd cell_6t
Xbit_r52_c57 bl_57 br_57 wl_52 vdd gnd cell_6t
Xbit_r53_c57 bl_57 br_57 wl_53 vdd gnd cell_6t
Xbit_r54_c57 bl_57 br_57 wl_54 vdd gnd cell_6t
Xbit_r55_c57 bl_57 br_57 wl_55 vdd gnd cell_6t
Xbit_r56_c57 bl_57 br_57 wl_56 vdd gnd cell_6t
Xbit_r57_c57 bl_57 br_57 wl_57 vdd gnd cell_6t
Xbit_r58_c57 bl_57 br_57 wl_58 vdd gnd cell_6t
Xbit_r59_c57 bl_57 br_57 wl_59 vdd gnd cell_6t
Xbit_r60_c57 bl_57 br_57 wl_60 vdd gnd cell_6t
Xbit_r61_c57 bl_57 br_57 wl_61 vdd gnd cell_6t
Xbit_r62_c57 bl_57 br_57 wl_62 vdd gnd cell_6t
Xbit_r63_c57 bl_57 br_57 wl_63 vdd gnd cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd cell_6t
Xbit_r1_c58 bl_58 br_58 wl_1 vdd gnd cell_6t
Xbit_r2_c58 bl_58 br_58 wl_2 vdd gnd cell_6t
Xbit_r3_c58 bl_58 br_58 wl_3 vdd gnd cell_6t
Xbit_r4_c58 bl_58 br_58 wl_4 vdd gnd cell_6t
Xbit_r5_c58 bl_58 br_58 wl_5 vdd gnd cell_6t
Xbit_r6_c58 bl_58 br_58 wl_6 vdd gnd cell_6t
Xbit_r7_c58 bl_58 br_58 wl_7 vdd gnd cell_6t
Xbit_r8_c58 bl_58 br_58 wl_8 vdd gnd cell_6t
Xbit_r9_c58 bl_58 br_58 wl_9 vdd gnd cell_6t
Xbit_r10_c58 bl_58 br_58 wl_10 vdd gnd cell_6t
Xbit_r11_c58 bl_58 br_58 wl_11 vdd gnd cell_6t
Xbit_r12_c58 bl_58 br_58 wl_12 vdd gnd cell_6t
Xbit_r13_c58 bl_58 br_58 wl_13 vdd gnd cell_6t
Xbit_r14_c58 bl_58 br_58 wl_14 vdd gnd cell_6t
Xbit_r15_c58 bl_58 br_58 wl_15 vdd gnd cell_6t
Xbit_r16_c58 bl_58 br_58 wl_16 vdd gnd cell_6t
Xbit_r17_c58 bl_58 br_58 wl_17 vdd gnd cell_6t
Xbit_r18_c58 bl_58 br_58 wl_18 vdd gnd cell_6t
Xbit_r19_c58 bl_58 br_58 wl_19 vdd gnd cell_6t
Xbit_r20_c58 bl_58 br_58 wl_20 vdd gnd cell_6t
Xbit_r21_c58 bl_58 br_58 wl_21 vdd gnd cell_6t
Xbit_r22_c58 bl_58 br_58 wl_22 vdd gnd cell_6t
Xbit_r23_c58 bl_58 br_58 wl_23 vdd gnd cell_6t
Xbit_r24_c58 bl_58 br_58 wl_24 vdd gnd cell_6t
Xbit_r25_c58 bl_58 br_58 wl_25 vdd gnd cell_6t
Xbit_r26_c58 bl_58 br_58 wl_26 vdd gnd cell_6t
Xbit_r27_c58 bl_58 br_58 wl_27 vdd gnd cell_6t
Xbit_r28_c58 bl_58 br_58 wl_28 vdd gnd cell_6t
Xbit_r29_c58 bl_58 br_58 wl_29 vdd gnd cell_6t
Xbit_r30_c58 bl_58 br_58 wl_30 vdd gnd cell_6t
Xbit_r31_c58 bl_58 br_58 wl_31 vdd gnd cell_6t
Xbit_r32_c58 bl_58 br_58 wl_32 vdd gnd cell_6t
Xbit_r33_c58 bl_58 br_58 wl_33 vdd gnd cell_6t
Xbit_r34_c58 bl_58 br_58 wl_34 vdd gnd cell_6t
Xbit_r35_c58 bl_58 br_58 wl_35 vdd gnd cell_6t
Xbit_r36_c58 bl_58 br_58 wl_36 vdd gnd cell_6t
Xbit_r37_c58 bl_58 br_58 wl_37 vdd gnd cell_6t
Xbit_r38_c58 bl_58 br_58 wl_38 vdd gnd cell_6t
Xbit_r39_c58 bl_58 br_58 wl_39 vdd gnd cell_6t
Xbit_r40_c58 bl_58 br_58 wl_40 vdd gnd cell_6t
Xbit_r41_c58 bl_58 br_58 wl_41 vdd gnd cell_6t
Xbit_r42_c58 bl_58 br_58 wl_42 vdd gnd cell_6t
Xbit_r43_c58 bl_58 br_58 wl_43 vdd gnd cell_6t
Xbit_r44_c58 bl_58 br_58 wl_44 vdd gnd cell_6t
Xbit_r45_c58 bl_58 br_58 wl_45 vdd gnd cell_6t
Xbit_r46_c58 bl_58 br_58 wl_46 vdd gnd cell_6t
Xbit_r47_c58 bl_58 br_58 wl_47 vdd gnd cell_6t
Xbit_r48_c58 bl_58 br_58 wl_48 vdd gnd cell_6t
Xbit_r49_c58 bl_58 br_58 wl_49 vdd gnd cell_6t
Xbit_r50_c58 bl_58 br_58 wl_50 vdd gnd cell_6t
Xbit_r51_c58 bl_58 br_58 wl_51 vdd gnd cell_6t
Xbit_r52_c58 bl_58 br_58 wl_52 vdd gnd cell_6t
Xbit_r53_c58 bl_58 br_58 wl_53 vdd gnd cell_6t
Xbit_r54_c58 bl_58 br_58 wl_54 vdd gnd cell_6t
Xbit_r55_c58 bl_58 br_58 wl_55 vdd gnd cell_6t
Xbit_r56_c58 bl_58 br_58 wl_56 vdd gnd cell_6t
Xbit_r57_c58 bl_58 br_58 wl_57 vdd gnd cell_6t
Xbit_r58_c58 bl_58 br_58 wl_58 vdd gnd cell_6t
Xbit_r59_c58 bl_58 br_58 wl_59 vdd gnd cell_6t
Xbit_r60_c58 bl_58 br_58 wl_60 vdd gnd cell_6t
Xbit_r61_c58 bl_58 br_58 wl_61 vdd gnd cell_6t
Xbit_r62_c58 bl_58 br_58 wl_62 vdd gnd cell_6t
Xbit_r63_c58 bl_58 br_58 wl_63 vdd gnd cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd cell_6t
Xbit_r1_c59 bl_59 br_59 wl_1 vdd gnd cell_6t
Xbit_r2_c59 bl_59 br_59 wl_2 vdd gnd cell_6t
Xbit_r3_c59 bl_59 br_59 wl_3 vdd gnd cell_6t
Xbit_r4_c59 bl_59 br_59 wl_4 vdd gnd cell_6t
Xbit_r5_c59 bl_59 br_59 wl_5 vdd gnd cell_6t
Xbit_r6_c59 bl_59 br_59 wl_6 vdd gnd cell_6t
Xbit_r7_c59 bl_59 br_59 wl_7 vdd gnd cell_6t
Xbit_r8_c59 bl_59 br_59 wl_8 vdd gnd cell_6t
Xbit_r9_c59 bl_59 br_59 wl_9 vdd gnd cell_6t
Xbit_r10_c59 bl_59 br_59 wl_10 vdd gnd cell_6t
Xbit_r11_c59 bl_59 br_59 wl_11 vdd gnd cell_6t
Xbit_r12_c59 bl_59 br_59 wl_12 vdd gnd cell_6t
Xbit_r13_c59 bl_59 br_59 wl_13 vdd gnd cell_6t
Xbit_r14_c59 bl_59 br_59 wl_14 vdd gnd cell_6t
Xbit_r15_c59 bl_59 br_59 wl_15 vdd gnd cell_6t
Xbit_r16_c59 bl_59 br_59 wl_16 vdd gnd cell_6t
Xbit_r17_c59 bl_59 br_59 wl_17 vdd gnd cell_6t
Xbit_r18_c59 bl_59 br_59 wl_18 vdd gnd cell_6t
Xbit_r19_c59 bl_59 br_59 wl_19 vdd gnd cell_6t
Xbit_r20_c59 bl_59 br_59 wl_20 vdd gnd cell_6t
Xbit_r21_c59 bl_59 br_59 wl_21 vdd gnd cell_6t
Xbit_r22_c59 bl_59 br_59 wl_22 vdd gnd cell_6t
Xbit_r23_c59 bl_59 br_59 wl_23 vdd gnd cell_6t
Xbit_r24_c59 bl_59 br_59 wl_24 vdd gnd cell_6t
Xbit_r25_c59 bl_59 br_59 wl_25 vdd gnd cell_6t
Xbit_r26_c59 bl_59 br_59 wl_26 vdd gnd cell_6t
Xbit_r27_c59 bl_59 br_59 wl_27 vdd gnd cell_6t
Xbit_r28_c59 bl_59 br_59 wl_28 vdd gnd cell_6t
Xbit_r29_c59 bl_59 br_59 wl_29 vdd gnd cell_6t
Xbit_r30_c59 bl_59 br_59 wl_30 vdd gnd cell_6t
Xbit_r31_c59 bl_59 br_59 wl_31 vdd gnd cell_6t
Xbit_r32_c59 bl_59 br_59 wl_32 vdd gnd cell_6t
Xbit_r33_c59 bl_59 br_59 wl_33 vdd gnd cell_6t
Xbit_r34_c59 bl_59 br_59 wl_34 vdd gnd cell_6t
Xbit_r35_c59 bl_59 br_59 wl_35 vdd gnd cell_6t
Xbit_r36_c59 bl_59 br_59 wl_36 vdd gnd cell_6t
Xbit_r37_c59 bl_59 br_59 wl_37 vdd gnd cell_6t
Xbit_r38_c59 bl_59 br_59 wl_38 vdd gnd cell_6t
Xbit_r39_c59 bl_59 br_59 wl_39 vdd gnd cell_6t
Xbit_r40_c59 bl_59 br_59 wl_40 vdd gnd cell_6t
Xbit_r41_c59 bl_59 br_59 wl_41 vdd gnd cell_6t
Xbit_r42_c59 bl_59 br_59 wl_42 vdd gnd cell_6t
Xbit_r43_c59 bl_59 br_59 wl_43 vdd gnd cell_6t
Xbit_r44_c59 bl_59 br_59 wl_44 vdd gnd cell_6t
Xbit_r45_c59 bl_59 br_59 wl_45 vdd gnd cell_6t
Xbit_r46_c59 bl_59 br_59 wl_46 vdd gnd cell_6t
Xbit_r47_c59 bl_59 br_59 wl_47 vdd gnd cell_6t
Xbit_r48_c59 bl_59 br_59 wl_48 vdd gnd cell_6t
Xbit_r49_c59 bl_59 br_59 wl_49 vdd gnd cell_6t
Xbit_r50_c59 bl_59 br_59 wl_50 vdd gnd cell_6t
Xbit_r51_c59 bl_59 br_59 wl_51 vdd gnd cell_6t
Xbit_r52_c59 bl_59 br_59 wl_52 vdd gnd cell_6t
Xbit_r53_c59 bl_59 br_59 wl_53 vdd gnd cell_6t
Xbit_r54_c59 bl_59 br_59 wl_54 vdd gnd cell_6t
Xbit_r55_c59 bl_59 br_59 wl_55 vdd gnd cell_6t
Xbit_r56_c59 bl_59 br_59 wl_56 vdd gnd cell_6t
Xbit_r57_c59 bl_59 br_59 wl_57 vdd gnd cell_6t
Xbit_r58_c59 bl_59 br_59 wl_58 vdd gnd cell_6t
Xbit_r59_c59 bl_59 br_59 wl_59 vdd gnd cell_6t
Xbit_r60_c59 bl_59 br_59 wl_60 vdd gnd cell_6t
Xbit_r61_c59 bl_59 br_59 wl_61 vdd gnd cell_6t
Xbit_r62_c59 bl_59 br_59 wl_62 vdd gnd cell_6t
Xbit_r63_c59 bl_59 br_59 wl_63 vdd gnd cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd cell_6t
Xbit_r1_c60 bl_60 br_60 wl_1 vdd gnd cell_6t
Xbit_r2_c60 bl_60 br_60 wl_2 vdd gnd cell_6t
Xbit_r3_c60 bl_60 br_60 wl_3 vdd gnd cell_6t
Xbit_r4_c60 bl_60 br_60 wl_4 vdd gnd cell_6t
Xbit_r5_c60 bl_60 br_60 wl_5 vdd gnd cell_6t
Xbit_r6_c60 bl_60 br_60 wl_6 vdd gnd cell_6t
Xbit_r7_c60 bl_60 br_60 wl_7 vdd gnd cell_6t
Xbit_r8_c60 bl_60 br_60 wl_8 vdd gnd cell_6t
Xbit_r9_c60 bl_60 br_60 wl_9 vdd gnd cell_6t
Xbit_r10_c60 bl_60 br_60 wl_10 vdd gnd cell_6t
Xbit_r11_c60 bl_60 br_60 wl_11 vdd gnd cell_6t
Xbit_r12_c60 bl_60 br_60 wl_12 vdd gnd cell_6t
Xbit_r13_c60 bl_60 br_60 wl_13 vdd gnd cell_6t
Xbit_r14_c60 bl_60 br_60 wl_14 vdd gnd cell_6t
Xbit_r15_c60 bl_60 br_60 wl_15 vdd gnd cell_6t
Xbit_r16_c60 bl_60 br_60 wl_16 vdd gnd cell_6t
Xbit_r17_c60 bl_60 br_60 wl_17 vdd gnd cell_6t
Xbit_r18_c60 bl_60 br_60 wl_18 vdd gnd cell_6t
Xbit_r19_c60 bl_60 br_60 wl_19 vdd gnd cell_6t
Xbit_r20_c60 bl_60 br_60 wl_20 vdd gnd cell_6t
Xbit_r21_c60 bl_60 br_60 wl_21 vdd gnd cell_6t
Xbit_r22_c60 bl_60 br_60 wl_22 vdd gnd cell_6t
Xbit_r23_c60 bl_60 br_60 wl_23 vdd gnd cell_6t
Xbit_r24_c60 bl_60 br_60 wl_24 vdd gnd cell_6t
Xbit_r25_c60 bl_60 br_60 wl_25 vdd gnd cell_6t
Xbit_r26_c60 bl_60 br_60 wl_26 vdd gnd cell_6t
Xbit_r27_c60 bl_60 br_60 wl_27 vdd gnd cell_6t
Xbit_r28_c60 bl_60 br_60 wl_28 vdd gnd cell_6t
Xbit_r29_c60 bl_60 br_60 wl_29 vdd gnd cell_6t
Xbit_r30_c60 bl_60 br_60 wl_30 vdd gnd cell_6t
Xbit_r31_c60 bl_60 br_60 wl_31 vdd gnd cell_6t
Xbit_r32_c60 bl_60 br_60 wl_32 vdd gnd cell_6t
Xbit_r33_c60 bl_60 br_60 wl_33 vdd gnd cell_6t
Xbit_r34_c60 bl_60 br_60 wl_34 vdd gnd cell_6t
Xbit_r35_c60 bl_60 br_60 wl_35 vdd gnd cell_6t
Xbit_r36_c60 bl_60 br_60 wl_36 vdd gnd cell_6t
Xbit_r37_c60 bl_60 br_60 wl_37 vdd gnd cell_6t
Xbit_r38_c60 bl_60 br_60 wl_38 vdd gnd cell_6t
Xbit_r39_c60 bl_60 br_60 wl_39 vdd gnd cell_6t
Xbit_r40_c60 bl_60 br_60 wl_40 vdd gnd cell_6t
Xbit_r41_c60 bl_60 br_60 wl_41 vdd gnd cell_6t
Xbit_r42_c60 bl_60 br_60 wl_42 vdd gnd cell_6t
Xbit_r43_c60 bl_60 br_60 wl_43 vdd gnd cell_6t
Xbit_r44_c60 bl_60 br_60 wl_44 vdd gnd cell_6t
Xbit_r45_c60 bl_60 br_60 wl_45 vdd gnd cell_6t
Xbit_r46_c60 bl_60 br_60 wl_46 vdd gnd cell_6t
Xbit_r47_c60 bl_60 br_60 wl_47 vdd gnd cell_6t
Xbit_r48_c60 bl_60 br_60 wl_48 vdd gnd cell_6t
Xbit_r49_c60 bl_60 br_60 wl_49 vdd gnd cell_6t
Xbit_r50_c60 bl_60 br_60 wl_50 vdd gnd cell_6t
Xbit_r51_c60 bl_60 br_60 wl_51 vdd gnd cell_6t
Xbit_r52_c60 bl_60 br_60 wl_52 vdd gnd cell_6t
Xbit_r53_c60 bl_60 br_60 wl_53 vdd gnd cell_6t
Xbit_r54_c60 bl_60 br_60 wl_54 vdd gnd cell_6t
Xbit_r55_c60 bl_60 br_60 wl_55 vdd gnd cell_6t
Xbit_r56_c60 bl_60 br_60 wl_56 vdd gnd cell_6t
Xbit_r57_c60 bl_60 br_60 wl_57 vdd gnd cell_6t
Xbit_r58_c60 bl_60 br_60 wl_58 vdd gnd cell_6t
Xbit_r59_c60 bl_60 br_60 wl_59 vdd gnd cell_6t
Xbit_r60_c60 bl_60 br_60 wl_60 vdd gnd cell_6t
Xbit_r61_c60 bl_60 br_60 wl_61 vdd gnd cell_6t
Xbit_r62_c60 bl_60 br_60 wl_62 vdd gnd cell_6t
Xbit_r63_c60 bl_60 br_60 wl_63 vdd gnd cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd cell_6t
Xbit_r1_c61 bl_61 br_61 wl_1 vdd gnd cell_6t
Xbit_r2_c61 bl_61 br_61 wl_2 vdd gnd cell_6t
Xbit_r3_c61 bl_61 br_61 wl_3 vdd gnd cell_6t
Xbit_r4_c61 bl_61 br_61 wl_4 vdd gnd cell_6t
Xbit_r5_c61 bl_61 br_61 wl_5 vdd gnd cell_6t
Xbit_r6_c61 bl_61 br_61 wl_6 vdd gnd cell_6t
Xbit_r7_c61 bl_61 br_61 wl_7 vdd gnd cell_6t
Xbit_r8_c61 bl_61 br_61 wl_8 vdd gnd cell_6t
Xbit_r9_c61 bl_61 br_61 wl_9 vdd gnd cell_6t
Xbit_r10_c61 bl_61 br_61 wl_10 vdd gnd cell_6t
Xbit_r11_c61 bl_61 br_61 wl_11 vdd gnd cell_6t
Xbit_r12_c61 bl_61 br_61 wl_12 vdd gnd cell_6t
Xbit_r13_c61 bl_61 br_61 wl_13 vdd gnd cell_6t
Xbit_r14_c61 bl_61 br_61 wl_14 vdd gnd cell_6t
Xbit_r15_c61 bl_61 br_61 wl_15 vdd gnd cell_6t
Xbit_r16_c61 bl_61 br_61 wl_16 vdd gnd cell_6t
Xbit_r17_c61 bl_61 br_61 wl_17 vdd gnd cell_6t
Xbit_r18_c61 bl_61 br_61 wl_18 vdd gnd cell_6t
Xbit_r19_c61 bl_61 br_61 wl_19 vdd gnd cell_6t
Xbit_r20_c61 bl_61 br_61 wl_20 vdd gnd cell_6t
Xbit_r21_c61 bl_61 br_61 wl_21 vdd gnd cell_6t
Xbit_r22_c61 bl_61 br_61 wl_22 vdd gnd cell_6t
Xbit_r23_c61 bl_61 br_61 wl_23 vdd gnd cell_6t
Xbit_r24_c61 bl_61 br_61 wl_24 vdd gnd cell_6t
Xbit_r25_c61 bl_61 br_61 wl_25 vdd gnd cell_6t
Xbit_r26_c61 bl_61 br_61 wl_26 vdd gnd cell_6t
Xbit_r27_c61 bl_61 br_61 wl_27 vdd gnd cell_6t
Xbit_r28_c61 bl_61 br_61 wl_28 vdd gnd cell_6t
Xbit_r29_c61 bl_61 br_61 wl_29 vdd gnd cell_6t
Xbit_r30_c61 bl_61 br_61 wl_30 vdd gnd cell_6t
Xbit_r31_c61 bl_61 br_61 wl_31 vdd gnd cell_6t
Xbit_r32_c61 bl_61 br_61 wl_32 vdd gnd cell_6t
Xbit_r33_c61 bl_61 br_61 wl_33 vdd gnd cell_6t
Xbit_r34_c61 bl_61 br_61 wl_34 vdd gnd cell_6t
Xbit_r35_c61 bl_61 br_61 wl_35 vdd gnd cell_6t
Xbit_r36_c61 bl_61 br_61 wl_36 vdd gnd cell_6t
Xbit_r37_c61 bl_61 br_61 wl_37 vdd gnd cell_6t
Xbit_r38_c61 bl_61 br_61 wl_38 vdd gnd cell_6t
Xbit_r39_c61 bl_61 br_61 wl_39 vdd gnd cell_6t
Xbit_r40_c61 bl_61 br_61 wl_40 vdd gnd cell_6t
Xbit_r41_c61 bl_61 br_61 wl_41 vdd gnd cell_6t
Xbit_r42_c61 bl_61 br_61 wl_42 vdd gnd cell_6t
Xbit_r43_c61 bl_61 br_61 wl_43 vdd gnd cell_6t
Xbit_r44_c61 bl_61 br_61 wl_44 vdd gnd cell_6t
Xbit_r45_c61 bl_61 br_61 wl_45 vdd gnd cell_6t
Xbit_r46_c61 bl_61 br_61 wl_46 vdd gnd cell_6t
Xbit_r47_c61 bl_61 br_61 wl_47 vdd gnd cell_6t
Xbit_r48_c61 bl_61 br_61 wl_48 vdd gnd cell_6t
Xbit_r49_c61 bl_61 br_61 wl_49 vdd gnd cell_6t
Xbit_r50_c61 bl_61 br_61 wl_50 vdd gnd cell_6t
Xbit_r51_c61 bl_61 br_61 wl_51 vdd gnd cell_6t
Xbit_r52_c61 bl_61 br_61 wl_52 vdd gnd cell_6t
Xbit_r53_c61 bl_61 br_61 wl_53 vdd gnd cell_6t
Xbit_r54_c61 bl_61 br_61 wl_54 vdd gnd cell_6t
Xbit_r55_c61 bl_61 br_61 wl_55 vdd gnd cell_6t
Xbit_r56_c61 bl_61 br_61 wl_56 vdd gnd cell_6t
Xbit_r57_c61 bl_61 br_61 wl_57 vdd gnd cell_6t
Xbit_r58_c61 bl_61 br_61 wl_58 vdd gnd cell_6t
Xbit_r59_c61 bl_61 br_61 wl_59 vdd gnd cell_6t
Xbit_r60_c61 bl_61 br_61 wl_60 vdd gnd cell_6t
Xbit_r61_c61 bl_61 br_61 wl_61 vdd gnd cell_6t
Xbit_r62_c61 bl_61 br_61 wl_62 vdd gnd cell_6t
Xbit_r63_c61 bl_61 br_61 wl_63 vdd gnd cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd cell_6t
Xbit_r1_c62 bl_62 br_62 wl_1 vdd gnd cell_6t
Xbit_r2_c62 bl_62 br_62 wl_2 vdd gnd cell_6t
Xbit_r3_c62 bl_62 br_62 wl_3 vdd gnd cell_6t
Xbit_r4_c62 bl_62 br_62 wl_4 vdd gnd cell_6t
Xbit_r5_c62 bl_62 br_62 wl_5 vdd gnd cell_6t
Xbit_r6_c62 bl_62 br_62 wl_6 vdd gnd cell_6t
Xbit_r7_c62 bl_62 br_62 wl_7 vdd gnd cell_6t
Xbit_r8_c62 bl_62 br_62 wl_8 vdd gnd cell_6t
Xbit_r9_c62 bl_62 br_62 wl_9 vdd gnd cell_6t
Xbit_r10_c62 bl_62 br_62 wl_10 vdd gnd cell_6t
Xbit_r11_c62 bl_62 br_62 wl_11 vdd gnd cell_6t
Xbit_r12_c62 bl_62 br_62 wl_12 vdd gnd cell_6t
Xbit_r13_c62 bl_62 br_62 wl_13 vdd gnd cell_6t
Xbit_r14_c62 bl_62 br_62 wl_14 vdd gnd cell_6t
Xbit_r15_c62 bl_62 br_62 wl_15 vdd gnd cell_6t
Xbit_r16_c62 bl_62 br_62 wl_16 vdd gnd cell_6t
Xbit_r17_c62 bl_62 br_62 wl_17 vdd gnd cell_6t
Xbit_r18_c62 bl_62 br_62 wl_18 vdd gnd cell_6t
Xbit_r19_c62 bl_62 br_62 wl_19 vdd gnd cell_6t
Xbit_r20_c62 bl_62 br_62 wl_20 vdd gnd cell_6t
Xbit_r21_c62 bl_62 br_62 wl_21 vdd gnd cell_6t
Xbit_r22_c62 bl_62 br_62 wl_22 vdd gnd cell_6t
Xbit_r23_c62 bl_62 br_62 wl_23 vdd gnd cell_6t
Xbit_r24_c62 bl_62 br_62 wl_24 vdd gnd cell_6t
Xbit_r25_c62 bl_62 br_62 wl_25 vdd gnd cell_6t
Xbit_r26_c62 bl_62 br_62 wl_26 vdd gnd cell_6t
Xbit_r27_c62 bl_62 br_62 wl_27 vdd gnd cell_6t
Xbit_r28_c62 bl_62 br_62 wl_28 vdd gnd cell_6t
Xbit_r29_c62 bl_62 br_62 wl_29 vdd gnd cell_6t
Xbit_r30_c62 bl_62 br_62 wl_30 vdd gnd cell_6t
Xbit_r31_c62 bl_62 br_62 wl_31 vdd gnd cell_6t
Xbit_r32_c62 bl_62 br_62 wl_32 vdd gnd cell_6t
Xbit_r33_c62 bl_62 br_62 wl_33 vdd gnd cell_6t
Xbit_r34_c62 bl_62 br_62 wl_34 vdd gnd cell_6t
Xbit_r35_c62 bl_62 br_62 wl_35 vdd gnd cell_6t
Xbit_r36_c62 bl_62 br_62 wl_36 vdd gnd cell_6t
Xbit_r37_c62 bl_62 br_62 wl_37 vdd gnd cell_6t
Xbit_r38_c62 bl_62 br_62 wl_38 vdd gnd cell_6t
Xbit_r39_c62 bl_62 br_62 wl_39 vdd gnd cell_6t
Xbit_r40_c62 bl_62 br_62 wl_40 vdd gnd cell_6t
Xbit_r41_c62 bl_62 br_62 wl_41 vdd gnd cell_6t
Xbit_r42_c62 bl_62 br_62 wl_42 vdd gnd cell_6t
Xbit_r43_c62 bl_62 br_62 wl_43 vdd gnd cell_6t
Xbit_r44_c62 bl_62 br_62 wl_44 vdd gnd cell_6t
Xbit_r45_c62 bl_62 br_62 wl_45 vdd gnd cell_6t
Xbit_r46_c62 bl_62 br_62 wl_46 vdd gnd cell_6t
Xbit_r47_c62 bl_62 br_62 wl_47 vdd gnd cell_6t
Xbit_r48_c62 bl_62 br_62 wl_48 vdd gnd cell_6t
Xbit_r49_c62 bl_62 br_62 wl_49 vdd gnd cell_6t
Xbit_r50_c62 bl_62 br_62 wl_50 vdd gnd cell_6t
Xbit_r51_c62 bl_62 br_62 wl_51 vdd gnd cell_6t
Xbit_r52_c62 bl_62 br_62 wl_52 vdd gnd cell_6t
Xbit_r53_c62 bl_62 br_62 wl_53 vdd gnd cell_6t
Xbit_r54_c62 bl_62 br_62 wl_54 vdd gnd cell_6t
Xbit_r55_c62 bl_62 br_62 wl_55 vdd gnd cell_6t
Xbit_r56_c62 bl_62 br_62 wl_56 vdd gnd cell_6t
Xbit_r57_c62 bl_62 br_62 wl_57 vdd gnd cell_6t
Xbit_r58_c62 bl_62 br_62 wl_58 vdd gnd cell_6t
Xbit_r59_c62 bl_62 br_62 wl_59 vdd gnd cell_6t
Xbit_r60_c62 bl_62 br_62 wl_60 vdd gnd cell_6t
Xbit_r61_c62 bl_62 br_62 wl_61 vdd gnd cell_6t
Xbit_r62_c62 bl_62 br_62 wl_62 vdd gnd cell_6t
Xbit_r63_c62 bl_62 br_62 wl_63 vdd gnd cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd cell_6t
Xbit_r1_c63 bl_63 br_63 wl_1 vdd gnd cell_6t
Xbit_r2_c63 bl_63 br_63 wl_2 vdd gnd cell_6t
Xbit_r3_c63 bl_63 br_63 wl_3 vdd gnd cell_6t
Xbit_r4_c63 bl_63 br_63 wl_4 vdd gnd cell_6t
Xbit_r5_c63 bl_63 br_63 wl_5 vdd gnd cell_6t
Xbit_r6_c63 bl_63 br_63 wl_6 vdd gnd cell_6t
Xbit_r7_c63 bl_63 br_63 wl_7 vdd gnd cell_6t
Xbit_r8_c63 bl_63 br_63 wl_8 vdd gnd cell_6t
Xbit_r9_c63 bl_63 br_63 wl_9 vdd gnd cell_6t
Xbit_r10_c63 bl_63 br_63 wl_10 vdd gnd cell_6t
Xbit_r11_c63 bl_63 br_63 wl_11 vdd gnd cell_6t
Xbit_r12_c63 bl_63 br_63 wl_12 vdd gnd cell_6t
Xbit_r13_c63 bl_63 br_63 wl_13 vdd gnd cell_6t
Xbit_r14_c63 bl_63 br_63 wl_14 vdd gnd cell_6t
Xbit_r15_c63 bl_63 br_63 wl_15 vdd gnd cell_6t
Xbit_r16_c63 bl_63 br_63 wl_16 vdd gnd cell_6t
Xbit_r17_c63 bl_63 br_63 wl_17 vdd gnd cell_6t
Xbit_r18_c63 bl_63 br_63 wl_18 vdd gnd cell_6t
Xbit_r19_c63 bl_63 br_63 wl_19 vdd gnd cell_6t
Xbit_r20_c63 bl_63 br_63 wl_20 vdd gnd cell_6t
Xbit_r21_c63 bl_63 br_63 wl_21 vdd gnd cell_6t
Xbit_r22_c63 bl_63 br_63 wl_22 vdd gnd cell_6t
Xbit_r23_c63 bl_63 br_63 wl_23 vdd gnd cell_6t
Xbit_r24_c63 bl_63 br_63 wl_24 vdd gnd cell_6t
Xbit_r25_c63 bl_63 br_63 wl_25 vdd gnd cell_6t
Xbit_r26_c63 bl_63 br_63 wl_26 vdd gnd cell_6t
Xbit_r27_c63 bl_63 br_63 wl_27 vdd gnd cell_6t
Xbit_r28_c63 bl_63 br_63 wl_28 vdd gnd cell_6t
Xbit_r29_c63 bl_63 br_63 wl_29 vdd gnd cell_6t
Xbit_r30_c63 bl_63 br_63 wl_30 vdd gnd cell_6t
Xbit_r31_c63 bl_63 br_63 wl_31 vdd gnd cell_6t
Xbit_r32_c63 bl_63 br_63 wl_32 vdd gnd cell_6t
Xbit_r33_c63 bl_63 br_63 wl_33 vdd gnd cell_6t
Xbit_r34_c63 bl_63 br_63 wl_34 vdd gnd cell_6t
Xbit_r35_c63 bl_63 br_63 wl_35 vdd gnd cell_6t
Xbit_r36_c63 bl_63 br_63 wl_36 vdd gnd cell_6t
Xbit_r37_c63 bl_63 br_63 wl_37 vdd gnd cell_6t
Xbit_r38_c63 bl_63 br_63 wl_38 vdd gnd cell_6t
Xbit_r39_c63 bl_63 br_63 wl_39 vdd gnd cell_6t
Xbit_r40_c63 bl_63 br_63 wl_40 vdd gnd cell_6t
Xbit_r41_c63 bl_63 br_63 wl_41 vdd gnd cell_6t
Xbit_r42_c63 bl_63 br_63 wl_42 vdd gnd cell_6t
Xbit_r43_c63 bl_63 br_63 wl_43 vdd gnd cell_6t
Xbit_r44_c63 bl_63 br_63 wl_44 vdd gnd cell_6t
Xbit_r45_c63 bl_63 br_63 wl_45 vdd gnd cell_6t
Xbit_r46_c63 bl_63 br_63 wl_46 vdd gnd cell_6t
Xbit_r47_c63 bl_63 br_63 wl_47 vdd gnd cell_6t
Xbit_r48_c63 bl_63 br_63 wl_48 vdd gnd cell_6t
Xbit_r49_c63 bl_63 br_63 wl_49 vdd gnd cell_6t
Xbit_r50_c63 bl_63 br_63 wl_50 vdd gnd cell_6t
Xbit_r51_c63 bl_63 br_63 wl_51 vdd gnd cell_6t
Xbit_r52_c63 bl_63 br_63 wl_52 vdd gnd cell_6t
Xbit_r53_c63 bl_63 br_63 wl_53 vdd gnd cell_6t
Xbit_r54_c63 bl_63 br_63 wl_54 vdd gnd cell_6t
Xbit_r55_c63 bl_63 br_63 wl_55 vdd gnd cell_6t
Xbit_r56_c63 bl_63 br_63 wl_56 vdd gnd cell_6t
Xbit_r57_c63 bl_63 br_63 wl_57 vdd gnd cell_6t
Xbit_r58_c63 bl_63 br_63 wl_58 vdd gnd cell_6t
Xbit_r59_c63 bl_63 br_63 wl_59 vdd gnd cell_6t
Xbit_r60_c63 bl_63 br_63 wl_60 vdd gnd cell_6t
Xbit_r61_c63 bl_63 br_63 wl_61 vdd gnd cell_6t
Xbit_r62_c63 bl_63 br_63 wl_62 vdd gnd cell_6t
Xbit_r63_c63 bl_63 br_63 wl_63 vdd gnd cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd cell_6t
Xbit_r1_c64 bl_64 br_64 wl_1 vdd gnd cell_6t
Xbit_r2_c64 bl_64 br_64 wl_2 vdd gnd cell_6t
Xbit_r3_c64 bl_64 br_64 wl_3 vdd gnd cell_6t
Xbit_r4_c64 bl_64 br_64 wl_4 vdd gnd cell_6t
Xbit_r5_c64 bl_64 br_64 wl_5 vdd gnd cell_6t
Xbit_r6_c64 bl_64 br_64 wl_6 vdd gnd cell_6t
Xbit_r7_c64 bl_64 br_64 wl_7 vdd gnd cell_6t
Xbit_r8_c64 bl_64 br_64 wl_8 vdd gnd cell_6t
Xbit_r9_c64 bl_64 br_64 wl_9 vdd gnd cell_6t
Xbit_r10_c64 bl_64 br_64 wl_10 vdd gnd cell_6t
Xbit_r11_c64 bl_64 br_64 wl_11 vdd gnd cell_6t
Xbit_r12_c64 bl_64 br_64 wl_12 vdd gnd cell_6t
Xbit_r13_c64 bl_64 br_64 wl_13 vdd gnd cell_6t
Xbit_r14_c64 bl_64 br_64 wl_14 vdd gnd cell_6t
Xbit_r15_c64 bl_64 br_64 wl_15 vdd gnd cell_6t
Xbit_r16_c64 bl_64 br_64 wl_16 vdd gnd cell_6t
Xbit_r17_c64 bl_64 br_64 wl_17 vdd gnd cell_6t
Xbit_r18_c64 bl_64 br_64 wl_18 vdd gnd cell_6t
Xbit_r19_c64 bl_64 br_64 wl_19 vdd gnd cell_6t
Xbit_r20_c64 bl_64 br_64 wl_20 vdd gnd cell_6t
Xbit_r21_c64 bl_64 br_64 wl_21 vdd gnd cell_6t
Xbit_r22_c64 bl_64 br_64 wl_22 vdd gnd cell_6t
Xbit_r23_c64 bl_64 br_64 wl_23 vdd gnd cell_6t
Xbit_r24_c64 bl_64 br_64 wl_24 vdd gnd cell_6t
Xbit_r25_c64 bl_64 br_64 wl_25 vdd gnd cell_6t
Xbit_r26_c64 bl_64 br_64 wl_26 vdd gnd cell_6t
Xbit_r27_c64 bl_64 br_64 wl_27 vdd gnd cell_6t
Xbit_r28_c64 bl_64 br_64 wl_28 vdd gnd cell_6t
Xbit_r29_c64 bl_64 br_64 wl_29 vdd gnd cell_6t
Xbit_r30_c64 bl_64 br_64 wl_30 vdd gnd cell_6t
Xbit_r31_c64 bl_64 br_64 wl_31 vdd gnd cell_6t
Xbit_r32_c64 bl_64 br_64 wl_32 vdd gnd cell_6t
Xbit_r33_c64 bl_64 br_64 wl_33 vdd gnd cell_6t
Xbit_r34_c64 bl_64 br_64 wl_34 vdd gnd cell_6t
Xbit_r35_c64 bl_64 br_64 wl_35 vdd gnd cell_6t
Xbit_r36_c64 bl_64 br_64 wl_36 vdd gnd cell_6t
Xbit_r37_c64 bl_64 br_64 wl_37 vdd gnd cell_6t
Xbit_r38_c64 bl_64 br_64 wl_38 vdd gnd cell_6t
Xbit_r39_c64 bl_64 br_64 wl_39 vdd gnd cell_6t
Xbit_r40_c64 bl_64 br_64 wl_40 vdd gnd cell_6t
Xbit_r41_c64 bl_64 br_64 wl_41 vdd gnd cell_6t
Xbit_r42_c64 bl_64 br_64 wl_42 vdd gnd cell_6t
Xbit_r43_c64 bl_64 br_64 wl_43 vdd gnd cell_6t
Xbit_r44_c64 bl_64 br_64 wl_44 vdd gnd cell_6t
Xbit_r45_c64 bl_64 br_64 wl_45 vdd gnd cell_6t
Xbit_r46_c64 bl_64 br_64 wl_46 vdd gnd cell_6t
Xbit_r47_c64 bl_64 br_64 wl_47 vdd gnd cell_6t
Xbit_r48_c64 bl_64 br_64 wl_48 vdd gnd cell_6t
Xbit_r49_c64 bl_64 br_64 wl_49 vdd gnd cell_6t
Xbit_r50_c64 bl_64 br_64 wl_50 vdd gnd cell_6t
Xbit_r51_c64 bl_64 br_64 wl_51 vdd gnd cell_6t
Xbit_r52_c64 bl_64 br_64 wl_52 vdd gnd cell_6t
Xbit_r53_c64 bl_64 br_64 wl_53 vdd gnd cell_6t
Xbit_r54_c64 bl_64 br_64 wl_54 vdd gnd cell_6t
Xbit_r55_c64 bl_64 br_64 wl_55 vdd gnd cell_6t
Xbit_r56_c64 bl_64 br_64 wl_56 vdd gnd cell_6t
Xbit_r57_c64 bl_64 br_64 wl_57 vdd gnd cell_6t
Xbit_r58_c64 bl_64 br_64 wl_58 vdd gnd cell_6t
Xbit_r59_c64 bl_64 br_64 wl_59 vdd gnd cell_6t
Xbit_r60_c64 bl_64 br_64 wl_60 vdd gnd cell_6t
Xbit_r61_c64 bl_64 br_64 wl_61 vdd gnd cell_6t
Xbit_r62_c64 bl_64 br_64 wl_62 vdd gnd cell_6t
Xbit_r63_c64 bl_64 br_64 wl_63 vdd gnd cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd cell_6t
Xbit_r1_c65 bl_65 br_65 wl_1 vdd gnd cell_6t
Xbit_r2_c65 bl_65 br_65 wl_2 vdd gnd cell_6t
Xbit_r3_c65 bl_65 br_65 wl_3 vdd gnd cell_6t
Xbit_r4_c65 bl_65 br_65 wl_4 vdd gnd cell_6t
Xbit_r5_c65 bl_65 br_65 wl_5 vdd gnd cell_6t
Xbit_r6_c65 bl_65 br_65 wl_6 vdd gnd cell_6t
Xbit_r7_c65 bl_65 br_65 wl_7 vdd gnd cell_6t
Xbit_r8_c65 bl_65 br_65 wl_8 vdd gnd cell_6t
Xbit_r9_c65 bl_65 br_65 wl_9 vdd gnd cell_6t
Xbit_r10_c65 bl_65 br_65 wl_10 vdd gnd cell_6t
Xbit_r11_c65 bl_65 br_65 wl_11 vdd gnd cell_6t
Xbit_r12_c65 bl_65 br_65 wl_12 vdd gnd cell_6t
Xbit_r13_c65 bl_65 br_65 wl_13 vdd gnd cell_6t
Xbit_r14_c65 bl_65 br_65 wl_14 vdd gnd cell_6t
Xbit_r15_c65 bl_65 br_65 wl_15 vdd gnd cell_6t
Xbit_r16_c65 bl_65 br_65 wl_16 vdd gnd cell_6t
Xbit_r17_c65 bl_65 br_65 wl_17 vdd gnd cell_6t
Xbit_r18_c65 bl_65 br_65 wl_18 vdd gnd cell_6t
Xbit_r19_c65 bl_65 br_65 wl_19 vdd gnd cell_6t
Xbit_r20_c65 bl_65 br_65 wl_20 vdd gnd cell_6t
Xbit_r21_c65 bl_65 br_65 wl_21 vdd gnd cell_6t
Xbit_r22_c65 bl_65 br_65 wl_22 vdd gnd cell_6t
Xbit_r23_c65 bl_65 br_65 wl_23 vdd gnd cell_6t
Xbit_r24_c65 bl_65 br_65 wl_24 vdd gnd cell_6t
Xbit_r25_c65 bl_65 br_65 wl_25 vdd gnd cell_6t
Xbit_r26_c65 bl_65 br_65 wl_26 vdd gnd cell_6t
Xbit_r27_c65 bl_65 br_65 wl_27 vdd gnd cell_6t
Xbit_r28_c65 bl_65 br_65 wl_28 vdd gnd cell_6t
Xbit_r29_c65 bl_65 br_65 wl_29 vdd gnd cell_6t
Xbit_r30_c65 bl_65 br_65 wl_30 vdd gnd cell_6t
Xbit_r31_c65 bl_65 br_65 wl_31 vdd gnd cell_6t
Xbit_r32_c65 bl_65 br_65 wl_32 vdd gnd cell_6t
Xbit_r33_c65 bl_65 br_65 wl_33 vdd gnd cell_6t
Xbit_r34_c65 bl_65 br_65 wl_34 vdd gnd cell_6t
Xbit_r35_c65 bl_65 br_65 wl_35 vdd gnd cell_6t
Xbit_r36_c65 bl_65 br_65 wl_36 vdd gnd cell_6t
Xbit_r37_c65 bl_65 br_65 wl_37 vdd gnd cell_6t
Xbit_r38_c65 bl_65 br_65 wl_38 vdd gnd cell_6t
Xbit_r39_c65 bl_65 br_65 wl_39 vdd gnd cell_6t
Xbit_r40_c65 bl_65 br_65 wl_40 vdd gnd cell_6t
Xbit_r41_c65 bl_65 br_65 wl_41 vdd gnd cell_6t
Xbit_r42_c65 bl_65 br_65 wl_42 vdd gnd cell_6t
Xbit_r43_c65 bl_65 br_65 wl_43 vdd gnd cell_6t
Xbit_r44_c65 bl_65 br_65 wl_44 vdd gnd cell_6t
Xbit_r45_c65 bl_65 br_65 wl_45 vdd gnd cell_6t
Xbit_r46_c65 bl_65 br_65 wl_46 vdd gnd cell_6t
Xbit_r47_c65 bl_65 br_65 wl_47 vdd gnd cell_6t
Xbit_r48_c65 bl_65 br_65 wl_48 vdd gnd cell_6t
Xbit_r49_c65 bl_65 br_65 wl_49 vdd gnd cell_6t
Xbit_r50_c65 bl_65 br_65 wl_50 vdd gnd cell_6t
Xbit_r51_c65 bl_65 br_65 wl_51 vdd gnd cell_6t
Xbit_r52_c65 bl_65 br_65 wl_52 vdd gnd cell_6t
Xbit_r53_c65 bl_65 br_65 wl_53 vdd gnd cell_6t
Xbit_r54_c65 bl_65 br_65 wl_54 vdd gnd cell_6t
Xbit_r55_c65 bl_65 br_65 wl_55 vdd gnd cell_6t
Xbit_r56_c65 bl_65 br_65 wl_56 vdd gnd cell_6t
Xbit_r57_c65 bl_65 br_65 wl_57 vdd gnd cell_6t
Xbit_r58_c65 bl_65 br_65 wl_58 vdd gnd cell_6t
Xbit_r59_c65 bl_65 br_65 wl_59 vdd gnd cell_6t
Xbit_r60_c65 bl_65 br_65 wl_60 vdd gnd cell_6t
Xbit_r61_c65 bl_65 br_65 wl_61 vdd gnd cell_6t
Xbit_r62_c65 bl_65 br_65 wl_62 vdd gnd cell_6t
Xbit_r63_c65 bl_65 br_65 wl_63 vdd gnd cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd cell_6t
Xbit_r1_c66 bl_66 br_66 wl_1 vdd gnd cell_6t
Xbit_r2_c66 bl_66 br_66 wl_2 vdd gnd cell_6t
Xbit_r3_c66 bl_66 br_66 wl_3 vdd gnd cell_6t
Xbit_r4_c66 bl_66 br_66 wl_4 vdd gnd cell_6t
Xbit_r5_c66 bl_66 br_66 wl_5 vdd gnd cell_6t
Xbit_r6_c66 bl_66 br_66 wl_6 vdd gnd cell_6t
Xbit_r7_c66 bl_66 br_66 wl_7 vdd gnd cell_6t
Xbit_r8_c66 bl_66 br_66 wl_8 vdd gnd cell_6t
Xbit_r9_c66 bl_66 br_66 wl_9 vdd gnd cell_6t
Xbit_r10_c66 bl_66 br_66 wl_10 vdd gnd cell_6t
Xbit_r11_c66 bl_66 br_66 wl_11 vdd gnd cell_6t
Xbit_r12_c66 bl_66 br_66 wl_12 vdd gnd cell_6t
Xbit_r13_c66 bl_66 br_66 wl_13 vdd gnd cell_6t
Xbit_r14_c66 bl_66 br_66 wl_14 vdd gnd cell_6t
Xbit_r15_c66 bl_66 br_66 wl_15 vdd gnd cell_6t
Xbit_r16_c66 bl_66 br_66 wl_16 vdd gnd cell_6t
Xbit_r17_c66 bl_66 br_66 wl_17 vdd gnd cell_6t
Xbit_r18_c66 bl_66 br_66 wl_18 vdd gnd cell_6t
Xbit_r19_c66 bl_66 br_66 wl_19 vdd gnd cell_6t
Xbit_r20_c66 bl_66 br_66 wl_20 vdd gnd cell_6t
Xbit_r21_c66 bl_66 br_66 wl_21 vdd gnd cell_6t
Xbit_r22_c66 bl_66 br_66 wl_22 vdd gnd cell_6t
Xbit_r23_c66 bl_66 br_66 wl_23 vdd gnd cell_6t
Xbit_r24_c66 bl_66 br_66 wl_24 vdd gnd cell_6t
Xbit_r25_c66 bl_66 br_66 wl_25 vdd gnd cell_6t
Xbit_r26_c66 bl_66 br_66 wl_26 vdd gnd cell_6t
Xbit_r27_c66 bl_66 br_66 wl_27 vdd gnd cell_6t
Xbit_r28_c66 bl_66 br_66 wl_28 vdd gnd cell_6t
Xbit_r29_c66 bl_66 br_66 wl_29 vdd gnd cell_6t
Xbit_r30_c66 bl_66 br_66 wl_30 vdd gnd cell_6t
Xbit_r31_c66 bl_66 br_66 wl_31 vdd gnd cell_6t
Xbit_r32_c66 bl_66 br_66 wl_32 vdd gnd cell_6t
Xbit_r33_c66 bl_66 br_66 wl_33 vdd gnd cell_6t
Xbit_r34_c66 bl_66 br_66 wl_34 vdd gnd cell_6t
Xbit_r35_c66 bl_66 br_66 wl_35 vdd gnd cell_6t
Xbit_r36_c66 bl_66 br_66 wl_36 vdd gnd cell_6t
Xbit_r37_c66 bl_66 br_66 wl_37 vdd gnd cell_6t
Xbit_r38_c66 bl_66 br_66 wl_38 vdd gnd cell_6t
Xbit_r39_c66 bl_66 br_66 wl_39 vdd gnd cell_6t
Xbit_r40_c66 bl_66 br_66 wl_40 vdd gnd cell_6t
Xbit_r41_c66 bl_66 br_66 wl_41 vdd gnd cell_6t
Xbit_r42_c66 bl_66 br_66 wl_42 vdd gnd cell_6t
Xbit_r43_c66 bl_66 br_66 wl_43 vdd gnd cell_6t
Xbit_r44_c66 bl_66 br_66 wl_44 vdd gnd cell_6t
Xbit_r45_c66 bl_66 br_66 wl_45 vdd gnd cell_6t
Xbit_r46_c66 bl_66 br_66 wl_46 vdd gnd cell_6t
Xbit_r47_c66 bl_66 br_66 wl_47 vdd gnd cell_6t
Xbit_r48_c66 bl_66 br_66 wl_48 vdd gnd cell_6t
Xbit_r49_c66 bl_66 br_66 wl_49 vdd gnd cell_6t
Xbit_r50_c66 bl_66 br_66 wl_50 vdd gnd cell_6t
Xbit_r51_c66 bl_66 br_66 wl_51 vdd gnd cell_6t
Xbit_r52_c66 bl_66 br_66 wl_52 vdd gnd cell_6t
Xbit_r53_c66 bl_66 br_66 wl_53 vdd gnd cell_6t
Xbit_r54_c66 bl_66 br_66 wl_54 vdd gnd cell_6t
Xbit_r55_c66 bl_66 br_66 wl_55 vdd gnd cell_6t
Xbit_r56_c66 bl_66 br_66 wl_56 vdd gnd cell_6t
Xbit_r57_c66 bl_66 br_66 wl_57 vdd gnd cell_6t
Xbit_r58_c66 bl_66 br_66 wl_58 vdd gnd cell_6t
Xbit_r59_c66 bl_66 br_66 wl_59 vdd gnd cell_6t
Xbit_r60_c66 bl_66 br_66 wl_60 vdd gnd cell_6t
Xbit_r61_c66 bl_66 br_66 wl_61 vdd gnd cell_6t
Xbit_r62_c66 bl_66 br_66 wl_62 vdd gnd cell_6t
Xbit_r63_c66 bl_66 br_66 wl_63 vdd gnd cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd cell_6t
Xbit_r1_c67 bl_67 br_67 wl_1 vdd gnd cell_6t
Xbit_r2_c67 bl_67 br_67 wl_2 vdd gnd cell_6t
Xbit_r3_c67 bl_67 br_67 wl_3 vdd gnd cell_6t
Xbit_r4_c67 bl_67 br_67 wl_4 vdd gnd cell_6t
Xbit_r5_c67 bl_67 br_67 wl_5 vdd gnd cell_6t
Xbit_r6_c67 bl_67 br_67 wl_6 vdd gnd cell_6t
Xbit_r7_c67 bl_67 br_67 wl_7 vdd gnd cell_6t
Xbit_r8_c67 bl_67 br_67 wl_8 vdd gnd cell_6t
Xbit_r9_c67 bl_67 br_67 wl_9 vdd gnd cell_6t
Xbit_r10_c67 bl_67 br_67 wl_10 vdd gnd cell_6t
Xbit_r11_c67 bl_67 br_67 wl_11 vdd gnd cell_6t
Xbit_r12_c67 bl_67 br_67 wl_12 vdd gnd cell_6t
Xbit_r13_c67 bl_67 br_67 wl_13 vdd gnd cell_6t
Xbit_r14_c67 bl_67 br_67 wl_14 vdd gnd cell_6t
Xbit_r15_c67 bl_67 br_67 wl_15 vdd gnd cell_6t
Xbit_r16_c67 bl_67 br_67 wl_16 vdd gnd cell_6t
Xbit_r17_c67 bl_67 br_67 wl_17 vdd gnd cell_6t
Xbit_r18_c67 bl_67 br_67 wl_18 vdd gnd cell_6t
Xbit_r19_c67 bl_67 br_67 wl_19 vdd gnd cell_6t
Xbit_r20_c67 bl_67 br_67 wl_20 vdd gnd cell_6t
Xbit_r21_c67 bl_67 br_67 wl_21 vdd gnd cell_6t
Xbit_r22_c67 bl_67 br_67 wl_22 vdd gnd cell_6t
Xbit_r23_c67 bl_67 br_67 wl_23 vdd gnd cell_6t
Xbit_r24_c67 bl_67 br_67 wl_24 vdd gnd cell_6t
Xbit_r25_c67 bl_67 br_67 wl_25 vdd gnd cell_6t
Xbit_r26_c67 bl_67 br_67 wl_26 vdd gnd cell_6t
Xbit_r27_c67 bl_67 br_67 wl_27 vdd gnd cell_6t
Xbit_r28_c67 bl_67 br_67 wl_28 vdd gnd cell_6t
Xbit_r29_c67 bl_67 br_67 wl_29 vdd gnd cell_6t
Xbit_r30_c67 bl_67 br_67 wl_30 vdd gnd cell_6t
Xbit_r31_c67 bl_67 br_67 wl_31 vdd gnd cell_6t
Xbit_r32_c67 bl_67 br_67 wl_32 vdd gnd cell_6t
Xbit_r33_c67 bl_67 br_67 wl_33 vdd gnd cell_6t
Xbit_r34_c67 bl_67 br_67 wl_34 vdd gnd cell_6t
Xbit_r35_c67 bl_67 br_67 wl_35 vdd gnd cell_6t
Xbit_r36_c67 bl_67 br_67 wl_36 vdd gnd cell_6t
Xbit_r37_c67 bl_67 br_67 wl_37 vdd gnd cell_6t
Xbit_r38_c67 bl_67 br_67 wl_38 vdd gnd cell_6t
Xbit_r39_c67 bl_67 br_67 wl_39 vdd gnd cell_6t
Xbit_r40_c67 bl_67 br_67 wl_40 vdd gnd cell_6t
Xbit_r41_c67 bl_67 br_67 wl_41 vdd gnd cell_6t
Xbit_r42_c67 bl_67 br_67 wl_42 vdd gnd cell_6t
Xbit_r43_c67 bl_67 br_67 wl_43 vdd gnd cell_6t
Xbit_r44_c67 bl_67 br_67 wl_44 vdd gnd cell_6t
Xbit_r45_c67 bl_67 br_67 wl_45 vdd gnd cell_6t
Xbit_r46_c67 bl_67 br_67 wl_46 vdd gnd cell_6t
Xbit_r47_c67 bl_67 br_67 wl_47 vdd gnd cell_6t
Xbit_r48_c67 bl_67 br_67 wl_48 vdd gnd cell_6t
Xbit_r49_c67 bl_67 br_67 wl_49 vdd gnd cell_6t
Xbit_r50_c67 bl_67 br_67 wl_50 vdd gnd cell_6t
Xbit_r51_c67 bl_67 br_67 wl_51 vdd gnd cell_6t
Xbit_r52_c67 bl_67 br_67 wl_52 vdd gnd cell_6t
Xbit_r53_c67 bl_67 br_67 wl_53 vdd gnd cell_6t
Xbit_r54_c67 bl_67 br_67 wl_54 vdd gnd cell_6t
Xbit_r55_c67 bl_67 br_67 wl_55 vdd gnd cell_6t
Xbit_r56_c67 bl_67 br_67 wl_56 vdd gnd cell_6t
Xbit_r57_c67 bl_67 br_67 wl_57 vdd gnd cell_6t
Xbit_r58_c67 bl_67 br_67 wl_58 vdd gnd cell_6t
Xbit_r59_c67 bl_67 br_67 wl_59 vdd gnd cell_6t
Xbit_r60_c67 bl_67 br_67 wl_60 vdd gnd cell_6t
Xbit_r61_c67 bl_67 br_67 wl_61 vdd gnd cell_6t
Xbit_r62_c67 bl_67 br_67 wl_62 vdd gnd cell_6t
Xbit_r63_c67 bl_67 br_67 wl_63 vdd gnd cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd cell_6t
Xbit_r1_c68 bl_68 br_68 wl_1 vdd gnd cell_6t
Xbit_r2_c68 bl_68 br_68 wl_2 vdd gnd cell_6t
Xbit_r3_c68 bl_68 br_68 wl_3 vdd gnd cell_6t
Xbit_r4_c68 bl_68 br_68 wl_4 vdd gnd cell_6t
Xbit_r5_c68 bl_68 br_68 wl_5 vdd gnd cell_6t
Xbit_r6_c68 bl_68 br_68 wl_6 vdd gnd cell_6t
Xbit_r7_c68 bl_68 br_68 wl_7 vdd gnd cell_6t
Xbit_r8_c68 bl_68 br_68 wl_8 vdd gnd cell_6t
Xbit_r9_c68 bl_68 br_68 wl_9 vdd gnd cell_6t
Xbit_r10_c68 bl_68 br_68 wl_10 vdd gnd cell_6t
Xbit_r11_c68 bl_68 br_68 wl_11 vdd gnd cell_6t
Xbit_r12_c68 bl_68 br_68 wl_12 vdd gnd cell_6t
Xbit_r13_c68 bl_68 br_68 wl_13 vdd gnd cell_6t
Xbit_r14_c68 bl_68 br_68 wl_14 vdd gnd cell_6t
Xbit_r15_c68 bl_68 br_68 wl_15 vdd gnd cell_6t
Xbit_r16_c68 bl_68 br_68 wl_16 vdd gnd cell_6t
Xbit_r17_c68 bl_68 br_68 wl_17 vdd gnd cell_6t
Xbit_r18_c68 bl_68 br_68 wl_18 vdd gnd cell_6t
Xbit_r19_c68 bl_68 br_68 wl_19 vdd gnd cell_6t
Xbit_r20_c68 bl_68 br_68 wl_20 vdd gnd cell_6t
Xbit_r21_c68 bl_68 br_68 wl_21 vdd gnd cell_6t
Xbit_r22_c68 bl_68 br_68 wl_22 vdd gnd cell_6t
Xbit_r23_c68 bl_68 br_68 wl_23 vdd gnd cell_6t
Xbit_r24_c68 bl_68 br_68 wl_24 vdd gnd cell_6t
Xbit_r25_c68 bl_68 br_68 wl_25 vdd gnd cell_6t
Xbit_r26_c68 bl_68 br_68 wl_26 vdd gnd cell_6t
Xbit_r27_c68 bl_68 br_68 wl_27 vdd gnd cell_6t
Xbit_r28_c68 bl_68 br_68 wl_28 vdd gnd cell_6t
Xbit_r29_c68 bl_68 br_68 wl_29 vdd gnd cell_6t
Xbit_r30_c68 bl_68 br_68 wl_30 vdd gnd cell_6t
Xbit_r31_c68 bl_68 br_68 wl_31 vdd gnd cell_6t
Xbit_r32_c68 bl_68 br_68 wl_32 vdd gnd cell_6t
Xbit_r33_c68 bl_68 br_68 wl_33 vdd gnd cell_6t
Xbit_r34_c68 bl_68 br_68 wl_34 vdd gnd cell_6t
Xbit_r35_c68 bl_68 br_68 wl_35 vdd gnd cell_6t
Xbit_r36_c68 bl_68 br_68 wl_36 vdd gnd cell_6t
Xbit_r37_c68 bl_68 br_68 wl_37 vdd gnd cell_6t
Xbit_r38_c68 bl_68 br_68 wl_38 vdd gnd cell_6t
Xbit_r39_c68 bl_68 br_68 wl_39 vdd gnd cell_6t
Xbit_r40_c68 bl_68 br_68 wl_40 vdd gnd cell_6t
Xbit_r41_c68 bl_68 br_68 wl_41 vdd gnd cell_6t
Xbit_r42_c68 bl_68 br_68 wl_42 vdd gnd cell_6t
Xbit_r43_c68 bl_68 br_68 wl_43 vdd gnd cell_6t
Xbit_r44_c68 bl_68 br_68 wl_44 vdd gnd cell_6t
Xbit_r45_c68 bl_68 br_68 wl_45 vdd gnd cell_6t
Xbit_r46_c68 bl_68 br_68 wl_46 vdd gnd cell_6t
Xbit_r47_c68 bl_68 br_68 wl_47 vdd gnd cell_6t
Xbit_r48_c68 bl_68 br_68 wl_48 vdd gnd cell_6t
Xbit_r49_c68 bl_68 br_68 wl_49 vdd gnd cell_6t
Xbit_r50_c68 bl_68 br_68 wl_50 vdd gnd cell_6t
Xbit_r51_c68 bl_68 br_68 wl_51 vdd gnd cell_6t
Xbit_r52_c68 bl_68 br_68 wl_52 vdd gnd cell_6t
Xbit_r53_c68 bl_68 br_68 wl_53 vdd gnd cell_6t
Xbit_r54_c68 bl_68 br_68 wl_54 vdd gnd cell_6t
Xbit_r55_c68 bl_68 br_68 wl_55 vdd gnd cell_6t
Xbit_r56_c68 bl_68 br_68 wl_56 vdd gnd cell_6t
Xbit_r57_c68 bl_68 br_68 wl_57 vdd gnd cell_6t
Xbit_r58_c68 bl_68 br_68 wl_58 vdd gnd cell_6t
Xbit_r59_c68 bl_68 br_68 wl_59 vdd gnd cell_6t
Xbit_r60_c68 bl_68 br_68 wl_60 vdd gnd cell_6t
Xbit_r61_c68 bl_68 br_68 wl_61 vdd gnd cell_6t
Xbit_r62_c68 bl_68 br_68 wl_62 vdd gnd cell_6t
Xbit_r63_c68 bl_68 br_68 wl_63 vdd gnd cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd cell_6t
Xbit_r1_c69 bl_69 br_69 wl_1 vdd gnd cell_6t
Xbit_r2_c69 bl_69 br_69 wl_2 vdd gnd cell_6t
Xbit_r3_c69 bl_69 br_69 wl_3 vdd gnd cell_6t
Xbit_r4_c69 bl_69 br_69 wl_4 vdd gnd cell_6t
Xbit_r5_c69 bl_69 br_69 wl_5 vdd gnd cell_6t
Xbit_r6_c69 bl_69 br_69 wl_6 vdd gnd cell_6t
Xbit_r7_c69 bl_69 br_69 wl_7 vdd gnd cell_6t
Xbit_r8_c69 bl_69 br_69 wl_8 vdd gnd cell_6t
Xbit_r9_c69 bl_69 br_69 wl_9 vdd gnd cell_6t
Xbit_r10_c69 bl_69 br_69 wl_10 vdd gnd cell_6t
Xbit_r11_c69 bl_69 br_69 wl_11 vdd gnd cell_6t
Xbit_r12_c69 bl_69 br_69 wl_12 vdd gnd cell_6t
Xbit_r13_c69 bl_69 br_69 wl_13 vdd gnd cell_6t
Xbit_r14_c69 bl_69 br_69 wl_14 vdd gnd cell_6t
Xbit_r15_c69 bl_69 br_69 wl_15 vdd gnd cell_6t
Xbit_r16_c69 bl_69 br_69 wl_16 vdd gnd cell_6t
Xbit_r17_c69 bl_69 br_69 wl_17 vdd gnd cell_6t
Xbit_r18_c69 bl_69 br_69 wl_18 vdd gnd cell_6t
Xbit_r19_c69 bl_69 br_69 wl_19 vdd gnd cell_6t
Xbit_r20_c69 bl_69 br_69 wl_20 vdd gnd cell_6t
Xbit_r21_c69 bl_69 br_69 wl_21 vdd gnd cell_6t
Xbit_r22_c69 bl_69 br_69 wl_22 vdd gnd cell_6t
Xbit_r23_c69 bl_69 br_69 wl_23 vdd gnd cell_6t
Xbit_r24_c69 bl_69 br_69 wl_24 vdd gnd cell_6t
Xbit_r25_c69 bl_69 br_69 wl_25 vdd gnd cell_6t
Xbit_r26_c69 bl_69 br_69 wl_26 vdd gnd cell_6t
Xbit_r27_c69 bl_69 br_69 wl_27 vdd gnd cell_6t
Xbit_r28_c69 bl_69 br_69 wl_28 vdd gnd cell_6t
Xbit_r29_c69 bl_69 br_69 wl_29 vdd gnd cell_6t
Xbit_r30_c69 bl_69 br_69 wl_30 vdd gnd cell_6t
Xbit_r31_c69 bl_69 br_69 wl_31 vdd gnd cell_6t
Xbit_r32_c69 bl_69 br_69 wl_32 vdd gnd cell_6t
Xbit_r33_c69 bl_69 br_69 wl_33 vdd gnd cell_6t
Xbit_r34_c69 bl_69 br_69 wl_34 vdd gnd cell_6t
Xbit_r35_c69 bl_69 br_69 wl_35 vdd gnd cell_6t
Xbit_r36_c69 bl_69 br_69 wl_36 vdd gnd cell_6t
Xbit_r37_c69 bl_69 br_69 wl_37 vdd gnd cell_6t
Xbit_r38_c69 bl_69 br_69 wl_38 vdd gnd cell_6t
Xbit_r39_c69 bl_69 br_69 wl_39 vdd gnd cell_6t
Xbit_r40_c69 bl_69 br_69 wl_40 vdd gnd cell_6t
Xbit_r41_c69 bl_69 br_69 wl_41 vdd gnd cell_6t
Xbit_r42_c69 bl_69 br_69 wl_42 vdd gnd cell_6t
Xbit_r43_c69 bl_69 br_69 wl_43 vdd gnd cell_6t
Xbit_r44_c69 bl_69 br_69 wl_44 vdd gnd cell_6t
Xbit_r45_c69 bl_69 br_69 wl_45 vdd gnd cell_6t
Xbit_r46_c69 bl_69 br_69 wl_46 vdd gnd cell_6t
Xbit_r47_c69 bl_69 br_69 wl_47 vdd gnd cell_6t
Xbit_r48_c69 bl_69 br_69 wl_48 vdd gnd cell_6t
Xbit_r49_c69 bl_69 br_69 wl_49 vdd gnd cell_6t
Xbit_r50_c69 bl_69 br_69 wl_50 vdd gnd cell_6t
Xbit_r51_c69 bl_69 br_69 wl_51 vdd gnd cell_6t
Xbit_r52_c69 bl_69 br_69 wl_52 vdd gnd cell_6t
Xbit_r53_c69 bl_69 br_69 wl_53 vdd gnd cell_6t
Xbit_r54_c69 bl_69 br_69 wl_54 vdd gnd cell_6t
Xbit_r55_c69 bl_69 br_69 wl_55 vdd gnd cell_6t
Xbit_r56_c69 bl_69 br_69 wl_56 vdd gnd cell_6t
Xbit_r57_c69 bl_69 br_69 wl_57 vdd gnd cell_6t
Xbit_r58_c69 bl_69 br_69 wl_58 vdd gnd cell_6t
Xbit_r59_c69 bl_69 br_69 wl_59 vdd gnd cell_6t
Xbit_r60_c69 bl_69 br_69 wl_60 vdd gnd cell_6t
Xbit_r61_c69 bl_69 br_69 wl_61 vdd gnd cell_6t
Xbit_r62_c69 bl_69 br_69 wl_62 vdd gnd cell_6t
Xbit_r63_c69 bl_69 br_69 wl_63 vdd gnd cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd cell_6t
Xbit_r1_c70 bl_70 br_70 wl_1 vdd gnd cell_6t
Xbit_r2_c70 bl_70 br_70 wl_2 vdd gnd cell_6t
Xbit_r3_c70 bl_70 br_70 wl_3 vdd gnd cell_6t
Xbit_r4_c70 bl_70 br_70 wl_4 vdd gnd cell_6t
Xbit_r5_c70 bl_70 br_70 wl_5 vdd gnd cell_6t
Xbit_r6_c70 bl_70 br_70 wl_6 vdd gnd cell_6t
Xbit_r7_c70 bl_70 br_70 wl_7 vdd gnd cell_6t
Xbit_r8_c70 bl_70 br_70 wl_8 vdd gnd cell_6t
Xbit_r9_c70 bl_70 br_70 wl_9 vdd gnd cell_6t
Xbit_r10_c70 bl_70 br_70 wl_10 vdd gnd cell_6t
Xbit_r11_c70 bl_70 br_70 wl_11 vdd gnd cell_6t
Xbit_r12_c70 bl_70 br_70 wl_12 vdd gnd cell_6t
Xbit_r13_c70 bl_70 br_70 wl_13 vdd gnd cell_6t
Xbit_r14_c70 bl_70 br_70 wl_14 vdd gnd cell_6t
Xbit_r15_c70 bl_70 br_70 wl_15 vdd gnd cell_6t
Xbit_r16_c70 bl_70 br_70 wl_16 vdd gnd cell_6t
Xbit_r17_c70 bl_70 br_70 wl_17 vdd gnd cell_6t
Xbit_r18_c70 bl_70 br_70 wl_18 vdd gnd cell_6t
Xbit_r19_c70 bl_70 br_70 wl_19 vdd gnd cell_6t
Xbit_r20_c70 bl_70 br_70 wl_20 vdd gnd cell_6t
Xbit_r21_c70 bl_70 br_70 wl_21 vdd gnd cell_6t
Xbit_r22_c70 bl_70 br_70 wl_22 vdd gnd cell_6t
Xbit_r23_c70 bl_70 br_70 wl_23 vdd gnd cell_6t
Xbit_r24_c70 bl_70 br_70 wl_24 vdd gnd cell_6t
Xbit_r25_c70 bl_70 br_70 wl_25 vdd gnd cell_6t
Xbit_r26_c70 bl_70 br_70 wl_26 vdd gnd cell_6t
Xbit_r27_c70 bl_70 br_70 wl_27 vdd gnd cell_6t
Xbit_r28_c70 bl_70 br_70 wl_28 vdd gnd cell_6t
Xbit_r29_c70 bl_70 br_70 wl_29 vdd gnd cell_6t
Xbit_r30_c70 bl_70 br_70 wl_30 vdd gnd cell_6t
Xbit_r31_c70 bl_70 br_70 wl_31 vdd gnd cell_6t
Xbit_r32_c70 bl_70 br_70 wl_32 vdd gnd cell_6t
Xbit_r33_c70 bl_70 br_70 wl_33 vdd gnd cell_6t
Xbit_r34_c70 bl_70 br_70 wl_34 vdd gnd cell_6t
Xbit_r35_c70 bl_70 br_70 wl_35 vdd gnd cell_6t
Xbit_r36_c70 bl_70 br_70 wl_36 vdd gnd cell_6t
Xbit_r37_c70 bl_70 br_70 wl_37 vdd gnd cell_6t
Xbit_r38_c70 bl_70 br_70 wl_38 vdd gnd cell_6t
Xbit_r39_c70 bl_70 br_70 wl_39 vdd gnd cell_6t
Xbit_r40_c70 bl_70 br_70 wl_40 vdd gnd cell_6t
Xbit_r41_c70 bl_70 br_70 wl_41 vdd gnd cell_6t
Xbit_r42_c70 bl_70 br_70 wl_42 vdd gnd cell_6t
Xbit_r43_c70 bl_70 br_70 wl_43 vdd gnd cell_6t
Xbit_r44_c70 bl_70 br_70 wl_44 vdd gnd cell_6t
Xbit_r45_c70 bl_70 br_70 wl_45 vdd gnd cell_6t
Xbit_r46_c70 bl_70 br_70 wl_46 vdd gnd cell_6t
Xbit_r47_c70 bl_70 br_70 wl_47 vdd gnd cell_6t
Xbit_r48_c70 bl_70 br_70 wl_48 vdd gnd cell_6t
Xbit_r49_c70 bl_70 br_70 wl_49 vdd gnd cell_6t
Xbit_r50_c70 bl_70 br_70 wl_50 vdd gnd cell_6t
Xbit_r51_c70 bl_70 br_70 wl_51 vdd gnd cell_6t
Xbit_r52_c70 bl_70 br_70 wl_52 vdd gnd cell_6t
Xbit_r53_c70 bl_70 br_70 wl_53 vdd gnd cell_6t
Xbit_r54_c70 bl_70 br_70 wl_54 vdd gnd cell_6t
Xbit_r55_c70 bl_70 br_70 wl_55 vdd gnd cell_6t
Xbit_r56_c70 bl_70 br_70 wl_56 vdd gnd cell_6t
Xbit_r57_c70 bl_70 br_70 wl_57 vdd gnd cell_6t
Xbit_r58_c70 bl_70 br_70 wl_58 vdd gnd cell_6t
Xbit_r59_c70 bl_70 br_70 wl_59 vdd gnd cell_6t
Xbit_r60_c70 bl_70 br_70 wl_60 vdd gnd cell_6t
Xbit_r61_c70 bl_70 br_70 wl_61 vdd gnd cell_6t
Xbit_r62_c70 bl_70 br_70 wl_62 vdd gnd cell_6t
Xbit_r63_c70 bl_70 br_70 wl_63 vdd gnd cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd cell_6t
Xbit_r1_c71 bl_71 br_71 wl_1 vdd gnd cell_6t
Xbit_r2_c71 bl_71 br_71 wl_2 vdd gnd cell_6t
Xbit_r3_c71 bl_71 br_71 wl_3 vdd gnd cell_6t
Xbit_r4_c71 bl_71 br_71 wl_4 vdd gnd cell_6t
Xbit_r5_c71 bl_71 br_71 wl_5 vdd gnd cell_6t
Xbit_r6_c71 bl_71 br_71 wl_6 vdd gnd cell_6t
Xbit_r7_c71 bl_71 br_71 wl_7 vdd gnd cell_6t
Xbit_r8_c71 bl_71 br_71 wl_8 vdd gnd cell_6t
Xbit_r9_c71 bl_71 br_71 wl_9 vdd gnd cell_6t
Xbit_r10_c71 bl_71 br_71 wl_10 vdd gnd cell_6t
Xbit_r11_c71 bl_71 br_71 wl_11 vdd gnd cell_6t
Xbit_r12_c71 bl_71 br_71 wl_12 vdd gnd cell_6t
Xbit_r13_c71 bl_71 br_71 wl_13 vdd gnd cell_6t
Xbit_r14_c71 bl_71 br_71 wl_14 vdd gnd cell_6t
Xbit_r15_c71 bl_71 br_71 wl_15 vdd gnd cell_6t
Xbit_r16_c71 bl_71 br_71 wl_16 vdd gnd cell_6t
Xbit_r17_c71 bl_71 br_71 wl_17 vdd gnd cell_6t
Xbit_r18_c71 bl_71 br_71 wl_18 vdd gnd cell_6t
Xbit_r19_c71 bl_71 br_71 wl_19 vdd gnd cell_6t
Xbit_r20_c71 bl_71 br_71 wl_20 vdd gnd cell_6t
Xbit_r21_c71 bl_71 br_71 wl_21 vdd gnd cell_6t
Xbit_r22_c71 bl_71 br_71 wl_22 vdd gnd cell_6t
Xbit_r23_c71 bl_71 br_71 wl_23 vdd gnd cell_6t
Xbit_r24_c71 bl_71 br_71 wl_24 vdd gnd cell_6t
Xbit_r25_c71 bl_71 br_71 wl_25 vdd gnd cell_6t
Xbit_r26_c71 bl_71 br_71 wl_26 vdd gnd cell_6t
Xbit_r27_c71 bl_71 br_71 wl_27 vdd gnd cell_6t
Xbit_r28_c71 bl_71 br_71 wl_28 vdd gnd cell_6t
Xbit_r29_c71 bl_71 br_71 wl_29 vdd gnd cell_6t
Xbit_r30_c71 bl_71 br_71 wl_30 vdd gnd cell_6t
Xbit_r31_c71 bl_71 br_71 wl_31 vdd gnd cell_6t
Xbit_r32_c71 bl_71 br_71 wl_32 vdd gnd cell_6t
Xbit_r33_c71 bl_71 br_71 wl_33 vdd gnd cell_6t
Xbit_r34_c71 bl_71 br_71 wl_34 vdd gnd cell_6t
Xbit_r35_c71 bl_71 br_71 wl_35 vdd gnd cell_6t
Xbit_r36_c71 bl_71 br_71 wl_36 vdd gnd cell_6t
Xbit_r37_c71 bl_71 br_71 wl_37 vdd gnd cell_6t
Xbit_r38_c71 bl_71 br_71 wl_38 vdd gnd cell_6t
Xbit_r39_c71 bl_71 br_71 wl_39 vdd gnd cell_6t
Xbit_r40_c71 bl_71 br_71 wl_40 vdd gnd cell_6t
Xbit_r41_c71 bl_71 br_71 wl_41 vdd gnd cell_6t
Xbit_r42_c71 bl_71 br_71 wl_42 vdd gnd cell_6t
Xbit_r43_c71 bl_71 br_71 wl_43 vdd gnd cell_6t
Xbit_r44_c71 bl_71 br_71 wl_44 vdd gnd cell_6t
Xbit_r45_c71 bl_71 br_71 wl_45 vdd gnd cell_6t
Xbit_r46_c71 bl_71 br_71 wl_46 vdd gnd cell_6t
Xbit_r47_c71 bl_71 br_71 wl_47 vdd gnd cell_6t
Xbit_r48_c71 bl_71 br_71 wl_48 vdd gnd cell_6t
Xbit_r49_c71 bl_71 br_71 wl_49 vdd gnd cell_6t
Xbit_r50_c71 bl_71 br_71 wl_50 vdd gnd cell_6t
Xbit_r51_c71 bl_71 br_71 wl_51 vdd gnd cell_6t
Xbit_r52_c71 bl_71 br_71 wl_52 vdd gnd cell_6t
Xbit_r53_c71 bl_71 br_71 wl_53 vdd gnd cell_6t
Xbit_r54_c71 bl_71 br_71 wl_54 vdd gnd cell_6t
Xbit_r55_c71 bl_71 br_71 wl_55 vdd gnd cell_6t
Xbit_r56_c71 bl_71 br_71 wl_56 vdd gnd cell_6t
Xbit_r57_c71 bl_71 br_71 wl_57 vdd gnd cell_6t
Xbit_r58_c71 bl_71 br_71 wl_58 vdd gnd cell_6t
Xbit_r59_c71 bl_71 br_71 wl_59 vdd gnd cell_6t
Xbit_r60_c71 bl_71 br_71 wl_60 vdd gnd cell_6t
Xbit_r61_c71 bl_71 br_71 wl_61 vdd gnd cell_6t
Xbit_r62_c71 bl_71 br_71 wl_62 vdd gnd cell_6t
Xbit_r63_c71 bl_71 br_71 wl_63 vdd gnd cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd cell_6t
Xbit_r1_c72 bl_72 br_72 wl_1 vdd gnd cell_6t
Xbit_r2_c72 bl_72 br_72 wl_2 vdd gnd cell_6t
Xbit_r3_c72 bl_72 br_72 wl_3 vdd gnd cell_6t
Xbit_r4_c72 bl_72 br_72 wl_4 vdd gnd cell_6t
Xbit_r5_c72 bl_72 br_72 wl_5 vdd gnd cell_6t
Xbit_r6_c72 bl_72 br_72 wl_6 vdd gnd cell_6t
Xbit_r7_c72 bl_72 br_72 wl_7 vdd gnd cell_6t
Xbit_r8_c72 bl_72 br_72 wl_8 vdd gnd cell_6t
Xbit_r9_c72 bl_72 br_72 wl_9 vdd gnd cell_6t
Xbit_r10_c72 bl_72 br_72 wl_10 vdd gnd cell_6t
Xbit_r11_c72 bl_72 br_72 wl_11 vdd gnd cell_6t
Xbit_r12_c72 bl_72 br_72 wl_12 vdd gnd cell_6t
Xbit_r13_c72 bl_72 br_72 wl_13 vdd gnd cell_6t
Xbit_r14_c72 bl_72 br_72 wl_14 vdd gnd cell_6t
Xbit_r15_c72 bl_72 br_72 wl_15 vdd gnd cell_6t
Xbit_r16_c72 bl_72 br_72 wl_16 vdd gnd cell_6t
Xbit_r17_c72 bl_72 br_72 wl_17 vdd gnd cell_6t
Xbit_r18_c72 bl_72 br_72 wl_18 vdd gnd cell_6t
Xbit_r19_c72 bl_72 br_72 wl_19 vdd gnd cell_6t
Xbit_r20_c72 bl_72 br_72 wl_20 vdd gnd cell_6t
Xbit_r21_c72 bl_72 br_72 wl_21 vdd gnd cell_6t
Xbit_r22_c72 bl_72 br_72 wl_22 vdd gnd cell_6t
Xbit_r23_c72 bl_72 br_72 wl_23 vdd gnd cell_6t
Xbit_r24_c72 bl_72 br_72 wl_24 vdd gnd cell_6t
Xbit_r25_c72 bl_72 br_72 wl_25 vdd gnd cell_6t
Xbit_r26_c72 bl_72 br_72 wl_26 vdd gnd cell_6t
Xbit_r27_c72 bl_72 br_72 wl_27 vdd gnd cell_6t
Xbit_r28_c72 bl_72 br_72 wl_28 vdd gnd cell_6t
Xbit_r29_c72 bl_72 br_72 wl_29 vdd gnd cell_6t
Xbit_r30_c72 bl_72 br_72 wl_30 vdd gnd cell_6t
Xbit_r31_c72 bl_72 br_72 wl_31 vdd gnd cell_6t
Xbit_r32_c72 bl_72 br_72 wl_32 vdd gnd cell_6t
Xbit_r33_c72 bl_72 br_72 wl_33 vdd gnd cell_6t
Xbit_r34_c72 bl_72 br_72 wl_34 vdd gnd cell_6t
Xbit_r35_c72 bl_72 br_72 wl_35 vdd gnd cell_6t
Xbit_r36_c72 bl_72 br_72 wl_36 vdd gnd cell_6t
Xbit_r37_c72 bl_72 br_72 wl_37 vdd gnd cell_6t
Xbit_r38_c72 bl_72 br_72 wl_38 vdd gnd cell_6t
Xbit_r39_c72 bl_72 br_72 wl_39 vdd gnd cell_6t
Xbit_r40_c72 bl_72 br_72 wl_40 vdd gnd cell_6t
Xbit_r41_c72 bl_72 br_72 wl_41 vdd gnd cell_6t
Xbit_r42_c72 bl_72 br_72 wl_42 vdd gnd cell_6t
Xbit_r43_c72 bl_72 br_72 wl_43 vdd gnd cell_6t
Xbit_r44_c72 bl_72 br_72 wl_44 vdd gnd cell_6t
Xbit_r45_c72 bl_72 br_72 wl_45 vdd gnd cell_6t
Xbit_r46_c72 bl_72 br_72 wl_46 vdd gnd cell_6t
Xbit_r47_c72 bl_72 br_72 wl_47 vdd gnd cell_6t
Xbit_r48_c72 bl_72 br_72 wl_48 vdd gnd cell_6t
Xbit_r49_c72 bl_72 br_72 wl_49 vdd gnd cell_6t
Xbit_r50_c72 bl_72 br_72 wl_50 vdd gnd cell_6t
Xbit_r51_c72 bl_72 br_72 wl_51 vdd gnd cell_6t
Xbit_r52_c72 bl_72 br_72 wl_52 vdd gnd cell_6t
Xbit_r53_c72 bl_72 br_72 wl_53 vdd gnd cell_6t
Xbit_r54_c72 bl_72 br_72 wl_54 vdd gnd cell_6t
Xbit_r55_c72 bl_72 br_72 wl_55 vdd gnd cell_6t
Xbit_r56_c72 bl_72 br_72 wl_56 vdd gnd cell_6t
Xbit_r57_c72 bl_72 br_72 wl_57 vdd gnd cell_6t
Xbit_r58_c72 bl_72 br_72 wl_58 vdd gnd cell_6t
Xbit_r59_c72 bl_72 br_72 wl_59 vdd gnd cell_6t
Xbit_r60_c72 bl_72 br_72 wl_60 vdd gnd cell_6t
Xbit_r61_c72 bl_72 br_72 wl_61 vdd gnd cell_6t
Xbit_r62_c72 bl_72 br_72 wl_62 vdd gnd cell_6t
Xbit_r63_c72 bl_72 br_72 wl_63 vdd gnd cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd cell_6t
Xbit_r1_c73 bl_73 br_73 wl_1 vdd gnd cell_6t
Xbit_r2_c73 bl_73 br_73 wl_2 vdd gnd cell_6t
Xbit_r3_c73 bl_73 br_73 wl_3 vdd gnd cell_6t
Xbit_r4_c73 bl_73 br_73 wl_4 vdd gnd cell_6t
Xbit_r5_c73 bl_73 br_73 wl_5 vdd gnd cell_6t
Xbit_r6_c73 bl_73 br_73 wl_6 vdd gnd cell_6t
Xbit_r7_c73 bl_73 br_73 wl_7 vdd gnd cell_6t
Xbit_r8_c73 bl_73 br_73 wl_8 vdd gnd cell_6t
Xbit_r9_c73 bl_73 br_73 wl_9 vdd gnd cell_6t
Xbit_r10_c73 bl_73 br_73 wl_10 vdd gnd cell_6t
Xbit_r11_c73 bl_73 br_73 wl_11 vdd gnd cell_6t
Xbit_r12_c73 bl_73 br_73 wl_12 vdd gnd cell_6t
Xbit_r13_c73 bl_73 br_73 wl_13 vdd gnd cell_6t
Xbit_r14_c73 bl_73 br_73 wl_14 vdd gnd cell_6t
Xbit_r15_c73 bl_73 br_73 wl_15 vdd gnd cell_6t
Xbit_r16_c73 bl_73 br_73 wl_16 vdd gnd cell_6t
Xbit_r17_c73 bl_73 br_73 wl_17 vdd gnd cell_6t
Xbit_r18_c73 bl_73 br_73 wl_18 vdd gnd cell_6t
Xbit_r19_c73 bl_73 br_73 wl_19 vdd gnd cell_6t
Xbit_r20_c73 bl_73 br_73 wl_20 vdd gnd cell_6t
Xbit_r21_c73 bl_73 br_73 wl_21 vdd gnd cell_6t
Xbit_r22_c73 bl_73 br_73 wl_22 vdd gnd cell_6t
Xbit_r23_c73 bl_73 br_73 wl_23 vdd gnd cell_6t
Xbit_r24_c73 bl_73 br_73 wl_24 vdd gnd cell_6t
Xbit_r25_c73 bl_73 br_73 wl_25 vdd gnd cell_6t
Xbit_r26_c73 bl_73 br_73 wl_26 vdd gnd cell_6t
Xbit_r27_c73 bl_73 br_73 wl_27 vdd gnd cell_6t
Xbit_r28_c73 bl_73 br_73 wl_28 vdd gnd cell_6t
Xbit_r29_c73 bl_73 br_73 wl_29 vdd gnd cell_6t
Xbit_r30_c73 bl_73 br_73 wl_30 vdd gnd cell_6t
Xbit_r31_c73 bl_73 br_73 wl_31 vdd gnd cell_6t
Xbit_r32_c73 bl_73 br_73 wl_32 vdd gnd cell_6t
Xbit_r33_c73 bl_73 br_73 wl_33 vdd gnd cell_6t
Xbit_r34_c73 bl_73 br_73 wl_34 vdd gnd cell_6t
Xbit_r35_c73 bl_73 br_73 wl_35 vdd gnd cell_6t
Xbit_r36_c73 bl_73 br_73 wl_36 vdd gnd cell_6t
Xbit_r37_c73 bl_73 br_73 wl_37 vdd gnd cell_6t
Xbit_r38_c73 bl_73 br_73 wl_38 vdd gnd cell_6t
Xbit_r39_c73 bl_73 br_73 wl_39 vdd gnd cell_6t
Xbit_r40_c73 bl_73 br_73 wl_40 vdd gnd cell_6t
Xbit_r41_c73 bl_73 br_73 wl_41 vdd gnd cell_6t
Xbit_r42_c73 bl_73 br_73 wl_42 vdd gnd cell_6t
Xbit_r43_c73 bl_73 br_73 wl_43 vdd gnd cell_6t
Xbit_r44_c73 bl_73 br_73 wl_44 vdd gnd cell_6t
Xbit_r45_c73 bl_73 br_73 wl_45 vdd gnd cell_6t
Xbit_r46_c73 bl_73 br_73 wl_46 vdd gnd cell_6t
Xbit_r47_c73 bl_73 br_73 wl_47 vdd gnd cell_6t
Xbit_r48_c73 bl_73 br_73 wl_48 vdd gnd cell_6t
Xbit_r49_c73 bl_73 br_73 wl_49 vdd gnd cell_6t
Xbit_r50_c73 bl_73 br_73 wl_50 vdd gnd cell_6t
Xbit_r51_c73 bl_73 br_73 wl_51 vdd gnd cell_6t
Xbit_r52_c73 bl_73 br_73 wl_52 vdd gnd cell_6t
Xbit_r53_c73 bl_73 br_73 wl_53 vdd gnd cell_6t
Xbit_r54_c73 bl_73 br_73 wl_54 vdd gnd cell_6t
Xbit_r55_c73 bl_73 br_73 wl_55 vdd gnd cell_6t
Xbit_r56_c73 bl_73 br_73 wl_56 vdd gnd cell_6t
Xbit_r57_c73 bl_73 br_73 wl_57 vdd gnd cell_6t
Xbit_r58_c73 bl_73 br_73 wl_58 vdd gnd cell_6t
Xbit_r59_c73 bl_73 br_73 wl_59 vdd gnd cell_6t
Xbit_r60_c73 bl_73 br_73 wl_60 vdd gnd cell_6t
Xbit_r61_c73 bl_73 br_73 wl_61 vdd gnd cell_6t
Xbit_r62_c73 bl_73 br_73 wl_62 vdd gnd cell_6t
Xbit_r63_c73 bl_73 br_73 wl_63 vdd gnd cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd cell_6t
Xbit_r1_c74 bl_74 br_74 wl_1 vdd gnd cell_6t
Xbit_r2_c74 bl_74 br_74 wl_2 vdd gnd cell_6t
Xbit_r3_c74 bl_74 br_74 wl_3 vdd gnd cell_6t
Xbit_r4_c74 bl_74 br_74 wl_4 vdd gnd cell_6t
Xbit_r5_c74 bl_74 br_74 wl_5 vdd gnd cell_6t
Xbit_r6_c74 bl_74 br_74 wl_6 vdd gnd cell_6t
Xbit_r7_c74 bl_74 br_74 wl_7 vdd gnd cell_6t
Xbit_r8_c74 bl_74 br_74 wl_8 vdd gnd cell_6t
Xbit_r9_c74 bl_74 br_74 wl_9 vdd gnd cell_6t
Xbit_r10_c74 bl_74 br_74 wl_10 vdd gnd cell_6t
Xbit_r11_c74 bl_74 br_74 wl_11 vdd gnd cell_6t
Xbit_r12_c74 bl_74 br_74 wl_12 vdd gnd cell_6t
Xbit_r13_c74 bl_74 br_74 wl_13 vdd gnd cell_6t
Xbit_r14_c74 bl_74 br_74 wl_14 vdd gnd cell_6t
Xbit_r15_c74 bl_74 br_74 wl_15 vdd gnd cell_6t
Xbit_r16_c74 bl_74 br_74 wl_16 vdd gnd cell_6t
Xbit_r17_c74 bl_74 br_74 wl_17 vdd gnd cell_6t
Xbit_r18_c74 bl_74 br_74 wl_18 vdd gnd cell_6t
Xbit_r19_c74 bl_74 br_74 wl_19 vdd gnd cell_6t
Xbit_r20_c74 bl_74 br_74 wl_20 vdd gnd cell_6t
Xbit_r21_c74 bl_74 br_74 wl_21 vdd gnd cell_6t
Xbit_r22_c74 bl_74 br_74 wl_22 vdd gnd cell_6t
Xbit_r23_c74 bl_74 br_74 wl_23 vdd gnd cell_6t
Xbit_r24_c74 bl_74 br_74 wl_24 vdd gnd cell_6t
Xbit_r25_c74 bl_74 br_74 wl_25 vdd gnd cell_6t
Xbit_r26_c74 bl_74 br_74 wl_26 vdd gnd cell_6t
Xbit_r27_c74 bl_74 br_74 wl_27 vdd gnd cell_6t
Xbit_r28_c74 bl_74 br_74 wl_28 vdd gnd cell_6t
Xbit_r29_c74 bl_74 br_74 wl_29 vdd gnd cell_6t
Xbit_r30_c74 bl_74 br_74 wl_30 vdd gnd cell_6t
Xbit_r31_c74 bl_74 br_74 wl_31 vdd gnd cell_6t
Xbit_r32_c74 bl_74 br_74 wl_32 vdd gnd cell_6t
Xbit_r33_c74 bl_74 br_74 wl_33 vdd gnd cell_6t
Xbit_r34_c74 bl_74 br_74 wl_34 vdd gnd cell_6t
Xbit_r35_c74 bl_74 br_74 wl_35 vdd gnd cell_6t
Xbit_r36_c74 bl_74 br_74 wl_36 vdd gnd cell_6t
Xbit_r37_c74 bl_74 br_74 wl_37 vdd gnd cell_6t
Xbit_r38_c74 bl_74 br_74 wl_38 vdd gnd cell_6t
Xbit_r39_c74 bl_74 br_74 wl_39 vdd gnd cell_6t
Xbit_r40_c74 bl_74 br_74 wl_40 vdd gnd cell_6t
Xbit_r41_c74 bl_74 br_74 wl_41 vdd gnd cell_6t
Xbit_r42_c74 bl_74 br_74 wl_42 vdd gnd cell_6t
Xbit_r43_c74 bl_74 br_74 wl_43 vdd gnd cell_6t
Xbit_r44_c74 bl_74 br_74 wl_44 vdd gnd cell_6t
Xbit_r45_c74 bl_74 br_74 wl_45 vdd gnd cell_6t
Xbit_r46_c74 bl_74 br_74 wl_46 vdd gnd cell_6t
Xbit_r47_c74 bl_74 br_74 wl_47 vdd gnd cell_6t
Xbit_r48_c74 bl_74 br_74 wl_48 vdd gnd cell_6t
Xbit_r49_c74 bl_74 br_74 wl_49 vdd gnd cell_6t
Xbit_r50_c74 bl_74 br_74 wl_50 vdd gnd cell_6t
Xbit_r51_c74 bl_74 br_74 wl_51 vdd gnd cell_6t
Xbit_r52_c74 bl_74 br_74 wl_52 vdd gnd cell_6t
Xbit_r53_c74 bl_74 br_74 wl_53 vdd gnd cell_6t
Xbit_r54_c74 bl_74 br_74 wl_54 vdd gnd cell_6t
Xbit_r55_c74 bl_74 br_74 wl_55 vdd gnd cell_6t
Xbit_r56_c74 bl_74 br_74 wl_56 vdd gnd cell_6t
Xbit_r57_c74 bl_74 br_74 wl_57 vdd gnd cell_6t
Xbit_r58_c74 bl_74 br_74 wl_58 vdd gnd cell_6t
Xbit_r59_c74 bl_74 br_74 wl_59 vdd gnd cell_6t
Xbit_r60_c74 bl_74 br_74 wl_60 vdd gnd cell_6t
Xbit_r61_c74 bl_74 br_74 wl_61 vdd gnd cell_6t
Xbit_r62_c74 bl_74 br_74 wl_62 vdd gnd cell_6t
Xbit_r63_c74 bl_74 br_74 wl_63 vdd gnd cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd cell_6t
Xbit_r1_c75 bl_75 br_75 wl_1 vdd gnd cell_6t
Xbit_r2_c75 bl_75 br_75 wl_2 vdd gnd cell_6t
Xbit_r3_c75 bl_75 br_75 wl_3 vdd gnd cell_6t
Xbit_r4_c75 bl_75 br_75 wl_4 vdd gnd cell_6t
Xbit_r5_c75 bl_75 br_75 wl_5 vdd gnd cell_6t
Xbit_r6_c75 bl_75 br_75 wl_6 vdd gnd cell_6t
Xbit_r7_c75 bl_75 br_75 wl_7 vdd gnd cell_6t
Xbit_r8_c75 bl_75 br_75 wl_8 vdd gnd cell_6t
Xbit_r9_c75 bl_75 br_75 wl_9 vdd gnd cell_6t
Xbit_r10_c75 bl_75 br_75 wl_10 vdd gnd cell_6t
Xbit_r11_c75 bl_75 br_75 wl_11 vdd gnd cell_6t
Xbit_r12_c75 bl_75 br_75 wl_12 vdd gnd cell_6t
Xbit_r13_c75 bl_75 br_75 wl_13 vdd gnd cell_6t
Xbit_r14_c75 bl_75 br_75 wl_14 vdd gnd cell_6t
Xbit_r15_c75 bl_75 br_75 wl_15 vdd gnd cell_6t
Xbit_r16_c75 bl_75 br_75 wl_16 vdd gnd cell_6t
Xbit_r17_c75 bl_75 br_75 wl_17 vdd gnd cell_6t
Xbit_r18_c75 bl_75 br_75 wl_18 vdd gnd cell_6t
Xbit_r19_c75 bl_75 br_75 wl_19 vdd gnd cell_6t
Xbit_r20_c75 bl_75 br_75 wl_20 vdd gnd cell_6t
Xbit_r21_c75 bl_75 br_75 wl_21 vdd gnd cell_6t
Xbit_r22_c75 bl_75 br_75 wl_22 vdd gnd cell_6t
Xbit_r23_c75 bl_75 br_75 wl_23 vdd gnd cell_6t
Xbit_r24_c75 bl_75 br_75 wl_24 vdd gnd cell_6t
Xbit_r25_c75 bl_75 br_75 wl_25 vdd gnd cell_6t
Xbit_r26_c75 bl_75 br_75 wl_26 vdd gnd cell_6t
Xbit_r27_c75 bl_75 br_75 wl_27 vdd gnd cell_6t
Xbit_r28_c75 bl_75 br_75 wl_28 vdd gnd cell_6t
Xbit_r29_c75 bl_75 br_75 wl_29 vdd gnd cell_6t
Xbit_r30_c75 bl_75 br_75 wl_30 vdd gnd cell_6t
Xbit_r31_c75 bl_75 br_75 wl_31 vdd gnd cell_6t
Xbit_r32_c75 bl_75 br_75 wl_32 vdd gnd cell_6t
Xbit_r33_c75 bl_75 br_75 wl_33 vdd gnd cell_6t
Xbit_r34_c75 bl_75 br_75 wl_34 vdd gnd cell_6t
Xbit_r35_c75 bl_75 br_75 wl_35 vdd gnd cell_6t
Xbit_r36_c75 bl_75 br_75 wl_36 vdd gnd cell_6t
Xbit_r37_c75 bl_75 br_75 wl_37 vdd gnd cell_6t
Xbit_r38_c75 bl_75 br_75 wl_38 vdd gnd cell_6t
Xbit_r39_c75 bl_75 br_75 wl_39 vdd gnd cell_6t
Xbit_r40_c75 bl_75 br_75 wl_40 vdd gnd cell_6t
Xbit_r41_c75 bl_75 br_75 wl_41 vdd gnd cell_6t
Xbit_r42_c75 bl_75 br_75 wl_42 vdd gnd cell_6t
Xbit_r43_c75 bl_75 br_75 wl_43 vdd gnd cell_6t
Xbit_r44_c75 bl_75 br_75 wl_44 vdd gnd cell_6t
Xbit_r45_c75 bl_75 br_75 wl_45 vdd gnd cell_6t
Xbit_r46_c75 bl_75 br_75 wl_46 vdd gnd cell_6t
Xbit_r47_c75 bl_75 br_75 wl_47 vdd gnd cell_6t
Xbit_r48_c75 bl_75 br_75 wl_48 vdd gnd cell_6t
Xbit_r49_c75 bl_75 br_75 wl_49 vdd gnd cell_6t
Xbit_r50_c75 bl_75 br_75 wl_50 vdd gnd cell_6t
Xbit_r51_c75 bl_75 br_75 wl_51 vdd gnd cell_6t
Xbit_r52_c75 bl_75 br_75 wl_52 vdd gnd cell_6t
Xbit_r53_c75 bl_75 br_75 wl_53 vdd gnd cell_6t
Xbit_r54_c75 bl_75 br_75 wl_54 vdd gnd cell_6t
Xbit_r55_c75 bl_75 br_75 wl_55 vdd gnd cell_6t
Xbit_r56_c75 bl_75 br_75 wl_56 vdd gnd cell_6t
Xbit_r57_c75 bl_75 br_75 wl_57 vdd gnd cell_6t
Xbit_r58_c75 bl_75 br_75 wl_58 vdd gnd cell_6t
Xbit_r59_c75 bl_75 br_75 wl_59 vdd gnd cell_6t
Xbit_r60_c75 bl_75 br_75 wl_60 vdd gnd cell_6t
Xbit_r61_c75 bl_75 br_75 wl_61 vdd gnd cell_6t
Xbit_r62_c75 bl_75 br_75 wl_62 vdd gnd cell_6t
Xbit_r63_c75 bl_75 br_75 wl_63 vdd gnd cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd cell_6t
Xbit_r1_c76 bl_76 br_76 wl_1 vdd gnd cell_6t
Xbit_r2_c76 bl_76 br_76 wl_2 vdd gnd cell_6t
Xbit_r3_c76 bl_76 br_76 wl_3 vdd gnd cell_6t
Xbit_r4_c76 bl_76 br_76 wl_4 vdd gnd cell_6t
Xbit_r5_c76 bl_76 br_76 wl_5 vdd gnd cell_6t
Xbit_r6_c76 bl_76 br_76 wl_6 vdd gnd cell_6t
Xbit_r7_c76 bl_76 br_76 wl_7 vdd gnd cell_6t
Xbit_r8_c76 bl_76 br_76 wl_8 vdd gnd cell_6t
Xbit_r9_c76 bl_76 br_76 wl_9 vdd gnd cell_6t
Xbit_r10_c76 bl_76 br_76 wl_10 vdd gnd cell_6t
Xbit_r11_c76 bl_76 br_76 wl_11 vdd gnd cell_6t
Xbit_r12_c76 bl_76 br_76 wl_12 vdd gnd cell_6t
Xbit_r13_c76 bl_76 br_76 wl_13 vdd gnd cell_6t
Xbit_r14_c76 bl_76 br_76 wl_14 vdd gnd cell_6t
Xbit_r15_c76 bl_76 br_76 wl_15 vdd gnd cell_6t
Xbit_r16_c76 bl_76 br_76 wl_16 vdd gnd cell_6t
Xbit_r17_c76 bl_76 br_76 wl_17 vdd gnd cell_6t
Xbit_r18_c76 bl_76 br_76 wl_18 vdd gnd cell_6t
Xbit_r19_c76 bl_76 br_76 wl_19 vdd gnd cell_6t
Xbit_r20_c76 bl_76 br_76 wl_20 vdd gnd cell_6t
Xbit_r21_c76 bl_76 br_76 wl_21 vdd gnd cell_6t
Xbit_r22_c76 bl_76 br_76 wl_22 vdd gnd cell_6t
Xbit_r23_c76 bl_76 br_76 wl_23 vdd gnd cell_6t
Xbit_r24_c76 bl_76 br_76 wl_24 vdd gnd cell_6t
Xbit_r25_c76 bl_76 br_76 wl_25 vdd gnd cell_6t
Xbit_r26_c76 bl_76 br_76 wl_26 vdd gnd cell_6t
Xbit_r27_c76 bl_76 br_76 wl_27 vdd gnd cell_6t
Xbit_r28_c76 bl_76 br_76 wl_28 vdd gnd cell_6t
Xbit_r29_c76 bl_76 br_76 wl_29 vdd gnd cell_6t
Xbit_r30_c76 bl_76 br_76 wl_30 vdd gnd cell_6t
Xbit_r31_c76 bl_76 br_76 wl_31 vdd gnd cell_6t
Xbit_r32_c76 bl_76 br_76 wl_32 vdd gnd cell_6t
Xbit_r33_c76 bl_76 br_76 wl_33 vdd gnd cell_6t
Xbit_r34_c76 bl_76 br_76 wl_34 vdd gnd cell_6t
Xbit_r35_c76 bl_76 br_76 wl_35 vdd gnd cell_6t
Xbit_r36_c76 bl_76 br_76 wl_36 vdd gnd cell_6t
Xbit_r37_c76 bl_76 br_76 wl_37 vdd gnd cell_6t
Xbit_r38_c76 bl_76 br_76 wl_38 vdd gnd cell_6t
Xbit_r39_c76 bl_76 br_76 wl_39 vdd gnd cell_6t
Xbit_r40_c76 bl_76 br_76 wl_40 vdd gnd cell_6t
Xbit_r41_c76 bl_76 br_76 wl_41 vdd gnd cell_6t
Xbit_r42_c76 bl_76 br_76 wl_42 vdd gnd cell_6t
Xbit_r43_c76 bl_76 br_76 wl_43 vdd gnd cell_6t
Xbit_r44_c76 bl_76 br_76 wl_44 vdd gnd cell_6t
Xbit_r45_c76 bl_76 br_76 wl_45 vdd gnd cell_6t
Xbit_r46_c76 bl_76 br_76 wl_46 vdd gnd cell_6t
Xbit_r47_c76 bl_76 br_76 wl_47 vdd gnd cell_6t
Xbit_r48_c76 bl_76 br_76 wl_48 vdd gnd cell_6t
Xbit_r49_c76 bl_76 br_76 wl_49 vdd gnd cell_6t
Xbit_r50_c76 bl_76 br_76 wl_50 vdd gnd cell_6t
Xbit_r51_c76 bl_76 br_76 wl_51 vdd gnd cell_6t
Xbit_r52_c76 bl_76 br_76 wl_52 vdd gnd cell_6t
Xbit_r53_c76 bl_76 br_76 wl_53 vdd gnd cell_6t
Xbit_r54_c76 bl_76 br_76 wl_54 vdd gnd cell_6t
Xbit_r55_c76 bl_76 br_76 wl_55 vdd gnd cell_6t
Xbit_r56_c76 bl_76 br_76 wl_56 vdd gnd cell_6t
Xbit_r57_c76 bl_76 br_76 wl_57 vdd gnd cell_6t
Xbit_r58_c76 bl_76 br_76 wl_58 vdd gnd cell_6t
Xbit_r59_c76 bl_76 br_76 wl_59 vdd gnd cell_6t
Xbit_r60_c76 bl_76 br_76 wl_60 vdd gnd cell_6t
Xbit_r61_c76 bl_76 br_76 wl_61 vdd gnd cell_6t
Xbit_r62_c76 bl_76 br_76 wl_62 vdd gnd cell_6t
Xbit_r63_c76 bl_76 br_76 wl_63 vdd gnd cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd cell_6t
Xbit_r1_c77 bl_77 br_77 wl_1 vdd gnd cell_6t
Xbit_r2_c77 bl_77 br_77 wl_2 vdd gnd cell_6t
Xbit_r3_c77 bl_77 br_77 wl_3 vdd gnd cell_6t
Xbit_r4_c77 bl_77 br_77 wl_4 vdd gnd cell_6t
Xbit_r5_c77 bl_77 br_77 wl_5 vdd gnd cell_6t
Xbit_r6_c77 bl_77 br_77 wl_6 vdd gnd cell_6t
Xbit_r7_c77 bl_77 br_77 wl_7 vdd gnd cell_6t
Xbit_r8_c77 bl_77 br_77 wl_8 vdd gnd cell_6t
Xbit_r9_c77 bl_77 br_77 wl_9 vdd gnd cell_6t
Xbit_r10_c77 bl_77 br_77 wl_10 vdd gnd cell_6t
Xbit_r11_c77 bl_77 br_77 wl_11 vdd gnd cell_6t
Xbit_r12_c77 bl_77 br_77 wl_12 vdd gnd cell_6t
Xbit_r13_c77 bl_77 br_77 wl_13 vdd gnd cell_6t
Xbit_r14_c77 bl_77 br_77 wl_14 vdd gnd cell_6t
Xbit_r15_c77 bl_77 br_77 wl_15 vdd gnd cell_6t
Xbit_r16_c77 bl_77 br_77 wl_16 vdd gnd cell_6t
Xbit_r17_c77 bl_77 br_77 wl_17 vdd gnd cell_6t
Xbit_r18_c77 bl_77 br_77 wl_18 vdd gnd cell_6t
Xbit_r19_c77 bl_77 br_77 wl_19 vdd gnd cell_6t
Xbit_r20_c77 bl_77 br_77 wl_20 vdd gnd cell_6t
Xbit_r21_c77 bl_77 br_77 wl_21 vdd gnd cell_6t
Xbit_r22_c77 bl_77 br_77 wl_22 vdd gnd cell_6t
Xbit_r23_c77 bl_77 br_77 wl_23 vdd gnd cell_6t
Xbit_r24_c77 bl_77 br_77 wl_24 vdd gnd cell_6t
Xbit_r25_c77 bl_77 br_77 wl_25 vdd gnd cell_6t
Xbit_r26_c77 bl_77 br_77 wl_26 vdd gnd cell_6t
Xbit_r27_c77 bl_77 br_77 wl_27 vdd gnd cell_6t
Xbit_r28_c77 bl_77 br_77 wl_28 vdd gnd cell_6t
Xbit_r29_c77 bl_77 br_77 wl_29 vdd gnd cell_6t
Xbit_r30_c77 bl_77 br_77 wl_30 vdd gnd cell_6t
Xbit_r31_c77 bl_77 br_77 wl_31 vdd gnd cell_6t
Xbit_r32_c77 bl_77 br_77 wl_32 vdd gnd cell_6t
Xbit_r33_c77 bl_77 br_77 wl_33 vdd gnd cell_6t
Xbit_r34_c77 bl_77 br_77 wl_34 vdd gnd cell_6t
Xbit_r35_c77 bl_77 br_77 wl_35 vdd gnd cell_6t
Xbit_r36_c77 bl_77 br_77 wl_36 vdd gnd cell_6t
Xbit_r37_c77 bl_77 br_77 wl_37 vdd gnd cell_6t
Xbit_r38_c77 bl_77 br_77 wl_38 vdd gnd cell_6t
Xbit_r39_c77 bl_77 br_77 wl_39 vdd gnd cell_6t
Xbit_r40_c77 bl_77 br_77 wl_40 vdd gnd cell_6t
Xbit_r41_c77 bl_77 br_77 wl_41 vdd gnd cell_6t
Xbit_r42_c77 bl_77 br_77 wl_42 vdd gnd cell_6t
Xbit_r43_c77 bl_77 br_77 wl_43 vdd gnd cell_6t
Xbit_r44_c77 bl_77 br_77 wl_44 vdd gnd cell_6t
Xbit_r45_c77 bl_77 br_77 wl_45 vdd gnd cell_6t
Xbit_r46_c77 bl_77 br_77 wl_46 vdd gnd cell_6t
Xbit_r47_c77 bl_77 br_77 wl_47 vdd gnd cell_6t
Xbit_r48_c77 bl_77 br_77 wl_48 vdd gnd cell_6t
Xbit_r49_c77 bl_77 br_77 wl_49 vdd gnd cell_6t
Xbit_r50_c77 bl_77 br_77 wl_50 vdd gnd cell_6t
Xbit_r51_c77 bl_77 br_77 wl_51 vdd gnd cell_6t
Xbit_r52_c77 bl_77 br_77 wl_52 vdd gnd cell_6t
Xbit_r53_c77 bl_77 br_77 wl_53 vdd gnd cell_6t
Xbit_r54_c77 bl_77 br_77 wl_54 vdd gnd cell_6t
Xbit_r55_c77 bl_77 br_77 wl_55 vdd gnd cell_6t
Xbit_r56_c77 bl_77 br_77 wl_56 vdd gnd cell_6t
Xbit_r57_c77 bl_77 br_77 wl_57 vdd gnd cell_6t
Xbit_r58_c77 bl_77 br_77 wl_58 vdd gnd cell_6t
Xbit_r59_c77 bl_77 br_77 wl_59 vdd gnd cell_6t
Xbit_r60_c77 bl_77 br_77 wl_60 vdd gnd cell_6t
Xbit_r61_c77 bl_77 br_77 wl_61 vdd gnd cell_6t
Xbit_r62_c77 bl_77 br_77 wl_62 vdd gnd cell_6t
Xbit_r63_c77 bl_77 br_77 wl_63 vdd gnd cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd cell_6t
Xbit_r1_c78 bl_78 br_78 wl_1 vdd gnd cell_6t
Xbit_r2_c78 bl_78 br_78 wl_2 vdd gnd cell_6t
Xbit_r3_c78 bl_78 br_78 wl_3 vdd gnd cell_6t
Xbit_r4_c78 bl_78 br_78 wl_4 vdd gnd cell_6t
Xbit_r5_c78 bl_78 br_78 wl_5 vdd gnd cell_6t
Xbit_r6_c78 bl_78 br_78 wl_6 vdd gnd cell_6t
Xbit_r7_c78 bl_78 br_78 wl_7 vdd gnd cell_6t
Xbit_r8_c78 bl_78 br_78 wl_8 vdd gnd cell_6t
Xbit_r9_c78 bl_78 br_78 wl_9 vdd gnd cell_6t
Xbit_r10_c78 bl_78 br_78 wl_10 vdd gnd cell_6t
Xbit_r11_c78 bl_78 br_78 wl_11 vdd gnd cell_6t
Xbit_r12_c78 bl_78 br_78 wl_12 vdd gnd cell_6t
Xbit_r13_c78 bl_78 br_78 wl_13 vdd gnd cell_6t
Xbit_r14_c78 bl_78 br_78 wl_14 vdd gnd cell_6t
Xbit_r15_c78 bl_78 br_78 wl_15 vdd gnd cell_6t
Xbit_r16_c78 bl_78 br_78 wl_16 vdd gnd cell_6t
Xbit_r17_c78 bl_78 br_78 wl_17 vdd gnd cell_6t
Xbit_r18_c78 bl_78 br_78 wl_18 vdd gnd cell_6t
Xbit_r19_c78 bl_78 br_78 wl_19 vdd gnd cell_6t
Xbit_r20_c78 bl_78 br_78 wl_20 vdd gnd cell_6t
Xbit_r21_c78 bl_78 br_78 wl_21 vdd gnd cell_6t
Xbit_r22_c78 bl_78 br_78 wl_22 vdd gnd cell_6t
Xbit_r23_c78 bl_78 br_78 wl_23 vdd gnd cell_6t
Xbit_r24_c78 bl_78 br_78 wl_24 vdd gnd cell_6t
Xbit_r25_c78 bl_78 br_78 wl_25 vdd gnd cell_6t
Xbit_r26_c78 bl_78 br_78 wl_26 vdd gnd cell_6t
Xbit_r27_c78 bl_78 br_78 wl_27 vdd gnd cell_6t
Xbit_r28_c78 bl_78 br_78 wl_28 vdd gnd cell_6t
Xbit_r29_c78 bl_78 br_78 wl_29 vdd gnd cell_6t
Xbit_r30_c78 bl_78 br_78 wl_30 vdd gnd cell_6t
Xbit_r31_c78 bl_78 br_78 wl_31 vdd gnd cell_6t
Xbit_r32_c78 bl_78 br_78 wl_32 vdd gnd cell_6t
Xbit_r33_c78 bl_78 br_78 wl_33 vdd gnd cell_6t
Xbit_r34_c78 bl_78 br_78 wl_34 vdd gnd cell_6t
Xbit_r35_c78 bl_78 br_78 wl_35 vdd gnd cell_6t
Xbit_r36_c78 bl_78 br_78 wl_36 vdd gnd cell_6t
Xbit_r37_c78 bl_78 br_78 wl_37 vdd gnd cell_6t
Xbit_r38_c78 bl_78 br_78 wl_38 vdd gnd cell_6t
Xbit_r39_c78 bl_78 br_78 wl_39 vdd gnd cell_6t
Xbit_r40_c78 bl_78 br_78 wl_40 vdd gnd cell_6t
Xbit_r41_c78 bl_78 br_78 wl_41 vdd gnd cell_6t
Xbit_r42_c78 bl_78 br_78 wl_42 vdd gnd cell_6t
Xbit_r43_c78 bl_78 br_78 wl_43 vdd gnd cell_6t
Xbit_r44_c78 bl_78 br_78 wl_44 vdd gnd cell_6t
Xbit_r45_c78 bl_78 br_78 wl_45 vdd gnd cell_6t
Xbit_r46_c78 bl_78 br_78 wl_46 vdd gnd cell_6t
Xbit_r47_c78 bl_78 br_78 wl_47 vdd gnd cell_6t
Xbit_r48_c78 bl_78 br_78 wl_48 vdd gnd cell_6t
Xbit_r49_c78 bl_78 br_78 wl_49 vdd gnd cell_6t
Xbit_r50_c78 bl_78 br_78 wl_50 vdd gnd cell_6t
Xbit_r51_c78 bl_78 br_78 wl_51 vdd gnd cell_6t
Xbit_r52_c78 bl_78 br_78 wl_52 vdd gnd cell_6t
Xbit_r53_c78 bl_78 br_78 wl_53 vdd gnd cell_6t
Xbit_r54_c78 bl_78 br_78 wl_54 vdd gnd cell_6t
Xbit_r55_c78 bl_78 br_78 wl_55 vdd gnd cell_6t
Xbit_r56_c78 bl_78 br_78 wl_56 vdd gnd cell_6t
Xbit_r57_c78 bl_78 br_78 wl_57 vdd gnd cell_6t
Xbit_r58_c78 bl_78 br_78 wl_58 vdd gnd cell_6t
Xbit_r59_c78 bl_78 br_78 wl_59 vdd gnd cell_6t
Xbit_r60_c78 bl_78 br_78 wl_60 vdd gnd cell_6t
Xbit_r61_c78 bl_78 br_78 wl_61 vdd gnd cell_6t
Xbit_r62_c78 bl_78 br_78 wl_62 vdd gnd cell_6t
Xbit_r63_c78 bl_78 br_78 wl_63 vdd gnd cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd cell_6t
Xbit_r1_c79 bl_79 br_79 wl_1 vdd gnd cell_6t
Xbit_r2_c79 bl_79 br_79 wl_2 vdd gnd cell_6t
Xbit_r3_c79 bl_79 br_79 wl_3 vdd gnd cell_6t
Xbit_r4_c79 bl_79 br_79 wl_4 vdd gnd cell_6t
Xbit_r5_c79 bl_79 br_79 wl_5 vdd gnd cell_6t
Xbit_r6_c79 bl_79 br_79 wl_6 vdd gnd cell_6t
Xbit_r7_c79 bl_79 br_79 wl_7 vdd gnd cell_6t
Xbit_r8_c79 bl_79 br_79 wl_8 vdd gnd cell_6t
Xbit_r9_c79 bl_79 br_79 wl_9 vdd gnd cell_6t
Xbit_r10_c79 bl_79 br_79 wl_10 vdd gnd cell_6t
Xbit_r11_c79 bl_79 br_79 wl_11 vdd gnd cell_6t
Xbit_r12_c79 bl_79 br_79 wl_12 vdd gnd cell_6t
Xbit_r13_c79 bl_79 br_79 wl_13 vdd gnd cell_6t
Xbit_r14_c79 bl_79 br_79 wl_14 vdd gnd cell_6t
Xbit_r15_c79 bl_79 br_79 wl_15 vdd gnd cell_6t
Xbit_r16_c79 bl_79 br_79 wl_16 vdd gnd cell_6t
Xbit_r17_c79 bl_79 br_79 wl_17 vdd gnd cell_6t
Xbit_r18_c79 bl_79 br_79 wl_18 vdd gnd cell_6t
Xbit_r19_c79 bl_79 br_79 wl_19 vdd gnd cell_6t
Xbit_r20_c79 bl_79 br_79 wl_20 vdd gnd cell_6t
Xbit_r21_c79 bl_79 br_79 wl_21 vdd gnd cell_6t
Xbit_r22_c79 bl_79 br_79 wl_22 vdd gnd cell_6t
Xbit_r23_c79 bl_79 br_79 wl_23 vdd gnd cell_6t
Xbit_r24_c79 bl_79 br_79 wl_24 vdd gnd cell_6t
Xbit_r25_c79 bl_79 br_79 wl_25 vdd gnd cell_6t
Xbit_r26_c79 bl_79 br_79 wl_26 vdd gnd cell_6t
Xbit_r27_c79 bl_79 br_79 wl_27 vdd gnd cell_6t
Xbit_r28_c79 bl_79 br_79 wl_28 vdd gnd cell_6t
Xbit_r29_c79 bl_79 br_79 wl_29 vdd gnd cell_6t
Xbit_r30_c79 bl_79 br_79 wl_30 vdd gnd cell_6t
Xbit_r31_c79 bl_79 br_79 wl_31 vdd gnd cell_6t
Xbit_r32_c79 bl_79 br_79 wl_32 vdd gnd cell_6t
Xbit_r33_c79 bl_79 br_79 wl_33 vdd gnd cell_6t
Xbit_r34_c79 bl_79 br_79 wl_34 vdd gnd cell_6t
Xbit_r35_c79 bl_79 br_79 wl_35 vdd gnd cell_6t
Xbit_r36_c79 bl_79 br_79 wl_36 vdd gnd cell_6t
Xbit_r37_c79 bl_79 br_79 wl_37 vdd gnd cell_6t
Xbit_r38_c79 bl_79 br_79 wl_38 vdd gnd cell_6t
Xbit_r39_c79 bl_79 br_79 wl_39 vdd gnd cell_6t
Xbit_r40_c79 bl_79 br_79 wl_40 vdd gnd cell_6t
Xbit_r41_c79 bl_79 br_79 wl_41 vdd gnd cell_6t
Xbit_r42_c79 bl_79 br_79 wl_42 vdd gnd cell_6t
Xbit_r43_c79 bl_79 br_79 wl_43 vdd gnd cell_6t
Xbit_r44_c79 bl_79 br_79 wl_44 vdd gnd cell_6t
Xbit_r45_c79 bl_79 br_79 wl_45 vdd gnd cell_6t
Xbit_r46_c79 bl_79 br_79 wl_46 vdd gnd cell_6t
Xbit_r47_c79 bl_79 br_79 wl_47 vdd gnd cell_6t
Xbit_r48_c79 bl_79 br_79 wl_48 vdd gnd cell_6t
Xbit_r49_c79 bl_79 br_79 wl_49 vdd gnd cell_6t
Xbit_r50_c79 bl_79 br_79 wl_50 vdd gnd cell_6t
Xbit_r51_c79 bl_79 br_79 wl_51 vdd gnd cell_6t
Xbit_r52_c79 bl_79 br_79 wl_52 vdd gnd cell_6t
Xbit_r53_c79 bl_79 br_79 wl_53 vdd gnd cell_6t
Xbit_r54_c79 bl_79 br_79 wl_54 vdd gnd cell_6t
Xbit_r55_c79 bl_79 br_79 wl_55 vdd gnd cell_6t
Xbit_r56_c79 bl_79 br_79 wl_56 vdd gnd cell_6t
Xbit_r57_c79 bl_79 br_79 wl_57 vdd gnd cell_6t
Xbit_r58_c79 bl_79 br_79 wl_58 vdd gnd cell_6t
Xbit_r59_c79 bl_79 br_79 wl_59 vdd gnd cell_6t
Xbit_r60_c79 bl_79 br_79 wl_60 vdd gnd cell_6t
Xbit_r61_c79 bl_79 br_79 wl_61 vdd gnd cell_6t
Xbit_r62_c79 bl_79 br_79 wl_62 vdd gnd cell_6t
Xbit_r63_c79 bl_79 br_79 wl_63 vdd gnd cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd cell_6t
Xbit_r1_c80 bl_80 br_80 wl_1 vdd gnd cell_6t
Xbit_r2_c80 bl_80 br_80 wl_2 vdd gnd cell_6t
Xbit_r3_c80 bl_80 br_80 wl_3 vdd gnd cell_6t
Xbit_r4_c80 bl_80 br_80 wl_4 vdd gnd cell_6t
Xbit_r5_c80 bl_80 br_80 wl_5 vdd gnd cell_6t
Xbit_r6_c80 bl_80 br_80 wl_6 vdd gnd cell_6t
Xbit_r7_c80 bl_80 br_80 wl_7 vdd gnd cell_6t
Xbit_r8_c80 bl_80 br_80 wl_8 vdd gnd cell_6t
Xbit_r9_c80 bl_80 br_80 wl_9 vdd gnd cell_6t
Xbit_r10_c80 bl_80 br_80 wl_10 vdd gnd cell_6t
Xbit_r11_c80 bl_80 br_80 wl_11 vdd gnd cell_6t
Xbit_r12_c80 bl_80 br_80 wl_12 vdd gnd cell_6t
Xbit_r13_c80 bl_80 br_80 wl_13 vdd gnd cell_6t
Xbit_r14_c80 bl_80 br_80 wl_14 vdd gnd cell_6t
Xbit_r15_c80 bl_80 br_80 wl_15 vdd gnd cell_6t
Xbit_r16_c80 bl_80 br_80 wl_16 vdd gnd cell_6t
Xbit_r17_c80 bl_80 br_80 wl_17 vdd gnd cell_6t
Xbit_r18_c80 bl_80 br_80 wl_18 vdd gnd cell_6t
Xbit_r19_c80 bl_80 br_80 wl_19 vdd gnd cell_6t
Xbit_r20_c80 bl_80 br_80 wl_20 vdd gnd cell_6t
Xbit_r21_c80 bl_80 br_80 wl_21 vdd gnd cell_6t
Xbit_r22_c80 bl_80 br_80 wl_22 vdd gnd cell_6t
Xbit_r23_c80 bl_80 br_80 wl_23 vdd gnd cell_6t
Xbit_r24_c80 bl_80 br_80 wl_24 vdd gnd cell_6t
Xbit_r25_c80 bl_80 br_80 wl_25 vdd gnd cell_6t
Xbit_r26_c80 bl_80 br_80 wl_26 vdd gnd cell_6t
Xbit_r27_c80 bl_80 br_80 wl_27 vdd gnd cell_6t
Xbit_r28_c80 bl_80 br_80 wl_28 vdd gnd cell_6t
Xbit_r29_c80 bl_80 br_80 wl_29 vdd gnd cell_6t
Xbit_r30_c80 bl_80 br_80 wl_30 vdd gnd cell_6t
Xbit_r31_c80 bl_80 br_80 wl_31 vdd gnd cell_6t
Xbit_r32_c80 bl_80 br_80 wl_32 vdd gnd cell_6t
Xbit_r33_c80 bl_80 br_80 wl_33 vdd gnd cell_6t
Xbit_r34_c80 bl_80 br_80 wl_34 vdd gnd cell_6t
Xbit_r35_c80 bl_80 br_80 wl_35 vdd gnd cell_6t
Xbit_r36_c80 bl_80 br_80 wl_36 vdd gnd cell_6t
Xbit_r37_c80 bl_80 br_80 wl_37 vdd gnd cell_6t
Xbit_r38_c80 bl_80 br_80 wl_38 vdd gnd cell_6t
Xbit_r39_c80 bl_80 br_80 wl_39 vdd gnd cell_6t
Xbit_r40_c80 bl_80 br_80 wl_40 vdd gnd cell_6t
Xbit_r41_c80 bl_80 br_80 wl_41 vdd gnd cell_6t
Xbit_r42_c80 bl_80 br_80 wl_42 vdd gnd cell_6t
Xbit_r43_c80 bl_80 br_80 wl_43 vdd gnd cell_6t
Xbit_r44_c80 bl_80 br_80 wl_44 vdd gnd cell_6t
Xbit_r45_c80 bl_80 br_80 wl_45 vdd gnd cell_6t
Xbit_r46_c80 bl_80 br_80 wl_46 vdd gnd cell_6t
Xbit_r47_c80 bl_80 br_80 wl_47 vdd gnd cell_6t
Xbit_r48_c80 bl_80 br_80 wl_48 vdd gnd cell_6t
Xbit_r49_c80 bl_80 br_80 wl_49 vdd gnd cell_6t
Xbit_r50_c80 bl_80 br_80 wl_50 vdd gnd cell_6t
Xbit_r51_c80 bl_80 br_80 wl_51 vdd gnd cell_6t
Xbit_r52_c80 bl_80 br_80 wl_52 vdd gnd cell_6t
Xbit_r53_c80 bl_80 br_80 wl_53 vdd gnd cell_6t
Xbit_r54_c80 bl_80 br_80 wl_54 vdd gnd cell_6t
Xbit_r55_c80 bl_80 br_80 wl_55 vdd gnd cell_6t
Xbit_r56_c80 bl_80 br_80 wl_56 vdd gnd cell_6t
Xbit_r57_c80 bl_80 br_80 wl_57 vdd gnd cell_6t
Xbit_r58_c80 bl_80 br_80 wl_58 vdd gnd cell_6t
Xbit_r59_c80 bl_80 br_80 wl_59 vdd gnd cell_6t
Xbit_r60_c80 bl_80 br_80 wl_60 vdd gnd cell_6t
Xbit_r61_c80 bl_80 br_80 wl_61 vdd gnd cell_6t
Xbit_r62_c80 bl_80 br_80 wl_62 vdd gnd cell_6t
Xbit_r63_c80 bl_80 br_80 wl_63 vdd gnd cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd cell_6t
Xbit_r1_c81 bl_81 br_81 wl_1 vdd gnd cell_6t
Xbit_r2_c81 bl_81 br_81 wl_2 vdd gnd cell_6t
Xbit_r3_c81 bl_81 br_81 wl_3 vdd gnd cell_6t
Xbit_r4_c81 bl_81 br_81 wl_4 vdd gnd cell_6t
Xbit_r5_c81 bl_81 br_81 wl_5 vdd gnd cell_6t
Xbit_r6_c81 bl_81 br_81 wl_6 vdd gnd cell_6t
Xbit_r7_c81 bl_81 br_81 wl_7 vdd gnd cell_6t
Xbit_r8_c81 bl_81 br_81 wl_8 vdd gnd cell_6t
Xbit_r9_c81 bl_81 br_81 wl_9 vdd gnd cell_6t
Xbit_r10_c81 bl_81 br_81 wl_10 vdd gnd cell_6t
Xbit_r11_c81 bl_81 br_81 wl_11 vdd gnd cell_6t
Xbit_r12_c81 bl_81 br_81 wl_12 vdd gnd cell_6t
Xbit_r13_c81 bl_81 br_81 wl_13 vdd gnd cell_6t
Xbit_r14_c81 bl_81 br_81 wl_14 vdd gnd cell_6t
Xbit_r15_c81 bl_81 br_81 wl_15 vdd gnd cell_6t
Xbit_r16_c81 bl_81 br_81 wl_16 vdd gnd cell_6t
Xbit_r17_c81 bl_81 br_81 wl_17 vdd gnd cell_6t
Xbit_r18_c81 bl_81 br_81 wl_18 vdd gnd cell_6t
Xbit_r19_c81 bl_81 br_81 wl_19 vdd gnd cell_6t
Xbit_r20_c81 bl_81 br_81 wl_20 vdd gnd cell_6t
Xbit_r21_c81 bl_81 br_81 wl_21 vdd gnd cell_6t
Xbit_r22_c81 bl_81 br_81 wl_22 vdd gnd cell_6t
Xbit_r23_c81 bl_81 br_81 wl_23 vdd gnd cell_6t
Xbit_r24_c81 bl_81 br_81 wl_24 vdd gnd cell_6t
Xbit_r25_c81 bl_81 br_81 wl_25 vdd gnd cell_6t
Xbit_r26_c81 bl_81 br_81 wl_26 vdd gnd cell_6t
Xbit_r27_c81 bl_81 br_81 wl_27 vdd gnd cell_6t
Xbit_r28_c81 bl_81 br_81 wl_28 vdd gnd cell_6t
Xbit_r29_c81 bl_81 br_81 wl_29 vdd gnd cell_6t
Xbit_r30_c81 bl_81 br_81 wl_30 vdd gnd cell_6t
Xbit_r31_c81 bl_81 br_81 wl_31 vdd gnd cell_6t
Xbit_r32_c81 bl_81 br_81 wl_32 vdd gnd cell_6t
Xbit_r33_c81 bl_81 br_81 wl_33 vdd gnd cell_6t
Xbit_r34_c81 bl_81 br_81 wl_34 vdd gnd cell_6t
Xbit_r35_c81 bl_81 br_81 wl_35 vdd gnd cell_6t
Xbit_r36_c81 bl_81 br_81 wl_36 vdd gnd cell_6t
Xbit_r37_c81 bl_81 br_81 wl_37 vdd gnd cell_6t
Xbit_r38_c81 bl_81 br_81 wl_38 vdd gnd cell_6t
Xbit_r39_c81 bl_81 br_81 wl_39 vdd gnd cell_6t
Xbit_r40_c81 bl_81 br_81 wl_40 vdd gnd cell_6t
Xbit_r41_c81 bl_81 br_81 wl_41 vdd gnd cell_6t
Xbit_r42_c81 bl_81 br_81 wl_42 vdd gnd cell_6t
Xbit_r43_c81 bl_81 br_81 wl_43 vdd gnd cell_6t
Xbit_r44_c81 bl_81 br_81 wl_44 vdd gnd cell_6t
Xbit_r45_c81 bl_81 br_81 wl_45 vdd gnd cell_6t
Xbit_r46_c81 bl_81 br_81 wl_46 vdd gnd cell_6t
Xbit_r47_c81 bl_81 br_81 wl_47 vdd gnd cell_6t
Xbit_r48_c81 bl_81 br_81 wl_48 vdd gnd cell_6t
Xbit_r49_c81 bl_81 br_81 wl_49 vdd gnd cell_6t
Xbit_r50_c81 bl_81 br_81 wl_50 vdd gnd cell_6t
Xbit_r51_c81 bl_81 br_81 wl_51 vdd gnd cell_6t
Xbit_r52_c81 bl_81 br_81 wl_52 vdd gnd cell_6t
Xbit_r53_c81 bl_81 br_81 wl_53 vdd gnd cell_6t
Xbit_r54_c81 bl_81 br_81 wl_54 vdd gnd cell_6t
Xbit_r55_c81 bl_81 br_81 wl_55 vdd gnd cell_6t
Xbit_r56_c81 bl_81 br_81 wl_56 vdd gnd cell_6t
Xbit_r57_c81 bl_81 br_81 wl_57 vdd gnd cell_6t
Xbit_r58_c81 bl_81 br_81 wl_58 vdd gnd cell_6t
Xbit_r59_c81 bl_81 br_81 wl_59 vdd gnd cell_6t
Xbit_r60_c81 bl_81 br_81 wl_60 vdd gnd cell_6t
Xbit_r61_c81 bl_81 br_81 wl_61 vdd gnd cell_6t
Xbit_r62_c81 bl_81 br_81 wl_62 vdd gnd cell_6t
Xbit_r63_c81 bl_81 br_81 wl_63 vdd gnd cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd cell_6t
Xbit_r1_c82 bl_82 br_82 wl_1 vdd gnd cell_6t
Xbit_r2_c82 bl_82 br_82 wl_2 vdd gnd cell_6t
Xbit_r3_c82 bl_82 br_82 wl_3 vdd gnd cell_6t
Xbit_r4_c82 bl_82 br_82 wl_4 vdd gnd cell_6t
Xbit_r5_c82 bl_82 br_82 wl_5 vdd gnd cell_6t
Xbit_r6_c82 bl_82 br_82 wl_6 vdd gnd cell_6t
Xbit_r7_c82 bl_82 br_82 wl_7 vdd gnd cell_6t
Xbit_r8_c82 bl_82 br_82 wl_8 vdd gnd cell_6t
Xbit_r9_c82 bl_82 br_82 wl_9 vdd gnd cell_6t
Xbit_r10_c82 bl_82 br_82 wl_10 vdd gnd cell_6t
Xbit_r11_c82 bl_82 br_82 wl_11 vdd gnd cell_6t
Xbit_r12_c82 bl_82 br_82 wl_12 vdd gnd cell_6t
Xbit_r13_c82 bl_82 br_82 wl_13 vdd gnd cell_6t
Xbit_r14_c82 bl_82 br_82 wl_14 vdd gnd cell_6t
Xbit_r15_c82 bl_82 br_82 wl_15 vdd gnd cell_6t
Xbit_r16_c82 bl_82 br_82 wl_16 vdd gnd cell_6t
Xbit_r17_c82 bl_82 br_82 wl_17 vdd gnd cell_6t
Xbit_r18_c82 bl_82 br_82 wl_18 vdd gnd cell_6t
Xbit_r19_c82 bl_82 br_82 wl_19 vdd gnd cell_6t
Xbit_r20_c82 bl_82 br_82 wl_20 vdd gnd cell_6t
Xbit_r21_c82 bl_82 br_82 wl_21 vdd gnd cell_6t
Xbit_r22_c82 bl_82 br_82 wl_22 vdd gnd cell_6t
Xbit_r23_c82 bl_82 br_82 wl_23 vdd gnd cell_6t
Xbit_r24_c82 bl_82 br_82 wl_24 vdd gnd cell_6t
Xbit_r25_c82 bl_82 br_82 wl_25 vdd gnd cell_6t
Xbit_r26_c82 bl_82 br_82 wl_26 vdd gnd cell_6t
Xbit_r27_c82 bl_82 br_82 wl_27 vdd gnd cell_6t
Xbit_r28_c82 bl_82 br_82 wl_28 vdd gnd cell_6t
Xbit_r29_c82 bl_82 br_82 wl_29 vdd gnd cell_6t
Xbit_r30_c82 bl_82 br_82 wl_30 vdd gnd cell_6t
Xbit_r31_c82 bl_82 br_82 wl_31 vdd gnd cell_6t
Xbit_r32_c82 bl_82 br_82 wl_32 vdd gnd cell_6t
Xbit_r33_c82 bl_82 br_82 wl_33 vdd gnd cell_6t
Xbit_r34_c82 bl_82 br_82 wl_34 vdd gnd cell_6t
Xbit_r35_c82 bl_82 br_82 wl_35 vdd gnd cell_6t
Xbit_r36_c82 bl_82 br_82 wl_36 vdd gnd cell_6t
Xbit_r37_c82 bl_82 br_82 wl_37 vdd gnd cell_6t
Xbit_r38_c82 bl_82 br_82 wl_38 vdd gnd cell_6t
Xbit_r39_c82 bl_82 br_82 wl_39 vdd gnd cell_6t
Xbit_r40_c82 bl_82 br_82 wl_40 vdd gnd cell_6t
Xbit_r41_c82 bl_82 br_82 wl_41 vdd gnd cell_6t
Xbit_r42_c82 bl_82 br_82 wl_42 vdd gnd cell_6t
Xbit_r43_c82 bl_82 br_82 wl_43 vdd gnd cell_6t
Xbit_r44_c82 bl_82 br_82 wl_44 vdd gnd cell_6t
Xbit_r45_c82 bl_82 br_82 wl_45 vdd gnd cell_6t
Xbit_r46_c82 bl_82 br_82 wl_46 vdd gnd cell_6t
Xbit_r47_c82 bl_82 br_82 wl_47 vdd gnd cell_6t
Xbit_r48_c82 bl_82 br_82 wl_48 vdd gnd cell_6t
Xbit_r49_c82 bl_82 br_82 wl_49 vdd gnd cell_6t
Xbit_r50_c82 bl_82 br_82 wl_50 vdd gnd cell_6t
Xbit_r51_c82 bl_82 br_82 wl_51 vdd gnd cell_6t
Xbit_r52_c82 bl_82 br_82 wl_52 vdd gnd cell_6t
Xbit_r53_c82 bl_82 br_82 wl_53 vdd gnd cell_6t
Xbit_r54_c82 bl_82 br_82 wl_54 vdd gnd cell_6t
Xbit_r55_c82 bl_82 br_82 wl_55 vdd gnd cell_6t
Xbit_r56_c82 bl_82 br_82 wl_56 vdd gnd cell_6t
Xbit_r57_c82 bl_82 br_82 wl_57 vdd gnd cell_6t
Xbit_r58_c82 bl_82 br_82 wl_58 vdd gnd cell_6t
Xbit_r59_c82 bl_82 br_82 wl_59 vdd gnd cell_6t
Xbit_r60_c82 bl_82 br_82 wl_60 vdd gnd cell_6t
Xbit_r61_c82 bl_82 br_82 wl_61 vdd gnd cell_6t
Xbit_r62_c82 bl_82 br_82 wl_62 vdd gnd cell_6t
Xbit_r63_c82 bl_82 br_82 wl_63 vdd gnd cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd cell_6t
Xbit_r1_c83 bl_83 br_83 wl_1 vdd gnd cell_6t
Xbit_r2_c83 bl_83 br_83 wl_2 vdd gnd cell_6t
Xbit_r3_c83 bl_83 br_83 wl_3 vdd gnd cell_6t
Xbit_r4_c83 bl_83 br_83 wl_4 vdd gnd cell_6t
Xbit_r5_c83 bl_83 br_83 wl_5 vdd gnd cell_6t
Xbit_r6_c83 bl_83 br_83 wl_6 vdd gnd cell_6t
Xbit_r7_c83 bl_83 br_83 wl_7 vdd gnd cell_6t
Xbit_r8_c83 bl_83 br_83 wl_8 vdd gnd cell_6t
Xbit_r9_c83 bl_83 br_83 wl_9 vdd gnd cell_6t
Xbit_r10_c83 bl_83 br_83 wl_10 vdd gnd cell_6t
Xbit_r11_c83 bl_83 br_83 wl_11 vdd gnd cell_6t
Xbit_r12_c83 bl_83 br_83 wl_12 vdd gnd cell_6t
Xbit_r13_c83 bl_83 br_83 wl_13 vdd gnd cell_6t
Xbit_r14_c83 bl_83 br_83 wl_14 vdd gnd cell_6t
Xbit_r15_c83 bl_83 br_83 wl_15 vdd gnd cell_6t
Xbit_r16_c83 bl_83 br_83 wl_16 vdd gnd cell_6t
Xbit_r17_c83 bl_83 br_83 wl_17 vdd gnd cell_6t
Xbit_r18_c83 bl_83 br_83 wl_18 vdd gnd cell_6t
Xbit_r19_c83 bl_83 br_83 wl_19 vdd gnd cell_6t
Xbit_r20_c83 bl_83 br_83 wl_20 vdd gnd cell_6t
Xbit_r21_c83 bl_83 br_83 wl_21 vdd gnd cell_6t
Xbit_r22_c83 bl_83 br_83 wl_22 vdd gnd cell_6t
Xbit_r23_c83 bl_83 br_83 wl_23 vdd gnd cell_6t
Xbit_r24_c83 bl_83 br_83 wl_24 vdd gnd cell_6t
Xbit_r25_c83 bl_83 br_83 wl_25 vdd gnd cell_6t
Xbit_r26_c83 bl_83 br_83 wl_26 vdd gnd cell_6t
Xbit_r27_c83 bl_83 br_83 wl_27 vdd gnd cell_6t
Xbit_r28_c83 bl_83 br_83 wl_28 vdd gnd cell_6t
Xbit_r29_c83 bl_83 br_83 wl_29 vdd gnd cell_6t
Xbit_r30_c83 bl_83 br_83 wl_30 vdd gnd cell_6t
Xbit_r31_c83 bl_83 br_83 wl_31 vdd gnd cell_6t
Xbit_r32_c83 bl_83 br_83 wl_32 vdd gnd cell_6t
Xbit_r33_c83 bl_83 br_83 wl_33 vdd gnd cell_6t
Xbit_r34_c83 bl_83 br_83 wl_34 vdd gnd cell_6t
Xbit_r35_c83 bl_83 br_83 wl_35 vdd gnd cell_6t
Xbit_r36_c83 bl_83 br_83 wl_36 vdd gnd cell_6t
Xbit_r37_c83 bl_83 br_83 wl_37 vdd gnd cell_6t
Xbit_r38_c83 bl_83 br_83 wl_38 vdd gnd cell_6t
Xbit_r39_c83 bl_83 br_83 wl_39 vdd gnd cell_6t
Xbit_r40_c83 bl_83 br_83 wl_40 vdd gnd cell_6t
Xbit_r41_c83 bl_83 br_83 wl_41 vdd gnd cell_6t
Xbit_r42_c83 bl_83 br_83 wl_42 vdd gnd cell_6t
Xbit_r43_c83 bl_83 br_83 wl_43 vdd gnd cell_6t
Xbit_r44_c83 bl_83 br_83 wl_44 vdd gnd cell_6t
Xbit_r45_c83 bl_83 br_83 wl_45 vdd gnd cell_6t
Xbit_r46_c83 bl_83 br_83 wl_46 vdd gnd cell_6t
Xbit_r47_c83 bl_83 br_83 wl_47 vdd gnd cell_6t
Xbit_r48_c83 bl_83 br_83 wl_48 vdd gnd cell_6t
Xbit_r49_c83 bl_83 br_83 wl_49 vdd gnd cell_6t
Xbit_r50_c83 bl_83 br_83 wl_50 vdd gnd cell_6t
Xbit_r51_c83 bl_83 br_83 wl_51 vdd gnd cell_6t
Xbit_r52_c83 bl_83 br_83 wl_52 vdd gnd cell_6t
Xbit_r53_c83 bl_83 br_83 wl_53 vdd gnd cell_6t
Xbit_r54_c83 bl_83 br_83 wl_54 vdd gnd cell_6t
Xbit_r55_c83 bl_83 br_83 wl_55 vdd gnd cell_6t
Xbit_r56_c83 bl_83 br_83 wl_56 vdd gnd cell_6t
Xbit_r57_c83 bl_83 br_83 wl_57 vdd gnd cell_6t
Xbit_r58_c83 bl_83 br_83 wl_58 vdd gnd cell_6t
Xbit_r59_c83 bl_83 br_83 wl_59 vdd gnd cell_6t
Xbit_r60_c83 bl_83 br_83 wl_60 vdd gnd cell_6t
Xbit_r61_c83 bl_83 br_83 wl_61 vdd gnd cell_6t
Xbit_r62_c83 bl_83 br_83 wl_62 vdd gnd cell_6t
Xbit_r63_c83 bl_83 br_83 wl_63 vdd gnd cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd cell_6t
Xbit_r1_c84 bl_84 br_84 wl_1 vdd gnd cell_6t
Xbit_r2_c84 bl_84 br_84 wl_2 vdd gnd cell_6t
Xbit_r3_c84 bl_84 br_84 wl_3 vdd gnd cell_6t
Xbit_r4_c84 bl_84 br_84 wl_4 vdd gnd cell_6t
Xbit_r5_c84 bl_84 br_84 wl_5 vdd gnd cell_6t
Xbit_r6_c84 bl_84 br_84 wl_6 vdd gnd cell_6t
Xbit_r7_c84 bl_84 br_84 wl_7 vdd gnd cell_6t
Xbit_r8_c84 bl_84 br_84 wl_8 vdd gnd cell_6t
Xbit_r9_c84 bl_84 br_84 wl_9 vdd gnd cell_6t
Xbit_r10_c84 bl_84 br_84 wl_10 vdd gnd cell_6t
Xbit_r11_c84 bl_84 br_84 wl_11 vdd gnd cell_6t
Xbit_r12_c84 bl_84 br_84 wl_12 vdd gnd cell_6t
Xbit_r13_c84 bl_84 br_84 wl_13 vdd gnd cell_6t
Xbit_r14_c84 bl_84 br_84 wl_14 vdd gnd cell_6t
Xbit_r15_c84 bl_84 br_84 wl_15 vdd gnd cell_6t
Xbit_r16_c84 bl_84 br_84 wl_16 vdd gnd cell_6t
Xbit_r17_c84 bl_84 br_84 wl_17 vdd gnd cell_6t
Xbit_r18_c84 bl_84 br_84 wl_18 vdd gnd cell_6t
Xbit_r19_c84 bl_84 br_84 wl_19 vdd gnd cell_6t
Xbit_r20_c84 bl_84 br_84 wl_20 vdd gnd cell_6t
Xbit_r21_c84 bl_84 br_84 wl_21 vdd gnd cell_6t
Xbit_r22_c84 bl_84 br_84 wl_22 vdd gnd cell_6t
Xbit_r23_c84 bl_84 br_84 wl_23 vdd gnd cell_6t
Xbit_r24_c84 bl_84 br_84 wl_24 vdd gnd cell_6t
Xbit_r25_c84 bl_84 br_84 wl_25 vdd gnd cell_6t
Xbit_r26_c84 bl_84 br_84 wl_26 vdd gnd cell_6t
Xbit_r27_c84 bl_84 br_84 wl_27 vdd gnd cell_6t
Xbit_r28_c84 bl_84 br_84 wl_28 vdd gnd cell_6t
Xbit_r29_c84 bl_84 br_84 wl_29 vdd gnd cell_6t
Xbit_r30_c84 bl_84 br_84 wl_30 vdd gnd cell_6t
Xbit_r31_c84 bl_84 br_84 wl_31 vdd gnd cell_6t
Xbit_r32_c84 bl_84 br_84 wl_32 vdd gnd cell_6t
Xbit_r33_c84 bl_84 br_84 wl_33 vdd gnd cell_6t
Xbit_r34_c84 bl_84 br_84 wl_34 vdd gnd cell_6t
Xbit_r35_c84 bl_84 br_84 wl_35 vdd gnd cell_6t
Xbit_r36_c84 bl_84 br_84 wl_36 vdd gnd cell_6t
Xbit_r37_c84 bl_84 br_84 wl_37 vdd gnd cell_6t
Xbit_r38_c84 bl_84 br_84 wl_38 vdd gnd cell_6t
Xbit_r39_c84 bl_84 br_84 wl_39 vdd gnd cell_6t
Xbit_r40_c84 bl_84 br_84 wl_40 vdd gnd cell_6t
Xbit_r41_c84 bl_84 br_84 wl_41 vdd gnd cell_6t
Xbit_r42_c84 bl_84 br_84 wl_42 vdd gnd cell_6t
Xbit_r43_c84 bl_84 br_84 wl_43 vdd gnd cell_6t
Xbit_r44_c84 bl_84 br_84 wl_44 vdd gnd cell_6t
Xbit_r45_c84 bl_84 br_84 wl_45 vdd gnd cell_6t
Xbit_r46_c84 bl_84 br_84 wl_46 vdd gnd cell_6t
Xbit_r47_c84 bl_84 br_84 wl_47 vdd gnd cell_6t
Xbit_r48_c84 bl_84 br_84 wl_48 vdd gnd cell_6t
Xbit_r49_c84 bl_84 br_84 wl_49 vdd gnd cell_6t
Xbit_r50_c84 bl_84 br_84 wl_50 vdd gnd cell_6t
Xbit_r51_c84 bl_84 br_84 wl_51 vdd gnd cell_6t
Xbit_r52_c84 bl_84 br_84 wl_52 vdd gnd cell_6t
Xbit_r53_c84 bl_84 br_84 wl_53 vdd gnd cell_6t
Xbit_r54_c84 bl_84 br_84 wl_54 vdd gnd cell_6t
Xbit_r55_c84 bl_84 br_84 wl_55 vdd gnd cell_6t
Xbit_r56_c84 bl_84 br_84 wl_56 vdd gnd cell_6t
Xbit_r57_c84 bl_84 br_84 wl_57 vdd gnd cell_6t
Xbit_r58_c84 bl_84 br_84 wl_58 vdd gnd cell_6t
Xbit_r59_c84 bl_84 br_84 wl_59 vdd gnd cell_6t
Xbit_r60_c84 bl_84 br_84 wl_60 vdd gnd cell_6t
Xbit_r61_c84 bl_84 br_84 wl_61 vdd gnd cell_6t
Xbit_r62_c84 bl_84 br_84 wl_62 vdd gnd cell_6t
Xbit_r63_c84 bl_84 br_84 wl_63 vdd gnd cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd cell_6t
Xbit_r1_c85 bl_85 br_85 wl_1 vdd gnd cell_6t
Xbit_r2_c85 bl_85 br_85 wl_2 vdd gnd cell_6t
Xbit_r3_c85 bl_85 br_85 wl_3 vdd gnd cell_6t
Xbit_r4_c85 bl_85 br_85 wl_4 vdd gnd cell_6t
Xbit_r5_c85 bl_85 br_85 wl_5 vdd gnd cell_6t
Xbit_r6_c85 bl_85 br_85 wl_6 vdd gnd cell_6t
Xbit_r7_c85 bl_85 br_85 wl_7 vdd gnd cell_6t
Xbit_r8_c85 bl_85 br_85 wl_8 vdd gnd cell_6t
Xbit_r9_c85 bl_85 br_85 wl_9 vdd gnd cell_6t
Xbit_r10_c85 bl_85 br_85 wl_10 vdd gnd cell_6t
Xbit_r11_c85 bl_85 br_85 wl_11 vdd gnd cell_6t
Xbit_r12_c85 bl_85 br_85 wl_12 vdd gnd cell_6t
Xbit_r13_c85 bl_85 br_85 wl_13 vdd gnd cell_6t
Xbit_r14_c85 bl_85 br_85 wl_14 vdd gnd cell_6t
Xbit_r15_c85 bl_85 br_85 wl_15 vdd gnd cell_6t
Xbit_r16_c85 bl_85 br_85 wl_16 vdd gnd cell_6t
Xbit_r17_c85 bl_85 br_85 wl_17 vdd gnd cell_6t
Xbit_r18_c85 bl_85 br_85 wl_18 vdd gnd cell_6t
Xbit_r19_c85 bl_85 br_85 wl_19 vdd gnd cell_6t
Xbit_r20_c85 bl_85 br_85 wl_20 vdd gnd cell_6t
Xbit_r21_c85 bl_85 br_85 wl_21 vdd gnd cell_6t
Xbit_r22_c85 bl_85 br_85 wl_22 vdd gnd cell_6t
Xbit_r23_c85 bl_85 br_85 wl_23 vdd gnd cell_6t
Xbit_r24_c85 bl_85 br_85 wl_24 vdd gnd cell_6t
Xbit_r25_c85 bl_85 br_85 wl_25 vdd gnd cell_6t
Xbit_r26_c85 bl_85 br_85 wl_26 vdd gnd cell_6t
Xbit_r27_c85 bl_85 br_85 wl_27 vdd gnd cell_6t
Xbit_r28_c85 bl_85 br_85 wl_28 vdd gnd cell_6t
Xbit_r29_c85 bl_85 br_85 wl_29 vdd gnd cell_6t
Xbit_r30_c85 bl_85 br_85 wl_30 vdd gnd cell_6t
Xbit_r31_c85 bl_85 br_85 wl_31 vdd gnd cell_6t
Xbit_r32_c85 bl_85 br_85 wl_32 vdd gnd cell_6t
Xbit_r33_c85 bl_85 br_85 wl_33 vdd gnd cell_6t
Xbit_r34_c85 bl_85 br_85 wl_34 vdd gnd cell_6t
Xbit_r35_c85 bl_85 br_85 wl_35 vdd gnd cell_6t
Xbit_r36_c85 bl_85 br_85 wl_36 vdd gnd cell_6t
Xbit_r37_c85 bl_85 br_85 wl_37 vdd gnd cell_6t
Xbit_r38_c85 bl_85 br_85 wl_38 vdd gnd cell_6t
Xbit_r39_c85 bl_85 br_85 wl_39 vdd gnd cell_6t
Xbit_r40_c85 bl_85 br_85 wl_40 vdd gnd cell_6t
Xbit_r41_c85 bl_85 br_85 wl_41 vdd gnd cell_6t
Xbit_r42_c85 bl_85 br_85 wl_42 vdd gnd cell_6t
Xbit_r43_c85 bl_85 br_85 wl_43 vdd gnd cell_6t
Xbit_r44_c85 bl_85 br_85 wl_44 vdd gnd cell_6t
Xbit_r45_c85 bl_85 br_85 wl_45 vdd gnd cell_6t
Xbit_r46_c85 bl_85 br_85 wl_46 vdd gnd cell_6t
Xbit_r47_c85 bl_85 br_85 wl_47 vdd gnd cell_6t
Xbit_r48_c85 bl_85 br_85 wl_48 vdd gnd cell_6t
Xbit_r49_c85 bl_85 br_85 wl_49 vdd gnd cell_6t
Xbit_r50_c85 bl_85 br_85 wl_50 vdd gnd cell_6t
Xbit_r51_c85 bl_85 br_85 wl_51 vdd gnd cell_6t
Xbit_r52_c85 bl_85 br_85 wl_52 vdd gnd cell_6t
Xbit_r53_c85 bl_85 br_85 wl_53 vdd gnd cell_6t
Xbit_r54_c85 bl_85 br_85 wl_54 vdd gnd cell_6t
Xbit_r55_c85 bl_85 br_85 wl_55 vdd gnd cell_6t
Xbit_r56_c85 bl_85 br_85 wl_56 vdd gnd cell_6t
Xbit_r57_c85 bl_85 br_85 wl_57 vdd gnd cell_6t
Xbit_r58_c85 bl_85 br_85 wl_58 vdd gnd cell_6t
Xbit_r59_c85 bl_85 br_85 wl_59 vdd gnd cell_6t
Xbit_r60_c85 bl_85 br_85 wl_60 vdd gnd cell_6t
Xbit_r61_c85 bl_85 br_85 wl_61 vdd gnd cell_6t
Xbit_r62_c85 bl_85 br_85 wl_62 vdd gnd cell_6t
Xbit_r63_c85 bl_85 br_85 wl_63 vdd gnd cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd cell_6t
Xbit_r1_c86 bl_86 br_86 wl_1 vdd gnd cell_6t
Xbit_r2_c86 bl_86 br_86 wl_2 vdd gnd cell_6t
Xbit_r3_c86 bl_86 br_86 wl_3 vdd gnd cell_6t
Xbit_r4_c86 bl_86 br_86 wl_4 vdd gnd cell_6t
Xbit_r5_c86 bl_86 br_86 wl_5 vdd gnd cell_6t
Xbit_r6_c86 bl_86 br_86 wl_6 vdd gnd cell_6t
Xbit_r7_c86 bl_86 br_86 wl_7 vdd gnd cell_6t
Xbit_r8_c86 bl_86 br_86 wl_8 vdd gnd cell_6t
Xbit_r9_c86 bl_86 br_86 wl_9 vdd gnd cell_6t
Xbit_r10_c86 bl_86 br_86 wl_10 vdd gnd cell_6t
Xbit_r11_c86 bl_86 br_86 wl_11 vdd gnd cell_6t
Xbit_r12_c86 bl_86 br_86 wl_12 vdd gnd cell_6t
Xbit_r13_c86 bl_86 br_86 wl_13 vdd gnd cell_6t
Xbit_r14_c86 bl_86 br_86 wl_14 vdd gnd cell_6t
Xbit_r15_c86 bl_86 br_86 wl_15 vdd gnd cell_6t
Xbit_r16_c86 bl_86 br_86 wl_16 vdd gnd cell_6t
Xbit_r17_c86 bl_86 br_86 wl_17 vdd gnd cell_6t
Xbit_r18_c86 bl_86 br_86 wl_18 vdd gnd cell_6t
Xbit_r19_c86 bl_86 br_86 wl_19 vdd gnd cell_6t
Xbit_r20_c86 bl_86 br_86 wl_20 vdd gnd cell_6t
Xbit_r21_c86 bl_86 br_86 wl_21 vdd gnd cell_6t
Xbit_r22_c86 bl_86 br_86 wl_22 vdd gnd cell_6t
Xbit_r23_c86 bl_86 br_86 wl_23 vdd gnd cell_6t
Xbit_r24_c86 bl_86 br_86 wl_24 vdd gnd cell_6t
Xbit_r25_c86 bl_86 br_86 wl_25 vdd gnd cell_6t
Xbit_r26_c86 bl_86 br_86 wl_26 vdd gnd cell_6t
Xbit_r27_c86 bl_86 br_86 wl_27 vdd gnd cell_6t
Xbit_r28_c86 bl_86 br_86 wl_28 vdd gnd cell_6t
Xbit_r29_c86 bl_86 br_86 wl_29 vdd gnd cell_6t
Xbit_r30_c86 bl_86 br_86 wl_30 vdd gnd cell_6t
Xbit_r31_c86 bl_86 br_86 wl_31 vdd gnd cell_6t
Xbit_r32_c86 bl_86 br_86 wl_32 vdd gnd cell_6t
Xbit_r33_c86 bl_86 br_86 wl_33 vdd gnd cell_6t
Xbit_r34_c86 bl_86 br_86 wl_34 vdd gnd cell_6t
Xbit_r35_c86 bl_86 br_86 wl_35 vdd gnd cell_6t
Xbit_r36_c86 bl_86 br_86 wl_36 vdd gnd cell_6t
Xbit_r37_c86 bl_86 br_86 wl_37 vdd gnd cell_6t
Xbit_r38_c86 bl_86 br_86 wl_38 vdd gnd cell_6t
Xbit_r39_c86 bl_86 br_86 wl_39 vdd gnd cell_6t
Xbit_r40_c86 bl_86 br_86 wl_40 vdd gnd cell_6t
Xbit_r41_c86 bl_86 br_86 wl_41 vdd gnd cell_6t
Xbit_r42_c86 bl_86 br_86 wl_42 vdd gnd cell_6t
Xbit_r43_c86 bl_86 br_86 wl_43 vdd gnd cell_6t
Xbit_r44_c86 bl_86 br_86 wl_44 vdd gnd cell_6t
Xbit_r45_c86 bl_86 br_86 wl_45 vdd gnd cell_6t
Xbit_r46_c86 bl_86 br_86 wl_46 vdd gnd cell_6t
Xbit_r47_c86 bl_86 br_86 wl_47 vdd gnd cell_6t
Xbit_r48_c86 bl_86 br_86 wl_48 vdd gnd cell_6t
Xbit_r49_c86 bl_86 br_86 wl_49 vdd gnd cell_6t
Xbit_r50_c86 bl_86 br_86 wl_50 vdd gnd cell_6t
Xbit_r51_c86 bl_86 br_86 wl_51 vdd gnd cell_6t
Xbit_r52_c86 bl_86 br_86 wl_52 vdd gnd cell_6t
Xbit_r53_c86 bl_86 br_86 wl_53 vdd gnd cell_6t
Xbit_r54_c86 bl_86 br_86 wl_54 vdd gnd cell_6t
Xbit_r55_c86 bl_86 br_86 wl_55 vdd gnd cell_6t
Xbit_r56_c86 bl_86 br_86 wl_56 vdd gnd cell_6t
Xbit_r57_c86 bl_86 br_86 wl_57 vdd gnd cell_6t
Xbit_r58_c86 bl_86 br_86 wl_58 vdd gnd cell_6t
Xbit_r59_c86 bl_86 br_86 wl_59 vdd gnd cell_6t
Xbit_r60_c86 bl_86 br_86 wl_60 vdd gnd cell_6t
Xbit_r61_c86 bl_86 br_86 wl_61 vdd gnd cell_6t
Xbit_r62_c86 bl_86 br_86 wl_62 vdd gnd cell_6t
Xbit_r63_c86 bl_86 br_86 wl_63 vdd gnd cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd cell_6t
Xbit_r1_c87 bl_87 br_87 wl_1 vdd gnd cell_6t
Xbit_r2_c87 bl_87 br_87 wl_2 vdd gnd cell_6t
Xbit_r3_c87 bl_87 br_87 wl_3 vdd gnd cell_6t
Xbit_r4_c87 bl_87 br_87 wl_4 vdd gnd cell_6t
Xbit_r5_c87 bl_87 br_87 wl_5 vdd gnd cell_6t
Xbit_r6_c87 bl_87 br_87 wl_6 vdd gnd cell_6t
Xbit_r7_c87 bl_87 br_87 wl_7 vdd gnd cell_6t
Xbit_r8_c87 bl_87 br_87 wl_8 vdd gnd cell_6t
Xbit_r9_c87 bl_87 br_87 wl_9 vdd gnd cell_6t
Xbit_r10_c87 bl_87 br_87 wl_10 vdd gnd cell_6t
Xbit_r11_c87 bl_87 br_87 wl_11 vdd gnd cell_6t
Xbit_r12_c87 bl_87 br_87 wl_12 vdd gnd cell_6t
Xbit_r13_c87 bl_87 br_87 wl_13 vdd gnd cell_6t
Xbit_r14_c87 bl_87 br_87 wl_14 vdd gnd cell_6t
Xbit_r15_c87 bl_87 br_87 wl_15 vdd gnd cell_6t
Xbit_r16_c87 bl_87 br_87 wl_16 vdd gnd cell_6t
Xbit_r17_c87 bl_87 br_87 wl_17 vdd gnd cell_6t
Xbit_r18_c87 bl_87 br_87 wl_18 vdd gnd cell_6t
Xbit_r19_c87 bl_87 br_87 wl_19 vdd gnd cell_6t
Xbit_r20_c87 bl_87 br_87 wl_20 vdd gnd cell_6t
Xbit_r21_c87 bl_87 br_87 wl_21 vdd gnd cell_6t
Xbit_r22_c87 bl_87 br_87 wl_22 vdd gnd cell_6t
Xbit_r23_c87 bl_87 br_87 wl_23 vdd gnd cell_6t
Xbit_r24_c87 bl_87 br_87 wl_24 vdd gnd cell_6t
Xbit_r25_c87 bl_87 br_87 wl_25 vdd gnd cell_6t
Xbit_r26_c87 bl_87 br_87 wl_26 vdd gnd cell_6t
Xbit_r27_c87 bl_87 br_87 wl_27 vdd gnd cell_6t
Xbit_r28_c87 bl_87 br_87 wl_28 vdd gnd cell_6t
Xbit_r29_c87 bl_87 br_87 wl_29 vdd gnd cell_6t
Xbit_r30_c87 bl_87 br_87 wl_30 vdd gnd cell_6t
Xbit_r31_c87 bl_87 br_87 wl_31 vdd gnd cell_6t
Xbit_r32_c87 bl_87 br_87 wl_32 vdd gnd cell_6t
Xbit_r33_c87 bl_87 br_87 wl_33 vdd gnd cell_6t
Xbit_r34_c87 bl_87 br_87 wl_34 vdd gnd cell_6t
Xbit_r35_c87 bl_87 br_87 wl_35 vdd gnd cell_6t
Xbit_r36_c87 bl_87 br_87 wl_36 vdd gnd cell_6t
Xbit_r37_c87 bl_87 br_87 wl_37 vdd gnd cell_6t
Xbit_r38_c87 bl_87 br_87 wl_38 vdd gnd cell_6t
Xbit_r39_c87 bl_87 br_87 wl_39 vdd gnd cell_6t
Xbit_r40_c87 bl_87 br_87 wl_40 vdd gnd cell_6t
Xbit_r41_c87 bl_87 br_87 wl_41 vdd gnd cell_6t
Xbit_r42_c87 bl_87 br_87 wl_42 vdd gnd cell_6t
Xbit_r43_c87 bl_87 br_87 wl_43 vdd gnd cell_6t
Xbit_r44_c87 bl_87 br_87 wl_44 vdd gnd cell_6t
Xbit_r45_c87 bl_87 br_87 wl_45 vdd gnd cell_6t
Xbit_r46_c87 bl_87 br_87 wl_46 vdd gnd cell_6t
Xbit_r47_c87 bl_87 br_87 wl_47 vdd gnd cell_6t
Xbit_r48_c87 bl_87 br_87 wl_48 vdd gnd cell_6t
Xbit_r49_c87 bl_87 br_87 wl_49 vdd gnd cell_6t
Xbit_r50_c87 bl_87 br_87 wl_50 vdd gnd cell_6t
Xbit_r51_c87 bl_87 br_87 wl_51 vdd gnd cell_6t
Xbit_r52_c87 bl_87 br_87 wl_52 vdd gnd cell_6t
Xbit_r53_c87 bl_87 br_87 wl_53 vdd gnd cell_6t
Xbit_r54_c87 bl_87 br_87 wl_54 vdd gnd cell_6t
Xbit_r55_c87 bl_87 br_87 wl_55 vdd gnd cell_6t
Xbit_r56_c87 bl_87 br_87 wl_56 vdd gnd cell_6t
Xbit_r57_c87 bl_87 br_87 wl_57 vdd gnd cell_6t
Xbit_r58_c87 bl_87 br_87 wl_58 vdd gnd cell_6t
Xbit_r59_c87 bl_87 br_87 wl_59 vdd gnd cell_6t
Xbit_r60_c87 bl_87 br_87 wl_60 vdd gnd cell_6t
Xbit_r61_c87 bl_87 br_87 wl_61 vdd gnd cell_6t
Xbit_r62_c87 bl_87 br_87 wl_62 vdd gnd cell_6t
Xbit_r63_c87 bl_87 br_87 wl_63 vdd gnd cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd cell_6t
Xbit_r1_c88 bl_88 br_88 wl_1 vdd gnd cell_6t
Xbit_r2_c88 bl_88 br_88 wl_2 vdd gnd cell_6t
Xbit_r3_c88 bl_88 br_88 wl_3 vdd gnd cell_6t
Xbit_r4_c88 bl_88 br_88 wl_4 vdd gnd cell_6t
Xbit_r5_c88 bl_88 br_88 wl_5 vdd gnd cell_6t
Xbit_r6_c88 bl_88 br_88 wl_6 vdd gnd cell_6t
Xbit_r7_c88 bl_88 br_88 wl_7 vdd gnd cell_6t
Xbit_r8_c88 bl_88 br_88 wl_8 vdd gnd cell_6t
Xbit_r9_c88 bl_88 br_88 wl_9 vdd gnd cell_6t
Xbit_r10_c88 bl_88 br_88 wl_10 vdd gnd cell_6t
Xbit_r11_c88 bl_88 br_88 wl_11 vdd gnd cell_6t
Xbit_r12_c88 bl_88 br_88 wl_12 vdd gnd cell_6t
Xbit_r13_c88 bl_88 br_88 wl_13 vdd gnd cell_6t
Xbit_r14_c88 bl_88 br_88 wl_14 vdd gnd cell_6t
Xbit_r15_c88 bl_88 br_88 wl_15 vdd gnd cell_6t
Xbit_r16_c88 bl_88 br_88 wl_16 vdd gnd cell_6t
Xbit_r17_c88 bl_88 br_88 wl_17 vdd gnd cell_6t
Xbit_r18_c88 bl_88 br_88 wl_18 vdd gnd cell_6t
Xbit_r19_c88 bl_88 br_88 wl_19 vdd gnd cell_6t
Xbit_r20_c88 bl_88 br_88 wl_20 vdd gnd cell_6t
Xbit_r21_c88 bl_88 br_88 wl_21 vdd gnd cell_6t
Xbit_r22_c88 bl_88 br_88 wl_22 vdd gnd cell_6t
Xbit_r23_c88 bl_88 br_88 wl_23 vdd gnd cell_6t
Xbit_r24_c88 bl_88 br_88 wl_24 vdd gnd cell_6t
Xbit_r25_c88 bl_88 br_88 wl_25 vdd gnd cell_6t
Xbit_r26_c88 bl_88 br_88 wl_26 vdd gnd cell_6t
Xbit_r27_c88 bl_88 br_88 wl_27 vdd gnd cell_6t
Xbit_r28_c88 bl_88 br_88 wl_28 vdd gnd cell_6t
Xbit_r29_c88 bl_88 br_88 wl_29 vdd gnd cell_6t
Xbit_r30_c88 bl_88 br_88 wl_30 vdd gnd cell_6t
Xbit_r31_c88 bl_88 br_88 wl_31 vdd gnd cell_6t
Xbit_r32_c88 bl_88 br_88 wl_32 vdd gnd cell_6t
Xbit_r33_c88 bl_88 br_88 wl_33 vdd gnd cell_6t
Xbit_r34_c88 bl_88 br_88 wl_34 vdd gnd cell_6t
Xbit_r35_c88 bl_88 br_88 wl_35 vdd gnd cell_6t
Xbit_r36_c88 bl_88 br_88 wl_36 vdd gnd cell_6t
Xbit_r37_c88 bl_88 br_88 wl_37 vdd gnd cell_6t
Xbit_r38_c88 bl_88 br_88 wl_38 vdd gnd cell_6t
Xbit_r39_c88 bl_88 br_88 wl_39 vdd gnd cell_6t
Xbit_r40_c88 bl_88 br_88 wl_40 vdd gnd cell_6t
Xbit_r41_c88 bl_88 br_88 wl_41 vdd gnd cell_6t
Xbit_r42_c88 bl_88 br_88 wl_42 vdd gnd cell_6t
Xbit_r43_c88 bl_88 br_88 wl_43 vdd gnd cell_6t
Xbit_r44_c88 bl_88 br_88 wl_44 vdd gnd cell_6t
Xbit_r45_c88 bl_88 br_88 wl_45 vdd gnd cell_6t
Xbit_r46_c88 bl_88 br_88 wl_46 vdd gnd cell_6t
Xbit_r47_c88 bl_88 br_88 wl_47 vdd gnd cell_6t
Xbit_r48_c88 bl_88 br_88 wl_48 vdd gnd cell_6t
Xbit_r49_c88 bl_88 br_88 wl_49 vdd gnd cell_6t
Xbit_r50_c88 bl_88 br_88 wl_50 vdd gnd cell_6t
Xbit_r51_c88 bl_88 br_88 wl_51 vdd gnd cell_6t
Xbit_r52_c88 bl_88 br_88 wl_52 vdd gnd cell_6t
Xbit_r53_c88 bl_88 br_88 wl_53 vdd gnd cell_6t
Xbit_r54_c88 bl_88 br_88 wl_54 vdd gnd cell_6t
Xbit_r55_c88 bl_88 br_88 wl_55 vdd gnd cell_6t
Xbit_r56_c88 bl_88 br_88 wl_56 vdd gnd cell_6t
Xbit_r57_c88 bl_88 br_88 wl_57 vdd gnd cell_6t
Xbit_r58_c88 bl_88 br_88 wl_58 vdd gnd cell_6t
Xbit_r59_c88 bl_88 br_88 wl_59 vdd gnd cell_6t
Xbit_r60_c88 bl_88 br_88 wl_60 vdd gnd cell_6t
Xbit_r61_c88 bl_88 br_88 wl_61 vdd gnd cell_6t
Xbit_r62_c88 bl_88 br_88 wl_62 vdd gnd cell_6t
Xbit_r63_c88 bl_88 br_88 wl_63 vdd gnd cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd cell_6t
Xbit_r1_c89 bl_89 br_89 wl_1 vdd gnd cell_6t
Xbit_r2_c89 bl_89 br_89 wl_2 vdd gnd cell_6t
Xbit_r3_c89 bl_89 br_89 wl_3 vdd gnd cell_6t
Xbit_r4_c89 bl_89 br_89 wl_4 vdd gnd cell_6t
Xbit_r5_c89 bl_89 br_89 wl_5 vdd gnd cell_6t
Xbit_r6_c89 bl_89 br_89 wl_6 vdd gnd cell_6t
Xbit_r7_c89 bl_89 br_89 wl_7 vdd gnd cell_6t
Xbit_r8_c89 bl_89 br_89 wl_8 vdd gnd cell_6t
Xbit_r9_c89 bl_89 br_89 wl_9 vdd gnd cell_6t
Xbit_r10_c89 bl_89 br_89 wl_10 vdd gnd cell_6t
Xbit_r11_c89 bl_89 br_89 wl_11 vdd gnd cell_6t
Xbit_r12_c89 bl_89 br_89 wl_12 vdd gnd cell_6t
Xbit_r13_c89 bl_89 br_89 wl_13 vdd gnd cell_6t
Xbit_r14_c89 bl_89 br_89 wl_14 vdd gnd cell_6t
Xbit_r15_c89 bl_89 br_89 wl_15 vdd gnd cell_6t
Xbit_r16_c89 bl_89 br_89 wl_16 vdd gnd cell_6t
Xbit_r17_c89 bl_89 br_89 wl_17 vdd gnd cell_6t
Xbit_r18_c89 bl_89 br_89 wl_18 vdd gnd cell_6t
Xbit_r19_c89 bl_89 br_89 wl_19 vdd gnd cell_6t
Xbit_r20_c89 bl_89 br_89 wl_20 vdd gnd cell_6t
Xbit_r21_c89 bl_89 br_89 wl_21 vdd gnd cell_6t
Xbit_r22_c89 bl_89 br_89 wl_22 vdd gnd cell_6t
Xbit_r23_c89 bl_89 br_89 wl_23 vdd gnd cell_6t
Xbit_r24_c89 bl_89 br_89 wl_24 vdd gnd cell_6t
Xbit_r25_c89 bl_89 br_89 wl_25 vdd gnd cell_6t
Xbit_r26_c89 bl_89 br_89 wl_26 vdd gnd cell_6t
Xbit_r27_c89 bl_89 br_89 wl_27 vdd gnd cell_6t
Xbit_r28_c89 bl_89 br_89 wl_28 vdd gnd cell_6t
Xbit_r29_c89 bl_89 br_89 wl_29 vdd gnd cell_6t
Xbit_r30_c89 bl_89 br_89 wl_30 vdd gnd cell_6t
Xbit_r31_c89 bl_89 br_89 wl_31 vdd gnd cell_6t
Xbit_r32_c89 bl_89 br_89 wl_32 vdd gnd cell_6t
Xbit_r33_c89 bl_89 br_89 wl_33 vdd gnd cell_6t
Xbit_r34_c89 bl_89 br_89 wl_34 vdd gnd cell_6t
Xbit_r35_c89 bl_89 br_89 wl_35 vdd gnd cell_6t
Xbit_r36_c89 bl_89 br_89 wl_36 vdd gnd cell_6t
Xbit_r37_c89 bl_89 br_89 wl_37 vdd gnd cell_6t
Xbit_r38_c89 bl_89 br_89 wl_38 vdd gnd cell_6t
Xbit_r39_c89 bl_89 br_89 wl_39 vdd gnd cell_6t
Xbit_r40_c89 bl_89 br_89 wl_40 vdd gnd cell_6t
Xbit_r41_c89 bl_89 br_89 wl_41 vdd gnd cell_6t
Xbit_r42_c89 bl_89 br_89 wl_42 vdd gnd cell_6t
Xbit_r43_c89 bl_89 br_89 wl_43 vdd gnd cell_6t
Xbit_r44_c89 bl_89 br_89 wl_44 vdd gnd cell_6t
Xbit_r45_c89 bl_89 br_89 wl_45 vdd gnd cell_6t
Xbit_r46_c89 bl_89 br_89 wl_46 vdd gnd cell_6t
Xbit_r47_c89 bl_89 br_89 wl_47 vdd gnd cell_6t
Xbit_r48_c89 bl_89 br_89 wl_48 vdd gnd cell_6t
Xbit_r49_c89 bl_89 br_89 wl_49 vdd gnd cell_6t
Xbit_r50_c89 bl_89 br_89 wl_50 vdd gnd cell_6t
Xbit_r51_c89 bl_89 br_89 wl_51 vdd gnd cell_6t
Xbit_r52_c89 bl_89 br_89 wl_52 vdd gnd cell_6t
Xbit_r53_c89 bl_89 br_89 wl_53 vdd gnd cell_6t
Xbit_r54_c89 bl_89 br_89 wl_54 vdd gnd cell_6t
Xbit_r55_c89 bl_89 br_89 wl_55 vdd gnd cell_6t
Xbit_r56_c89 bl_89 br_89 wl_56 vdd gnd cell_6t
Xbit_r57_c89 bl_89 br_89 wl_57 vdd gnd cell_6t
Xbit_r58_c89 bl_89 br_89 wl_58 vdd gnd cell_6t
Xbit_r59_c89 bl_89 br_89 wl_59 vdd gnd cell_6t
Xbit_r60_c89 bl_89 br_89 wl_60 vdd gnd cell_6t
Xbit_r61_c89 bl_89 br_89 wl_61 vdd gnd cell_6t
Xbit_r62_c89 bl_89 br_89 wl_62 vdd gnd cell_6t
Xbit_r63_c89 bl_89 br_89 wl_63 vdd gnd cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd cell_6t
Xbit_r1_c90 bl_90 br_90 wl_1 vdd gnd cell_6t
Xbit_r2_c90 bl_90 br_90 wl_2 vdd gnd cell_6t
Xbit_r3_c90 bl_90 br_90 wl_3 vdd gnd cell_6t
Xbit_r4_c90 bl_90 br_90 wl_4 vdd gnd cell_6t
Xbit_r5_c90 bl_90 br_90 wl_5 vdd gnd cell_6t
Xbit_r6_c90 bl_90 br_90 wl_6 vdd gnd cell_6t
Xbit_r7_c90 bl_90 br_90 wl_7 vdd gnd cell_6t
Xbit_r8_c90 bl_90 br_90 wl_8 vdd gnd cell_6t
Xbit_r9_c90 bl_90 br_90 wl_9 vdd gnd cell_6t
Xbit_r10_c90 bl_90 br_90 wl_10 vdd gnd cell_6t
Xbit_r11_c90 bl_90 br_90 wl_11 vdd gnd cell_6t
Xbit_r12_c90 bl_90 br_90 wl_12 vdd gnd cell_6t
Xbit_r13_c90 bl_90 br_90 wl_13 vdd gnd cell_6t
Xbit_r14_c90 bl_90 br_90 wl_14 vdd gnd cell_6t
Xbit_r15_c90 bl_90 br_90 wl_15 vdd gnd cell_6t
Xbit_r16_c90 bl_90 br_90 wl_16 vdd gnd cell_6t
Xbit_r17_c90 bl_90 br_90 wl_17 vdd gnd cell_6t
Xbit_r18_c90 bl_90 br_90 wl_18 vdd gnd cell_6t
Xbit_r19_c90 bl_90 br_90 wl_19 vdd gnd cell_6t
Xbit_r20_c90 bl_90 br_90 wl_20 vdd gnd cell_6t
Xbit_r21_c90 bl_90 br_90 wl_21 vdd gnd cell_6t
Xbit_r22_c90 bl_90 br_90 wl_22 vdd gnd cell_6t
Xbit_r23_c90 bl_90 br_90 wl_23 vdd gnd cell_6t
Xbit_r24_c90 bl_90 br_90 wl_24 vdd gnd cell_6t
Xbit_r25_c90 bl_90 br_90 wl_25 vdd gnd cell_6t
Xbit_r26_c90 bl_90 br_90 wl_26 vdd gnd cell_6t
Xbit_r27_c90 bl_90 br_90 wl_27 vdd gnd cell_6t
Xbit_r28_c90 bl_90 br_90 wl_28 vdd gnd cell_6t
Xbit_r29_c90 bl_90 br_90 wl_29 vdd gnd cell_6t
Xbit_r30_c90 bl_90 br_90 wl_30 vdd gnd cell_6t
Xbit_r31_c90 bl_90 br_90 wl_31 vdd gnd cell_6t
Xbit_r32_c90 bl_90 br_90 wl_32 vdd gnd cell_6t
Xbit_r33_c90 bl_90 br_90 wl_33 vdd gnd cell_6t
Xbit_r34_c90 bl_90 br_90 wl_34 vdd gnd cell_6t
Xbit_r35_c90 bl_90 br_90 wl_35 vdd gnd cell_6t
Xbit_r36_c90 bl_90 br_90 wl_36 vdd gnd cell_6t
Xbit_r37_c90 bl_90 br_90 wl_37 vdd gnd cell_6t
Xbit_r38_c90 bl_90 br_90 wl_38 vdd gnd cell_6t
Xbit_r39_c90 bl_90 br_90 wl_39 vdd gnd cell_6t
Xbit_r40_c90 bl_90 br_90 wl_40 vdd gnd cell_6t
Xbit_r41_c90 bl_90 br_90 wl_41 vdd gnd cell_6t
Xbit_r42_c90 bl_90 br_90 wl_42 vdd gnd cell_6t
Xbit_r43_c90 bl_90 br_90 wl_43 vdd gnd cell_6t
Xbit_r44_c90 bl_90 br_90 wl_44 vdd gnd cell_6t
Xbit_r45_c90 bl_90 br_90 wl_45 vdd gnd cell_6t
Xbit_r46_c90 bl_90 br_90 wl_46 vdd gnd cell_6t
Xbit_r47_c90 bl_90 br_90 wl_47 vdd gnd cell_6t
Xbit_r48_c90 bl_90 br_90 wl_48 vdd gnd cell_6t
Xbit_r49_c90 bl_90 br_90 wl_49 vdd gnd cell_6t
Xbit_r50_c90 bl_90 br_90 wl_50 vdd gnd cell_6t
Xbit_r51_c90 bl_90 br_90 wl_51 vdd gnd cell_6t
Xbit_r52_c90 bl_90 br_90 wl_52 vdd gnd cell_6t
Xbit_r53_c90 bl_90 br_90 wl_53 vdd gnd cell_6t
Xbit_r54_c90 bl_90 br_90 wl_54 vdd gnd cell_6t
Xbit_r55_c90 bl_90 br_90 wl_55 vdd gnd cell_6t
Xbit_r56_c90 bl_90 br_90 wl_56 vdd gnd cell_6t
Xbit_r57_c90 bl_90 br_90 wl_57 vdd gnd cell_6t
Xbit_r58_c90 bl_90 br_90 wl_58 vdd gnd cell_6t
Xbit_r59_c90 bl_90 br_90 wl_59 vdd gnd cell_6t
Xbit_r60_c90 bl_90 br_90 wl_60 vdd gnd cell_6t
Xbit_r61_c90 bl_90 br_90 wl_61 vdd gnd cell_6t
Xbit_r62_c90 bl_90 br_90 wl_62 vdd gnd cell_6t
Xbit_r63_c90 bl_90 br_90 wl_63 vdd gnd cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd cell_6t
Xbit_r1_c91 bl_91 br_91 wl_1 vdd gnd cell_6t
Xbit_r2_c91 bl_91 br_91 wl_2 vdd gnd cell_6t
Xbit_r3_c91 bl_91 br_91 wl_3 vdd gnd cell_6t
Xbit_r4_c91 bl_91 br_91 wl_4 vdd gnd cell_6t
Xbit_r5_c91 bl_91 br_91 wl_5 vdd gnd cell_6t
Xbit_r6_c91 bl_91 br_91 wl_6 vdd gnd cell_6t
Xbit_r7_c91 bl_91 br_91 wl_7 vdd gnd cell_6t
Xbit_r8_c91 bl_91 br_91 wl_8 vdd gnd cell_6t
Xbit_r9_c91 bl_91 br_91 wl_9 vdd gnd cell_6t
Xbit_r10_c91 bl_91 br_91 wl_10 vdd gnd cell_6t
Xbit_r11_c91 bl_91 br_91 wl_11 vdd gnd cell_6t
Xbit_r12_c91 bl_91 br_91 wl_12 vdd gnd cell_6t
Xbit_r13_c91 bl_91 br_91 wl_13 vdd gnd cell_6t
Xbit_r14_c91 bl_91 br_91 wl_14 vdd gnd cell_6t
Xbit_r15_c91 bl_91 br_91 wl_15 vdd gnd cell_6t
Xbit_r16_c91 bl_91 br_91 wl_16 vdd gnd cell_6t
Xbit_r17_c91 bl_91 br_91 wl_17 vdd gnd cell_6t
Xbit_r18_c91 bl_91 br_91 wl_18 vdd gnd cell_6t
Xbit_r19_c91 bl_91 br_91 wl_19 vdd gnd cell_6t
Xbit_r20_c91 bl_91 br_91 wl_20 vdd gnd cell_6t
Xbit_r21_c91 bl_91 br_91 wl_21 vdd gnd cell_6t
Xbit_r22_c91 bl_91 br_91 wl_22 vdd gnd cell_6t
Xbit_r23_c91 bl_91 br_91 wl_23 vdd gnd cell_6t
Xbit_r24_c91 bl_91 br_91 wl_24 vdd gnd cell_6t
Xbit_r25_c91 bl_91 br_91 wl_25 vdd gnd cell_6t
Xbit_r26_c91 bl_91 br_91 wl_26 vdd gnd cell_6t
Xbit_r27_c91 bl_91 br_91 wl_27 vdd gnd cell_6t
Xbit_r28_c91 bl_91 br_91 wl_28 vdd gnd cell_6t
Xbit_r29_c91 bl_91 br_91 wl_29 vdd gnd cell_6t
Xbit_r30_c91 bl_91 br_91 wl_30 vdd gnd cell_6t
Xbit_r31_c91 bl_91 br_91 wl_31 vdd gnd cell_6t
Xbit_r32_c91 bl_91 br_91 wl_32 vdd gnd cell_6t
Xbit_r33_c91 bl_91 br_91 wl_33 vdd gnd cell_6t
Xbit_r34_c91 bl_91 br_91 wl_34 vdd gnd cell_6t
Xbit_r35_c91 bl_91 br_91 wl_35 vdd gnd cell_6t
Xbit_r36_c91 bl_91 br_91 wl_36 vdd gnd cell_6t
Xbit_r37_c91 bl_91 br_91 wl_37 vdd gnd cell_6t
Xbit_r38_c91 bl_91 br_91 wl_38 vdd gnd cell_6t
Xbit_r39_c91 bl_91 br_91 wl_39 vdd gnd cell_6t
Xbit_r40_c91 bl_91 br_91 wl_40 vdd gnd cell_6t
Xbit_r41_c91 bl_91 br_91 wl_41 vdd gnd cell_6t
Xbit_r42_c91 bl_91 br_91 wl_42 vdd gnd cell_6t
Xbit_r43_c91 bl_91 br_91 wl_43 vdd gnd cell_6t
Xbit_r44_c91 bl_91 br_91 wl_44 vdd gnd cell_6t
Xbit_r45_c91 bl_91 br_91 wl_45 vdd gnd cell_6t
Xbit_r46_c91 bl_91 br_91 wl_46 vdd gnd cell_6t
Xbit_r47_c91 bl_91 br_91 wl_47 vdd gnd cell_6t
Xbit_r48_c91 bl_91 br_91 wl_48 vdd gnd cell_6t
Xbit_r49_c91 bl_91 br_91 wl_49 vdd gnd cell_6t
Xbit_r50_c91 bl_91 br_91 wl_50 vdd gnd cell_6t
Xbit_r51_c91 bl_91 br_91 wl_51 vdd gnd cell_6t
Xbit_r52_c91 bl_91 br_91 wl_52 vdd gnd cell_6t
Xbit_r53_c91 bl_91 br_91 wl_53 vdd gnd cell_6t
Xbit_r54_c91 bl_91 br_91 wl_54 vdd gnd cell_6t
Xbit_r55_c91 bl_91 br_91 wl_55 vdd gnd cell_6t
Xbit_r56_c91 bl_91 br_91 wl_56 vdd gnd cell_6t
Xbit_r57_c91 bl_91 br_91 wl_57 vdd gnd cell_6t
Xbit_r58_c91 bl_91 br_91 wl_58 vdd gnd cell_6t
Xbit_r59_c91 bl_91 br_91 wl_59 vdd gnd cell_6t
Xbit_r60_c91 bl_91 br_91 wl_60 vdd gnd cell_6t
Xbit_r61_c91 bl_91 br_91 wl_61 vdd gnd cell_6t
Xbit_r62_c91 bl_91 br_91 wl_62 vdd gnd cell_6t
Xbit_r63_c91 bl_91 br_91 wl_63 vdd gnd cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd cell_6t
Xbit_r1_c92 bl_92 br_92 wl_1 vdd gnd cell_6t
Xbit_r2_c92 bl_92 br_92 wl_2 vdd gnd cell_6t
Xbit_r3_c92 bl_92 br_92 wl_3 vdd gnd cell_6t
Xbit_r4_c92 bl_92 br_92 wl_4 vdd gnd cell_6t
Xbit_r5_c92 bl_92 br_92 wl_5 vdd gnd cell_6t
Xbit_r6_c92 bl_92 br_92 wl_6 vdd gnd cell_6t
Xbit_r7_c92 bl_92 br_92 wl_7 vdd gnd cell_6t
Xbit_r8_c92 bl_92 br_92 wl_8 vdd gnd cell_6t
Xbit_r9_c92 bl_92 br_92 wl_9 vdd gnd cell_6t
Xbit_r10_c92 bl_92 br_92 wl_10 vdd gnd cell_6t
Xbit_r11_c92 bl_92 br_92 wl_11 vdd gnd cell_6t
Xbit_r12_c92 bl_92 br_92 wl_12 vdd gnd cell_6t
Xbit_r13_c92 bl_92 br_92 wl_13 vdd gnd cell_6t
Xbit_r14_c92 bl_92 br_92 wl_14 vdd gnd cell_6t
Xbit_r15_c92 bl_92 br_92 wl_15 vdd gnd cell_6t
Xbit_r16_c92 bl_92 br_92 wl_16 vdd gnd cell_6t
Xbit_r17_c92 bl_92 br_92 wl_17 vdd gnd cell_6t
Xbit_r18_c92 bl_92 br_92 wl_18 vdd gnd cell_6t
Xbit_r19_c92 bl_92 br_92 wl_19 vdd gnd cell_6t
Xbit_r20_c92 bl_92 br_92 wl_20 vdd gnd cell_6t
Xbit_r21_c92 bl_92 br_92 wl_21 vdd gnd cell_6t
Xbit_r22_c92 bl_92 br_92 wl_22 vdd gnd cell_6t
Xbit_r23_c92 bl_92 br_92 wl_23 vdd gnd cell_6t
Xbit_r24_c92 bl_92 br_92 wl_24 vdd gnd cell_6t
Xbit_r25_c92 bl_92 br_92 wl_25 vdd gnd cell_6t
Xbit_r26_c92 bl_92 br_92 wl_26 vdd gnd cell_6t
Xbit_r27_c92 bl_92 br_92 wl_27 vdd gnd cell_6t
Xbit_r28_c92 bl_92 br_92 wl_28 vdd gnd cell_6t
Xbit_r29_c92 bl_92 br_92 wl_29 vdd gnd cell_6t
Xbit_r30_c92 bl_92 br_92 wl_30 vdd gnd cell_6t
Xbit_r31_c92 bl_92 br_92 wl_31 vdd gnd cell_6t
Xbit_r32_c92 bl_92 br_92 wl_32 vdd gnd cell_6t
Xbit_r33_c92 bl_92 br_92 wl_33 vdd gnd cell_6t
Xbit_r34_c92 bl_92 br_92 wl_34 vdd gnd cell_6t
Xbit_r35_c92 bl_92 br_92 wl_35 vdd gnd cell_6t
Xbit_r36_c92 bl_92 br_92 wl_36 vdd gnd cell_6t
Xbit_r37_c92 bl_92 br_92 wl_37 vdd gnd cell_6t
Xbit_r38_c92 bl_92 br_92 wl_38 vdd gnd cell_6t
Xbit_r39_c92 bl_92 br_92 wl_39 vdd gnd cell_6t
Xbit_r40_c92 bl_92 br_92 wl_40 vdd gnd cell_6t
Xbit_r41_c92 bl_92 br_92 wl_41 vdd gnd cell_6t
Xbit_r42_c92 bl_92 br_92 wl_42 vdd gnd cell_6t
Xbit_r43_c92 bl_92 br_92 wl_43 vdd gnd cell_6t
Xbit_r44_c92 bl_92 br_92 wl_44 vdd gnd cell_6t
Xbit_r45_c92 bl_92 br_92 wl_45 vdd gnd cell_6t
Xbit_r46_c92 bl_92 br_92 wl_46 vdd gnd cell_6t
Xbit_r47_c92 bl_92 br_92 wl_47 vdd gnd cell_6t
Xbit_r48_c92 bl_92 br_92 wl_48 vdd gnd cell_6t
Xbit_r49_c92 bl_92 br_92 wl_49 vdd gnd cell_6t
Xbit_r50_c92 bl_92 br_92 wl_50 vdd gnd cell_6t
Xbit_r51_c92 bl_92 br_92 wl_51 vdd gnd cell_6t
Xbit_r52_c92 bl_92 br_92 wl_52 vdd gnd cell_6t
Xbit_r53_c92 bl_92 br_92 wl_53 vdd gnd cell_6t
Xbit_r54_c92 bl_92 br_92 wl_54 vdd gnd cell_6t
Xbit_r55_c92 bl_92 br_92 wl_55 vdd gnd cell_6t
Xbit_r56_c92 bl_92 br_92 wl_56 vdd gnd cell_6t
Xbit_r57_c92 bl_92 br_92 wl_57 vdd gnd cell_6t
Xbit_r58_c92 bl_92 br_92 wl_58 vdd gnd cell_6t
Xbit_r59_c92 bl_92 br_92 wl_59 vdd gnd cell_6t
Xbit_r60_c92 bl_92 br_92 wl_60 vdd gnd cell_6t
Xbit_r61_c92 bl_92 br_92 wl_61 vdd gnd cell_6t
Xbit_r62_c92 bl_92 br_92 wl_62 vdd gnd cell_6t
Xbit_r63_c92 bl_92 br_92 wl_63 vdd gnd cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd cell_6t
Xbit_r1_c93 bl_93 br_93 wl_1 vdd gnd cell_6t
Xbit_r2_c93 bl_93 br_93 wl_2 vdd gnd cell_6t
Xbit_r3_c93 bl_93 br_93 wl_3 vdd gnd cell_6t
Xbit_r4_c93 bl_93 br_93 wl_4 vdd gnd cell_6t
Xbit_r5_c93 bl_93 br_93 wl_5 vdd gnd cell_6t
Xbit_r6_c93 bl_93 br_93 wl_6 vdd gnd cell_6t
Xbit_r7_c93 bl_93 br_93 wl_7 vdd gnd cell_6t
Xbit_r8_c93 bl_93 br_93 wl_8 vdd gnd cell_6t
Xbit_r9_c93 bl_93 br_93 wl_9 vdd gnd cell_6t
Xbit_r10_c93 bl_93 br_93 wl_10 vdd gnd cell_6t
Xbit_r11_c93 bl_93 br_93 wl_11 vdd gnd cell_6t
Xbit_r12_c93 bl_93 br_93 wl_12 vdd gnd cell_6t
Xbit_r13_c93 bl_93 br_93 wl_13 vdd gnd cell_6t
Xbit_r14_c93 bl_93 br_93 wl_14 vdd gnd cell_6t
Xbit_r15_c93 bl_93 br_93 wl_15 vdd gnd cell_6t
Xbit_r16_c93 bl_93 br_93 wl_16 vdd gnd cell_6t
Xbit_r17_c93 bl_93 br_93 wl_17 vdd gnd cell_6t
Xbit_r18_c93 bl_93 br_93 wl_18 vdd gnd cell_6t
Xbit_r19_c93 bl_93 br_93 wl_19 vdd gnd cell_6t
Xbit_r20_c93 bl_93 br_93 wl_20 vdd gnd cell_6t
Xbit_r21_c93 bl_93 br_93 wl_21 vdd gnd cell_6t
Xbit_r22_c93 bl_93 br_93 wl_22 vdd gnd cell_6t
Xbit_r23_c93 bl_93 br_93 wl_23 vdd gnd cell_6t
Xbit_r24_c93 bl_93 br_93 wl_24 vdd gnd cell_6t
Xbit_r25_c93 bl_93 br_93 wl_25 vdd gnd cell_6t
Xbit_r26_c93 bl_93 br_93 wl_26 vdd gnd cell_6t
Xbit_r27_c93 bl_93 br_93 wl_27 vdd gnd cell_6t
Xbit_r28_c93 bl_93 br_93 wl_28 vdd gnd cell_6t
Xbit_r29_c93 bl_93 br_93 wl_29 vdd gnd cell_6t
Xbit_r30_c93 bl_93 br_93 wl_30 vdd gnd cell_6t
Xbit_r31_c93 bl_93 br_93 wl_31 vdd gnd cell_6t
Xbit_r32_c93 bl_93 br_93 wl_32 vdd gnd cell_6t
Xbit_r33_c93 bl_93 br_93 wl_33 vdd gnd cell_6t
Xbit_r34_c93 bl_93 br_93 wl_34 vdd gnd cell_6t
Xbit_r35_c93 bl_93 br_93 wl_35 vdd gnd cell_6t
Xbit_r36_c93 bl_93 br_93 wl_36 vdd gnd cell_6t
Xbit_r37_c93 bl_93 br_93 wl_37 vdd gnd cell_6t
Xbit_r38_c93 bl_93 br_93 wl_38 vdd gnd cell_6t
Xbit_r39_c93 bl_93 br_93 wl_39 vdd gnd cell_6t
Xbit_r40_c93 bl_93 br_93 wl_40 vdd gnd cell_6t
Xbit_r41_c93 bl_93 br_93 wl_41 vdd gnd cell_6t
Xbit_r42_c93 bl_93 br_93 wl_42 vdd gnd cell_6t
Xbit_r43_c93 bl_93 br_93 wl_43 vdd gnd cell_6t
Xbit_r44_c93 bl_93 br_93 wl_44 vdd gnd cell_6t
Xbit_r45_c93 bl_93 br_93 wl_45 vdd gnd cell_6t
Xbit_r46_c93 bl_93 br_93 wl_46 vdd gnd cell_6t
Xbit_r47_c93 bl_93 br_93 wl_47 vdd gnd cell_6t
Xbit_r48_c93 bl_93 br_93 wl_48 vdd gnd cell_6t
Xbit_r49_c93 bl_93 br_93 wl_49 vdd gnd cell_6t
Xbit_r50_c93 bl_93 br_93 wl_50 vdd gnd cell_6t
Xbit_r51_c93 bl_93 br_93 wl_51 vdd gnd cell_6t
Xbit_r52_c93 bl_93 br_93 wl_52 vdd gnd cell_6t
Xbit_r53_c93 bl_93 br_93 wl_53 vdd gnd cell_6t
Xbit_r54_c93 bl_93 br_93 wl_54 vdd gnd cell_6t
Xbit_r55_c93 bl_93 br_93 wl_55 vdd gnd cell_6t
Xbit_r56_c93 bl_93 br_93 wl_56 vdd gnd cell_6t
Xbit_r57_c93 bl_93 br_93 wl_57 vdd gnd cell_6t
Xbit_r58_c93 bl_93 br_93 wl_58 vdd gnd cell_6t
Xbit_r59_c93 bl_93 br_93 wl_59 vdd gnd cell_6t
Xbit_r60_c93 bl_93 br_93 wl_60 vdd gnd cell_6t
Xbit_r61_c93 bl_93 br_93 wl_61 vdd gnd cell_6t
Xbit_r62_c93 bl_93 br_93 wl_62 vdd gnd cell_6t
Xbit_r63_c93 bl_93 br_93 wl_63 vdd gnd cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd cell_6t
Xbit_r1_c94 bl_94 br_94 wl_1 vdd gnd cell_6t
Xbit_r2_c94 bl_94 br_94 wl_2 vdd gnd cell_6t
Xbit_r3_c94 bl_94 br_94 wl_3 vdd gnd cell_6t
Xbit_r4_c94 bl_94 br_94 wl_4 vdd gnd cell_6t
Xbit_r5_c94 bl_94 br_94 wl_5 vdd gnd cell_6t
Xbit_r6_c94 bl_94 br_94 wl_6 vdd gnd cell_6t
Xbit_r7_c94 bl_94 br_94 wl_7 vdd gnd cell_6t
Xbit_r8_c94 bl_94 br_94 wl_8 vdd gnd cell_6t
Xbit_r9_c94 bl_94 br_94 wl_9 vdd gnd cell_6t
Xbit_r10_c94 bl_94 br_94 wl_10 vdd gnd cell_6t
Xbit_r11_c94 bl_94 br_94 wl_11 vdd gnd cell_6t
Xbit_r12_c94 bl_94 br_94 wl_12 vdd gnd cell_6t
Xbit_r13_c94 bl_94 br_94 wl_13 vdd gnd cell_6t
Xbit_r14_c94 bl_94 br_94 wl_14 vdd gnd cell_6t
Xbit_r15_c94 bl_94 br_94 wl_15 vdd gnd cell_6t
Xbit_r16_c94 bl_94 br_94 wl_16 vdd gnd cell_6t
Xbit_r17_c94 bl_94 br_94 wl_17 vdd gnd cell_6t
Xbit_r18_c94 bl_94 br_94 wl_18 vdd gnd cell_6t
Xbit_r19_c94 bl_94 br_94 wl_19 vdd gnd cell_6t
Xbit_r20_c94 bl_94 br_94 wl_20 vdd gnd cell_6t
Xbit_r21_c94 bl_94 br_94 wl_21 vdd gnd cell_6t
Xbit_r22_c94 bl_94 br_94 wl_22 vdd gnd cell_6t
Xbit_r23_c94 bl_94 br_94 wl_23 vdd gnd cell_6t
Xbit_r24_c94 bl_94 br_94 wl_24 vdd gnd cell_6t
Xbit_r25_c94 bl_94 br_94 wl_25 vdd gnd cell_6t
Xbit_r26_c94 bl_94 br_94 wl_26 vdd gnd cell_6t
Xbit_r27_c94 bl_94 br_94 wl_27 vdd gnd cell_6t
Xbit_r28_c94 bl_94 br_94 wl_28 vdd gnd cell_6t
Xbit_r29_c94 bl_94 br_94 wl_29 vdd gnd cell_6t
Xbit_r30_c94 bl_94 br_94 wl_30 vdd gnd cell_6t
Xbit_r31_c94 bl_94 br_94 wl_31 vdd gnd cell_6t
Xbit_r32_c94 bl_94 br_94 wl_32 vdd gnd cell_6t
Xbit_r33_c94 bl_94 br_94 wl_33 vdd gnd cell_6t
Xbit_r34_c94 bl_94 br_94 wl_34 vdd gnd cell_6t
Xbit_r35_c94 bl_94 br_94 wl_35 vdd gnd cell_6t
Xbit_r36_c94 bl_94 br_94 wl_36 vdd gnd cell_6t
Xbit_r37_c94 bl_94 br_94 wl_37 vdd gnd cell_6t
Xbit_r38_c94 bl_94 br_94 wl_38 vdd gnd cell_6t
Xbit_r39_c94 bl_94 br_94 wl_39 vdd gnd cell_6t
Xbit_r40_c94 bl_94 br_94 wl_40 vdd gnd cell_6t
Xbit_r41_c94 bl_94 br_94 wl_41 vdd gnd cell_6t
Xbit_r42_c94 bl_94 br_94 wl_42 vdd gnd cell_6t
Xbit_r43_c94 bl_94 br_94 wl_43 vdd gnd cell_6t
Xbit_r44_c94 bl_94 br_94 wl_44 vdd gnd cell_6t
Xbit_r45_c94 bl_94 br_94 wl_45 vdd gnd cell_6t
Xbit_r46_c94 bl_94 br_94 wl_46 vdd gnd cell_6t
Xbit_r47_c94 bl_94 br_94 wl_47 vdd gnd cell_6t
Xbit_r48_c94 bl_94 br_94 wl_48 vdd gnd cell_6t
Xbit_r49_c94 bl_94 br_94 wl_49 vdd gnd cell_6t
Xbit_r50_c94 bl_94 br_94 wl_50 vdd gnd cell_6t
Xbit_r51_c94 bl_94 br_94 wl_51 vdd gnd cell_6t
Xbit_r52_c94 bl_94 br_94 wl_52 vdd gnd cell_6t
Xbit_r53_c94 bl_94 br_94 wl_53 vdd gnd cell_6t
Xbit_r54_c94 bl_94 br_94 wl_54 vdd gnd cell_6t
Xbit_r55_c94 bl_94 br_94 wl_55 vdd gnd cell_6t
Xbit_r56_c94 bl_94 br_94 wl_56 vdd gnd cell_6t
Xbit_r57_c94 bl_94 br_94 wl_57 vdd gnd cell_6t
Xbit_r58_c94 bl_94 br_94 wl_58 vdd gnd cell_6t
Xbit_r59_c94 bl_94 br_94 wl_59 vdd gnd cell_6t
Xbit_r60_c94 bl_94 br_94 wl_60 vdd gnd cell_6t
Xbit_r61_c94 bl_94 br_94 wl_61 vdd gnd cell_6t
Xbit_r62_c94 bl_94 br_94 wl_62 vdd gnd cell_6t
Xbit_r63_c94 bl_94 br_94 wl_63 vdd gnd cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd cell_6t
Xbit_r1_c95 bl_95 br_95 wl_1 vdd gnd cell_6t
Xbit_r2_c95 bl_95 br_95 wl_2 vdd gnd cell_6t
Xbit_r3_c95 bl_95 br_95 wl_3 vdd gnd cell_6t
Xbit_r4_c95 bl_95 br_95 wl_4 vdd gnd cell_6t
Xbit_r5_c95 bl_95 br_95 wl_5 vdd gnd cell_6t
Xbit_r6_c95 bl_95 br_95 wl_6 vdd gnd cell_6t
Xbit_r7_c95 bl_95 br_95 wl_7 vdd gnd cell_6t
Xbit_r8_c95 bl_95 br_95 wl_8 vdd gnd cell_6t
Xbit_r9_c95 bl_95 br_95 wl_9 vdd gnd cell_6t
Xbit_r10_c95 bl_95 br_95 wl_10 vdd gnd cell_6t
Xbit_r11_c95 bl_95 br_95 wl_11 vdd gnd cell_6t
Xbit_r12_c95 bl_95 br_95 wl_12 vdd gnd cell_6t
Xbit_r13_c95 bl_95 br_95 wl_13 vdd gnd cell_6t
Xbit_r14_c95 bl_95 br_95 wl_14 vdd gnd cell_6t
Xbit_r15_c95 bl_95 br_95 wl_15 vdd gnd cell_6t
Xbit_r16_c95 bl_95 br_95 wl_16 vdd gnd cell_6t
Xbit_r17_c95 bl_95 br_95 wl_17 vdd gnd cell_6t
Xbit_r18_c95 bl_95 br_95 wl_18 vdd gnd cell_6t
Xbit_r19_c95 bl_95 br_95 wl_19 vdd gnd cell_6t
Xbit_r20_c95 bl_95 br_95 wl_20 vdd gnd cell_6t
Xbit_r21_c95 bl_95 br_95 wl_21 vdd gnd cell_6t
Xbit_r22_c95 bl_95 br_95 wl_22 vdd gnd cell_6t
Xbit_r23_c95 bl_95 br_95 wl_23 vdd gnd cell_6t
Xbit_r24_c95 bl_95 br_95 wl_24 vdd gnd cell_6t
Xbit_r25_c95 bl_95 br_95 wl_25 vdd gnd cell_6t
Xbit_r26_c95 bl_95 br_95 wl_26 vdd gnd cell_6t
Xbit_r27_c95 bl_95 br_95 wl_27 vdd gnd cell_6t
Xbit_r28_c95 bl_95 br_95 wl_28 vdd gnd cell_6t
Xbit_r29_c95 bl_95 br_95 wl_29 vdd gnd cell_6t
Xbit_r30_c95 bl_95 br_95 wl_30 vdd gnd cell_6t
Xbit_r31_c95 bl_95 br_95 wl_31 vdd gnd cell_6t
Xbit_r32_c95 bl_95 br_95 wl_32 vdd gnd cell_6t
Xbit_r33_c95 bl_95 br_95 wl_33 vdd gnd cell_6t
Xbit_r34_c95 bl_95 br_95 wl_34 vdd gnd cell_6t
Xbit_r35_c95 bl_95 br_95 wl_35 vdd gnd cell_6t
Xbit_r36_c95 bl_95 br_95 wl_36 vdd gnd cell_6t
Xbit_r37_c95 bl_95 br_95 wl_37 vdd gnd cell_6t
Xbit_r38_c95 bl_95 br_95 wl_38 vdd gnd cell_6t
Xbit_r39_c95 bl_95 br_95 wl_39 vdd gnd cell_6t
Xbit_r40_c95 bl_95 br_95 wl_40 vdd gnd cell_6t
Xbit_r41_c95 bl_95 br_95 wl_41 vdd gnd cell_6t
Xbit_r42_c95 bl_95 br_95 wl_42 vdd gnd cell_6t
Xbit_r43_c95 bl_95 br_95 wl_43 vdd gnd cell_6t
Xbit_r44_c95 bl_95 br_95 wl_44 vdd gnd cell_6t
Xbit_r45_c95 bl_95 br_95 wl_45 vdd gnd cell_6t
Xbit_r46_c95 bl_95 br_95 wl_46 vdd gnd cell_6t
Xbit_r47_c95 bl_95 br_95 wl_47 vdd gnd cell_6t
Xbit_r48_c95 bl_95 br_95 wl_48 vdd gnd cell_6t
Xbit_r49_c95 bl_95 br_95 wl_49 vdd gnd cell_6t
Xbit_r50_c95 bl_95 br_95 wl_50 vdd gnd cell_6t
Xbit_r51_c95 bl_95 br_95 wl_51 vdd gnd cell_6t
Xbit_r52_c95 bl_95 br_95 wl_52 vdd gnd cell_6t
Xbit_r53_c95 bl_95 br_95 wl_53 vdd gnd cell_6t
Xbit_r54_c95 bl_95 br_95 wl_54 vdd gnd cell_6t
Xbit_r55_c95 bl_95 br_95 wl_55 vdd gnd cell_6t
Xbit_r56_c95 bl_95 br_95 wl_56 vdd gnd cell_6t
Xbit_r57_c95 bl_95 br_95 wl_57 vdd gnd cell_6t
Xbit_r58_c95 bl_95 br_95 wl_58 vdd gnd cell_6t
Xbit_r59_c95 bl_95 br_95 wl_59 vdd gnd cell_6t
Xbit_r60_c95 bl_95 br_95 wl_60 vdd gnd cell_6t
Xbit_r61_c95 bl_95 br_95 wl_61 vdd gnd cell_6t
Xbit_r62_c95 bl_95 br_95 wl_62 vdd gnd cell_6t
Xbit_r63_c95 bl_95 br_95 wl_63 vdd gnd cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd cell_6t
Xbit_r1_c96 bl_96 br_96 wl_1 vdd gnd cell_6t
Xbit_r2_c96 bl_96 br_96 wl_2 vdd gnd cell_6t
Xbit_r3_c96 bl_96 br_96 wl_3 vdd gnd cell_6t
Xbit_r4_c96 bl_96 br_96 wl_4 vdd gnd cell_6t
Xbit_r5_c96 bl_96 br_96 wl_5 vdd gnd cell_6t
Xbit_r6_c96 bl_96 br_96 wl_6 vdd gnd cell_6t
Xbit_r7_c96 bl_96 br_96 wl_7 vdd gnd cell_6t
Xbit_r8_c96 bl_96 br_96 wl_8 vdd gnd cell_6t
Xbit_r9_c96 bl_96 br_96 wl_9 vdd gnd cell_6t
Xbit_r10_c96 bl_96 br_96 wl_10 vdd gnd cell_6t
Xbit_r11_c96 bl_96 br_96 wl_11 vdd gnd cell_6t
Xbit_r12_c96 bl_96 br_96 wl_12 vdd gnd cell_6t
Xbit_r13_c96 bl_96 br_96 wl_13 vdd gnd cell_6t
Xbit_r14_c96 bl_96 br_96 wl_14 vdd gnd cell_6t
Xbit_r15_c96 bl_96 br_96 wl_15 vdd gnd cell_6t
Xbit_r16_c96 bl_96 br_96 wl_16 vdd gnd cell_6t
Xbit_r17_c96 bl_96 br_96 wl_17 vdd gnd cell_6t
Xbit_r18_c96 bl_96 br_96 wl_18 vdd gnd cell_6t
Xbit_r19_c96 bl_96 br_96 wl_19 vdd gnd cell_6t
Xbit_r20_c96 bl_96 br_96 wl_20 vdd gnd cell_6t
Xbit_r21_c96 bl_96 br_96 wl_21 vdd gnd cell_6t
Xbit_r22_c96 bl_96 br_96 wl_22 vdd gnd cell_6t
Xbit_r23_c96 bl_96 br_96 wl_23 vdd gnd cell_6t
Xbit_r24_c96 bl_96 br_96 wl_24 vdd gnd cell_6t
Xbit_r25_c96 bl_96 br_96 wl_25 vdd gnd cell_6t
Xbit_r26_c96 bl_96 br_96 wl_26 vdd gnd cell_6t
Xbit_r27_c96 bl_96 br_96 wl_27 vdd gnd cell_6t
Xbit_r28_c96 bl_96 br_96 wl_28 vdd gnd cell_6t
Xbit_r29_c96 bl_96 br_96 wl_29 vdd gnd cell_6t
Xbit_r30_c96 bl_96 br_96 wl_30 vdd gnd cell_6t
Xbit_r31_c96 bl_96 br_96 wl_31 vdd gnd cell_6t
Xbit_r32_c96 bl_96 br_96 wl_32 vdd gnd cell_6t
Xbit_r33_c96 bl_96 br_96 wl_33 vdd gnd cell_6t
Xbit_r34_c96 bl_96 br_96 wl_34 vdd gnd cell_6t
Xbit_r35_c96 bl_96 br_96 wl_35 vdd gnd cell_6t
Xbit_r36_c96 bl_96 br_96 wl_36 vdd gnd cell_6t
Xbit_r37_c96 bl_96 br_96 wl_37 vdd gnd cell_6t
Xbit_r38_c96 bl_96 br_96 wl_38 vdd gnd cell_6t
Xbit_r39_c96 bl_96 br_96 wl_39 vdd gnd cell_6t
Xbit_r40_c96 bl_96 br_96 wl_40 vdd gnd cell_6t
Xbit_r41_c96 bl_96 br_96 wl_41 vdd gnd cell_6t
Xbit_r42_c96 bl_96 br_96 wl_42 vdd gnd cell_6t
Xbit_r43_c96 bl_96 br_96 wl_43 vdd gnd cell_6t
Xbit_r44_c96 bl_96 br_96 wl_44 vdd gnd cell_6t
Xbit_r45_c96 bl_96 br_96 wl_45 vdd gnd cell_6t
Xbit_r46_c96 bl_96 br_96 wl_46 vdd gnd cell_6t
Xbit_r47_c96 bl_96 br_96 wl_47 vdd gnd cell_6t
Xbit_r48_c96 bl_96 br_96 wl_48 vdd gnd cell_6t
Xbit_r49_c96 bl_96 br_96 wl_49 vdd gnd cell_6t
Xbit_r50_c96 bl_96 br_96 wl_50 vdd gnd cell_6t
Xbit_r51_c96 bl_96 br_96 wl_51 vdd gnd cell_6t
Xbit_r52_c96 bl_96 br_96 wl_52 vdd gnd cell_6t
Xbit_r53_c96 bl_96 br_96 wl_53 vdd gnd cell_6t
Xbit_r54_c96 bl_96 br_96 wl_54 vdd gnd cell_6t
Xbit_r55_c96 bl_96 br_96 wl_55 vdd gnd cell_6t
Xbit_r56_c96 bl_96 br_96 wl_56 vdd gnd cell_6t
Xbit_r57_c96 bl_96 br_96 wl_57 vdd gnd cell_6t
Xbit_r58_c96 bl_96 br_96 wl_58 vdd gnd cell_6t
Xbit_r59_c96 bl_96 br_96 wl_59 vdd gnd cell_6t
Xbit_r60_c96 bl_96 br_96 wl_60 vdd gnd cell_6t
Xbit_r61_c96 bl_96 br_96 wl_61 vdd gnd cell_6t
Xbit_r62_c96 bl_96 br_96 wl_62 vdd gnd cell_6t
Xbit_r63_c96 bl_96 br_96 wl_63 vdd gnd cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd cell_6t
Xbit_r1_c97 bl_97 br_97 wl_1 vdd gnd cell_6t
Xbit_r2_c97 bl_97 br_97 wl_2 vdd gnd cell_6t
Xbit_r3_c97 bl_97 br_97 wl_3 vdd gnd cell_6t
Xbit_r4_c97 bl_97 br_97 wl_4 vdd gnd cell_6t
Xbit_r5_c97 bl_97 br_97 wl_5 vdd gnd cell_6t
Xbit_r6_c97 bl_97 br_97 wl_6 vdd gnd cell_6t
Xbit_r7_c97 bl_97 br_97 wl_7 vdd gnd cell_6t
Xbit_r8_c97 bl_97 br_97 wl_8 vdd gnd cell_6t
Xbit_r9_c97 bl_97 br_97 wl_9 vdd gnd cell_6t
Xbit_r10_c97 bl_97 br_97 wl_10 vdd gnd cell_6t
Xbit_r11_c97 bl_97 br_97 wl_11 vdd gnd cell_6t
Xbit_r12_c97 bl_97 br_97 wl_12 vdd gnd cell_6t
Xbit_r13_c97 bl_97 br_97 wl_13 vdd gnd cell_6t
Xbit_r14_c97 bl_97 br_97 wl_14 vdd gnd cell_6t
Xbit_r15_c97 bl_97 br_97 wl_15 vdd gnd cell_6t
Xbit_r16_c97 bl_97 br_97 wl_16 vdd gnd cell_6t
Xbit_r17_c97 bl_97 br_97 wl_17 vdd gnd cell_6t
Xbit_r18_c97 bl_97 br_97 wl_18 vdd gnd cell_6t
Xbit_r19_c97 bl_97 br_97 wl_19 vdd gnd cell_6t
Xbit_r20_c97 bl_97 br_97 wl_20 vdd gnd cell_6t
Xbit_r21_c97 bl_97 br_97 wl_21 vdd gnd cell_6t
Xbit_r22_c97 bl_97 br_97 wl_22 vdd gnd cell_6t
Xbit_r23_c97 bl_97 br_97 wl_23 vdd gnd cell_6t
Xbit_r24_c97 bl_97 br_97 wl_24 vdd gnd cell_6t
Xbit_r25_c97 bl_97 br_97 wl_25 vdd gnd cell_6t
Xbit_r26_c97 bl_97 br_97 wl_26 vdd gnd cell_6t
Xbit_r27_c97 bl_97 br_97 wl_27 vdd gnd cell_6t
Xbit_r28_c97 bl_97 br_97 wl_28 vdd gnd cell_6t
Xbit_r29_c97 bl_97 br_97 wl_29 vdd gnd cell_6t
Xbit_r30_c97 bl_97 br_97 wl_30 vdd gnd cell_6t
Xbit_r31_c97 bl_97 br_97 wl_31 vdd gnd cell_6t
Xbit_r32_c97 bl_97 br_97 wl_32 vdd gnd cell_6t
Xbit_r33_c97 bl_97 br_97 wl_33 vdd gnd cell_6t
Xbit_r34_c97 bl_97 br_97 wl_34 vdd gnd cell_6t
Xbit_r35_c97 bl_97 br_97 wl_35 vdd gnd cell_6t
Xbit_r36_c97 bl_97 br_97 wl_36 vdd gnd cell_6t
Xbit_r37_c97 bl_97 br_97 wl_37 vdd gnd cell_6t
Xbit_r38_c97 bl_97 br_97 wl_38 vdd gnd cell_6t
Xbit_r39_c97 bl_97 br_97 wl_39 vdd gnd cell_6t
Xbit_r40_c97 bl_97 br_97 wl_40 vdd gnd cell_6t
Xbit_r41_c97 bl_97 br_97 wl_41 vdd gnd cell_6t
Xbit_r42_c97 bl_97 br_97 wl_42 vdd gnd cell_6t
Xbit_r43_c97 bl_97 br_97 wl_43 vdd gnd cell_6t
Xbit_r44_c97 bl_97 br_97 wl_44 vdd gnd cell_6t
Xbit_r45_c97 bl_97 br_97 wl_45 vdd gnd cell_6t
Xbit_r46_c97 bl_97 br_97 wl_46 vdd gnd cell_6t
Xbit_r47_c97 bl_97 br_97 wl_47 vdd gnd cell_6t
Xbit_r48_c97 bl_97 br_97 wl_48 vdd gnd cell_6t
Xbit_r49_c97 bl_97 br_97 wl_49 vdd gnd cell_6t
Xbit_r50_c97 bl_97 br_97 wl_50 vdd gnd cell_6t
Xbit_r51_c97 bl_97 br_97 wl_51 vdd gnd cell_6t
Xbit_r52_c97 bl_97 br_97 wl_52 vdd gnd cell_6t
Xbit_r53_c97 bl_97 br_97 wl_53 vdd gnd cell_6t
Xbit_r54_c97 bl_97 br_97 wl_54 vdd gnd cell_6t
Xbit_r55_c97 bl_97 br_97 wl_55 vdd gnd cell_6t
Xbit_r56_c97 bl_97 br_97 wl_56 vdd gnd cell_6t
Xbit_r57_c97 bl_97 br_97 wl_57 vdd gnd cell_6t
Xbit_r58_c97 bl_97 br_97 wl_58 vdd gnd cell_6t
Xbit_r59_c97 bl_97 br_97 wl_59 vdd gnd cell_6t
Xbit_r60_c97 bl_97 br_97 wl_60 vdd gnd cell_6t
Xbit_r61_c97 bl_97 br_97 wl_61 vdd gnd cell_6t
Xbit_r62_c97 bl_97 br_97 wl_62 vdd gnd cell_6t
Xbit_r63_c97 bl_97 br_97 wl_63 vdd gnd cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd cell_6t
Xbit_r1_c98 bl_98 br_98 wl_1 vdd gnd cell_6t
Xbit_r2_c98 bl_98 br_98 wl_2 vdd gnd cell_6t
Xbit_r3_c98 bl_98 br_98 wl_3 vdd gnd cell_6t
Xbit_r4_c98 bl_98 br_98 wl_4 vdd gnd cell_6t
Xbit_r5_c98 bl_98 br_98 wl_5 vdd gnd cell_6t
Xbit_r6_c98 bl_98 br_98 wl_6 vdd gnd cell_6t
Xbit_r7_c98 bl_98 br_98 wl_7 vdd gnd cell_6t
Xbit_r8_c98 bl_98 br_98 wl_8 vdd gnd cell_6t
Xbit_r9_c98 bl_98 br_98 wl_9 vdd gnd cell_6t
Xbit_r10_c98 bl_98 br_98 wl_10 vdd gnd cell_6t
Xbit_r11_c98 bl_98 br_98 wl_11 vdd gnd cell_6t
Xbit_r12_c98 bl_98 br_98 wl_12 vdd gnd cell_6t
Xbit_r13_c98 bl_98 br_98 wl_13 vdd gnd cell_6t
Xbit_r14_c98 bl_98 br_98 wl_14 vdd gnd cell_6t
Xbit_r15_c98 bl_98 br_98 wl_15 vdd gnd cell_6t
Xbit_r16_c98 bl_98 br_98 wl_16 vdd gnd cell_6t
Xbit_r17_c98 bl_98 br_98 wl_17 vdd gnd cell_6t
Xbit_r18_c98 bl_98 br_98 wl_18 vdd gnd cell_6t
Xbit_r19_c98 bl_98 br_98 wl_19 vdd gnd cell_6t
Xbit_r20_c98 bl_98 br_98 wl_20 vdd gnd cell_6t
Xbit_r21_c98 bl_98 br_98 wl_21 vdd gnd cell_6t
Xbit_r22_c98 bl_98 br_98 wl_22 vdd gnd cell_6t
Xbit_r23_c98 bl_98 br_98 wl_23 vdd gnd cell_6t
Xbit_r24_c98 bl_98 br_98 wl_24 vdd gnd cell_6t
Xbit_r25_c98 bl_98 br_98 wl_25 vdd gnd cell_6t
Xbit_r26_c98 bl_98 br_98 wl_26 vdd gnd cell_6t
Xbit_r27_c98 bl_98 br_98 wl_27 vdd gnd cell_6t
Xbit_r28_c98 bl_98 br_98 wl_28 vdd gnd cell_6t
Xbit_r29_c98 bl_98 br_98 wl_29 vdd gnd cell_6t
Xbit_r30_c98 bl_98 br_98 wl_30 vdd gnd cell_6t
Xbit_r31_c98 bl_98 br_98 wl_31 vdd gnd cell_6t
Xbit_r32_c98 bl_98 br_98 wl_32 vdd gnd cell_6t
Xbit_r33_c98 bl_98 br_98 wl_33 vdd gnd cell_6t
Xbit_r34_c98 bl_98 br_98 wl_34 vdd gnd cell_6t
Xbit_r35_c98 bl_98 br_98 wl_35 vdd gnd cell_6t
Xbit_r36_c98 bl_98 br_98 wl_36 vdd gnd cell_6t
Xbit_r37_c98 bl_98 br_98 wl_37 vdd gnd cell_6t
Xbit_r38_c98 bl_98 br_98 wl_38 vdd gnd cell_6t
Xbit_r39_c98 bl_98 br_98 wl_39 vdd gnd cell_6t
Xbit_r40_c98 bl_98 br_98 wl_40 vdd gnd cell_6t
Xbit_r41_c98 bl_98 br_98 wl_41 vdd gnd cell_6t
Xbit_r42_c98 bl_98 br_98 wl_42 vdd gnd cell_6t
Xbit_r43_c98 bl_98 br_98 wl_43 vdd gnd cell_6t
Xbit_r44_c98 bl_98 br_98 wl_44 vdd gnd cell_6t
Xbit_r45_c98 bl_98 br_98 wl_45 vdd gnd cell_6t
Xbit_r46_c98 bl_98 br_98 wl_46 vdd gnd cell_6t
Xbit_r47_c98 bl_98 br_98 wl_47 vdd gnd cell_6t
Xbit_r48_c98 bl_98 br_98 wl_48 vdd gnd cell_6t
Xbit_r49_c98 bl_98 br_98 wl_49 vdd gnd cell_6t
Xbit_r50_c98 bl_98 br_98 wl_50 vdd gnd cell_6t
Xbit_r51_c98 bl_98 br_98 wl_51 vdd gnd cell_6t
Xbit_r52_c98 bl_98 br_98 wl_52 vdd gnd cell_6t
Xbit_r53_c98 bl_98 br_98 wl_53 vdd gnd cell_6t
Xbit_r54_c98 bl_98 br_98 wl_54 vdd gnd cell_6t
Xbit_r55_c98 bl_98 br_98 wl_55 vdd gnd cell_6t
Xbit_r56_c98 bl_98 br_98 wl_56 vdd gnd cell_6t
Xbit_r57_c98 bl_98 br_98 wl_57 vdd gnd cell_6t
Xbit_r58_c98 bl_98 br_98 wl_58 vdd gnd cell_6t
Xbit_r59_c98 bl_98 br_98 wl_59 vdd gnd cell_6t
Xbit_r60_c98 bl_98 br_98 wl_60 vdd gnd cell_6t
Xbit_r61_c98 bl_98 br_98 wl_61 vdd gnd cell_6t
Xbit_r62_c98 bl_98 br_98 wl_62 vdd gnd cell_6t
Xbit_r63_c98 bl_98 br_98 wl_63 vdd gnd cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd cell_6t
Xbit_r1_c99 bl_99 br_99 wl_1 vdd gnd cell_6t
Xbit_r2_c99 bl_99 br_99 wl_2 vdd gnd cell_6t
Xbit_r3_c99 bl_99 br_99 wl_3 vdd gnd cell_6t
Xbit_r4_c99 bl_99 br_99 wl_4 vdd gnd cell_6t
Xbit_r5_c99 bl_99 br_99 wl_5 vdd gnd cell_6t
Xbit_r6_c99 bl_99 br_99 wl_6 vdd gnd cell_6t
Xbit_r7_c99 bl_99 br_99 wl_7 vdd gnd cell_6t
Xbit_r8_c99 bl_99 br_99 wl_8 vdd gnd cell_6t
Xbit_r9_c99 bl_99 br_99 wl_9 vdd gnd cell_6t
Xbit_r10_c99 bl_99 br_99 wl_10 vdd gnd cell_6t
Xbit_r11_c99 bl_99 br_99 wl_11 vdd gnd cell_6t
Xbit_r12_c99 bl_99 br_99 wl_12 vdd gnd cell_6t
Xbit_r13_c99 bl_99 br_99 wl_13 vdd gnd cell_6t
Xbit_r14_c99 bl_99 br_99 wl_14 vdd gnd cell_6t
Xbit_r15_c99 bl_99 br_99 wl_15 vdd gnd cell_6t
Xbit_r16_c99 bl_99 br_99 wl_16 vdd gnd cell_6t
Xbit_r17_c99 bl_99 br_99 wl_17 vdd gnd cell_6t
Xbit_r18_c99 bl_99 br_99 wl_18 vdd gnd cell_6t
Xbit_r19_c99 bl_99 br_99 wl_19 vdd gnd cell_6t
Xbit_r20_c99 bl_99 br_99 wl_20 vdd gnd cell_6t
Xbit_r21_c99 bl_99 br_99 wl_21 vdd gnd cell_6t
Xbit_r22_c99 bl_99 br_99 wl_22 vdd gnd cell_6t
Xbit_r23_c99 bl_99 br_99 wl_23 vdd gnd cell_6t
Xbit_r24_c99 bl_99 br_99 wl_24 vdd gnd cell_6t
Xbit_r25_c99 bl_99 br_99 wl_25 vdd gnd cell_6t
Xbit_r26_c99 bl_99 br_99 wl_26 vdd gnd cell_6t
Xbit_r27_c99 bl_99 br_99 wl_27 vdd gnd cell_6t
Xbit_r28_c99 bl_99 br_99 wl_28 vdd gnd cell_6t
Xbit_r29_c99 bl_99 br_99 wl_29 vdd gnd cell_6t
Xbit_r30_c99 bl_99 br_99 wl_30 vdd gnd cell_6t
Xbit_r31_c99 bl_99 br_99 wl_31 vdd gnd cell_6t
Xbit_r32_c99 bl_99 br_99 wl_32 vdd gnd cell_6t
Xbit_r33_c99 bl_99 br_99 wl_33 vdd gnd cell_6t
Xbit_r34_c99 bl_99 br_99 wl_34 vdd gnd cell_6t
Xbit_r35_c99 bl_99 br_99 wl_35 vdd gnd cell_6t
Xbit_r36_c99 bl_99 br_99 wl_36 vdd gnd cell_6t
Xbit_r37_c99 bl_99 br_99 wl_37 vdd gnd cell_6t
Xbit_r38_c99 bl_99 br_99 wl_38 vdd gnd cell_6t
Xbit_r39_c99 bl_99 br_99 wl_39 vdd gnd cell_6t
Xbit_r40_c99 bl_99 br_99 wl_40 vdd gnd cell_6t
Xbit_r41_c99 bl_99 br_99 wl_41 vdd gnd cell_6t
Xbit_r42_c99 bl_99 br_99 wl_42 vdd gnd cell_6t
Xbit_r43_c99 bl_99 br_99 wl_43 vdd gnd cell_6t
Xbit_r44_c99 bl_99 br_99 wl_44 vdd gnd cell_6t
Xbit_r45_c99 bl_99 br_99 wl_45 vdd gnd cell_6t
Xbit_r46_c99 bl_99 br_99 wl_46 vdd gnd cell_6t
Xbit_r47_c99 bl_99 br_99 wl_47 vdd gnd cell_6t
Xbit_r48_c99 bl_99 br_99 wl_48 vdd gnd cell_6t
Xbit_r49_c99 bl_99 br_99 wl_49 vdd gnd cell_6t
Xbit_r50_c99 bl_99 br_99 wl_50 vdd gnd cell_6t
Xbit_r51_c99 bl_99 br_99 wl_51 vdd gnd cell_6t
Xbit_r52_c99 bl_99 br_99 wl_52 vdd gnd cell_6t
Xbit_r53_c99 bl_99 br_99 wl_53 vdd gnd cell_6t
Xbit_r54_c99 bl_99 br_99 wl_54 vdd gnd cell_6t
Xbit_r55_c99 bl_99 br_99 wl_55 vdd gnd cell_6t
Xbit_r56_c99 bl_99 br_99 wl_56 vdd gnd cell_6t
Xbit_r57_c99 bl_99 br_99 wl_57 vdd gnd cell_6t
Xbit_r58_c99 bl_99 br_99 wl_58 vdd gnd cell_6t
Xbit_r59_c99 bl_99 br_99 wl_59 vdd gnd cell_6t
Xbit_r60_c99 bl_99 br_99 wl_60 vdd gnd cell_6t
Xbit_r61_c99 bl_99 br_99 wl_61 vdd gnd cell_6t
Xbit_r62_c99 bl_99 br_99 wl_62 vdd gnd cell_6t
Xbit_r63_c99 bl_99 br_99 wl_63 vdd gnd cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd cell_6t
Xbit_r1_c100 bl_100 br_100 wl_1 vdd gnd cell_6t
Xbit_r2_c100 bl_100 br_100 wl_2 vdd gnd cell_6t
Xbit_r3_c100 bl_100 br_100 wl_3 vdd gnd cell_6t
Xbit_r4_c100 bl_100 br_100 wl_4 vdd gnd cell_6t
Xbit_r5_c100 bl_100 br_100 wl_5 vdd gnd cell_6t
Xbit_r6_c100 bl_100 br_100 wl_6 vdd gnd cell_6t
Xbit_r7_c100 bl_100 br_100 wl_7 vdd gnd cell_6t
Xbit_r8_c100 bl_100 br_100 wl_8 vdd gnd cell_6t
Xbit_r9_c100 bl_100 br_100 wl_9 vdd gnd cell_6t
Xbit_r10_c100 bl_100 br_100 wl_10 vdd gnd cell_6t
Xbit_r11_c100 bl_100 br_100 wl_11 vdd gnd cell_6t
Xbit_r12_c100 bl_100 br_100 wl_12 vdd gnd cell_6t
Xbit_r13_c100 bl_100 br_100 wl_13 vdd gnd cell_6t
Xbit_r14_c100 bl_100 br_100 wl_14 vdd gnd cell_6t
Xbit_r15_c100 bl_100 br_100 wl_15 vdd gnd cell_6t
Xbit_r16_c100 bl_100 br_100 wl_16 vdd gnd cell_6t
Xbit_r17_c100 bl_100 br_100 wl_17 vdd gnd cell_6t
Xbit_r18_c100 bl_100 br_100 wl_18 vdd gnd cell_6t
Xbit_r19_c100 bl_100 br_100 wl_19 vdd gnd cell_6t
Xbit_r20_c100 bl_100 br_100 wl_20 vdd gnd cell_6t
Xbit_r21_c100 bl_100 br_100 wl_21 vdd gnd cell_6t
Xbit_r22_c100 bl_100 br_100 wl_22 vdd gnd cell_6t
Xbit_r23_c100 bl_100 br_100 wl_23 vdd gnd cell_6t
Xbit_r24_c100 bl_100 br_100 wl_24 vdd gnd cell_6t
Xbit_r25_c100 bl_100 br_100 wl_25 vdd gnd cell_6t
Xbit_r26_c100 bl_100 br_100 wl_26 vdd gnd cell_6t
Xbit_r27_c100 bl_100 br_100 wl_27 vdd gnd cell_6t
Xbit_r28_c100 bl_100 br_100 wl_28 vdd gnd cell_6t
Xbit_r29_c100 bl_100 br_100 wl_29 vdd gnd cell_6t
Xbit_r30_c100 bl_100 br_100 wl_30 vdd gnd cell_6t
Xbit_r31_c100 bl_100 br_100 wl_31 vdd gnd cell_6t
Xbit_r32_c100 bl_100 br_100 wl_32 vdd gnd cell_6t
Xbit_r33_c100 bl_100 br_100 wl_33 vdd gnd cell_6t
Xbit_r34_c100 bl_100 br_100 wl_34 vdd gnd cell_6t
Xbit_r35_c100 bl_100 br_100 wl_35 vdd gnd cell_6t
Xbit_r36_c100 bl_100 br_100 wl_36 vdd gnd cell_6t
Xbit_r37_c100 bl_100 br_100 wl_37 vdd gnd cell_6t
Xbit_r38_c100 bl_100 br_100 wl_38 vdd gnd cell_6t
Xbit_r39_c100 bl_100 br_100 wl_39 vdd gnd cell_6t
Xbit_r40_c100 bl_100 br_100 wl_40 vdd gnd cell_6t
Xbit_r41_c100 bl_100 br_100 wl_41 vdd gnd cell_6t
Xbit_r42_c100 bl_100 br_100 wl_42 vdd gnd cell_6t
Xbit_r43_c100 bl_100 br_100 wl_43 vdd gnd cell_6t
Xbit_r44_c100 bl_100 br_100 wl_44 vdd gnd cell_6t
Xbit_r45_c100 bl_100 br_100 wl_45 vdd gnd cell_6t
Xbit_r46_c100 bl_100 br_100 wl_46 vdd gnd cell_6t
Xbit_r47_c100 bl_100 br_100 wl_47 vdd gnd cell_6t
Xbit_r48_c100 bl_100 br_100 wl_48 vdd gnd cell_6t
Xbit_r49_c100 bl_100 br_100 wl_49 vdd gnd cell_6t
Xbit_r50_c100 bl_100 br_100 wl_50 vdd gnd cell_6t
Xbit_r51_c100 bl_100 br_100 wl_51 vdd gnd cell_6t
Xbit_r52_c100 bl_100 br_100 wl_52 vdd gnd cell_6t
Xbit_r53_c100 bl_100 br_100 wl_53 vdd gnd cell_6t
Xbit_r54_c100 bl_100 br_100 wl_54 vdd gnd cell_6t
Xbit_r55_c100 bl_100 br_100 wl_55 vdd gnd cell_6t
Xbit_r56_c100 bl_100 br_100 wl_56 vdd gnd cell_6t
Xbit_r57_c100 bl_100 br_100 wl_57 vdd gnd cell_6t
Xbit_r58_c100 bl_100 br_100 wl_58 vdd gnd cell_6t
Xbit_r59_c100 bl_100 br_100 wl_59 vdd gnd cell_6t
Xbit_r60_c100 bl_100 br_100 wl_60 vdd gnd cell_6t
Xbit_r61_c100 bl_100 br_100 wl_61 vdd gnd cell_6t
Xbit_r62_c100 bl_100 br_100 wl_62 vdd gnd cell_6t
Xbit_r63_c100 bl_100 br_100 wl_63 vdd gnd cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd cell_6t
Xbit_r1_c101 bl_101 br_101 wl_1 vdd gnd cell_6t
Xbit_r2_c101 bl_101 br_101 wl_2 vdd gnd cell_6t
Xbit_r3_c101 bl_101 br_101 wl_3 vdd gnd cell_6t
Xbit_r4_c101 bl_101 br_101 wl_4 vdd gnd cell_6t
Xbit_r5_c101 bl_101 br_101 wl_5 vdd gnd cell_6t
Xbit_r6_c101 bl_101 br_101 wl_6 vdd gnd cell_6t
Xbit_r7_c101 bl_101 br_101 wl_7 vdd gnd cell_6t
Xbit_r8_c101 bl_101 br_101 wl_8 vdd gnd cell_6t
Xbit_r9_c101 bl_101 br_101 wl_9 vdd gnd cell_6t
Xbit_r10_c101 bl_101 br_101 wl_10 vdd gnd cell_6t
Xbit_r11_c101 bl_101 br_101 wl_11 vdd gnd cell_6t
Xbit_r12_c101 bl_101 br_101 wl_12 vdd gnd cell_6t
Xbit_r13_c101 bl_101 br_101 wl_13 vdd gnd cell_6t
Xbit_r14_c101 bl_101 br_101 wl_14 vdd gnd cell_6t
Xbit_r15_c101 bl_101 br_101 wl_15 vdd gnd cell_6t
Xbit_r16_c101 bl_101 br_101 wl_16 vdd gnd cell_6t
Xbit_r17_c101 bl_101 br_101 wl_17 vdd gnd cell_6t
Xbit_r18_c101 bl_101 br_101 wl_18 vdd gnd cell_6t
Xbit_r19_c101 bl_101 br_101 wl_19 vdd gnd cell_6t
Xbit_r20_c101 bl_101 br_101 wl_20 vdd gnd cell_6t
Xbit_r21_c101 bl_101 br_101 wl_21 vdd gnd cell_6t
Xbit_r22_c101 bl_101 br_101 wl_22 vdd gnd cell_6t
Xbit_r23_c101 bl_101 br_101 wl_23 vdd gnd cell_6t
Xbit_r24_c101 bl_101 br_101 wl_24 vdd gnd cell_6t
Xbit_r25_c101 bl_101 br_101 wl_25 vdd gnd cell_6t
Xbit_r26_c101 bl_101 br_101 wl_26 vdd gnd cell_6t
Xbit_r27_c101 bl_101 br_101 wl_27 vdd gnd cell_6t
Xbit_r28_c101 bl_101 br_101 wl_28 vdd gnd cell_6t
Xbit_r29_c101 bl_101 br_101 wl_29 vdd gnd cell_6t
Xbit_r30_c101 bl_101 br_101 wl_30 vdd gnd cell_6t
Xbit_r31_c101 bl_101 br_101 wl_31 vdd gnd cell_6t
Xbit_r32_c101 bl_101 br_101 wl_32 vdd gnd cell_6t
Xbit_r33_c101 bl_101 br_101 wl_33 vdd gnd cell_6t
Xbit_r34_c101 bl_101 br_101 wl_34 vdd gnd cell_6t
Xbit_r35_c101 bl_101 br_101 wl_35 vdd gnd cell_6t
Xbit_r36_c101 bl_101 br_101 wl_36 vdd gnd cell_6t
Xbit_r37_c101 bl_101 br_101 wl_37 vdd gnd cell_6t
Xbit_r38_c101 bl_101 br_101 wl_38 vdd gnd cell_6t
Xbit_r39_c101 bl_101 br_101 wl_39 vdd gnd cell_6t
Xbit_r40_c101 bl_101 br_101 wl_40 vdd gnd cell_6t
Xbit_r41_c101 bl_101 br_101 wl_41 vdd gnd cell_6t
Xbit_r42_c101 bl_101 br_101 wl_42 vdd gnd cell_6t
Xbit_r43_c101 bl_101 br_101 wl_43 vdd gnd cell_6t
Xbit_r44_c101 bl_101 br_101 wl_44 vdd gnd cell_6t
Xbit_r45_c101 bl_101 br_101 wl_45 vdd gnd cell_6t
Xbit_r46_c101 bl_101 br_101 wl_46 vdd gnd cell_6t
Xbit_r47_c101 bl_101 br_101 wl_47 vdd gnd cell_6t
Xbit_r48_c101 bl_101 br_101 wl_48 vdd gnd cell_6t
Xbit_r49_c101 bl_101 br_101 wl_49 vdd gnd cell_6t
Xbit_r50_c101 bl_101 br_101 wl_50 vdd gnd cell_6t
Xbit_r51_c101 bl_101 br_101 wl_51 vdd gnd cell_6t
Xbit_r52_c101 bl_101 br_101 wl_52 vdd gnd cell_6t
Xbit_r53_c101 bl_101 br_101 wl_53 vdd gnd cell_6t
Xbit_r54_c101 bl_101 br_101 wl_54 vdd gnd cell_6t
Xbit_r55_c101 bl_101 br_101 wl_55 vdd gnd cell_6t
Xbit_r56_c101 bl_101 br_101 wl_56 vdd gnd cell_6t
Xbit_r57_c101 bl_101 br_101 wl_57 vdd gnd cell_6t
Xbit_r58_c101 bl_101 br_101 wl_58 vdd gnd cell_6t
Xbit_r59_c101 bl_101 br_101 wl_59 vdd gnd cell_6t
Xbit_r60_c101 bl_101 br_101 wl_60 vdd gnd cell_6t
Xbit_r61_c101 bl_101 br_101 wl_61 vdd gnd cell_6t
Xbit_r62_c101 bl_101 br_101 wl_62 vdd gnd cell_6t
Xbit_r63_c101 bl_101 br_101 wl_63 vdd gnd cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd cell_6t
Xbit_r1_c102 bl_102 br_102 wl_1 vdd gnd cell_6t
Xbit_r2_c102 bl_102 br_102 wl_2 vdd gnd cell_6t
Xbit_r3_c102 bl_102 br_102 wl_3 vdd gnd cell_6t
Xbit_r4_c102 bl_102 br_102 wl_4 vdd gnd cell_6t
Xbit_r5_c102 bl_102 br_102 wl_5 vdd gnd cell_6t
Xbit_r6_c102 bl_102 br_102 wl_6 vdd gnd cell_6t
Xbit_r7_c102 bl_102 br_102 wl_7 vdd gnd cell_6t
Xbit_r8_c102 bl_102 br_102 wl_8 vdd gnd cell_6t
Xbit_r9_c102 bl_102 br_102 wl_9 vdd gnd cell_6t
Xbit_r10_c102 bl_102 br_102 wl_10 vdd gnd cell_6t
Xbit_r11_c102 bl_102 br_102 wl_11 vdd gnd cell_6t
Xbit_r12_c102 bl_102 br_102 wl_12 vdd gnd cell_6t
Xbit_r13_c102 bl_102 br_102 wl_13 vdd gnd cell_6t
Xbit_r14_c102 bl_102 br_102 wl_14 vdd gnd cell_6t
Xbit_r15_c102 bl_102 br_102 wl_15 vdd gnd cell_6t
Xbit_r16_c102 bl_102 br_102 wl_16 vdd gnd cell_6t
Xbit_r17_c102 bl_102 br_102 wl_17 vdd gnd cell_6t
Xbit_r18_c102 bl_102 br_102 wl_18 vdd gnd cell_6t
Xbit_r19_c102 bl_102 br_102 wl_19 vdd gnd cell_6t
Xbit_r20_c102 bl_102 br_102 wl_20 vdd gnd cell_6t
Xbit_r21_c102 bl_102 br_102 wl_21 vdd gnd cell_6t
Xbit_r22_c102 bl_102 br_102 wl_22 vdd gnd cell_6t
Xbit_r23_c102 bl_102 br_102 wl_23 vdd gnd cell_6t
Xbit_r24_c102 bl_102 br_102 wl_24 vdd gnd cell_6t
Xbit_r25_c102 bl_102 br_102 wl_25 vdd gnd cell_6t
Xbit_r26_c102 bl_102 br_102 wl_26 vdd gnd cell_6t
Xbit_r27_c102 bl_102 br_102 wl_27 vdd gnd cell_6t
Xbit_r28_c102 bl_102 br_102 wl_28 vdd gnd cell_6t
Xbit_r29_c102 bl_102 br_102 wl_29 vdd gnd cell_6t
Xbit_r30_c102 bl_102 br_102 wl_30 vdd gnd cell_6t
Xbit_r31_c102 bl_102 br_102 wl_31 vdd gnd cell_6t
Xbit_r32_c102 bl_102 br_102 wl_32 vdd gnd cell_6t
Xbit_r33_c102 bl_102 br_102 wl_33 vdd gnd cell_6t
Xbit_r34_c102 bl_102 br_102 wl_34 vdd gnd cell_6t
Xbit_r35_c102 bl_102 br_102 wl_35 vdd gnd cell_6t
Xbit_r36_c102 bl_102 br_102 wl_36 vdd gnd cell_6t
Xbit_r37_c102 bl_102 br_102 wl_37 vdd gnd cell_6t
Xbit_r38_c102 bl_102 br_102 wl_38 vdd gnd cell_6t
Xbit_r39_c102 bl_102 br_102 wl_39 vdd gnd cell_6t
Xbit_r40_c102 bl_102 br_102 wl_40 vdd gnd cell_6t
Xbit_r41_c102 bl_102 br_102 wl_41 vdd gnd cell_6t
Xbit_r42_c102 bl_102 br_102 wl_42 vdd gnd cell_6t
Xbit_r43_c102 bl_102 br_102 wl_43 vdd gnd cell_6t
Xbit_r44_c102 bl_102 br_102 wl_44 vdd gnd cell_6t
Xbit_r45_c102 bl_102 br_102 wl_45 vdd gnd cell_6t
Xbit_r46_c102 bl_102 br_102 wl_46 vdd gnd cell_6t
Xbit_r47_c102 bl_102 br_102 wl_47 vdd gnd cell_6t
Xbit_r48_c102 bl_102 br_102 wl_48 vdd gnd cell_6t
Xbit_r49_c102 bl_102 br_102 wl_49 vdd gnd cell_6t
Xbit_r50_c102 bl_102 br_102 wl_50 vdd gnd cell_6t
Xbit_r51_c102 bl_102 br_102 wl_51 vdd gnd cell_6t
Xbit_r52_c102 bl_102 br_102 wl_52 vdd gnd cell_6t
Xbit_r53_c102 bl_102 br_102 wl_53 vdd gnd cell_6t
Xbit_r54_c102 bl_102 br_102 wl_54 vdd gnd cell_6t
Xbit_r55_c102 bl_102 br_102 wl_55 vdd gnd cell_6t
Xbit_r56_c102 bl_102 br_102 wl_56 vdd gnd cell_6t
Xbit_r57_c102 bl_102 br_102 wl_57 vdd gnd cell_6t
Xbit_r58_c102 bl_102 br_102 wl_58 vdd gnd cell_6t
Xbit_r59_c102 bl_102 br_102 wl_59 vdd gnd cell_6t
Xbit_r60_c102 bl_102 br_102 wl_60 vdd gnd cell_6t
Xbit_r61_c102 bl_102 br_102 wl_61 vdd gnd cell_6t
Xbit_r62_c102 bl_102 br_102 wl_62 vdd gnd cell_6t
Xbit_r63_c102 bl_102 br_102 wl_63 vdd gnd cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd cell_6t
Xbit_r1_c103 bl_103 br_103 wl_1 vdd gnd cell_6t
Xbit_r2_c103 bl_103 br_103 wl_2 vdd gnd cell_6t
Xbit_r3_c103 bl_103 br_103 wl_3 vdd gnd cell_6t
Xbit_r4_c103 bl_103 br_103 wl_4 vdd gnd cell_6t
Xbit_r5_c103 bl_103 br_103 wl_5 vdd gnd cell_6t
Xbit_r6_c103 bl_103 br_103 wl_6 vdd gnd cell_6t
Xbit_r7_c103 bl_103 br_103 wl_7 vdd gnd cell_6t
Xbit_r8_c103 bl_103 br_103 wl_8 vdd gnd cell_6t
Xbit_r9_c103 bl_103 br_103 wl_9 vdd gnd cell_6t
Xbit_r10_c103 bl_103 br_103 wl_10 vdd gnd cell_6t
Xbit_r11_c103 bl_103 br_103 wl_11 vdd gnd cell_6t
Xbit_r12_c103 bl_103 br_103 wl_12 vdd gnd cell_6t
Xbit_r13_c103 bl_103 br_103 wl_13 vdd gnd cell_6t
Xbit_r14_c103 bl_103 br_103 wl_14 vdd gnd cell_6t
Xbit_r15_c103 bl_103 br_103 wl_15 vdd gnd cell_6t
Xbit_r16_c103 bl_103 br_103 wl_16 vdd gnd cell_6t
Xbit_r17_c103 bl_103 br_103 wl_17 vdd gnd cell_6t
Xbit_r18_c103 bl_103 br_103 wl_18 vdd gnd cell_6t
Xbit_r19_c103 bl_103 br_103 wl_19 vdd gnd cell_6t
Xbit_r20_c103 bl_103 br_103 wl_20 vdd gnd cell_6t
Xbit_r21_c103 bl_103 br_103 wl_21 vdd gnd cell_6t
Xbit_r22_c103 bl_103 br_103 wl_22 vdd gnd cell_6t
Xbit_r23_c103 bl_103 br_103 wl_23 vdd gnd cell_6t
Xbit_r24_c103 bl_103 br_103 wl_24 vdd gnd cell_6t
Xbit_r25_c103 bl_103 br_103 wl_25 vdd gnd cell_6t
Xbit_r26_c103 bl_103 br_103 wl_26 vdd gnd cell_6t
Xbit_r27_c103 bl_103 br_103 wl_27 vdd gnd cell_6t
Xbit_r28_c103 bl_103 br_103 wl_28 vdd gnd cell_6t
Xbit_r29_c103 bl_103 br_103 wl_29 vdd gnd cell_6t
Xbit_r30_c103 bl_103 br_103 wl_30 vdd gnd cell_6t
Xbit_r31_c103 bl_103 br_103 wl_31 vdd gnd cell_6t
Xbit_r32_c103 bl_103 br_103 wl_32 vdd gnd cell_6t
Xbit_r33_c103 bl_103 br_103 wl_33 vdd gnd cell_6t
Xbit_r34_c103 bl_103 br_103 wl_34 vdd gnd cell_6t
Xbit_r35_c103 bl_103 br_103 wl_35 vdd gnd cell_6t
Xbit_r36_c103 bl_103 br_103 wl_36 vdd gnd cell_6t
Xbit_r37_c103 bl_103 br_103 wl_37 vdd gnd cell_6t
Xbit_r38_c103 bl_103 br_103 wl_38 vdd gnd cell_6t
Xbit_r39_c103 bl_103 br_103 wl_39 vdd gnd cell_6t
Xbit_r40_c103 bl_103 br_103 wl_40 vdd gnd cell_6t
Xbit_r41_c103 bl_103 br_103 wl_41 vdd gnd cell_6t
Xbit_r42_c103 bl_103 br_103 wl_42 vdd gnd cell_6t
Xbit_r43_c103 bl_103 br_103 wl_43 vdd gnd cell_6t
Xbit_r44_c103 bl_103 br_103 wl_44 vdd gnd cell_6t
Xbit_r45_c103 bl_103 br_103 wl_45 vdd gnd cell_6t
Xbit_r46_c103 bl_103 br_103 wl_46 vdd gnd cell_6t
Xbit_r47_c103 bl_103 br_103 wl_47 vdd gnd cell_6t
Xbit_r48_c103 bl_103 br_103 wl_48 vdd gnd cell_6t
Xbit_r49_c103 bl_103 br_103 wl_49 vdd gnd cell_6t
Xbit_r50_c103 bl_103 br_103 wl_50 vdd gnd cell_6t
Xbit_r51_c103 bl_103 br_103 wl_51 vdd gnd cell_6t
Xbit_r52_c103 bl_103 br_103 wl_52 vdd gnd cell_6t
Xbit_r53_c103 bl_103 br_103 wl_53 vdd gnd cell_6t
Xbit_r54_c103 bl_103 br_103 wl_54 vdd gnd cell_6t
Xbit_r55_c103 bl_103 br_103 wl_55 vdd gnd cell_6t
Xbit_r56_c103 bl_103 br_103 wl_56 vdd gnd cell_6t
Xbit_r57_c103 bl_103 br_103 wl_57 vdd gnd cell_6t
Xbit_r58_c103 bl_103 br_103 wl_58 vdd gnd cell_6t
Xbit_r59_c103 bl_103 br_103 wl_59 vdd gnd cell_6t
Xbit_r60_c103 bl_103 br_103 wl_60 vdd gnd cell_6t
Xbit_r61_c103 bl_103 br_103 wl_61 vdd gnd cell_6t
Xbit_r62_c103 bl_103 br_103 wl_62 vdd gnd cell_6t
Xbit_r63_c103 bl_103 br_103 wl_63 vdd gnd cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd cell_6t
Xbit_r1_c104 bl_104 br_104 wl_1 vdd gnd cell_6t
Xbit_r2_c104 bl_104 br_104 wl_2 vdd gnd cell_6t
Xbit_r3_c104 bl_104 br_104 wl_3 vdd gnd cell_6t
Xbit_r4_c104 bl_104 br_104 wl_4 vdd gnd cell_6t
Xbit_r5_c104 bl_104 br_104 wl_5 vdd gnd cell_6t
Xbit_r6_c104 bl_104 br_104 wl_6 vdd gnd cell_6t
Xbit_r7_c104 bl_104 br_104 wl_7 vdd gnd cell_6t
Xbit_r8_c104 bl_104 br_104 wl_8 vdd gnd cell_6t
Xbit_r9_c104 bl_104 br_104 wl_9 vdd gnd cell_6t
Xbit_r10_c104 bl_104 br_104 wl_10 vdd gnd cell_6t
Xbit_r11_c104 bl_104 br_104 wl_11 vdd gnd cell_6t
Xbit_r12_c104 bl_104 br_104 wl_12 vdd gnd cell_6t
Xbit_r13_c104 bl_104 br_104 wl_13 vdd gnd cell_6t
Xbit_r14_c104 bl_104 br_104 wl_14 vdd gnd cell_6t
Xbit_r15_c104 bl_104 br_104 wl_15 vdd gnd cell_6t
Xbit_r16_c104 bl_104 br_104 wl_16 vdd gnd cell_6t
Xbit_r17_c104 bl_104 br_104 wl_17 vdd gnd cell_6t
Xbit_r18_c104 bl_104 br_104 wl_18 vdd gnd cell_6t
Xbit_r19_c104 bl_104 br_104 wl_19 vdd gnd cell_6t
Xbit_r20_c104 bl_104 br_104 wl_20 vdd gnd cell_6t
Xbit_r21_c104 bl_104 br_104 wl_21 vdd gnd cell_6t
Xbit_r22_c104 bl_104 br_104 wl_22 vdd gnd cell_6t
Xbit_r23_c104 bl_104 br_104 wl_23 vdd gnd cell_6t
Xbit_r24_c104 bl_104 br_104 wl_24 vdd gnd cell_6t
Xbit_r25_c104 bl_104 br_104 wl_25 vdd gnd cell_6t
Xbit_r26_c104 bl_104 br_104 wl_26 vdd gnd cell_6t
Xbit_r27_c104 bl_104 br_104 wl_27 vdd gnd cell_6t
Xbit_r28_c104 bl_104 br_104 wl_28 vdd gnd cell_6t
Xbit_r29_c104 bl_104 br_104 wl_29 vdd gnd cell_6t
Xbit_r30_c104 bl_104 br_104 wl_30 vdd gnd cell_6t
Xbit_r31_c104 bl_104 br_104 wl_31 vdd gnd cell_6t
Xbit_r32_c104 bl_104 br_104 wl_32 vdd gnd cell_6t
Xbit_r33_c104 bl_104 br_104 wl_33 vdd gnd cell_6t
Xbit_r34_c104 bl_104 br_104 wl_34 vdd gnd cell_6t
Xbit_r35_c104 bl_104 br_104 wl_35 vdd gnd cell_6t
Xbit_r36_c104 bl_104 br_104 wl_36 vdd gnd cell_6t
Xbit_r37_c104 bl_104 br_104 wl_37 vdd gnd cell_6t
Xbit_r38_c104 bl_104 br_104 wl_38 vdd gnd cell_6t
Xbit_r39_c104 bl_104 br_104 wl_39 vdd gnd cell_6t
Xbit_r40_c104 bl_104 br_104 wl_40 vdd gnd cell_6t
Xbit_r41_c104 bl_104 br_104 wl_41 vdd gnd cell_6t
Xbit_r42_c104 bl_104 br_104 wl_42 vdd gnd cell_6t
Xbit_r43_c104 bl_104 br_104 wl_43 vdd gnd cell_6t
Xbit_r44_c104 bl_104 br_104 wl_44 vdd gnd cell_6t
Xbit_r45_c104 bl_104 br_104 wl_45 vdd gnd cell_6t
Xbit_r46_c104 bl_104 br_104 wl_46 vdd gnd cell_6t
Xbit_r47_c104 bl_104 br_104 wl_47 vdd gnd cell_6t
Xbit_r48_c104 bl_104 br_104 wl_48 vdd gnd cell_6t
Xbit_r49_c104 bl_104 br_104 wl_49 vdd gnd cell_6t
Xbit_r50_c104 bl_104 br_104 wl_50 vdd gnd cell_6t
Xbit_r51_c104 bl_104 br_104 wl_51 vdd gnd cell_6t
Xbit_r52_c104 bl_104 br_104 wl_52 vdd gnd cell_6t
Xbit_r53_c104 bl_104 br_104 wl_53 vdd gnd cell_6t
Xbit_r54_c104 bl_104 br_104 wl_54 vdd gnd cell_6t
Xbit_r55_c104 bl_104 br_104 wl_55 vdd gnd cell_6t
Xbit_r56_c104 bl_104 br_104 wl_56 vdd gnd cell_6t
Xbit_r57_c104 bl_104 br_104 wl_57 vdd gnd cell_6t
Xbit_r58_c104 bl_104 br_104 wl_58 vdd gnd cell_6t
Xbit_r59_c104 bl_104 br_104 wl_59 vdd gnd cell_6t
Xbit_r60_c104 bl_104 br_104 wl_60 vdd gnd cell_6t
Xbit_r61_c104 bl_104 br_104 wl_61 vdd gnd cell_6t
Xbit_r62_c104 bl_104 br_104 wl_62 vdd gnd cell_6t
Xbit_r63_c104 bl_104 br_104 wl_63 vdd gnd cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd cell_6t
Xbit_r1_c105 bl_105 br_105 wl_1 vdd gnd cell_6t
Xbit_r2_c105 bl_105 br_105 wl_2 vdd gnd cell_6t
Xbit_r3_c105 bl_105 br_105 wl_3 vdd gnd cell_6t
Xbit_r4_c105 bl_105 br_105 wl_4 vdd gnd cell_6t
Xbit_r5_c105 bl_105 br_105 wl_5 vdd gnd cell_6t
Xbit_r6_c105 bl_105 br_105 wl_6 vdd gnd cell_6t
Xbit_r7_c105 bl_105 br_105 wl_7 vdd gnd cell_6t
Xbit_r8_c105 bl_105 br_105 wl_8 vdd gnd cell_6t
Xbit_r9_c105 bl_105 br_105 wl_9 vdd gnd cell_6t
Xbit_r10_c105 bl_105 br_105 wl_10 vdd gnd cell_6t
Xbit_r11_c105 bl_105 br_105 wl_11 vdd gnd cell_6t
Xbit_r12_c105 bl_105 br_105 wl_12 vdd gnd cell_6t
Xbit_r13_c105 bl_105 br_105 wl_13 vdd gnd cell_6t
Xbit_r14_c105 bl_105 br_105 wl_14 vdd gnd cell_6t
Xbit_r15_c105 bl_105 br_105 wl_15 vdd gnd cell_6t
Xbit_r16_c105 bl_105 br_105 wl_16 vdd gnd cell_6t
Xbit_r17_c105 bl_105 br_105 wl_17 vdd gnd cell_6t
Xbit_r18_c105 bl_105 br_105 wl_18 vdd gnd cell_6t
Xbit_r19_c105 bl_105 br_105 wl_19 vdd gnd cell_6t
Xbit_r20_c105 bl_105 br_105 wl_20 vdd gnd cell_6t
Xbit_r21_c105 bl_105 br_105 wl_21 vdd gnd cell_6t
Xbit_r22_c105 bl_105 br_105 wl_22 vdd gnd cell_6t
Xbit_r23_c105 bl_105 br_105 wl_23 vdd gnd cell_6t
Xbit_r24_c105 bl_105 br_105 wl_24 vdd gnd cell_6t
Xbit_r25_c105 bl_105 br_105 wl_25 vdd gnd cell_6t
Xbit_r26_c105 bl_105 br_105 wl_26 vdd gnd cell_6t
Xbit_r27_c105 bl_105 br_105 wl_27 vdd gnd cell_6t
Xbit_r28_c105 bl_105 br_105 wl_28 vdd gnd cell_6t
Xbit_r29_c105 bl_105 br_105 wl_29 vdd gnd cell_6t
Xbit_r30_c105 bl_105 br_105 wl_30 vdd gnd cell_6t
Xbit_r31_c105 bl_105 br_105 wl_31 vdd gnd cell_6t
Xbit_r32_c105 bl_105 br_105 wl_32 vdd gnd cell_6t
Xbit_r33_c105 bl_105 br_105 wl_33 vdd gnd cell_6t
Xbit_r34_c105 bl_105 br_105 wl_34 vdd gnd cell_6t
Xbit_r35_c105 bl_105 br_105 wl_35 vdd gnd cell_6t
Xbit_r36_c105 bl_105 br_105 wl_36 vdd gnd cell_6t
Xbit_r37_c105 bl_105 br_105 wl_37 vdd gnd cell_6t
Xbit_r38_c105 bl_105 br_105 wl_38 vdd gnd cell_6t
Xbit_r39_c105 bl_105 br_105 wl_39 vdd gnd cell_6t
Xbit_r40_c105 bl_105 br_105 wl_40 vdd gnd cell_6t
Xbit_r41_c105 bl_105 br_105 wl_41 vdd gnd cell_6t
Xbit_r42_c105 bl_105 br_105 wl_42 vdd gnd cell_6t
Xbit_r43_c105 bl_105 br_105 wl_43 vdd gnd cell_6t
Xbit_r44_c105 bl_105 br_105 wl_44 vdd gnd cell_6t
Xbit_r45_c105 bl_105 br_105 wl_45 vdd gnd cell_6t
Xbit_r46_c105 bl_105 br_105 wl_46 vdd gnd cell_6t
Xbit_r47_c105 bl_105 br_105 wl_47 vdd gnd cell_6t
Xbit_r48_c105 bl_105 br_105 wl_48 vdd gnd cell_6t
Xbit_r49_c105 bl_105 br_105 wl_49 vdd gnd cell_6t
Xbit_r50_c105 bl_105 br_105 wl_50 vdd gnd cell_6t
Xbit_r51_c105 bl_105 br_105 wl_51 vdd gnd cell_6t
Xbit_r52_c105 bl_105 br_105 wl_52 vdd gnd cell_6t
Xbit_r53_c105 bl_105 br_105 wl_53 vdd gnd cell_6t
Xbit_r54_c105 bl_105 br_105 wl_54 vdd gnd cell_6t
Xbit_r55_c105 bl_105 br_105 wl_55 vdd gnd cell_6t
Xbit_r56_c105 bl_105 br_105 wl_56 vdd gnd cell_6t
Xbit_r57_c105 bl_105 br_105 wl_57 vdd gnd cell_6t
Xbit_r58_c105 bl_105 br_105 wl_58 vdd gnd cell_6t
Xbit_r59_c105 bl_105 br_105 wl_59 vdd gnd cell_6t
Xbit_r60_c105 bl_105 br_105 wl_60 vdd gnd cell_6t
Xbit_r61_c105 bl_105 br_105 wl_61 vdd gnd cell_6t
Xbit_r62_c105 bl_105 br_105 wl_62 vdd gnd cell_6t
Xbit_r63_c105 bl_105 br_105 wl_63 vdd gnd cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd cell_6t
Xbit_r1_c106 bl_106 br_106 wl_1 vdd gnd cell_6t
Xbit_r2_c106 bl_106 br_106 wl_2 vdd gnd cell_6t
Xbit_r3_c106 bl_106 br_106 wl_3 vdd gnd cell_6t
Xbit_r4_c106 bl_106 br_106 wl_4 vdd gnd cell_6t
Xbit_r5_c106 bl_106 br_106 wl_5 vdd gnd cell_6t
Xbit_r6_c106 bl_106 br_106 wl_6 vdd gnd cell_6t
Xbit_r7_c106 bl_106 br_106 wl_7 vdd gnd cell_6t
Xbit_r8_c106 bl_106 br_106 wl_8 vdd gnd cell_6t
Xbit_r9_c106 bl_106 br_106 wl_9 vdd gnd cell_6t
Xbit_r10_c106 bl_106 br_106 wl_10 vdd gnd cell_6t
Xbit_r11_c106 bl_106 br_106 wl_11 vdd gnd cell_6t
Xbit_r12_c106 bl_106 br_106 wl_12 vdd gnd cell_6t
Xbit_r13_c106 bl_106 br_106 wl_13 vdd gnd cell_6t
Xbit_r14_c106 bl_106 br_106 wl_14 vdd gnd cell_6t
Xbit_r15_c106 bl_106 br_106 wl_15 vdd gnd cell_6t
Xbit_r16_c106 bl_106 br_106 wl_16 vdd gnd cell_6t
Xbit_r17_c106 bl_106 br_106 wl_17 vdd gnd cell_6t
Xbit_r18_c106 bl_106 br_106 wl_18 vdd gnd cell_6t
Xbit_r19_c106 bl_106 br_106 wl_19 vdd gnd cell_6t
Xbit_r20_c106 bl_106 br_106 wl_20 vdd gnd cell_6t
Xbit_r21_c106 bl_106 br_106 wl_21 vdd gnd cell_6t
Xbit_r22_c106 bl_106 br_106 wl_22 vdd gnd cell_6t
Xbit_r23_c106 bl_106 br_106 wl_23 vdd gnd cell_6t
Xbit_r24_c106 bl_106 br_106 wl_24 vdd gnd cell_6t
Xbit_r25_c106 bl_106 br_106 wl_25 vdd gnd cell_6t
Xbit_r26_c106 bl_106 br_106 wl_26 vdd gnd cell_6t
Xbit_r27_c106 bl_106 br_106 wl_27 vdd gnd cell_6t
Xbit_r28_c106 bl_106 br_106 wl_28 vdd gnd cell_6t
Xbit_r29_c106 bl_106 br_106 wl_29 vdd gnd cell_6t
Xbit_r30_c106 bl_106 br_106 wl_30 vdd gnd cell_6t
Xbit_r31_c106 bl_106 br_106 wl_31 vdd gnd cell_6t
Xbit_r32_c106 bl_106 br_106 wl_32 vdd gnd cell_6t
Xbit_r33_c106 bl_106 br_106 wl_33 vdd gnd cell_6t
Xbit_r34_c106 bl_106 br_106 wl_34 vdd gnd cell_6t
Xbit_r35_c106 bl_106 br_106 wl_35 vdd gnd cell_6t
Xbit_r36_c106 bl_106 br_106 wl_36 vdd gnd cell_6t
Xbit_r37_c106 bl_106 br_106 wl_37 vdd gnd cell_6t
Xbit_r38_c106 bl_106 br_106 wl_38 vdd gnd cell_6t
Xbit_r39_c106 bl_106 br_106 wl_39 vdd gnd cell_6t
Xbit_r40_c106 bl_106 br_106 wl_40 vdd gnd cell_6t
Xbit_r41_c106 bl_106 br_106 wl_41 vdd gnd cell_6t
Xbit_r42_c106 bl_106 br_106 wl_42 vdd gnd cell_6t
Xbit_r43_c106 bl_106 br_106 wl_43 vdd gnd cell_6t
Xbit_r44_c106 bl_106 br_106 wl_44 vdd gnd cell_6t
Xbit_r45_c106 bl_106 br_106 wl_45 vdd gnd cell_6t
Xbit_r46_c106 bl_106 br_106 wl_46 vdd gnd cell_6t
Xbit_r47_c106 bl_106 br_106 wl_47 vdd gnd cell_6t
Xbit_r48_c106 bl_106 br_106 wl_48 vdd gnd cell_6t
Xbit_r49_c106 bl_106 br_106 wl_49 vdd gnd cell_6t
Xbit_r50_c106 bl_106 br_106 wl_50 vdd gnd cell_6t
Xbit_r51_c106 bl_106 br_106 wl_51 vdd gnd cell_6t
Xbit_r52_c106 bl_106 br_106 wl_52 vdd gnd cell_6t
Xbit_r53_c106 bl_106 br_106 wl_53 vdd gnd cell_6t
Xbit_r54_c106 bl_106 br_106 wl_54 vdd gnd cell_6t
Xbit_r55_c106 bl_106 br_106 wl_55 vdd gnd cell_6t
Xbit_r56_c106 bl_106 br_106 wl_56 vdd gnd cell_6t
Xbit_r57_c106 bl_106 br_106 wl_57 vdd gnd cell_6t
Xbit_r58_c106 bl_106 br_106 wl_58 vdd gnd cell_6t
Xbit_r59_c106 bl_106 br_106 wl_59 vdd gnd cell_6t
Xbit_r60_c106 bl_106 br_106 wl_60 vdd gnd cell_6t
Xbit_r61_c106 bl_106 br_106 wl_61 vdd gnd cell_6t
Xbit_r62_c106 bl_106 br_106 wl_62 vdd gnd cell_6t
Xbit_r63_c106 bl_106 br_106 wl_63 vdd gnd cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd cell_6t
Xbit_r1_c107 bl_107 br_107 wl_1 vdd gnd cell_6t
Xbit_r2_c107 bl_107 br_107 wl_2 vdd gnd cell_6t
Xbit_r3_c107 bl_107 br_107 wl_3 vdd gnd cell_6t
Xbit_r4_c107 bl_107 br_107 wl_4 vdd gnd cell_6t
Xbit_r5_c107 bl_107 br_107 wl_5 vdd gnd cell_6t
Xbit_r6_c107 bl_107 br_107 wl_6 vdd gnd cell_6t
Xbit_r7_c107 bl_107 br_107 wl_7 vdd gnd cell_6t
Xbit_r8_c107 bl_107 br_107 wl_8 vdd gnd cell_6t
Xbit_r9_c107 bl_107 br_107 wl_9 vdd gnd cell_6t
Xbit_r10_c107 bl_107 br_107 wl_10 vdd gnd cell_6t
Xbit_r11_c107 bl_107 br_107 wl_11 vdd gnd cell_6t
Xbit_r12_c107 bl_107 br_107 wl_12 vdd gnd cell_6t
Xbit_r13_c107 bl_107 br_107 wl_13 vdd gnd cell_6t
Xbit_r14_c107 bl_107 br_107 wl_14 vdd gnd cell_6t
Xbit_r15_c107 bl_107 br_107 wl_15 vdd gnd cell_6t
Xbit_r16_c107 bl_107 br_107 wl_16 vdd gnd cell_6t
Xbit_r17_c107 bl_107 br_107 wl_17 vdd gnd cell_6t
Xbit_r18_c107 bl_107 br_107 wl_18 vdd gnd cell_6t
Xbit_r19_c107 bl_107 br_107 wl_19 vdd gnd cell_6t
Xbit_r20_c107 bl_107 br_107 wl_20 vdd gnd cell_6t
Xbit_r21_c107 bl_107 br_107 wl_21 vdd gnd cell_6t
Xbit_r22_c107 bl_107 br_107 wl_22 vdd gnd cell_6t
Xbit_r23_c107 bl_107 br_107 wl_23 vdd gnd cell_6t
Xbit_r24_c107 bl_107 br_107 wl_24 vdd gnd cell_6t
Xbit_r25_c107 bl_107 br_107 wl_25 vdd gnd cell_6t
Xbit_r26_c107 bl_107 br_107 wl_26 vdd gnd cell_6t
Xbit_r27_c107 bl_107 br_107 wl_27 vdd gnd cell_6t
Xbit_r28_c107 bl_107 br_107 wl_28 vdd gnd cell_6t
Xbit_r29_c107 bl_107 br_107 wl_29 vdd gnd cell_6t
Xbit_r30_c107 bl_107 br_107 wl_30 vdd gnd cell_6t
Xbit_r31_c107 bl_107 br_107 wl_31 vdd gnd cell_6t
Xbit_r32_c107 bl_107 br_107 wl_32 vdd gnd cell_6t
Xbit_r33_c107 bl_107 br_107 wl_33 vdd gnd cell_6t
Xbit_r34_c107 bl_107 br_107 wl_34 vdd gnd cell_6t
Xbit_r35_c107 bl_107 br_107 wl_35 vdd gnd cell_6t
Xbit_r36_c107 bl_107 br_107 wl_36 vdd gnd cell_6t
Xbit_r37_c107 bl_107 br_107 wl_37 vdd gnd cell_6t
Xbit_r38_c107 bl_107 br_107 wl_38 vdd gnd cell_6t
Xbit_r39_c107 bl_107 br_107 wl_39 vdd gnd cell_6t
Xbit_r40_c107 bl_107 br_107 wl_40 vdd gnd cell_6t
Xbit_r41_c107 bl_107 br_107 wl_41 vdd gnd cell_6t
Xbit_r42_c107 bl_107 br_107 wl_42 vdd gnd cell_6t
Xbit_r43_c107 bl_107 br_107 wl_43 vdd gnd cell_6t
Xbit_r44_c107 bl_107 br_107 wl_44 vdd gnd cell_6t
Xbit_r45_c107 bl_107 br_107 wl_45 vdd gnd cell_6t
Xbit_r46_c107 bl_107 br_107 wl_46 vdd gnd cell_6t
Xbit_r47_c107 bl_107 br_107 wl_47 vdd gnd cell_6t
Xbit_r48_c107 bl_107 br_107 wl_48 vdd gnd cell_6t
Xbit_r49_c107 bl_107 br_107 wl_49 vdd gnd cell_6t
Xbit_r50_c107 bl_107 br_107 wl_50 vdd gnd cell_6t
Xbit_r51_c107 bl_107 br_107 wl_51 vdd gnd cell_6t
Xbit_r52_c107 bl_107 br_107 wl_52 vdd gnd cell_6t
Xbit_r53_c107 bl_107 br_107 wl_53 vdd gnd cell_6t
Xbit_r54_c107 bl_107 br_107 wl_54 vdd gnd cell_6t
Xbit_r55_c107 bl_107 br_107 wl_55 vdd gnd cell_6t
Xbit_r56_c107 bl_107 br_107 wl_56 vdd gnd cell_6t
Xbit_r57_c107 bl_107 br_107 wl_57 vdd gnd cell_6t
Xbit_r58_c107 bl_107 br_107 wl_58 vdd gnd cell_6t
Xbit_r59_c107 bl_107 br_107 wl_59 vdd gnd cell_6t
Xbit_r60_c107 bl_107 br_107 wl_60 vdd gnd cell_6t
Xbit_r61_c107 bl_107 br_107 wl_61 vdd gnd cell_6t
Xbit_r62_c107 bl_107 br_107 wl_62 vdd gnd cell_6t
Xbit_r63_c107 bl_107 br_107 wl_63 vdd gnd cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd cell_6t
Xbit_r1_c108 bl_108 br_108 wl_1 vdd gnd cell_6t
Xbit_r2_c108 bl_108 br_108 wl_2 vdd gnd cell_6t
Xbit_r3_c108 bl_108 br_108 wl_3 vdd gnd cell_6t
Xbit_r4_c108 bl_108 br_108 wl_4 vdd gnd cell_6t
Xbit_r5_c108 bl_108 br_108 wl_5 vdd gnd cell_6t
Xbit_r6_c108 bl_108 br_108 wl_6 vdd gnd cell_6t
Xbit_r7_c108 bl_108 br_108 wl_7 vdd gnd cell_6t
Xbit_r8_c108 bl_108 br_108 wl_8 vdd gnd cell_6t
Xbit_r9_c108 bl_108 br_108 wl_9 vdd gnd cell_6t
Xbit_r10_c108 bl_108 br_108 wl_10 vdd gnd cell_6t
Xbit_r11_c108 bl_108 br_108 wl_11 vdd gnd cell_6t
Xbit_r12_c108 bl_108 br_108 wl_12 vdd gnd cell_6t
Xbit_r13_c108 bl_108 br_108 wl_13 vdd gnd cell_6t
Xbit_r14_c108 bl_108 br_108 wl_14 vdd gnd cell_6t
Xbit_r15_c108 bl_108 br_108 wl_15 vdd gnd cell_6t
Xbit_r16_c108 bl_108 br_108 wl_16 vdd gnd cell_6t
Xbit_r17_c108 bl_108 br_108 wl_17 vdd gnd cell_6t
Xbit_r18_c108 bl_108 br_108 wl_18 vdd gnd cell_6t
Xbit_r19_c108 bl_108 br_108 wl_19 vdd gnd cell_6t
Xbit_r20_c108 bl_108 br_108 wl_20 vdd gnd cell_6t
Xbit_r21_c108 bl_108 br_108 wl_21 vdd gnd cell_6t
Xbit_r22_c108 bl_108 br_108 wl_22 vdd gnd cell_6t
Xbit_r23_c108 bl_108 br_108 wl_23 vdd gnd cell_6t
Xbit_r24_c108 bl_108 br_108 wl_24 vdd gnd cell_6t
Xbit_r25_c108 bl_108 br_108 wl_25 vdd gnd cell_6t
Xbit_r26_c108 bl_108 br_108 wl_26 vdd gnd cell_6t
Xbit_r27_c108 bl_108 br_108 wl_27 vdd gnd cell_6t
Xbit_r28_c108 bl_108 br_108 wl_28 vdd gnd cell_6t
Xbit_r29_c108 bl_108 br_108 wl_29 vdd gnd cell_6t
Xbit_r30_c108 bl_108 br_108 wl_30 vdd gnd cell_6t
Xbit_r31_c108 bl_108 br_108 wl_31 vdd gnd cell_6t
Xbit_r32_c108 bl_108 br_108 wl_32 vdd gnd cell_6t
Xbit_r33_c108 bl_108 br_108 wl_33 vdd gnd cell_6t
Xbit_r34_c108 bl_108 br_108 wl_34 vdd gnd cell_6t
Xbit_r35_c108 bl_108 br_108 wl_35 vdd gnd cell_6t
Xbit_r36_c108 bl_108 br_108 wl_36 vdd gnd cell_6t
Xbit_r37_c108 bl_108 br_108 wl_37 vdd gnd cell_6t
Xbit_r38_c108 bl_108 br_108 wl_38 vdd gnd cell_6t
Xbit_r39_c108 bl_108 br_108 wl_39 vdd gnd cell_6t
Xbit_r40_c108 bl_108 br_108 wl_40 vdd gnd cell_6t
Xbit_r41_c108 bl_108 br_108 wl_41 vdd gnd cell_6t
Xbit_r42_c108 bl_108 br_108 wl_42 vdd gnd cell_6t
Xbit_r43_c108 bl_108 br_108 wl_43 vdd gnd cell_6t
Xbit_r44_c108 bl_108 br_108 wl_44 vdd gnd cell_6t
Xbit_r45_c108 bl_108 br_108 wl_45 vdd gnd cell_6t
Xbit_r46_c108 bl_108 br_108 wl_46 vdd gnd cell_6t
Xbit_r47_c108 bl_108 br_108 wl_47 vdd gnd cell_6t
Xbit_r48_c108 bl_108 br_108 wl_48 vdd gnd cell_6t
Xbit_r49_c108 bl_108 br_108 wl_49 vdd gnd cell_6t
Xbit_r50_c108 bl_108 br_108 wl_50 vdd gnd cell_6t
Xbit_r51_c108 bl_108 br_108 wl_51 vdd gnd cell_6t
Xbit_r52_c108 bl_108 br_108 wl_52 vdd gnd cell_6t
Xbit_r53_c108 bl_108 br_108 wl_53 vdd gnd cell_6t
Xbit_r54_c108 bl_108 br_108 wl_54 vdd gnd cell_6t
Xbit_r55_c108 bl_108 br_108 wl_55 vdd gnd cell_6t
Xbit_r56_c108 bl_108 br_108 wl_56 vdd gnd cell_6t
Xbit_r57_c108 bl_108 br_108 wl_57 vdd gnd cell_6t
Xbit_r58_c108 bl_108 br_108 wl_58 vdd gnd cell_6t
Xbit_r59_c108 bl_108 br_108 wl_59 vdd gnd cell_6t
Xbit_r60_c108 bl_108 br_108 wl_60 vdd gnd cell_6t
Xbit_r61_c108 bl_108 br_108 wl_61 vdd gnd cell_6t
Xbit_r62_c108 bl_108 br_108 wl_62 vdd gnd cell_6t
Xbit_r63_c108 bl_108 br_108 wl_63 vdd gnd cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd cell_6t
Xbit_r1_c109 bl_109 br_109 wl_1 vdd gnd cell_6t
Xbit_r2_c109 bl_109 br_109 wl_2 vdd gnd cell_6t
Xbit_r3_c109 bl_109 br_109 wl_3 vdd gnd cell_6t
Xbit_r4_c109 bl_109 br_109 wl_4 vdd gnd cell_6t
Xbit_r5_c109 bl_109 br_109 wl_5 vdd gnd cell_6t
Xbit_r6_c109 bl_109 br_109 wl_6 vdd gnd cell_6t
Xbit_r7_c109 bl_109 br_109 wl_7 vdd gnd cell_6t
Xbit_r8_c109 bl_109 br_109 wl_8 vdd gnd cell_6t
Xbit_r9_c109 bl_109 br_109 wl_9 vdd gnd cell_6t
Xbit_r10_c109 bl_109 br_109 wl_10 vdd gnd cell_6t
Xbit_r11_c109 bl_109 br_109 wl_11 vdd gnd cell_6t
Xbit_r12_c109 bl_109 br_109 wl_12 vdd gnd cell_6t
Xbit_r13_c109 bl_109 br_109 wl_13 vdd gnd cell_6t
Xbit_r14_c109 bl_109 br_109 wl_14 vdd gnd cell_6t
Xbit_r15_c109 bl_109 br_109 wl_15 vdd gnd cell_6t
Xbit_r16_c109 bl_109 br_109 wl_16 vdd gnd cell_6t
Xbit_r17_c109 bl_109 br_109 wl_17 vdd gnd cell_6t
Xbit_r18_c109 bl_109 br_109 wl_18 vdd gnd cell_6t
Xbit_r19_c109 bl_109 br_109 wl_19 vdd gnd cell_6t
Xbit_r20_c109 bl_109 br_109 wl_20 vdd gnd cell_6t
Xbit_r21_c109 bl_109 br_109 wl_21 vdd gnd cell_6t
Xbit_r22_c109 bl_109 br_109 wl_22 vdd gnd cell_6t
Xbit_r23_c109 bl_109 br_109 wl_23 vdd gnd cell_6t
Xbit_r24_c109 bl_109 br_109 wl_24 vdd gnd cell_6t
Xbit_r25_c109 bl_109 br_109 wl_25 vdd gnd cell_6t
Xbit_r26_c109 bl_109 br_109 wl_26 vdd gnd cell_6t
Xbit_r27_c109 bl_109 br_109 wl_27 vdd gnd cell_6t
Xbit_r28_c109 bl_109 br_109 wl_28 vdd gnd cell_6t
Xbit_r29_c109 bl_109 br_109 wl_29 vdd gnd cell_6t
Xbit_r30_c109 bl_109 br_109 wl_30 vdd gnd cell_6t
Xbit_r31_c109 bl_109 br_109 wl_31 vdd gnd cell_6t
Xbit_r32_c109 bl_109 br_109 wl_32 vdd gnd cell_6t
Xbit_r33_c109 bl_109 br_109 wl_33 vdd gnd cell_6t
Xbit_r34_c109 bl_109 br_109 wl_34 vdd gnd cell_6t
Xbit_r35_c109 bl_109 br_109 wl_35 vdd gnd cell_6t
Xbit_r36_c109 bl_109 br_109 wl_36 vdd gnd cell_6t
Xbit_r37_c109 bl_109 br_109 wl_37 vdd gnd cell_6t
Xbit_r38_c109 bl_109 br_109 wl_38 vdd gnd cell_6t
Xbit_r39_c109 bl_109 br_109 wl_39 vdd gnd cell_6t
Xbit_r40_c109 bl_109 br_109 wl_40 vdd gnd cell_6t
Xbit_r41_c109 bl_109 br_109 wl_41 vdd gnd cell_6t
Xbit_r42_c109 bl_109 br_109 wl_42 vdd gnd cell_6t
Xbit_r43_c109 bl_109 br_109 wl_43 vdd gnd cell_6t
Xbit_r44_c109 bl_109 br_109 wl_44 vdd gnd cell_6t
Xbit_r45_c109 bl_109 br_109 wl_45 vdd gnd cell_6t
Xbit_r46_c109 bl_109 br_109 wl_46 vdd gnd cell_6t
Xbit_r47_c109 bl_109 br_109 wl_47 vdd gnd cell_6t
Xbit_r48_c109 bl_109 br_109 wl_48 vdd gnd cell_6t
Xbit_r49_c109 bl_109 br_109 wl_49 vdd gnd cell_6t
Xbit_r50_c109 bl_109 br_109 wl_50 vdd gnd cell_6t
Xbit_r51_c109 bl_109 br_109 wl_51 vdd gnd cell_6t
Xbit_r52_c109 bl_109 br_109 wl_52 vdd gnd cell_6t
Xbit_r53_c109 bl_109 br_109 wl_53 vdd gnd cell_6t
Xbit_r54_c109 bl_109 br_109 wl_54 vdd gnd cell_6t
Xbit_r55_c109 bl_109 br_109 wl_55 vdd gnd cell_6t
Xbit_r56_c109 bl_109 br_109 wl_56 vdd gnd cell_6t
Xbit_r57_c109 bl_109 br_109 wl_57 vdd gnd cell_6t
Xbit_r58_c109 bl_109 br_109 wl_58 vdd gnd cell_6t
Xbit_r59_c109 bl_109 br_109 wl_59 vdd gnd cell_6t
Xbit_r60_c109 bl_109 br_109 wl_60 vdd gnd cell_6t
Xbit_r61_c109 bl_109 br_109 wl_61 vdd gnd cell_6t
Xbit_r62_c109 bl_109 br_109 wl_62 vdd gnd cell_6t
Xbit_r63_c109 bl_109 br_109 wl_63 vdd gnd cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd cell_6t
Xbit_r1_c110 bl_110 br_110 wl_1 vdd gnd cell_6t
Xbit_r2_c110 bl_110 br_110 wl_2 vdd gnd cell_6t
Xbit_r3_c110 bl_110 br_110 wl_3 vdd gnd cell_6t
Xbit_r4_c110 bl_110 br_110 wl_4 vdd gnd cell_6t
Xbit_r5_c110 bl_110 br_110 wl_5 vdd gnd cell_6t
Xbit_r6_c110 bl_110 br_110 wl_6 vdd gnd cell_6t
Xbit_r7_c110 bl_110 br_110 wl_7 vdd gnd cell_6t
Xbit_r8_c110 bl_110 br_110 wl_8 vdd gnd cell_6t
Xbit_r9_c110 bl_110 br_110 wl_9 vdd gnd cell_6t
Xbit_r10_c110 bl_110 br_110 wl_10 vdd gnd cell_6t
Xbit_r11_c110 bl_110 br_110 wl_11 vdd gnd cell_6t
Xbit_r12_c110 bl_110 br_110 wl_12 vdd gnd cell_6t
Xbit_r13_c110 bl_110 br_110 wl_13 vdd gnd cell_6t
Xbit_r14_c110 bl_110 br_110 wl_14 vdd gnd cell_6t
Xbit_r15_c110 bl_110 br_110 wl_15 vdd gnd cell_6t
Xbit_r16_c110 bl_110 br_110 wl_16 vdd gnd cell_6t
Xbit_r17_c110 bl_110 br_110 wl_17 vdd gnd cell_6t
Xbit_r18_c110 bl_110 br_110 wl_18 vdd gnd cell_6t
Xbit_r19_c110 bl_110 br_110 wl_19 vdd gnd cell_6t
Xbit_r20_c110 bl_110 br_110 wl_20 vdd gnd cell_6t
Xbit_r21_c110 bl_110 br_110 wl_21 vdd gnd cell_6t
Xbit_r22_c110 bl_110 br_110 wl_22 vdd gnd cell_6t
Xbit_r23_c110 bl_110 br_110 wl_23 vdd gnd cell_6t
Xbit_r24_c110 bl_110 br_110 wl_24 vdd gnd cell_6t
Xbit_r25_c110 bl_110 br_110 wl_25 vdd gnd cell_6t
Xbit_r26_c110 bl_110 br_110 wl_26 vdd gnd cell_6t
Xbit_r27_c110 bl_110 br_110 wl_27 vdd gnd cell_6t
Xbit_r28_c110 bl_110 br_110 wl_28 vdd gnd cell_6t
Xbit_r29_c110 bl_110 br_110 wl_29 vdd gnd cell_6t
Xbit_r30_c110 bl_110 br_110 wl_30 vdd gnd cell_6t
Xbit_r31_c110 bl_110 br_110 wl_31 vdd gnd cell_6t
Xbit_r32_c110 bl_110 br_110 wl_32 vdd gnd cell_6t
Xbit_r33_c110 bl_110 br_110 wl_33 vdd gnd cell_6t
Xbit_r34_c110 bl_110 br_110 wl_34 vdd gnd cell_6t
Xbit_r35_c110 bl_110 br_110 wl_35 vdd gnd cell_6t
Xbit_r36_c110 bl_110 br_110 wl_36 vdd gnd cell_6t
Xbit_r37_c110 bl_110 br_110 wl_37 vdd gnd cell_6t
Xbit_r38_c110 bl_110 br_110 wl_38 vdd gnd cell_6t
Xbit_r39_c110 bl_110 br_110 wl_39 vdd gnd cell_6t
Xbit_r40_c110 bl_110 br_110 wl_40 vdd gnd cell_6t
Xbit_r41_c110 bl_110 br_110 wl_41 vdd gnd cell_6t
Xbit_r42_c110 bl_110 br_110 wl_42 vdd gnd cell_6t
Xbit_r43_c110 bl_110 br_110 wl_43 vdd gnd cell_6t
Xbit_r44_c110 bl_110 br_110 wl_44 vdd gnd cell_6t
Xbit_r45_c110 bl_110 br_110 wl_45 vdd gnd cell_6t
Xbit_r46_c110 bl_110 br_110 wl_46 vdd gnd cell_6t
Xbit_r47_c110 bl_110 br_110 wl_47 vdd gnd cell_6t
Xbit_r48_c110 bl_110 br_110 wl_48 vdd gnd cell_6t
Xbit_r49_c110 bl_110 br_110 wl_49 vdd gnd cell_6t
Xbit_r50_c110 bl_110 br_110 wl_50 vdd gnd cell_6t
Xbit_r51_c110 bl_110 br_110 wl_51 vdd gnd cell_6t
Xbit_r52_c110 bl_110 br_110 wl_52 vdd gnd cell_6t
Xbit_r53_c110 bl_110 br_110 wl_53 vdd gnd cell_6t
Xbit_r54_c110 bl_110 br_110 wl_54 vdd gnd cell_6t
Xbit_r55_c110 bl_110 br_110 wl_55 vdd gnd cell_6t
Xbit_r56_c110 bl_110 br_110 wl_56 vdd gnd cell_6t
Xbit_r57_c110 bl_110 br_110 wl_57 vdd gnd cell_6t
Xbit_r58_c110 bl_110 br_110 wl_58 vdd gnd cell_6t
Xbit_r59_c110 bl_110 br_110 wl_59 vdd gnd cell_6t
Xbit_r60_c110 bl_110 br_110 wl_60 vdd gnd cell_6t
Xbit_r61_c110 bl_110 br_110 wl_61 vdd gnd cell_6t
Xbit_r62_c110 bl_110 br_110 wl_62 vdd gnd cell_6t
Xbit_r63_c110 bl_110 br_110 wl_63 vdd gnd cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd cell_6t
Xbit_r1_c111 bl_111 br_111 wl_1 vdd gnd cell_6t
Xbit_r2_c111 bl_111 br_111 wl_2 vdd gnd cell_6t
Xbit_r3_c111 bl_111 br_111 wl_3 vdd gnd cell_6t
Xbit_r4_c111 bl_111 br_111 wl_4 vdd gnd cell_6t
Xbit_r5_c111 bl_111 br_111 wl_5 vdd gnd cell_6t
Xbit_r6_c111 bl_111 br_111 wl_6 vdd gnd cell_6t
Xbit_r7_c111 bl_111 br_111 wl_7 vdd gnd cell_6t
Xbit_r8_c111 bl_111 br_111 wl_8 vdd gnd cell_6t
Xbit_r9_c111 bl_111 br_111 wl_9 vdd gnd cell_6t
Xbit_r10_c111 bl_111 br_111 wl_10 vdd gnd cell_6t
Xbit_r11_c111 bl_111 br_111 wl_11 vdd gnd cell_6t
Xbit_r12_c111 bl_111 br_111 wl_12 vdd gnd cell_6t
Xbit_r13_c111 bl_111 br_111 wl_13 vdd gnd cell_6t
Xbit_r14_c111 bl_111 br_111 wl_14 vdd gnd cell_6t
Xbit_r15_c111 bl_111 br_111 wl_15 vdd gnd cell_6t
Xbit_r16_c111 bl_111 br_111 wl_16 vdd gnd cell_6t
Xbit_r17_c111 bl_111 br_111 wl_17 vdd gnd cell_6t
Xbit_r18_c111 bl_111 br_111 wl_18 vdd gnd cell_6t
Xbit_r19_c111 bl_111 br_111 wl_19 vdd gnd cell_6t
Xbit_r20_c111 bl_111 br_111 wl_20 vdd gnd cell_6t
Xbit_r21_c111 bl_111 br_111 wl_21 vdd gnd cell_6t
Xbit_r22_c111 bl_111 br_111 wl_22 vdd gnd cell_6t
Xbit_r23_c111 bl_111 br_111 wl_23 vdd gnd cell_6t
Xbit_r24_c111 bl_111 br_111 wl_24 vdd gnd cell_6t
Xbit_r25_c111 bl_111 br_111 wl_25 vdd gnd cell_6t
Xbit_r26_c111 bl_111 br_111 wl_26 vdd gnd cell_6t
Xbit_r27_c111 bl_111 br_111 wl_27 vdd gnd cell_6t
Xbit_r28_c111 bl_111 br_111 wl_28 vdd gnd cell_6t
Xbit_r29_c111 bl_111 br_111 wl_29 vdd gnd cell_6t
Xbit_r30_c111 bl_111 br_111 wl_30 vdd gnd cell_6t
Xbit_r31_c111 bl_111 br_111 wl_31 vdd gnd cell_6t
Xbit_r32_c111 bl_111 br_111 wl_32 vdd gnd cell_6t
Xbit_r33_c111 bl_111 br_111 wl_33 vdd gnd cell_6t
Xbit_r34_c111 bl_111 br_111 wl_34 vdd gnd cell_6t
Xbit_r35_c111 bl_111 br_111 wl_35 vdd gnd cell_6t
Xbit_r36_c111 bl_111 br_111 wl_36 vdd gnd cell_6t
Xbit_r37_c111 bl_111 br_111 wl_37 vdd gnd cell_6t
Xbit_r38_c111 bl_111 br_111 wl_38 vdd gnd cell_6t
Xbit_r39_c111 bl_111 br_111 wl_39 vdd gnd cell_6t
Xbit_r40_c111 bl_111 br_111 wl_40 vdd gnd cell_6t
Xbit_r41_c111 bl_111 br_111 wl_41 vdd gnd cell_6t
Xbit_r42_c111 bl_111 br_111 wl_42 vdd gnd cell_6t
Xbit_r43_c111 bl_111 br_111 wl_43 vdd gnd cell_6t
Xbit_r44_c111 bl_111 br_111 wl_44 vdd gnd cell_6t
Xbit_r45_c111 bl_111 br_111 wl_45 vdd gnd cell_6t
Xbit_r46_c111 bl_111 br_111 wl_46 vdd gnd cell_6t
Xbit_r47_c111 bl_111 br_111 wl_47 vdd gnd cell_6t
Xbit_r48_c111 bl_111 br_111 wl_48 vdd gnd cell_6t
Xbit_r49_c111 bl_111 br_111 wl_49 vdd gnd cell_6t
Xbit_r50_c111 bl_111 br_111 wl_50 vdd gnd cell_6t
Xbit_r51_c111 bl_111 br_111 wl_51 vdd gnd cell_6t
Xbit_r52_c111 bl_111 br_111 wl_52 vdd gnd cell_6t
Xbit_r53_c111 bl_111 br_111 wl_53 vdd gnd cell_6t
Xbit_r54_c111 bl_111 br_111 wl_54 vdd gnd cell_6t
Xbit_r55_c111 bl_111 br_111 wl_55 vdd gnd cell_6t
Xbit_r56_c111 bl_111 br_111 wl_56 vdd gnd cell_6t
Xbit_r57_c111 bl_111 br_111 wl_57 vdd gnd cell_6t
Xbit_r58_c111 bl_111 br_111 wl_58 vdd gnd cell_6t
Xbit_r59_c111 bl_111 br_111 wl_59 vdd gnd cell_6t
Xbit_r60_c111 bl_111 br_111 wl_60 vdd gnd cell_6t
Xbit_r61_c111 bl_111 br_111 wl_61 vdd gnd cell_6t
Xbit_r62_c111 bl_111 br_111 wl_62 vdd gnd cell_6t
Xbit_r63_c111 bl_111 br_111 wl_63 vdd gnd cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd cell_6t
Xbit_r1_c112 bl_112 br_112 wl_1 vdd gnd cell_6t
Xbit_r2_c112 bl_112 br_112 wl_2 vdd gnd cell_6t
Xbit_r3_c112 bl_112 br_112 wl_3 vdd gnd cell_6t
Xbit_r4_c112 bl_112 br_112 wl_4 vdd gnd cell_6t
Xbit_r5_c112 bl_112 br_112 wl_5 vdd gnd cell_6t
Xbit_r6_c112 bl_112 br_112 wl_6 vdd gnd cell_6t
Xbit_r7_c112 bl_112 br_112 wl_7 vdd gnd cell_6t
Xbit_r8_c112 bl_112 br_112 wl_8 vdd gnd cell_6t
Xbit_r9_c112 bl_112 br_112 wl_9 vdd gnd cell_6t
Xbit_r10_c112 bl_112 br_112 wl_10 vdd gnd cell_6t
Xbit_r11_c112 bl_112 br_112 wl_11 vdd gnd cell_6t
Xbit_r12_c112 bl_112 br_112 wl_12 vdd gnd cell_6t
Xbit_r13_c112 bl_112 br_112 wl_13 vdd gnd cell_6t
Xbit_r14_c112 bl_112 br_112 wl_14 vdd gnd cell_6t
Xbit_r15_c112 bl_112 br_112 wl_15 vdd gnd cell_6t
Xbit_r16_c112 bl_112 br_112 wl_16 vdd gnd cell_6t
Xbit_r17_c112 bl_112 br_112 wl_17 vdd gnd cell_6t
Xbit_r18_c112 bl_112 br_112 wl_18 vdd gnd cell_6t
Xbit_r19_c112 bl_112 br_112 wl_19 vdd gnd cell_6t
Xbit_r20_c112 bl_112 br_112 wl_20 vdd gnd cell_6t
Xbit_r21_c112 bl_112 br_112 wl_21 vdd gnd cell_6t
Xbit_r22_c112 bl_112 br_112 wl_22 vdd gnd cell_6t
Xbit_r23_c112 bl_112 br_112 wl_23 vdd gnd cell_6t
Xbit_r24_c112 bl_112 br_112 wl_24 vdd gnd cell_6t
Xbit_r25_c112 bl_112 br_112 wl_25 vdd gnd cell_6t
Xbit_r26_c112 bl_112 br_112 wl_26 vdd gnd cell_6t
Xbit_r27_c112 bl_112 br_112 wl_27 vdd gnd cell_6t
Xbit_r28_c112 bl_112 br_112 wl_28 vdd gnd cell_6t
Xbit_r29_c112 bl_112 br_112 wl_29 vdd gnd cell_6t
Xbit_r30_c112 bl_112 br_112 wl_30 vdd gnd cell_6t
Xbit_r31_c112 bl_112 br_112 wl_31 vdd gnd cell_6t
Xbit_r32_c112 bl_112 br_112 wl_32 vdd gnd cell_6t
Xbit_r33_c112 bl_112 br_112 wl_33 vdd gnd cell_6t
Xbit_r34_c112 bl_112 br_112 wl_34 vdd gnd cell_6t
Xbit_r35_c112 bl_112 br_112 wl_35 vdd gnd cell_6t
Xbit_r36_c112 bl_112 br_112 wl_36 vdd gnd cell_6t
Xbit_r37_c112 bl_112 br_112 wl_37 vdd gnd cell_6t
Xbit_r38_c112 bl_112 br_112 wl_38 vdd gnd cell_6t
Xbit_r39_c112 bl_112 br_112 wl_39 vdd gnd cell_6t
Xbit_r40_c112 bl_112 br_112 wl_40 vdd gnd cell_6t
Xbit_r41_c112 bl_112 br_112 wl_41 vdd gnd cell_6t
Xbit_r42_c112 bl_112 br_112 wl_42 vdd gnd cell_6t
Xbit_r43_c112 bl_112 br_112 wl_43 vdd gnd cell_6t
Xbit_r44_c112 bl_112 br_112 wl_44 vdd gnd cell_6t
Xbit_r45_c112 bl_112 br_112 wl_45 vdd gnd cell_6t
Xbit_r46_c112 bl_112 br_112 wl_46 vdd gnd cell_6t
Xbit_r47_c112 bl_112 br_112 wl_47 vdd gnd cell_6t
Xbit_r48_c112 bl_112 br_112 wl_48 vdd gnd cell_6t
Xbit_r49_c112 bl_112 br_112 wl_49 vdd gnd cell_6t
Xbit_r50_c112 bl_112 br_112 wl_50 vdd gnd cell_6t
Xbit_r51_c112 bl_112 br_112 wl_51 vdd gnd cell_6t
Xbit_r52_c112 bl_112 br_112 wl_52 vdd gnd cell_6t
Xbit_r53_c112 bl_112 br_112 wl_53 vdd gnd cell_6t
Xbit_r54_c112 bl_112 br_112 wl_54 vdd gnd cell_6t
Xbit_r55_c112 bl_112 br_112 wl_55 vdd gnd cell_6t
Xbit_r56_c112 bl_112 br_112 wl_56 vdd gnd cell_6t
Xbit_r57_c112 bl_112 br_112 wl_57 vdd gnd cell_6t
Xbit_r58_c112 bl_112 br_112 wl_58 vdd gnd cell_6t
Xbit_r59_c112 bl_112 br_112 wl_59 vdd gnd cell_6t
Xbit_r60_c112 bl_112 br_112 wl_60 vdd gnd cell_6t
Xbit_r61_c112 bl_112 br_112 wl_61 vdd gnd cell_6t
Xbit_r62_c112 bl_112 br_112 wl_62 vdd gnd cell_6t
Xbit_r63_c112 bl_112 br_112 wl_63 vdd gnd cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd cell_6t
Xbit_r1_c113 bl_113 br_113 wl_1 vdd gnd cell_6t
Xbit_r2_c113 bl_113 br_113 wl_2 vdd gnd cell_6t
Xbit_r3_c113 bl_113 br_113 wl_3 vdd gnd cell_6t
Xbit_r4_c113 bl_113 br_113 wl_4 vdd gnd cell_6t
Xbit_r5_c113 bl_113 br_113 wl_5 vdd gnd cell_6t
Xbit_r6_c113 bl_113 br_113 wl_6 vdd gnd cell_6t
Xbit_r7_c113 bl_113 br_113 wl_7 vdd gnd cell_6t
Xbit_r8_c113 bl_113 br_113 wl_8 vdd gnd cell_6t
Xbit_r9_c113 bl_113 br_113 wl_9 vdd gnd cell_6t
Xbit_r10_c113 bl_113 br_113 wl_10 vdd gnd cell_6t
Xbit_r11_c113 bl_113 br_113 wl_11 vdd gnd cell_6t
Xbit_r12_c113 bl_113 br_113 wl_12 vdd gnd cell_6t
Xbit_r13_c113 bl_113 br_113 wl_13 vdd gnd cell_6t
Xbit_r14_c113 bl_113 br_113 wl_14 vdd gnd cell_6t
Xbit_r15_c113 bl_113 br_113 wl_15 vdd gnd cell_6t
Xbit_r16_c113 bl_113 br_113 wl_16 vdd gnd cell_6t
Xbit_r17_c113 bl_113 br_113 wl_17 vdd gnd cell_6t
Xbit_r18_c113 bl_113 br_113 wl_18 vdd gnd cell_6t
Xbit_r19_c113 bl_113 br_113 wl_19 vdd gnd cell_6t
Xbit_r20_c113 bl_113 br_113 wl_20 vdd gnd cell_6t
Xbit_r21_c113 bl_113 br_113 wl_21 vdd gnd cell_6t
Xbit_r22_c113 bl_113 br_113 wl_22 vdd gnd cell_6t
Xbit_r23_c113 bl_113 br_113 wl_23 vdd gnd cell_6t
Xbit_r24_c113 bl_113 br_113 wl_24 vdd gnd cell_6t
Xbit_r25_c113 bl_113 br_113 wl_25 vdd gnd cell_6t
Xbit_r26_c113 bl_113 br_113 wl_26 vdd gnd cell_6t
Xbit_r27_c113 bl_113 br_113 wl_27 vdd gnd cell_6t
Xbit_r28_c113 bl_113 br_113 wl_28 vdd gnd cell_6t
Xbit_r29_c113 bl_113 br_113 wl_29 vdd gnd cell_6t
Xbit_r30_c113 bl_113 br_113 wl_30 vdd gnd cell_6t
Xbit_r31_c113 bl_113 br_113 wl_31 vdd gnd cell_6t
Xbit_r32_c113 bl_113 br_113 wl_32 vdd gnd cell_6t
Xbit_r33_c113 bl_113 br_113 wl_33 vdd gnd cell_6t
Xbit_r34_c113 bl_113 br_113 wl_34 vdd gnd cell_6t
Xbit_r35_c113 bl_113 br_113 wl_35 vdd gnd cell_6t
Xbit_r36_c113 bl_113 br_113 wl_36 vdd gnd cell_6t
Xbit_r37_c113 bl_113 br_113 wl_37 vdd gnd cell_6t
Xbit_r38_c113 bl_113 br_113 wl_38 vdd gnd cell_6t
Xbit_r39_c113 bl_113 br_113 wl_39 vdd gnd cell_6t
Xbit_r40_c113 bl_113 br_113 wl_40 vdd gnd cell_6t
Xbit_r41_c113 bl_113 br_113 wl_41 vdd gnd cell_6t
Xbit_r42_c113 bl_113 br_113 wl_42 vdd gnd cell_6t
Xbit_r43_c113 bl_113 br_113 wl_43 vdd gnd cell_6t
Xbit_r44_c113 bl_113 br_113 wl_44 vdd gnd cell_6t
Xbit_r45_c113 bl_113 br_113 wl_45 vdd gnd cell_6t
Xbit_r46_c113 bl_113 br_113 wl_46 vdd gnd cell_6t
Xbit_r47_c113 bl_113 br_113 wl_47 vdd gnd cell_6t
Xbit_r48_c113 bl_113 br_113 wl_48 vdd gnd cell_6t
Xbit_r49_c113 bl_113 br_113 wl_49 vdd gnd cell_6t
Xbit_r50_c113 bl_113 br_113 wl_50 vdd gnd cell_6t
Xbit_r51_c113 bl_113 br_113 wl_51 vdd gnd cell_6t
Xbit_r52_c113 bl_113 br_113 wl_52 vdd gnd cell_6t
Xbit_r53_c113 bl_113 br_113 wl_53 vdd gnd cell_6t
Xbit_r54_c113 bl_113 br_113 wl_54 vdd gnd cell_6t
Xbit_r55_c113 bl_113 br_113 wl_55 vdd gnd cell_6t
Xbit_r56_c113 bl_113 br_113 wl_56 vdd gnd cell_6t
Xbit_r57_c113 bl_113 br_113 wl_57 vdd gnd cell_6t
Xbit_r58_c113 bl_113 br_113 wl_58 vdd gnd cell_6t
Xbit_r59_c113 bl_113 br_113 wl_59 vdd gnd cell_6t
Xbit_r60_c113 bl_113 br_113 wl_60 vdd gnd cell_6t
Xbit_r61_c113 bl_113 br_113 wl_61 vdd gnd cell_6t
Xbit_r62_c113 bl_113 br_113 wl_62 vdd gnd cell_6t
Xbit_r63_c113 bl_113 br_113 wl_63 vdd gnd cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd cell_6t
Xbit_r1_c114 bl_114 br_114 wl_1 vdd gnd cell_6t
Xbit_r2_c114 bl_114 br_114 wl_2 vdd gnd cell_6t
Xbit_r3_c114 bl_114 br_114 wl_3 vdd gnd cell_6t
Xbit_r4_c114 bl_114 br_114 wl_4 vdd gnd cell_6t
Xbit_r5_c114 bl_114 br_114 wl_5 vdd gnd cell_6t
Xbit_r6_c114 bl_114 br_114 wl_6 vdd gnd cell_6t
Xbit_r7_c114 bl_114 br_114 wl_7 vdd gnd cell_6t
Xbit_r8_c114 bl_114 br_114 wl_8 vdd gnd cell_6t
Xbit_r9_c114 bl_114 br_114 wl_9 vdd gnd cell_6t
Xbit_r10_c114 bl_114 br_114 wl_10 vdd gnd cell_6t
Xbit_r11_c114 bl_114 br_114 wl_11 vdd gnd cell_6t
Xbit_r12_c114 bl_114 br_114 wl_12 vdd gnd cell_6t
Xbit_r13_c114 bl_114 br_114 wl_13 vdd gnd cell_6t
Xbit_r14_c114 bl_114 br_114 wl_14 vdd gnd cell_6t
Xbit_r15_c114 bl_114 br_114 wl_15 vdd gnd cell_6t
Xbit_r16_c114 bl_114 br_114 wl_16 vdd gnd cell_6t
Xbit_r17_c114 bl_114 br_114 wl_17 vdd gnd cell_6t
Xbit_r18_c114 bl_114 br_114 wl_18 vdd gnd cell_6t
Xbit_r19_c114 bl_114 br_114 wl_19 vdd gnd cell_6t
Xbit_r20_c114 bl_114 br_114 wl_20 vdd gnd cell_6t
Xbit_r21_c114 bl_114 br_114 wl_21 vdd gnd cell_6t
Xbit_r22_c114 bl_114 br_114 wl_22 vdd gnd cell_6t
Xbit_r23_c114 bl_114 br_114 wl_23 vdd gnd cell_6t
Xbit_r24_c114 bl_114 br_114 wl_24 vdd gnd cell_6t
Xbit_r25_c114 bl_114 br_114 wl_25 vdd gnd cell_6t
Xbit_r26_c114 bl_114 br_114 wl_26 vdd gnd cell_6t
Xbit_r27_c114 bl_114 br_114 wl_27 vdd gnd cell_6t
Xbit_r28_c114 bl_114 br_114 wl_28 vdd gnd cell_6t
Xbit_r29_c114 bl_114 br_114 wl_29 vdd gnd cell_6t
Xbit_r30_c114 bl_114 br_114 wl_30 vdd gnd cell_6t
Xbit_r31_c114 bl_114 br_114 wl_31 vdd gnd cell_6t
Xbit_r32_c114 bl_114 br_114 wl_32 vdd gnd cell_6t
Xbit_r33_c114 bl_114 br_114 wl_33 vdd gnd cell_6t
Xbit_r34_c114 bl_114 br_114 wl_34 vdd gnd cell_6t
Xbit_r35_c114 bl_114 br_114 wl_35 vdd gnd cell_6t
Xbit_r36_c114 bl_114 br_114 wl_36 vdd gnd cell_6t
Xbit_r37_c114 bl_114 br_114 wl_37 vdd gnd cell_6t
Xbit_r38_c114 bl_114 br_114 wl_38 vdd gnd cell_6t
Xbit_r39_c114 bl_114 br_114 wl_39 vdd gnd cell_6t
Xbit_r40_c114 bl_114 br_114 wl_40 vdd gnd cell_6t
Xbit_r41_c114 bl_114 br_114 wl_41 vdd gnd cell_6t
Xbit_r42_c114 bl_114 br_114 wl_42 vdd gnd cell_6t
Xbit_r43_c114 bl_114 br_114 wl_43 vdd gnd cell_6t
Xbit_r44_c114 bl_114 br_114 wl_44 vdd gnd cell_6t
Xbit_r45_c114 bl_114 br_114 wl_45 vdd gnd cell_6t
Xbit_r46_c114 bl_114 br_114 wl_46 vdd gnd cell_6t
Xbit_r47_c114 bl_114 br_114 wl_47 vdd gnd cell_6t
Xbit_r48_c114 bl_114 br_114 wl_48 vdd gnd cell_6t
Xbit_r49_c114 bl_114 br_114 wl_49 vdd gnd cell_6t
Xbit_r50_c114 bl_114 br_114 wl_50 vdd gnd cell_6t
Xbit_r51_c114 bl_114 br_114 wl_51 vdd gnd cell_6t
Xbit_r52_c114 bl_114 br_114 wl_52 vdd gnd cell_6t
Xbit_r53_c114 bl_114 br_114 wl_53 vdd gnd cell_6t
Xbit_r54_c114 bl_114 br_114 wl_54 vdd gnd cell_6t
Xbit_r55_c114 bl_114 br_114 wl_55 vdd gnd cell_6t
Xbit_r56_c114 bl_114 br_114 wl_56 vdd gnd cell_6t
Xbit_r57_c114 bl_114 br_114 wl_57 vdd gnd cell_6t
Xbit_r58_c114 bl_114 br_114 wl_58 vdd gnd cell_6t
Xbit_r59_c114 bl_114 br_114 wl_59 vdd gnd cell_6t
Xbit_r60_c114 bl_114 br_114 wl_60 vdd gnd cell_6t
Xbit_r61_c114 bl_114 br_114 wl_61 vdd gnd cell_6t
Xbit_r62_c114 bl_114 br_114 wl_62 vdd gnd cell_6t
Xbit_r63_c114 bl_114 br_114 wl_63 vdd gnd cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd cell_6t
Xbit_r1_c115 bl_115 br_115 wl_1 vdd gnd cell_6t
Xbit_r2_c115 bl_115 br_115 wl_2 vdd gnd cell_6t
Xbit_r3_c115 bl_115 br_115 wl_3 vdd gnd cell_6t
Xbit_r4_c115 bl_115 br_115 wl_4 vdd gnd cell_6t
Xbit_r5_c115 bl_115 br_115 wl_5 vdd gnd cell_6t
Xbit_r6_c115 bl_115 br_115 wl_6 vdd gnd cell_6t
Xbit_r7_c115 bl_115 br_115 wl_7 vdd gnd cell_6t
Xbit_r8_c115 bl_115 br_115 wl_8 vdd gnd cell_6t
Xbit_r9_c115 bl_115 br_115 wl_9 vdd gnd cell_6t
Xbit_r10_c115 bl_115 br_115 wl_10 vdd gnd cell_6t
Xbit_r11_c115 bl_115 br_115 wl_11 vdd gnd cell_6t
Xbit_r12_c115 bl_115 br_115 wl_12 vdd gnd cell_6t
Xbit_r13_c115 bl_115 br_115 wl_13 vdd gnd cell_6t
Xbit_r14_c115 bl_115 br_115 wl_14 vdd gnd cell_6t
Xbit_r15_c115 bl_115 br_115 wl_15 vdd gnd cell_6t
Xbit_r16_c115 bl_115 br_115 wl_16 vdd gnd cell_6t
Xbit_r17_c115 bl_115 br_115 wl_17 vdd gnd cell_6t
Xbit_r18_c115 bl_115 br_115 wl_18 vdd gnd cell_6t
Xbit_r19_c115 bl_115 br_115 wl_19 vdd gnd cell_6t
Xbit_r20_c115 bl_115 br_115 wl_20 vdd gnd cell_6t
Xbit_r21_c115 bl_115 br_115 wl_21 vdd gnd cell_6t
Xbit_r22_c115 bl_115 br_115 wl_22 vdd gnd cell_6t
Xbit_r23_c115 bl_115 br_115 wl_23 vdd gnd cell_6t
Xbit_r24_c115 bl_115 br_115 wl_24 vdd gnd cell_6t
Xbit_r25_c115 bl_115 br_115 wl_25 vdd gnd cell_6t
Xbit_r26_c115 bl_115 br_115 wl_26 vdd gnd cell_6t
Xbit_r27_c115 bl_115 br_115 wl_27 vdd gnd cell_6t
Xbit_r28_c115 bl_115 br_115 wl_28 vdd gnd cell_6t
Xbit_r29_c115 bl_115 br_115 wl_29 vdd gnd cell_6t
Xbit_r30_c115 bl_115 br_115 wl_30 vdd gnd cell_6t
Xbit_r31_c115 bl_115 br_115 wl_31 vdd gnd cell_6t
Xbit_r32_c115 bl_115 br_115 wl_32 vdd gnd cell_6t
Xbit_r33_c115 bl_115 br_115 wl_33 vdd gnd cell_6t
Xbit_r34_c115 bl_115 br_115 wl_34 vdd gnd cell_6t
Xbit_r35_c115 bl_115 br_115 wl_35 vdd gnd cell_6t
Xbit_r36_c115 bl_115 br_115 wl_36 vdd gnd cell_6t
Xbit_r37_c115 bl_115 br_115 wl_37 vdd gnd cell_6t
Xbit_r38_c115 bl_115 br_115 wl_38 vdd gnd cell_6t
Xbit_r39_c115 bl_115 br_115 wl_39 vdd gnd cell_6t
Xbit_r40_c115 bl_115 br_115 wl_40 vdd gnd cell_6t
Xbit_r41_c115 bl_115 br_115 wl_41 vdd gnd cell_6t
Xbit_r42_c115 bl_115 br_115 wl_42 vdd gnd cell_6t
Xbit_r43_c115 bl_115 br_115 wl_43 vdd gnd cell_6t
Xbit_r44_c115 bl_115 br_115 wl_44 vdd gnd cell_6t
Xbit_r45_c115 bl_115 br_115 wl_45 vdd gnd cell_6t
Xbit_r46_c115 bl_115 br_115 wl_46 vdd gnd cell_6t
Xbit_r47_c115 bl_115 br_115 wl_47 vdd gnd cell_6t
Xbit_r48_c115 bl_115 br_115 wl_48 vdd gnd cell_6t
Xbit_r49_c115 bl_115 br_115 wl_49 vdd gnd cell_6t
Xbit_r50_c115 bl_115 br_115 wl_50 vdd gnd cell_6t
Xbit_r51_c115 bl_115 br_115 wl_51 vdd gnd cell_6t
Xbit_r52_c115 bl_115 br_115 wl_52 vdd gnd cell_6t
Xbit_r53_c115 bl_115 br_115 wl_53 vdd gnd cell_6t
Xbit_r54_c115 bl_115 br_115 wl_54 vdd gnd cell_6t
Xbit_r55_c115 bl_115 br_115 wl_55 vdd gnd cell_6t
Xbit_r56_c115 bl_115 br_115 wl_56 vdd gnd cell_6t
Xbit_r57_c115 bl_115 br_115 wl_57 vdd gnd cell_6t
Xbit_r58_c115 bl_115 br_115 wl_58 vdd gnd cell_6t
Xbit_r59_c115 bl_115 br_115 wl_59 vdd gnd cell_6t
Xbit_r60_c115 bl_115 br_115 wl_60 vdd gnd cell_6t
Xbit_r61_c115 bl_115 br_115 wl_61 vdd gnd cell_6t
Xbit_r62_c115 bl_115 br_115 wl_62 vdd gnd cell_6t
Xbit_r63_c115 bl_115 br_115 wl_63 vdd gnd cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd cell_6t
Xbit_r1_c116 bl_116 br_116 wl_1 vdd gnd cell_6t
Xbit_r2_c116 bl_116 br_116 wl_2 vdd gnd cell_6t
Xbit_r3_c116 bl_116 br_116 wl_3 vdd gnd cell_6t
Xbit_r4_c116 bl_116 br_116 wl_4 vdd gnd cell_6t
Xbit_r5_c116 bl_116 br_116 wl_5 vdd gnd cell_6t
Xbit_r6_c116 bl_116 br_116 wl_6 vdd gnd cell_6t
Xbit_r7_c116 bl_116 br_116 wl_7 vdd gnd cell_6t
Xbit_r8_c116 bl_116 br_116 wl_8 vdd gnd cell_6t
Xbit_r9_c116 bl_116 br_116 wl_9 vdd gnd cell_6t
Xbit_r10_c116 bl_116 br_116 wl_10 vdd gnd cell_6t
Xbit_r11_c116 bl_116 br_116 wl_11 vdd gnd cell_6t
Xbit_r12_c116 bl_116 br_116 wl_12 vdd gnd cell_6t
Xbit_r13_c116 bl_116 br_116 wl_13 vdd gnd cell_6t
Xbit_r14_c116 bl_116 br_116 wl_14 vdd gnd cell_6t
Xbit_r15_c116 bl_116 br_116 wl_15 vdd gnd cell_6t
Xbit_r16_c116 bl_116 br_116 wl_16 vdd gnd cell_6t
Xbit_r17_c116 bl_116 br_116 wl_17 vdd gnd cell_6t
Xbit_r18_c116 bl_116 br_116 wl_18 vdd gnd cell_6t
Xbit_r19_c116 bl_116 br_116 wl_19 vdd gnd cell_6t
Xbit_r20_c116 bl_116 br_116 wl_20 vdd gnd cell_6t
Xbit_r21_c116 bl_116 br_116 wl_21 vdd gnd cell_6t
Xbit_r22_c116 bl_116 br_116 wl_22 vdd gnd cell_6t
Xbit_r23_c116 bl_116 br_116 wl_23 vdd gnd cell_6t
Xbit_r24_c116 bl_116 br_116 wl_24 vdd gnd cell_6t
Xbit_r25_c116 bl_116 br_116 wl_25 vdd gnd cell_6t
Xbit_r26_c116 bl_116 br_116 wl_26 vdd gnd cell_6t
Xbit_r27_c116 bl_116 br_116 wl_27 vdd gnd cell_6t
Xbit_r28_c116 bl_116 br_116 wl_28 vdd gnd cell_6t
Xbit_r29_c116 bl_116 br_116 wl_29 vdd gnd cell_6t
Xbit_r30_c116 bl_116 br_116 wl_30 vdd gnd cell_6t
Xbit_r31_c116 bl_116 br_116 wl_31 vdd gnd cell_6t
Xbit_r32_c116 bl_116 br_116 wl_32 vdd gnd cell_6t
Xbit_r33_c116 bl_116 br_116 wl_33 vdd gnd cell_6t
Xbit_r34_c116 bl_116 br_116 wl_34 vdd gnd cell_6t
Xbit_r35_c116 bl_116 br_116 wl_35 vdd gnd cell_6t
Xbit_r36_c116 bl_116 br_116 wl_36 vdd gnd cell_6t
Xbit_r37_c116 bl_116 br_116 wl_37 vdd gnd cell_6t
Xbit_r38_c116 bl_116 br_116 wl_38 vdd gnd cell_6t
Xbit_r39_c116 bl_116 br_116 wl_39 vdd gnd cell_6t
Xbit_r40_c116 bl_116 br_116 wl_40 vdd gnd cell_6t
Xbit_r41_c116 bl_116 br_116 wl_41 vdd gnd cell_6t
Xbit_r42_c116 bl_116 br_116 wl_42 vdd gnd cell_6t
Xbit_r43_c116 bl_116 br_116 wl_43 vdd gnd cell_6t
Xbit_r44_c116 bl_116 br_116 wl_44 vdd gnd cell_6t
Xbit_r45_c116 bl_116 br_116 wl_45 vdd gnd cell_6t
Xbit_r46_c116 bl_116 br_116 wl_46 vdd gnd cell_6t
Xbit_r47_c116 bl_116 br_116 wl_47 vdd gnd cell_6t
Xbit_r48_c116 bl_116 br_116 wl_48 vdd gnd cell_6t
Xbit_r49_c116 bl_116 br_116 wl_49 vdd gnd cell_6t
Xbit_r50_c116 bl_116 br_116 wl_50 vdd gnd cell_6t
Xbit_r51_c116 bl_116 br_116 wl_51 vdd gnd cell_6t
Xbit_r52_c116 bl_116 br_116 wl_52 vdd gnd cell_6t
Xbit_r53_c116 bl_116 br_116 wl_53 vdd gnd cell_6t
Xbit_r54_c116 bl_116 br_116 wl_54 vdd gnd cell_6t
Xbit_r55_c116 bl_116 br_116 wl_55 vdd gnd cell_6t
Xbit_r56_c116 bl_116 br_116 wl_56 vdd gnd cell_6t
Xbit_r57_c116 bl_116 br_116 wl_57 vdd gnd cell_6t
Xbit_r58_c116 bl_116 br_116 wl_58 vdd gnd cell_6t
Xbit_r59_c116 bl_116 br_116 wl_59 vdd gnd cell_6t
Xbit_r60_c116 bl_116 br_116 wl_60 vdd gnd cell_6t
Xbit_r61_c116 bl_116 br_116 wl_61 vdd gnd cell_6t
Xbit_r62_c116 bl_116 br_116 wl_62 vdd gnd cell_6t
Xbit_r63_c116 bl_116 br_116 wl_63 vdd gnd cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd cell_6t
Xbit_r1_c117 bl_117 br_117 wl_1 vdd gnd cell_6t
Xbit_r2_c117 bl_117 br_117 wl_2 vdd gnd cell_6t
Xbit_r3_c117 bl_117 br_117 wl_3 vdd gnd cell_6t
Xbit_r4_c117 bl_117 br_117 wl_4 vdd gnd cell_6t
Xbit_r5_c117 bl_117 br_117 wl_5 vdd gnd cell_6t
Xbit_r6_c117 bl_117 br_117 wl_6 vdd gnd cell_6t
Xbit_r7_c117 bl_117 br_117 wl_7 vdd gnd cell_6t
Xbit_r8_c117 bl_117 br_117 wl_8 vdd gnd cell_6t
Xbit_r9_c117 bl_117 br_117 wl_9 vdd gnd cell_6t
Xbit_r10_c117 bl_117 br_117 wl_10 vdd gnd cell_6t
Xbit_r11_c117 bl_117 br_117 wl_11 vdd gnd cell_6t
Xbit_r12_c117 bl_117 br_117 wl_12 vdd gnd cell_6t
Xbit_r13_c117 bl_117 br_117 wl_13 vdd gnd cell_6t
Xbit_r14_c117 bl_117 br_117 wl_14 vdd gnd cell_6t
Xbit_r15_c117 bl_117 br_117 wl_15 vdd gnd cell_6t
Xbit_r16_c117 bl_117 br_117 wl_16 vdd gnd cell_6t
Xbit_r17_c117 bl_117 br_117 wl_17 vdd gnd cell_6t
Xbit_r18_c117 bl_117 br_117 wl_18 vdd gnd cell_6t
Xbit_r19_c117 bl_117 br_117 wl_19 vdd gnd cell_6t
Xbit_r20_c117 bl_117 br_117 wl_20 vdd gnd cell_6t
Xbit_r21_c117 bl_117 br_117 wl_21 vdd gnd cell_6t
Xbit_r22_c117 bl_117 br_117 wl_22 vdd gnd cell_6t
Xbit_r23_c117 bl_117 br_117 wl_23 vdd gnd cell_6t
Xbit_r24_c117 bl_117 br_117 wl_24 vdd gnd cell_6t
Xbit_r25_c117 bl_117 br_117 wl_25 vdd gnd cell_6t
Xbit_r26_c117 bl_117 br_117 wl_26 vdd gnd cell_6t
Xbit_r27_c117 bl_117 br_117 wl_27 vdd gnd cell_6t
Xbit_r28_c117 bl_117 br_117 wl_28 vdd gnd cell_6t
Xbit_r29_c117 bl_117 br_117 wl_29 vdd gnd cell_6t
Xbit_r30_c117 bl_117 br_117 wl_30 vdd gnd cell_6t
Xbit_r31_c117 bl_117 br_117 wl_31 vdd gnd cell_6t
Xbit_r32_c117 bl_117 br_117 wl_32 vdd gnd cell_6t
Xbit_r33_c117 bl_117 br_117 wl_33 vdd gnd cell_6t
Xbit_r34_c117 bl_117 br_117 wl_34 vdd gnd cell_6t
Xbit_r35_c117 bl_117 br_117 wl_35 vdd gnd cell_6t
Xbit_r36_c117 bl_117 br_117 wl_36 vdd gnd cell_6t
Xbit_r37_c117 bl_117 br_117 wl_37 vdd gnd cell_6t
Xbit_r38_c117 bl_117 br_117 wl_38 vdd gnd cell_6t
Xbit_r39_c117 bl_117 br_117 wl_39 vdd gnd cell_6t
Xbit_r40_c117 bl_117 br_117 wl_40 vdd gnd cell_6t
Xbit_r41_c117 bl_117 br_117 wl_41 vdd gnd cell_6t
Xbit_r42_c117 bl_117 br_117 wl_42 vdd gnd cell_6t
Xbit_r43_c117 bl_117 br_117 wl_43 vdd gnd cell_6t
Xbit_r44_c117 bl_117 br_117 wl_44 vdd gnd cell_6t
Xbit_r45_c117 bl_117 br_117 wl_45 vdd gnd cell_6t
Xbit_r46_c117 bl_117 br_117 wl_46 vdd gnd cell_6t
Xbit_r47_c117 bl_117 br_117 wl_47 vdd gnd cell_6t
Xbit_r48_c117 bl_117 br_117 wl_48 vdd gnd cell_6t
Xbit_r49_c117 bl_117 br_117 wl_49 vdd gnd cell_6t
Xbit_r50_c117 bl_117 br_117 wl_50 vdd gnd cell_6t
Xbit_r51_c117 bl_117 br_117 wl_51 vdd gnd cell_6t
Xbit_r52_c117 bl_117 br_117 wl_52 vdd gnd cell_6t
Xbit_r53_c117 bl_117 br_117 wl_53 vdd gnd cell_6t
Xbit_r54_c117 bl_117 br_117 wl_54 vdd gnd cell_6t
Xbit_r55_c117 bl_117 br_117 wl_55 vdd gnd cell_6t
Xbit_r56_c117 bl_117 br_117 wl_56 vdd gnd cell_6t
Xbit_r57_c117 bl_117 br_117 wl_57 vdd gnd cell_6t
Xbit_r58_c117 bl_117 br_117 wl_58 vdd gnd cell_6t
Xbit_r59_c117 bl_117 br_117 wl_59 vdd gnd cell_6t
Xbit_r60_c117 bl_117 br_117 wl_60 vdd gnd cell_6t
Xbit_r61_c117 bl_117 br_117 wl_61 vdd gnd cell_6t
Xbit_r62_c117 bl_117 br_117 wl_62 vdd gnd cell_6t
Xbit_r63_c117 bl_117 br_117 wl_63 vdd gnd cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd cell_6t
Xbit_r1_c118 bl_118 br_118 wl_1 vdd gnd cell_6t
Xbit_r2_c118 bl_118 br_118 wl_2 vdd gnd cell_6t
Xbit_r3_c118 bl_118 br_118 wl_3 vdd gnd cell_6t
Xbit_r4_c118 bl_118 br_118 wl_4 vdd gnd cell_6t
Xbit_r5_c118 bl_118 br_118 wl_5 vdd gnd cell_6t
Xbit_r6_c118 bl_118 br_118 wl_6 vdd gnd cell_6t
Xbit_r7_c118 bl_118 br_118 wl_7 vdd gnd cell_6t
Xbit_r8_c118 bl_118 br_118 wl_8 vdd gnd cell_6t
Xbit_r9_c118 bl_118 br_118 wl_9 vdd gnd cell_6t
Xbit_r10_c118 bl_118 br_118 wl_10 vdd gnd cell_6t
Xbit_r11_c118 bl_118 br_118 wl_11 vdd gnd cell_6t
Xbit_r12_c118 bl_118 br_118 wl_12 vdd gnd cell_6t
Xbit_r13_c118 bl_118 br_118 wl_13 vdd gnd cell_6t
Xbit_r14_c118 bl_118 br_118 wl_14 vdd gnd cell_6t
Xbit_r15_c118 bl_118 br_118 wl_15 vdd gnd cell_6t
Xbit_r16_c118 bl_118 br_118 wl_16 vdd gnd cell_6t
Xbit_r17_c118 bl_118 br_118 wl_17 vdd gnd cell_6t
Xbit_r18_c118 bl_118 br_118 wl_18 vdd gnd cell_6t
Xbit_r19_c118 bl_118 br_118 wl_19 vdd gnd cell_6t
Xbit_r20_c118 bl_118 br_118 wl_20 vdd gnd cell_6t
Xbit_r21_c118 bl_118 br_118 wl_21 vdd gnd cell_6t
Xbit_r22_c118 bl_118 br_118 wl_22 vdd gnd cell_6t
Xbit_r23_c118 bl_118 br_118 wl_23 vdd gnd cell_6t
Xbit_r24_c118 bl_118 br_118 wl_24 vdd gnd cell_6t
Xbit_r25_c118 bl_118 br_118 wl_25 vdd gnd cell_6t
Xbit_r26_c118 bl_118 br_118 wl_26 vdd gnd cell_6t
Xbit_r27_c118 bl_118 br_118 wl_27 vdd gnd cell_6t
Xbit_r28_c118 bl_118 br_118 wl_28 vdd gnd cell_6t
Xbit_r29_c118 bl_118 br_118 wl_29 vdd gnd cell_6t
Xbit_r30_c118 bl_118 br_118 wl_30 vdd gnd cell_6t
Xbit_r31_c118 bl_118 br_118 wl_31 vdd gnd cell_6t
Xbit_r32_c118 bl_118 br_118 wl_32 vdd gnd cell_6t
Xbit_r33_c118 bl_118 br_118 wl_33 vdd gnd cell_6t
Xbit_r34_c118 bl_118 br_118 wl_34 vdd gnd cell_6t
Xbit_r35_c118 bl_118 br_118 wl_35 vdd gnd cell_6t
Xbit_r36_c118 bl_118 br_118 wl_36 vdd gnd cell_6t
Xbit_r37_c118 bl_118 br_118 wl_37 vdd gnd cell_6t
Xbit_r38_c118 bl_118 br_118 wl_38 vdd gnd cell_6t
Xbit_r39_c118 bl_118 br_118 wl_39 vdd gnd cell_6t
Xbit_r40_c118 bl_118 br_118 wl_40 vdd gnd cell_6t
Xbit_r41_c118 bl_118 br_118 wl_41 vdd gnd cell_6t
Xbit_r42_c118 bl_118 br_118 wl_42 vdd gnd cell_6t
Xbit_r43_c118 bl_118 br_118 wl_43 vdd gnd cell_6t
Xbit_r44_c118 bl_118 br_118 wl_44 vdd gnd cell_6t
Xbit_r45_c118 bl_118 br_118 wl_45 vdd gnd cell_6t
Xbit_r46_c118 bl_118 br_118 wl_46 vdd gnd cell_6t
Xbit_r47_c118 bl_118 br_118 wl_47 vdd gnd cell_6t
Xbit_r48_c118 bl_118 br_118 wl_48 vdd gnd cell_6t
Xbit_r49_c118 bl_118 br_118 wl_49 vdd gnd cell_6t
Xbit_r50_c118 bl_118 br_118 wl_50 vdd gnd cell_6t
Xbit_r51_c118 bl_118 br_118 wl_51 vdd gnd cell_6t
Xbit_r52_c118 bl_118 br_118 wl_52 vdd gnd cell_6t
Xbit_r53_c118 bl_118 br_118 wl_53 vdd gnd cell_6t
Xbit_r54_c118 bl_118 br_118 wl_54 vdd gnd cell_6t
Xbit_r55_c118 bl_118 br_118 wl_55 vdd gnd cell_6t
Xbit_r56_c118 bl_118 br_118 wl_56 vdd gnd cell_6t
Xbit_r57_c118 bl_118 br_118 wl_57 vdd gnd cell_6t
Xbit_r58_c118 bl_118 br_118 wl_58 vdd gnd cell_6t
Xbit_r59_c118 bl_118 br_118 wl_59 vdd gnd cell_6t
Xbit_r60_c118 bl_118 br_118 wl_60 vdd gnd cell_6t
Xbit_r61_c118 bl_118 br_118 wl_61 vdd gnd cell_6t
Xbit_r62_c118 bl_118 br_118 wl_62 vdd gnd cell_6t
Xbit_r63_c118 bl_118 br_118 wl_63 vdd gnd cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd cell_6t
Xbit_r1_c119 bl_119 br_119 wl_1 vdd gnd cell_6t
Xbit_r2_c119 bl_119 br_119 wl_2 vdd gnd cell_6t
Xbit_r3_c119 bl_119 br_119 wl_3 vdd gnd cell_6t
Xbit_r4_c119 bl_119 br_119 wl_4 vdd gnd cell_6t
Xbit_r5_c119 bl_119 br_119 wl_5 vdd gnd cell_6t
Xbit_r6_c119 bl_119 br_119 wl_6 vdd gnd cell_6t
Xbit_r7_c119 bl_119 br_119 wl_7 vdd gnd cell_6t
Xbit_r8_c119 bl_119 br_119 wl_8 vdd gnd cell_6t
Xbit_r9_c119 bl_119 br_119 wl_9 vdd gnd cell_6t
Xbit_r10_c119 bl_119 br_119 wl_10 vdd gnd cell_6t
Xbit_r11_c119 bl_119 br_119 wl_11 vdd gnd cell_6t
Xbit_r12_c119 bl_119 br_119 wl_12 vdd gnd cell_6t
Xbit_r13_c119 bl_119 br_119 wl_13 vdd gnd cell_6t
Xbit_r14_c119 bl_119 br_119 wl_14 vdd gnd cell_6t
Xbit_r15_c119 bl_119 br_119 wl_15 vdd gnd cell_6t
Xbit_r16_c119 bl_119 br_119 wl_16 vdd gnd cell_6t
Xbit_r17_c119 bl_119 br_119 wl_17 vdd gnd cell_6t
Xbit_r18_c119 bl_119 br_119 wl_18 vdd gnd cell_6t
Xbit_r19_c119 bl_119 br_119 wl_19 vdd gnd cell_6t
Xbit_r20_c119 bl_119 br_119 wl_20 vdd gnd cell_6t
Xbit_r21_c119 bl_119 br_119 wl_21 vdd gnd cell_6t
Xbit_r22_c119 bl_119 br_119 wl_22 vdd gnd cell_6t
Xbit_r23_c119 bl_119 br_119 wl_23 vdd gnd cell_6t
Xbit_r24_c119 bl_119 br_119 wl_24 vdd gnd cell_6t
Xbit_r25_c119 bl_119 br_119 wl_25 vdd gnd cell_6t
Xbit_r26_c119 bl_119 br_119 wl_26 vdd gnd cell_6t
Xbit_r27_c119 bl_119 br_119 wl_27 vdd gnd cell_6t
Xbit_r28_c119 bl_119 br_119 wl_28 vdd gnd cell_6t
Xbit_r29_c119 bl_119 br_119 wl_29 vdd gnd cell_6t
Xbit_r30_c119 bl_119 br_119 wl_30 vdd gnd cell_6t
Xbit_r31_c119 bl_119 br_119 wl_31 vdd gnd cell_6t
Xbit_r32_c119 bl_119 br_119 wl_32 vdd gnd cell_6t
Xbit_r33_c119 bl_119 br_119 wl_33 vdd gnd cell_6t
Xbit_r34_c119 bl_119 br_119 wl_34 vdd gnd cell_6t
Xbit_r35_c119 bl_119 br_119 wl_35 vdd gnd cell_6t
Xbit_r36_c119 bl_119 br_119 wl_36 vdd gnd cell_6t
Xbit_r37_c119 bl_119 br_119 wl_37 vdd gnd cell_6t
Xbit_r38_c119 bl_119 br_119 wl_38 vdd gnd cell_6t
Xbit_r39_c119 bl_119 br_119 wl_39 vdd gnd cell_6t
Xbit_r40_c119 bl_119 br_119 wl_40 vdd gnd cell_6t
Xbit_r41_c119 bl_119 br_119 wl_41 vdd gnd cell_6t
Xbit_r42_c119 bl_119 br_119 wl_42 vdd gnd cell_6t
Xbit_r43_c119 bl_119 br_119 wl_43 vdd gnd cell_6t
Xbit_r44_c119 bl_119 br_119 wl_44 vdd gnd cell_6t
Xbit_r45_c119 bl_119 br_119 wl_45 vdd gnd cell_6t
Xbit_r46_c119 bl_119 br_119 wl_46 vdd gnd cell_6t
Xbit_r47_c119 bl_119 br_119 wl_47 vdd gnd cell_6t
Xbit_r48_c119 bl_119 br_119 wl_48 vdd gnd cell_6t
Xbit_r49_c119 bl_119 br_119 wl_49 vdd gnd cell_6t
Xbit_r50_c119 bl_119 br_119 wl_50 vdd gnd cell_6t
Xbit_r51_c119 bl_119 br_119 wl_51 vdd gnd cell_6t
Xbit_r52_c119 bl_119 br_119 wl_52 vdd gnd cell_6t
Xbit_r53_c119 bl_119 br_119 wl_53 vdd gnd cell_6t
Xbit_r54_c119 bl_119 br_119 wl_54 vdd gnd cell_6t
Xbit_r55_c119 bl_119 br_119 wl_55 vdd gnd cell_6t
Xbit_r56_c119 bl_119 br_119 wl_56 vdd gnd cell_6t
Xbit_r57_c119 bl_119 br_119 wl_57 vdd gnd cell_6t
Xbit_r58_c119 bl_119 br_119 wl_58 vdd gnd cell_6t
Xbit_r59_c119 bl_119 br_119 wl_59 vdd gnd cell_6t
Xbit_r60_c119 bl_119 br_119 wl_60 vdd gnd cell_6t
Xbit_r61_c119 bl_119 br_119 wl_61 vdd gnd cell_6t
Xbit_r62_c119 bl_119 br_119 wl_62 vdd gnd cell_6t
Xbit_r63_c119 bl_119 br_119 wl_63 vdd gnd cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd cell_6t
Xbit_r1_c120 bl_120 br_120 wl_1 vdd gnd cell_6t
Xbit_r2_c120 bl_120 br_120 wl_2 vdd gnd cell_6t
Xbit_r3_c120 bl_120 br_120 wl_3 vdd gnd cell_6t
Xbit_r4_c120 bl_120 br_120 wl_4 vdd gnd cell_6t
Xbit_r5_c120 bl_120 br_120 wl_5 vdd gnd cell_6t
Xbit_r6_c120 bl_120 br_120 wl_6 vdd gnd cell_6t
Xbit_r7_c120 bl_120 br_120 wl_7 vdd gnd cell_6t
Xbit_r8_c120 bl_120 br_120 wl_8 vdd gnd cell_6t
Xbit_r9_c120 bl_120 br_120 wl_9 vdd gnd cell_6t
Xbit_r10_c120 bl_120 br_120 wl_10 vdd gnd cell_6t
Xbit_r11_c120 bl_120 br_120 wl_11 vdd gnd cell_6t
Xbit_r12_c120 bl_120 br_120 wl_12 vdd gnd cell_6t
Xbit_r13_c120 bl_120 br_120 wl_13 vdd gnd cell_6t
Xbit_r14_c120 bl_120 br_120 wl_14 vdd gnd cell_6t
Xbit_r15_c120 bl_120 br_120 wl_15 vdd gnd cell_6t
Xbit_r16_c120 bl_120 br_120 wl_16 vdd gnd cell_6t
Xbit_r17_c120 bl_120 br_120 wl_17 vdd gnd cell_6t
Xbit_r18_c120 bl_120 br_120 wl_18 vdd gnd cell_6t
Xbit_r19_c120 bl_120 br_120 wl_19 vdd gnd cell_6t
Xbit_r20_c120 bl_120 br_120 wl_20 vdd gnd cell_6t
Xbit_r21_c120 bl_120 br_120 wl_21 vdd gnd cell_6t
Xbit_r22_c120 bl_120 br_120 wl_22 vdd gnd cell_6t
Xbit_r23_c120 bl_120 br_120 wl_23 vdd gnd cell_6t
Xbit_r24_c120 bl_120 br_120 wl_24 vdd gnd cell_6t
Xbit_r25_c120 bl_120 br_120 wl_25 vdd gnd cell_6t
Xbit_r26_c120 bl_120 br_120 wl_26 vdd gnd cell_6t
Xbit_r27_c120 bl_120 br_120 wl_27 vdd gnd cell_6t
Xbit_r28_c120 bl_120 br_120 wl_28 vdd gnd cell_6t
Xbit_r29_c120 bl_120 br_120 wl_29 vdd gnd cell_6t
Xbit_r30_c120 bl_120 br_120 wl_30 vdd gnd cell_6t
Xbit_r31_c120 bl_120 br_120 wl_31 vdd gnd cell_6t
Xbit_r32_c120 bl_120 br_120 wl_32 vdd gnd cell_6t
Xbit_r33_c120 bl_120 br_120 wl_33 vdd gnd cell_6t
Xbit_r34_c120 bl_120 br_120 wl_34 vdd gnd cell_6t
Xbit_r35_c120 bl_120 br_120 wl_35 vdd gnd cell_6t
Xbit_r36_c120 bl_120 br_120 wl_36 vdd gnd cell_6t
Xbit_r37_c120 bl_120 br_120 wl_37 vdd gnd cell_6t
Xbit_r38_c120 bl_120 br_120 wl_38 vdd gnd cell_6t
Xbit_r39_c120 bl_120 br_120 wl_39 vdd gnd cell_6t
Xbit_r40_c120 bl_120 br_120 wl_40 vdd gnd cell_6t
Xbit_r41_c120 bl_120 br_120 wl_41 vdd gnd cell_6t
Xbit_r42_c120 bl_120 br_120 wl_42 vdd gnd cell_6t
Xbit_r43_c120 bl_120 br_120 wl_43 vdd gnd cell_6t
Xbit_r44_c120 bl_120 br_120 wl_44 vdd gnd cell_6t
Xbit_r45_c120 bl_120 br_120 wl_45 vdd gnd cell_6t
Xbit_r46_c120 bl_120 br_120 wl_46 vdd gnd cell_6t
Xbit_r47_c120 bl_120 br_120 wl_47 vdd gnd cell_6t
Xbit_r48_c120 bl_120 br_120 wl_48 vdd gnd cell_6t
Xbit_r49_c120 bl_120 br_120 wl_49 vdd gnd cell_6t
Xbit_r50_c120 bl_120 br_120 wl_50 vdd gnd cell_6t
Xbit_r51_c120 bl_120 br_120 wl_51 vdd gnd cell_6t
Xbit_r52_c120 bl_120 br_120 wl_52 vdd gnd cell_6t
Xbit_r53_c120 bl_120 br_120 wl_53 vdd gnd cell_6t
Xbit_r54_c120 bl_120 br_120 wl_54 vdd gnd cell_6t
Xbit_r55_c120 bl_120 br_120 wl_55 vdd gnd cell_6t
Xbit_r56_c120 bl_120 br_120 wl_56 vdd gnd cell_6t
Xbit_r57_c120 bl_120 br_120 wl_57 vdd gnd cell_6t
Xbit_r58_c120 bl_120 br_120 wl_58 vdd gnd cell_6t
Xbit_r59_c120 bl_120 br_120 wl_59 vdd gnd cell_6t
Xbit_r60_c120 bl_120 br_120 wl_60 vdd gnd cell_6t
Xbit_r61_c120 bl_120 br_120 wl_61 vdd gnd cell_6t
Xbit_r62_c120 bl_120 br_120 wl_62 vdd gnd cell_6t
Xbit_r63_c120 bl_120 br_120 wl_63 vdd gnd cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd cell_6t
Xbit_r1_c121 bl_121 br_121 wl_1 vdd gnd cell_6t
Xbit_r2_c121 bl_121 br_121 wl_2 vdd gnd cell_6t
Xbit_r3_c121 bl_121 br_121 wl_3 vdd gnd cell_6t
Xbit_r4_c121 bl_121 br_121 wl_4 vdd gnd cell_6t
Xbit_r5_c121 bl_121 br_121 wl_5 vdd gnd cell_6t
Xbit_r6_c121 bl_121 br_121 wl_6 vdd gnd cell_6t
Xbit_r7_c121 bl_121 br_121 wl_7 vdd gnd cell_6t
Xbit_r8_c121 bl_121 br_121 wl_8 vdd gnd cell_6t
Xbit_r9_c121 bl_121 br_121 wl_9 vdd gnd cell_6t
Xbit_r10_c121 bl_121 br_121 wl_10 vdd gnd cell_6t
Xbit_r11_c121 bl_121 br_121 wl_11 vdd gnd cell_6t
Xbit_r12_c121 bl_121 br_121 wl_12 vdd gnd cell_6t
Xbit_r13_c121 bl_121 br_121 wl_13 vdd gnd cell_6t
Xbit_r14_c121 bl_121 br_121 wl_14 vdd gnd cell_6t
Xbit_r15_c121 bl_121 br_121 wl_15 vdd gnd cell_6t
Xbit_r16_c121 bl_121 br_121 wl_16 vdd gnd cell_6t
Xbit_r17_c121 bl_121 br_121 wl_17 vdd gnd cell_6t
Xbit_r18_c121 bl_121 br_121 wl_18 vdd gnd cell_6t
Xbit_r19_c121 bl_121 br_121 wl_19 vdd gnd cell_6t
Xbit_r20_c121 bl_121 br_121 wl_20 vdd gnd cell_6t
Xbit_r21_c121 bl_121 br_121 wl_21 vdd gnd cell_6t
Xbit_r22_c121 bl_121 br_121 wl_22 vdd gnd cell_6t
Xbit_r23_c121 bl_121 br_121 wl_23 vdd gnd cell_6t
Xbit_r24_c121 bl_121 br_121 wl_24 vdd gnd cell_6t
Xbit_r25_c121 bl_121 br_121 wl_25 vdd gnd cell_6t
Xbit_r26_c121 bl_121 br_121 wl_26 vdd gnd cell_6t
Xbit_r27_c121 bl_121 br_121 wl_27 vdd gnd cell_6t
Xbit_r28_c121 bl_121 br_121 wl_28 vdd gnd cell_6t
Xbit_r29_c121 bl_121 br_121 wl_29 vdd gnd cell_6t
Xbit_r30_c121 bl_121 br_121 wl_30 vdd gnd cell_6t
Xbit_r31_c121 bl_121 br_121 wl_31 vdd gnd cell_6t
Xbit_r32_c121 bl_121 br_121 wl_32 vdd gnd cell_6t
Xbit_r33_c121 bl_121 br_121 wl_33 vdd gnd cell_6t
Xbit_r34_c121 bl_121 br_121 wl_34 vdd gnd cell_6t
Xbit_r35_c121 bl_121 br_121 wl_35 vdd gnd cell_6t
Xbit_r36_c121 bl_121 br_121 wl_36 vdd gnd cell_6t
Xbit_r37_c121 bl_121 br_121 wl_37 vdd gnd cell_6t
Xbit_r38_c121 bl_121 br_121 wl_38 vdd gnd cell_6t
Xbit_r39_c121 bl_121 br_121 wl_39 vdd gnd cell_6t
Xbit_r40_c121 bl_121 br_121 wl_40 vdd gnd cell_6t
Xbit_r41_c121 bl_121 br_121 wl_41 vdd gnd cell_6t
Xbit_r42_c121 bl_121 br_121 wl_42 vdd gnd cell_6t
Xbit_r43_c121 bl_121 br_121 wl_43 vdd gnd cell_6t
Xbit_r44_c121 bl_121 br_121 wl_44 vdd gnd cell_6t
Xbit_r45_c121 bl_121 br_121 wl_45 vdd gnd cell_6t
Xbit_r46_c121 bl_121 br_121 wl_46 vdd gnd cell_6t
Xbit_r47_c121 bl_121 br_121 wl_47 vdd gnd cell_6t
Xbit_r48_c121 bl_121 br_121 wl_48 vdd gnd cell_6t
Xbit_r49_c121 bl_121 br_121 wl_49 vdd gnd cell_6t
Xbit_r50_c121 bl_121 br_121 wl_50 vdd gnd cell_6t
Xbit_r51_c121 bl_121 br_121 wl_51 vdd gnd cell_6t
Xbit_r52_c121 bl_121 br_121 wl_52 vdd gnd cell_6t
Xbit_r53_c121 bl_121 br_121 wl_53 vdd gnd cell_6t
Xbit_r54_c121 bl_121 br_121 wl_54 vdd gnd cell_6t
Xbit_r55_c121 bl_121 br_121 wl_55 vdd gnd cell_6t
Xbit_r56_c121 bl_121 br_121 wl_56 vdd gnd cell_6t
Xbit_r57_c121 bl_121 br_121 wl_57 vdd gnd cell_6t
Xbit_r58_c121 bl_121 br_121 wl_58 vdd gnd cell_6t
Xbit_r59_c121 bl_121 br_121 wl_59 vdd gnd cell_6t
Xbit_r60_c121 bl_121 br_121 wl_60 vdd gnd cell_6t
Xbit_r61_c121 bl_121 br_121 wl_61 vdd gnd cell_6t
Xbit_r62_c121 bl_121 br_121 wl_62 vdd gnd cell_6t
Xbit_r63_c121 bl_121 br_121 wl_63 vdd gnd cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd cell_6t
Xbit_r1_c122 bl_122 br_122 wl_1 vdd gnd cell_6t
Xbit_r2_c122 bl_122 br_122 wl_2 vdd gnd cell_6t
Xbit_r3_c122 bl_122 br_122 wl_3 vdd gnd cell_6t
Xbit_r4_c122 bl_122 br_122 wl_4 vdd gnd cell_6t
Xbit_r5_c122 bl_122 br_122 wl_5 vdd gnd cell_6t
Xbit_r6_c122 bl_122 br_122 wl_6 vdd gnd cell_6t
Xbit_r7_c122 bl_122 br_122 wl_7 vdd gnd cell_6t
Xbit_r8_c122 bl_122 br_122 wl_8 vdd gnd cell_6t
Xbit_r9_c122 bl_122 br_122 wl_9 vdd gnd cell_6t
Xbit_r10_c122 bl_122 br_122 wl_10 vdd gnd cell_6t
Xbit_r11_c122 bl_122 br_122 wl_11 vdd gnd cell_6t
Xbit_r12_c122 bl_122 br_122 wl_12 vdd gnd cell_6t
Xbit_r13_c122 bl_122 br_122 wl_13 vdd gnd cell_6t
Xbit_r14_c122 bl_122 br_122 wl_14 vdd gnd cell_6t
Xbit_r15_c122 bl_122 br_122 wl_15 vdd gnd cell_6t
Xbit_r16_c122 bl_122 br_122 wl_16 vdd gnd cell_6t
Xbit_r17_c122 bl_122 br_122 wl_17 vdd gnd cell_6t
Xbit_r18_c122 bl_122 br_122 wl_18 vdd gnd cell_6t
Xbit_r19_c122 bl_122 br_122 wl_19 vdd gnd cell_6t
Xbit_r20_c122 bl_122 br_122 wl_20 vdd gnd cell_6t
Xbit_r21_c122 bl_122 br_122 wl_21 vdd gnd cell_6t
Xbit_r22_c122 bl_122 br_122 wl_22 vdd gnd cell_6t
Xbit_r23_c122 bl_122 br_122 wl_23 vdd gnd cell_6t
Xbit_r24_c122 bl_122 br_122 wl_24 vdd gnd cell_6t
Xbit_r25_c122 bl_122 br_122 wl_25 vdd gnd cell_6t
Xbit_r26_c122 bl_122 br_122 wl_26 vdd gnd cell_6t
Xbit_r27_c122 bl_122 br_122 wl_27 vdd gnd cell_6t
Xbit_r28_c122 bl_122 br_122 wl_28 vdd gnd cell_6t
Xbit_r29_c122 bl_122 br_122 wl_29 vdd gnd cell_6t
Xbit_r30_c122 bl_122 br_122 wl_30 vdd gnd cell_6t
Xbit_r31_c122 bl_122 br_122 wl_31 vdd gnd cell_6t
Xbit_r32_c122 bl_122 br_122 wl_32 vdd gnd cell_6t
Xbit_r33_c122 bl_122 br_122 wl_33 vdd gnd cell_6t
Xbit_r34_c122 bl_122 br_122 wl_34 vdd gnd cell_6t
Xbit_r35_c122 bl_122 br_122 wl_35 vdd gnd cell_6t
Xbit_r36_c122 bl_122 br_122 wl_36 vdd gnd cell_6t
Xbit_r37_c122 bl_122 br_122 wl_37 vdd gnd cell_6t
Xbit_r38_c122 bl_122 br_122 wl_38 vdd gnd cell_6t
Xbit_r39_c122 bl_122 br_122 wl_39 vdd gnd cell_6t
Xbit_r40_c122 bl_122 br_122 wl_40 vdd gnd cell_6t
Xbit_r41_c122 bl_122 br_122 wl_41 vdd gnd cell_6t
Xbit_r42_c122 bl_122 br_122 wl_42 vdd gnd cell_6t
Xbit_r43_c122 bl_122 br_122 wl_43 vdd gnd cell_6t
Xbit_r44_c122 bl_122 br_122 wl_44 vdd gnd cell_6t
Xbit_r45_c122 bl_122 br_122 wl_45 vdd gnd cell_6t
Xbit_r46_c122 bl_122 br_122 wl_46 vdd gnd cell_6t
Xbit_r47_c122 bl_122 br_122 wl_47 vdd gnd cell_6t
Xbit_r48_c122 bl_122 br_122 wl_48 vdd gnd cell_6t
Xbit_r49_c122 bl_122 br_122 wl_49 vdd gnd cell_6t
Xbit_r50_c122 bl_122 br_122 wl_50 vdd gnd cell_6t
Xbit_r51_c122 bl_122 br_122 wl_51 vdd gnd cell_6t
Xbit_r52_c122 bl_122 br_122 wl_52 vdd gnd cell_6t
Xbit_r53_c122 bl_122 br_122 wl_53 vdd gnd cell_6t
Xbit_r54_c122 bl_122 br_122 wl_54 vdd gnd cell_6t
Xbit_r55_c122 bl_122 br_122 wl_55 vdd gnd cell_6t
Xbit_r56_c122 bl_122 br_122 wl_56 vdd gnd cell_6t
Xbit_r57_c122 bl_122 br_122 wl_57 vdd gnd cell_6t
Xbit_r58_c122 bl_122 br_122 wl_58 vdd gnd cell_6t
Xbit_r59_c122 bl_122 br_122 wl_59 vdd gnd cell_6t
Xbit_r60_c122 bl_122 br_122 wl_60 vdd gnd cell_6t
Xbit_r61_c122 bl_122 br_122 wl_61 vdd gnd cell_6t
Xbit_r62_c122 bl_122 br_122 wl_62 vdd gnd cell_6t
Xbit_r63_c122 bl_122 br_122 wl_63 vdd gnd cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd cell_6t
Xbit_r1_c123 bl_123 br_123 wl_1 vdd gnd cell_6t
Xbit_r2_c123 bl_123 br_123 wl_2 vdd gnd cell_6t
Xbit_r3_c123 bl_123 br_123 wl_3 vdd gnd cell_6t
Xbit_r4_c123 bl_123 br_123 wl_4 vdd gnd cell_6t
Xbit_r5_c123 bl_123 br_123 wl_5 vdd gnd cell_6t
Xbit_r6_c123 bl_123 br_123 wl_6 vdd gnd cell_6t
Xbit_r7_c123 bl_123 br_123 wl_7 vdd gnd cell_6t
Xbit_r8_c123 bl_123 br_123 wl_8 vdd gnd cell_6t
Xbit_r9_c123 bl_123 br_123 wl_9 vdd gnd cell_6t
Xbit_r10_c123 bl_123 br_123 wl_10 vdd gnd cell_6t
Xbit_r11_c123 bl_123 br_123 wl_11 vdd gnd cell_6t
Xbit_r12_c123 bl_123 br_123 wl_12 vdd gnd cell_6t
Xbit_r13_c123 bl_123 br_123 wl_13 vdd gnd cell_6t
Xbit_r14_c123 bl_123 br_123 wl_14 vdd gnd cell_6t
Xbit_r15_c123 bl_123 br_123 wl_15 vdd gnd cell_6t
Xbit_r16_c123 bl_123 br_123 wl_16 vdd gnd cell_6t
Xbit_r17_c123 bl_123 br_123 wl_17 vdd gnd cell_6t
Xbit_r18_c123 bl_123 br_123 wl_18 vdd gnd cell_6t
Xbit_r19_c123 bl_123 br_123 wl_19 vdd gnd cell_6t
Xbit_r20_c123 bl_123 br_123 wl_20 vdd gnd cell_6t
Xbit_r21_c123 bl_123 br_123 wl_21 vdd gnd cell_6t
Xbit_r22_c123 bl_123 br_123 wl_22 vdd gnd cell_6t
Xbit_r23_c123 bl_123 br_123 wl_23 vdd gnd cell_6t
Xbit_r24_c123 bl_123 br_123 wl_24 vdd gnd cell_6t
Xbit_r25_c123 bl_123 br_123 wl_25 vdd gnd cell_6t
Xbit_r26_c123 bl_123 br_123 wl_26 vdd gnd cell_6t
Xbit_r27_c123 bl_123 br_123 wl_27 vdd gnd cell_6t
Xbit_r28_c123 bl_123 br_123 wl_28 vdd gnd cell_6t
Xbit_r29_c123 bl_123 br_123 wl_29 vdd gnd cell_6t
Xbit_r30_c123 bl_123 br_123 wl_30 vdd gnd cell_6t
Xbit_r31_c123 bl_123 br_123 wl_31 vdd gnd cell_6t
Xbit_r32_c123 bl_123 br_123 wl_32 vdd gnd cell_6t
Xbit_r33_c123 bl_123 br_123 wl_33 vdd gnd cell_6t
Xbit_r34_c123 bl_123 br_123 wl_34 vdd gnd cell_6t
Xbit_r35_c123 bl_123 br_123 wl_35 vdd gnd cell_6t
Xbit_r36_c123 bl_123 br_123 wl_36 vdd gnd cell_6t
Xbit_r37_c123 bl_123 br_123 wl_37 vdd gnd cell_6t
Xbit_r38_c123 bl_123 br_123 wl_38 vdd gnd cell_6t
Xbit_r39_c123 bl_123 br_123 wl_39 vdd gnd cell_6t
Xbit_r40_c123 bl_123 br_123 wl_40 vdd gnd cell_6t
Xbit_r41_c123 bl_123 br_123 wl_41 vdd gnd cell_6t
Xbit_r42_c123 bl_123 br_123 wl_42 vdd gnd cell_6t
Xbit_r43_c123 bl_123 br_123 wl_43 vdd gnd cell_6t
Xbit_r44_c123 bl_123 br_123 wl_44 vdd gnd cell_6t
Xbit_r45_c123 bl_123 br_123 wl_45 vdd gnd cell_6t
Xbit_r46_c123 bl_123 br_123 wl_46 vdd gnd cell_6t
Xbit_r47_c123 bl_123 br_123 wl_47 vdd gnd cell_6t
Xbit_r48_c123 bl_123 br_123 wl_48 vdd gnd cell_6t
Xbit_r49_c123 bl_123 br_123 wl_49 vdd gnd cell_6t
Xbit_r50_c123 bl_123 br_123 wl_50 vdd gnd cell_6t
Xbit_r51_c123 bl_123 br_123 wl_51 vdd gnd cell_6t
Xbit_r52_c123 bl_123 br_123 wl_52 vdd gnd cell_6t
Xbit_r53_c123 bl_123 br_123 wl_53 vdd gnd cell_6t
Xbit_r54_c123 bl_123 br_123 wl_54 vdd gnd cell_6t
Xbit_r55_c123 bl_123 br_123 wl_55 vdd gnd cell_6t
Xbit_r56_c123 bl_123 br_123 wl_56 vdd gnd cell_6t
Xbit_r57_c123 bl_123 br_123 wl_57 vdd gnd cell_6t
Xbit_r58_c123 bl_123 br_123 wl_58 vdd gnd cell_6t
Xbit_r59_c123 bl_123 br_123 wl_59 vdd gnd cell_6t
Xbit_r60_c123 bl_123 br_123 wl_60 vdd gnd cell_6t
Xbit_r61_c123 bl_123 br_123 wl_61 vdd gnd cell_6t
Xbit_r62_c123 bl_123 br_123 wl_62 vdd gnd cell_6t
Xbit_r63_c123 bl_123 br_123 wl_63 vdd gnd cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd cell_6t
Xbit_r1_c124 bl_124 br_124 wl_1 vdd gnd cell_6t
Xbit_r2_c124 bl_124 br_124 wl_2 vdd gnd cell_6t
Xbit_r3_c124 bl_124 br_124 wl_3 vdd gnd cell_6t
Xbit_r4_c124 bl_124 br_124 wl_4 vdd gnd cell_6t
Xbit_r5_c124 bl_124 br_124 wl_5 vdd gnd cell_6t
Xbit_r6_c124 bl_124 br_124 wl_6 vdd gnd cell_6t
Xbit_r7_c124 bl_124 br_124 wl_7 vdd gnd cell_6t
Xbit_r8_c124 bl_124 br_124 wl_8 vdd gnd cell_6t
Xbit_r9_c124 bl_124 br_124 wl_9 vdd gnd cell_6t
Xbit_r10_c124 bl_124 br_124 wl_10 vdd gnd cell_6t
Xbit_r11_c124 bl_124 br_124 wl_11 vdd gnd cell_6t
Xbit_r12_c124 bl_124 br_124 wl_12 vdd gnd cell_6t
Xbit_r13_c124 bl_124 br_124 wl_13 vdd gnd cell_6t
Xbit_r14_c124 bl_124 br_124 wl_14 vdd gnd cell_6t
Xbit_r15_c124 bl_124 br_124 wl_15 vdd gnd cell_6t
Xbit_r16_c124 bl_124 br_124 wl_16 vdd gnd cell_6t
Xbit_r17_c124 bl_124 br_124 wl_17 vdd gnd cell_6t
Xbit_r18_c124 bl_124 br_124 wl_18 vdd gnd cell_6t
Xbit_r19_c124 bl_124 br_124 wl_19 vdd gnd cell_6t
Xbit_r20_c124 bl_124 br_124 wl_20 vdd gnd cell_6t
Xbit_r21_c124 bl_124 br_124 wl_21 vdd gnd cell_6t
Xbit_r22_c124 bl_124 br_124 wl_22 vdd gnd cell_6t
Xbit_r23_c124 bl_124 br_124 wl_23 vdd gnd cell_6t
Xbit_r24_c124 bl_124 br_124 wl_24 vdd gnd cell_6t
Xbit_r25_c124 bl_124 br_124 wl_25 vdd gnd cell_6t
Xbit_r26_c124 bl_124 br_124 wl_26 vdd gnd cell_6t
Xbit_r27_c124 bl_124 br_124 wl_27 vdd gnd cell_6t
Xbit_r28_c124 bl_124 br_124 wl_28 vdd gnd cell_6t
Xbit_r29_c124 bl_124 br_124 wl_29 vdd gnd cell_6t
Xbit_r30_c124 bl_124 br_124 wl_30 vdd gnd cell_6t
Xbit_r31_c124 bl_124 br_124 wl_31 vdd gnd cell_6t
Xbit_r32_c124 bl_124 br_124 wl_32 vdd gnd cell_6t
Xbit_r33_c124 bl_124 br_124 wl_33 vdd gnd cell_6t
Xbit_r34_c124 bl_124 br_124 wl_34 vdd gnd cell_6t
Xbit_r35_c124 bl_124 br_124 wl_35 vdd gnd cell_6t
Xbit_r36_c124 bl_124 br_124 wl_36 vdd gnd cell_6t
Xbit_r37_c124 bl_124 br_124 wl_37 vdd gnd cell_6t
Xbit_r38_c124 bl_124 br_124 wl_38 vdd gnd cell_6t
Xbit_r39_c124 bl_124 br_124 wl_39 vdd gnd cell_6t
Xbit_r40_c124 bl_124 br_124 wl_40 vdd gnd cell_6t
Xbit_r41_c124 bl_124 br_124 wl_41 vdd gnd cell_6t
Xbit_r42_c124 bl_124 br_124 wl_42 vdd gnd cell_6t
Xbit_r43_c124 bl_124 br_124 wl_43 vdd gnd cell_6t
Xbit_r44_c124 bl_124 br_124 wl_44 vdd gnd cell_6t
Xbit_r45_c124 bl_124 br_124 wl_45 vdd gnd cell_6t
Xbit_r46_c124 bl_124 br_124 wl_46 vdd gnd cell_6t
Xbit_r47_c124 bl_124 br_124 wl_47 vdd gnd cell_6t
Xbit_r48_c124 bl_124 br_124 wl_48 vdd gnd cell_6t
Xbit_r49_c124 bl_124 br_124 wl_49 vdd gnd cell_6t
Xbit_r50_c124 bl_124 br_124 wl_50 vdd gnd cell_6t
Xbit_r51_c124 bl_124 br_124 wl_51 vdd gnd cell_6t
Xbit_r52_c124 bl_124 br_124 wl_52 vdd gnd cell_6t
Xbit_r53_c124 bl_124 br_124 wl_53 vdd gnd cell_6t
Xbit_r54_c124 bl_124 br_124 wl_54 vdd gnd cell_6t
Xbit_r55_c124 bl_124 br_124 wl_55 vdd gnd cell_6t
Xbit_r56_c124 bl_124 br_124 wl_56 vdd gnd cell_6t
Xbit_r57_c124 bl_124 br_124 wl_57 vdd gnd cell_6t
Xbit_r58_c124 bl_124 br_124 wl_58 vdd gnd cell_6t
Xbit_r59_c124 bl_124 br_124 wl_59 vdd gnd cell_6t
Xbit_r60_c124 bl_124 br_124 wl_60 vdd gnd cell_6t
Xbit_r61_c124 bl_124 br_124 wl_61 vdd gnd cell_6t
Xbit_r62_c124 bl_124 br_124 wl_62 vdd gnd cell_6t
Xbit_r63_c124 bl_124 br_124 wl_63 vdd gnd cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd cell_6t
Xbit_r1_c125 bl_125 br_125 wl_1 vdd gnd cell_6t
Xbit_r2_c125 bl_125 br_125 wl_2 vdd gnd cell_6t
Xbit_r3_c125 bl_125 br_125 wl_3 vdd gnd cell_6t
Xbit_r4_c125 bl_125 br_125 wl_4 vdd gnd cell_6t
Xbit_r5_c125 bl_125 br_125 wl_5 vdd gnd cell_6t
Xbit_r6_c125 bl_125 br_125 wl_6 vdd gnd cell_6t
Xbit_r7_c125 bl_125 br_125 wl_7 vdd gnd cell_6t
Xbit_r8_c125 bl_125 br_125 wl_8 vdd gnd cell_6t
Xbit_r9_c125 bl_125 br_125 wl_9 vdd gnd cell_6t
Xbit_r10_c125 bl_125 br_125 wl_10 vdd gnd cell_6t
Xbit_r11_c125 bl_125 br_125 wl_11 vdd gnd cell_6t
Xbit_r12_c125 bl_125 br_125 wl_12 vdd gnd cell_6t
Xbit_r13_c125 bl_125 br_125 wl_13 vdd gnd cell_6t
Xbit_r14_c125 bl_125 br_125 wl_14 vdd gnd cell_6t
Xbit_r15_c125 bl_125 br_125 wl_15 vdd gnd cell_6t
Xbit_r16_c125 bl_125 br_125 wl_16 vdd gnd cell_6t
Xbit_r17_c125 bl_125 br_125 wl_17 vdd gnd cell_6t
Xbit_r18_c125 bl_125 br_125 wl_18 vdd gnd cell_6t
Xbit_r19_c125 bl_125 br_125 wl_19 vdd gnd cell_6t
Xbit_r20_c125 bl_125 br_125 wl_20 vdd gnd cell_6t
Xbit_r21_c125 bl_125 br_125 wl_21 vdd gnd cell_6t
Xbit_r22_c125 bl_125 br_125 wl_22 vdd gnd cell_6t
Xbit_r23_c125 bl_125 br_125 wl_23 vdd gnd cell_6t
Xbit_r24_c125 bl_125 br_125 wl_24 vdd gnd cell_6t
Xbit_r25_c125 bl_125 br_125 wl_25 vdd gnd cell_6t
Xbit_r26_c125 bl_125 br_125 wl_26 vdd gnd cell_6t
Xbit_r27_c125 bl_125 br_125 wl_27 vdd gnd cell_6t
Xbit_r28_c125 bl_125 br_125 wl_28 vdd gnd cell_6t
Xbit_r29_c125 bl_125 br_125 wl_29 vdd gnd cell_6t
Xbit_r30_c125 bl_125 br_125 wl_30 vdd gnd cell_6t
Xbit_r31_c125 bl_125 br_125 wl_31 vdd gnd cell_6t
Xbit_r32_c125 bl_125 br_125 wl_32 vdd gnd cell_6t
Xbit_r33_c125 bl_125 br_125 wl_33 vdd gnd cell_6t
Xbit_r34_c125 bl_125 br_125 wl_34 vdd gnd cell_6t
Xbit_r35_c125 bl_125 br_125 wl_35 vdd gnd cell_6t
Xbit_r36_c125 bl_125 br_125 wl_36 vdd gnd cell_6t
Xbit_r37_c125 bl_125 br_125 wl_37 vdd gnd cell_6t
Xbit_r38_c125 bl_125 br_125 wl_38 vdd gnd cell_6t
Xbit_r39_c125 bl_125 br_125 wl_39 vdd gnd cell_6t
Xbit_r40_c125 bl_125 br_125 wl_40 vdd gnd cell_6t
Xbit_r41_c125 bl_125 br_125 wl_41 vdd gnd cell_6t
Xbit_r42_c125 bl_125 br_125 wl_42 vdd gnd cell_6t
Xbit_r43_c125 bl_125 br_125 wl_43 vdd gnd cell_6t
Xbit_r44_c125 bl_125 br_125 wl_44 vdd gnd cell_6t
Xbit_r45_c125 bl_125 br_125 wl_45 vdd gnd cell_6t
Xbit_r46_c125 bl_125 br_125 wl_46 vdd gnd cell_6t
Xbit_r47_c125 bl_125 br_125 wl_47 vdd gnd cell_6t
Xbit_r48_c125 bl_125 br_125 wl_48 vdd gnd cell_6t
Xbit_r49_c125 bl_125 br_125 wl_49 vdd gnd cell_6t
Xbit_r50_c125 bl_125 br_125 wl_50 vdd gnd cell_6t
Xbit_r51_c125 bl_125 br_125 wl_51 vdd gnd cell_6t
Xbit_r52_c125 bl_125 br_125 wl_52 vdd gnd cell_6t
Xbit_r53_c125 bl_125 br_125 wl_53 vdd gnd cell_6t
Xbit_r54_c125 bl_125 br_125 wl_54 vdd gnd cell_6t
Xbit_r55_c125 bl_125 br_125 wl_55 vdd gnd cell_6t
Xbit_r56_c125 bl_125 br_125 wl_56 vdd gnd cell_6t
Xbit_r57_c125 bl_125 br_125 wl_57 vdd gnd cell_6t
Xbit_r58_c125 bl_125 br_125 wl_58 vdd gnd cell_6t
Xbit_r59_c125 bl_125 br_125 wl_59 vdd gnd cell_6t
Xbit_r60_c125 bl_125 br_125 wl_60 vdd gnd cell_6t
Xbit_r61_c125 bl_125 br_125 wl_61 vdd gnd cell_6t
Xbit_r62_c125 bl_125 br_125 wl_62 vdd gnd cell_6t
Xbit_r63_c125 bl_125 br_125 wl_63 vdd gnd cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd cell_6t
Xbit_r1_c126 bl_126 br_126 wl_1 vdd gnd cell_6t
Xbit_r2_c126 bl_126 br_126 wl_2 vdd gnd cell_6t
Xbit_r3_c126 bl_126 br_126 wl_3 vdd gnd cell_6t
Xbit_r4_c126 bl_126 br_126 wl_4 vdd gnd cell_6t
Xbit_r5_c126 bl_126 br_126 wl_5 vdd gnd cell_6t
Xbit_r6_c126 bl_126 br_126 wl_6 vdd gnd cell_6t
Xbit_r7_c126 bl_126 br_126 wl_7 vdd gnd cell_6t
Xbit_r8_c126 bl_126 br_126 wl_8 vdd gnd cell_6t
Xbit_r9_c126 bl_126 br_126 wl_9 vdd gnd cell_6t
Xbit_r10_c126 bl_126 br_126 wl_10 vdd gnd cell_6t
Xbit_r11_c126 bl_126 br_126 wl_11 vdd gnd cell_6t
Xbit_r12_c126 bl_126 br_126 wl_12 vdd gnd cell_6t
Xbit_r13_c126 bl_126 br_126 wl_13 vdd gnd cell_6t
Xbit_r14_c126 bl_126 br_126 wl_14 vdd gnd cell_6t
Xbit_r15_c126 bl_126 br_126 wl_15 vdd gnd cell_6t
Xbit_r16_c126 bl_126 br_126 wl_16 vdd gnd cell_6t
Xbit_r17_c126 bl_126 br_126 wl_17 vdd gnd cell_6t
Xbit_r18_c126 bl_126 br_126 wl_18 vdd gnd cell_6t
Xbit_r19_c126 bl_126 br_126 wl_19 vdd gnd cell_6t
Xbit_r20_c126 bl_126 br_126 wl_20 vdd gnd cell_6t
Xbit_r21_c126 bl_126 br_126 wl_21 vdd gnd cell_6t
Xbit_r22_c126 bl_126 br_126 wl_22 vdd gnd cell_6t
Xbit_r23_c126 bl_126 br_126 wl_23 vdd gnd cell_6t
Xbit_r24_c126 bl_126 br_126 wl_24 vdd gnd cell_6t
Xbit_r25_c126 bl_126 br_126 wl_25 vdd gnd cell_6t
Xbit_r26_c126 bl_126 br_126 wl_26 vdd gnd cell_6t
Xbit_r27_c126 bl_126 br_126 wl_27 vdd gnd cell_6t
Xbit_r28_c126 bl_126 br_126 wl_28 vdd gnd cell_6t
Xbit_r29_c126 bl_126 br_126 wl_29 vdd gnd cell_6t
Xbit_r30_c126 bl_126 br_126 wl_30 vdd gnd cell_6t
Xbit_r31_c126 bl_126 br_126 wl_31 vdd gnd cell_6t
Xbit_r32_c126 bl_126 br_126 wl_32 vdd gnd cell_6t
Xbit_r33_c126 bl_126 br_126 wl_33 vdd gnd cell_6t
Xbit_r34_c126 bl_126 br_126 wl_34 vdd gnd cell_6t
Xbit_r35_c126 bl_126 br_126 wl_35 vdd gnd cell_6t
Xbit_r36_c126 bl_126 br_126 wl_36 vdd gnd cell_6t
Xbit_r37_c126 bl_126 br_126 wl_37 vdd gnd cell_6t
Xbit_r38_c126 bl_126 br_126 wl_38 vdd gnd cell_6t
Xbit_r39_c126 bl_126 br_126 wl_39 vdd gnd cell_6t
Xbit_r40_c126 bl_126 br_126 wl_40 vdd gnd cell_6t
Xbit_r41_c126 bl_126 br_126 wl_41 vdd gnd cell_6t
Xbit_r42_c126 bl_126 br_126 wl_42 vdd gnd cell_6t
Xbit_r43_c126 bl_126 br_126 wl_43 vdd gnd cell_6t
Xbit_r44_c126 bl_126 br_126 wl_44 vdd gnd cell_6t
Xbit_r45_c126 bl_126 br_126 wl_45 vdd gnd cell_6t
Xbit_r46_c126 bl_126 br_126 wl_46 vdd gnd cell_6t
Xbit_r47_c126 bl_126 br_126 wl_47 vdd gnd cell_6t
Xbit_r48_c126 bl_126 br_126 wl_48 vdd gnd cell_6t
Xbit_r49_c126 bl_126 br_126 wl_49 vdd gnd cell_6t
Xbit_r50_c126 bl_126 br_126 wl_50 vdd gnd cell_6t
Xbit_r51_c126 bl_126 br_126 wl_51 vdd gnd cell_6t
Xbit_r52_c126 bl_126 br_126 wl_52 vdd gnd cell_6t
Xbit_r53_c126 bl_126 br_126 wl_53 vdd gnd cell_6t
Xbit_r54_c126 bl_126 br_126 wl_54 vdd gnd cell_6t
Xbit_r55_c126 bl_126 br_126 wl_55 vdd gnd cell_6t
Xbit_r56_c126 bl_126 br_126 wl_56 vdd gnd cell_6t
Xbit_r57_c126 bl_126 br_126 wl_57 vdd gnd cell_6t
Xbit_r58_c126 bl_126 br_126 wl_58 vdd gnd cell_6t
Xbit_r59_c126 bl_126 br_126 wl_59 vdd gnd cell_6t
Xbit_r60_c126 bl_126 br_126 wl_60 vdd gnd cell_6t
Xbit_r61_c126 bl_126 br_126 wl_61 vdd gnd cell_6t
Xbit_r62_c126 bl_126 br_126 wl_62 vdd gnd cell_6t
Xbit_r63_c126 bl_126 br_126 wl_63 vdd gnd cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd cell_6t
Xbit_r1_c127 bl_127 br_127 wl_1 vdd gnd cell_6t
Xbit_r2_c127 bl_127 br_127 wl_2 vdd gnd cell_6t
Xbit_r3_c127 bl_127 br_127 wl_3 vdd gnd cell_6t
Xbit_r4_c127 bl_127 br_127 wl_4 vdd gnd cell_6t
Xbit_r5_c127 bl_127 br_127 wl_5 vdd gnd cell_6t
Xbit_r6_c127 bl_127 br_127 wl_6 vdd gnd cell_6t
Xbit_r7_c127 bl_127 br_127 wl_7 vdd gnd cell_6t
Xbit_r8_c127 bl_127 br_127 wl_8 vdd gnd cell_6t
Xbit_r9_c127 bl_127 br_127 wl_9 vdd gnd cell_6t
Xbit_r10_c127 bl_127 br_127 wl_10 vdd gnd cell_6t
Xbit_r11_c127 bl_127 br_127 wl_11 vdd gnd cell_6t
Xbit_r12_c127 bl_127 br_127 wl_12 vdd gnd cell_6t
Xbit_r13_c127 bl_127 br_127 wl_13 vdd gnd cell_6t
Xbit_r14_c127 bl_127 br_127 wl_14 vdd gnd cell_6t
Xbit_r15_c127 bl_127 br_127 wl_15 vdd gnd cell_6t
Xbit_r16_c127 bl_127 br_127 wl_16 vdd gnd cell_6t
Xbit_r17_c127 bl_127 br_127 wl_17 vdd gnd cell_6t
Xbit_r18_c127 bl_127 br_127 wl_18 vdd gnd cell_6t
Xbit_r19_c127 bl_127 br_127 wl_19 vdd gnd cell_6t
Xbit_r20_c127 bl_127 br_127 wl_20 vdd gnd cell_6t
Xbit_r21_c127 bl_127 br_127 wl_21 vdd gnd cell_6t
Xbit_r22_c127 bl_127 br_127 wl_22 vdd gnd cell_6t
Xbit_r23_c127 bl_127 br_127 wl_23 vdd gnd cell_6t
Xbit_r24_c127 bl_127 br_127 wl_24 vdd gnd cell_6t
Xbit_r25_c127 bl_127 br_127 wl_25 vdd gnd cell_6t
Xbit_r26_c127 bl_127 br_127 wl_26 vdd gnd cell_6t
Xbit_r27_c127 bl_127 br_127 wl_27 vdd gnd cell_6t
Xbit_r28_c127 bl_127 br_127 wl_28 vdd gnd cell_6t
Xbit_r29_c127 bl_127 br_127 wl_29 vdd gnd cell_6t
Xbit_r30_c127 bl_127 br_127 wl_30 vdd gnd cell_6t
Xbit_r31_c127 bl_127 br_127 wl_31 vdd gnd cell_6t
Xbit_r32_c127 bl_127 br_127 wl_32 vdd gnd cell_6t
Xbit_r33_c127 bl_127 br_127 wl_33 vdd gnd cell_6t
Xbit_r34_c127 bl_127 br_127 wl_34 vdd gnd cell_6t
Xbit_r35_c127 bl_127 br_127 wl_35 vdd gnd cell_6t
Xbit_r36_c127 bl_127 br_127 wl_36 vdd gnd cell_6t
Xbit_r37_c127 bl_127 br_127 wl_37 vdd gnd cell_6t
Xbit_r38_c127 bl_127 br_127 wl_38 vdd gnd cell_6t
Xbit_r39_c127 bl_127 br_127 wl_39 vdd gnd cell_6t
Xbit_r40_c127 bl_127 br_127 wl_40 vdd gnd cell_6t
Xbit_r41_c127 bl_127 br_127 wl_41 vdd gnd cell_6t
Xbit_r42_c127 bl_127 br_127 wl_42 vdd gnd cell_6t
Xbit_r43_c127 bl_127 br_127 wl_43 vdd gnd cell_6t
Xbit_r44_c127 bl_127 br_127 wl_44 vdd gnd cell_6t
Xbit_r45_c127 bl_127 br_127 wl_45 vdd gnd cell_6t
Xbit_r46_c127 bl_127 br_127 wl_46 vdd gnd cell_6t
Xbit_r47_c127 bl_127 br_127 wl_47 vdd gnd cell_6t
Xbit_r48_c127 bl_127 br_127 wl_48 vdd gnd cell_6t
Xbit_r49_c127 bl_127 br_127 wl_49 vdd gnd cell_6t
Xbit_r50_c127 bl_127 br_127 wl_50 vdd gnd cell_6t
Xbit_r51_c127 bl_127 br_127 wl_51 vdd gnd cell_6t
Xbit_r52_c127 bl_127 br_127 wl_52 vdd gnd cell_6t
Xbit_r53_c127 bl_127 br_127 wl_53 vdd gnd cell_6t
Xbit_r54_c127 bl_127 br_127 wl_54 vdd gnd cell_6t
Xbit_r55_c127 bl_127 br_127 wl_55 vdd gnd cell_6t
Xbit_r56_c127 bl_127 br_127 wl_56 vdd gnd cell_6t
Xbit_r57_c127 bl_127 br_127 wl_57 vdd gnd cell_6t
Xbit_r58_c127 bl_127 br_127 wl_58 vdd gnd cell_6t
Xbit_r59_c127 bl_127 br_127 wl_59 vdd gnd cell_6t
Xbit_r60_c127 bl_127 br_127 wl_60 vdd gnd cell_6t
Xbit_r61_c127 bl_127 br_127 wl_61 vdd gnd cell_6t
Xbit_r62_c127 bl_127 br_127 wl_62 vdd gnd cell_6t
Xbit_r63_c127 bl_127 br_127 wl_63 vdd gnd cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd cell_6t
Xbit_r1_c128 bl_128 br_128 wl_1 vdd gnd cell_6t
Xbit_r2_c128 bl_128 br_128 wl_2 vdd gnd cell_6t
Xbit_r3_c128 bl_128 br_128 wl_3 vdd gnd cell_6t
Xbit_r4_c128 bl_128 br_128 wl_4 vdd gnd cell_6t
Xbit_r5_c128 bl_128 br_128 wl_5 vdd gnd cell_6t
Xbit_r6_c128 bl_128 br_128 wl_6 vdd gnd cell_6t
Xbit_r7_c128 bl_128 br_128 wl_7 vdd gnd cell_6t
Xbit_r8_c128 bl_128 br_128 wl_8 vdd gnd cell_6t
Xbit_r9_c128 bl_128 br_128 wl_9 vdd gnd cell_6t
Xbit_r10_c128 bl_128 br_128 wl_10 vdd gnd cell_6t
Xbit_r11_c128 bl_128 br_128 wl_11 vdd gnd cell_6t
Xbit_r12_c128 bl_128 br_128 wl_12 vdd gnd cell_6t
Xbit_r13_c128 bl_128 br_128 wl_13 vdd gnd cell_6t
Xbit_r14_c128 bl_128 br_128 wl_14 vdd gnd cell_6t
Xbit_r15_c128 bl_128 br_128 wl_15 vdd gnd cell_6t
Xbit_r16_c128 bl_128 br_128 wl_16 vdd gnd cell_6t
Xbit_r17_c128 bl_128 br_128 wl_17 vdd gnd cell_6t
Xbit_r18_c128 bl_128 br_128 wl_18 vdd gnd cell_6t
Xbit_r19_c128 bl_128 br_128 wl_19 vdd gnd cell_6t
Xbit_r20_c128 bl_128 br_128 wl_20 vdd gnd cell_6t
Xbit_r21_c128 bl_128 br_128 wl_21 vdd gnd cell_6t
Xbit_r22_c128 bl_128 br_128 wl_22 vdd gnd cell_6t
Xbit_r23_c128 bl_128 br_128 wl_23 vdd gnd cell_6t
Xbit_r24_c128 bl_128 br_128 wl_24 vdd gnd cell_6t
Xbit_r25_c128 bl_128 br_128 wl_25 vdd gnd cell_6t
Xbit_r26_c128 bl_128 br_128 wl_26 vdd gnd cell_6t
Xbit_r27_c128 bl_128 br_128 wl_27 vdd gnd cell_6t
Xbit_r28_c128 bl_128 br_128 wl_28 vdd gnd cell_6t
Xbit_r29_c128 bl_128 br_128 wl_29 vdd gnd cell_6t
Xbit_r30_c128 bl_128 br_128 wl_30 vdd gnd cell_6t
Xbit_r31_c128 bl_128 br_128 wl_31 vdd gnd cell_6t
Xbit_r32_c128 bl_128 br_128 wl_32 vdd gnd cell_6t
Xbit_r33_c128 bl_128 br_128 wl_33 vdd gnd cell_6t
Xbit_r34_c128 bl_128 br_128 wl_34 vdd gnd cell_6t
Xbit_r35_c128 bl_128 br_128 wl_35 vdd gnd cell_6t
Xbit_r36_c128 bl_128 br_128 wl_36 vdd gnd cell_6t
Xbit_r37_c128 bl_128 br_128 wl_37 vdd gnd cell_6t
Xbit_r38_c128 bl_128 br_128 wl_38 vdd gnd cell_6t
Xbit_r39_c128 bl_128 br_128 wl_39 vdd gnd cell_6t
Xbit_r40_c128 bl_128 br_128 wl_40 vdd gnd cell_6t
Xbit_r41_c128 bl_128 br_128 wl_41 vdd gnd cell_6t
Xbit_r42_c128 bl_128 br_128 wl_42 vdd gnd cell_6t
Xbit_r43_c128 bl_128 br_128 wl_43 vdd gnd cell_6t
Xbit_r44_c128 bl_128 br_128 wl_44 vdd gnd cell_6t
Xbit_r45_c128 bl_128 br_128 wl_45 vdd gnd cell_6t
Xbit_r46_c128 bl_128 br_128 wl_46 vdd gnd cell_6t
Xbit_r47_c128 bl_128 br_128 wl_47 vdd gnd cell_6t
Xbit_r48_c128 bl_128 br_128 wl_48 vdd gnd cell_6t
Xbit_r49_c128 bl_128 br_128 wl_49 vdd gnd cell_6t
Xbit_r50_c128 bl_128 br_128 wl_50 vdd gnd cell_6t
Xbit_r51_c128 bl_128 br_128 wl_51 vdd gnd cell_6t
Xbit_r52_c128 bl_128 br_128 wl_52 vdd gnd cell_6t
Xbit_r53_c128 bl_128 br_128 wl_53 vdd gnd cell_6t
Xbit_r54_c128 bl_128 br_128 wl_54 vdd gnd cell_6t
Xbit_r55_c128 bl_128 br_128 wl_55 vdd gnd cell_6t
Xbit_r56_c128 bl_128 br_128 wl_56 vdd gnd cell_6t
Xbit_r57_c128 bl_128 br_128 wl_57 vdd gnd cell_6t
Xbit_r58_c128 bl_128 br_128 wl_58 vdd gnd cell_6t
Xbit_r59_c128 bl_128 br_128 wl_59 vdd gnd cell_6t
Xbit_r60_c128 bl_128 br_128 wl_60 vdd gnd cell_6t
Xbit_r61_c128 bl_128 br_128 wl_61 vdd gnd cell_6t
Xbit_r62_c128 bl_128 br_128 wl_62 vdd gnd cell_6t
Xbit_r63_c128 bl_128 br_128 wl_63 vdd gnd cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd cell_6t
Xbit_r1_c129 bl_129 br_129 wl_1 vdd gnd cell_6t
Xbit_r2_c129 bl_129 br_129 wl_2 vdd gnd cell_6t
Xbit_r3_c129 bl_129 br_129 wl_3 vdd gnd cell_6t
Xbit_r4_c129 bl_129 br_129 wl_4 vdd gnd cell_6t
Xbit_r5_c129 bl_129 br_129 wl_5 vdd gnd cell_6t
Xbit_r6_c129 bl_129 br_129 wl_6 vdd gnd cell_6t
Xbit_r7_c129 bl_129 br_129 wl_7 vdd gnd cell_6t
Xbit_r8_c129 bl_129 br_129 wl_8 vdd gnd cell_6t
Xbit_r9_c129 bl_129 br_129 wl_9 vdd gnd cell_6t
Xbit_r10_c129 bl_129 br_129 wl_10 vdd gnd cell_6t
Xbit_r11_c129 bl_129 br_129 wl_11 vdd gnd cell_6t
Xbit_r12_c129 bl_129 br_129 wl_12 vdd gnd cell_6t
Xbit_r13_c129 bl_129 br_129 wl_13 vdd gnd cell_6t
Xbit_r14_c129 bl_129 br_129 wl_14 vdd gnd cell_6t
Xbit_r15_c129 bl_129 br_129 wl_15 vdd gnd cell_6t
Xbit_r16_c129 bl_129 br_129 wl_16 vdd gnd cell_6t
Xbit_r17_c129 bl_129 br_129 wl_17 vdd gnd cell_6t
Xbit_r18_c129 bl_129 br_129 wl_18 vdd gnd cell_6t
Xbit_r19_c129 bl_129 br_129 wl_19 vdd gnd cell_6t
Xbit_r20_c129 bl_129 br_129 wl_20 vdd gnd cell_6t
Xbit_r21_c129 bl_129 br_129 wl_21 vdd gnd cell_6t
Xbit_r22_c129 bl_129 br_129 wl_22 vdd gnd cell_6t
Xbit_r23_c129 bl_129 br_129 wl_23 vdd gnd cell_6t
Xbit_r24_c129 bl_129 br_129 wl_24 vdd gnd cell_6t
Xbit_r25_c129 bl_129 br_129 wl_25 vdd gnd cell_6t
Xbit_r26_c129 bl_129 br_129 wl_26 vdd gnd cell_6t
Xbit_r27_c129 bl_129 br_129 wl_27 vdd gnd cell_6t
Xbit_r28_c129 bl_129 br_129 wl_28 vdd gnd cell_6t
Xbit_r29_c129 bl_129 br_129 wl_29 vdd gnd cell_6t
Xbit_r30_c129 bl_129 br_129 wl_30 vdd gnd cell_6t
Xbit_r31_c129 bl_129 br_129 wl_31 vdd gnd cell_6t
Xbit_r32_c129 bl_129 br_129 wl_32 vdd gnd cell_6t
Xbit_r33_c129 bl_129 br_129 wl_33 vdd gnd cell_6t
Xbit_r34_c129 bl_129 br_129 wl_34 vdd gnd cell_6t
Xbit_r35_c129 bl_129 br_129 wl_35 vdd gnd cell_6t
Xbit_r36_c129 bl_129 br_129 wl_36 vdd gnd cell_6t
Xbit_r37_c129 bl_129 br_129 wl_37 vdd gnd cell_6t
Xbit_r38_c129 bl_129 br_129 wl_38 vdd gnd cell_6t
Xbit_r39_c129 bl_129 br_129 wl_39 vdd gnd cell_6t
Xbit_r40_c129 bl_129 br_129 wl_40 vdd gnd cell_6t
Xbit_r41_c129 bl_129 br_129 wl_41 vdd gnd cell_6t
Xbit_r42_c129 bl_129 br_129 wl_42 vdd gnd cell_6t
Xbit_r43_c129 bl_129 br_129 wl_43 vdd gnd cell_6t
Xbit_r44_c129 bl_129 br_129 wl_44 vdd gnd cell_6t
Xbit_r45_c129 bl_129 br_129 wl_45 vdd gnd cell_6t
Xbit_r46_c129 bl_129 br_129 wl_46 vdd gnd cell_6t
Xbit_r47_c129 bl_129 br_129 wl_47 vdd gnd cell_6t
Xbit_r48_c129 bl_129 br_129 wl_48 vdd gnd cell_6t
Xbit_r49_c129 bl_129 br_129 wl_49 vdd gnd cell_6t
Xbit_r50_c129 bl_129 br_129 wl_50 vdd gnd cell_6t
Xbit_r51_c129 bl_129 br_129 wl_51 vdd gnd cell_6t
Xbit_r52_c129 bl_129 br_129 wl_52 vdd gnd cell_6t
Xbit_r53_c129 bl_129 br_129 wl_53 vdd gnd cell_6t
Xbit_r54_c129 bl_129 br_129 wl_54 vdd gnd cell_6t
Xbit_r55_c129 bl_129 br_129 wl_55 vdd gnd cell_6t
Xbit_r56_c129 bl_129 br_129 wl_56 vdd gnd cell_6t
Xbit_r57_c129 bl_129 br_129 wl_57 vdd gnd cell_6t
Xbit_r58_c129 bl_129 br_129 wl_58 vdd gnd cell_6t
Xbit_r59_c129 bl_129 br_129 wl_59 vdd gnd cell_6t
Xbit_r60_c129 bl_129 br_129 wl_60 vdd gnd cell_6t
Xbit_r61_c129 bl_129 br_129 wl_61 vdd gnd cell_6t
Xbit_r62_c129 bl_129 br_129 wl_62 vdd gnd cell_6t
Xbit_r63_c129 bl_129 br_129 wl_63 vdd gnd cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd cell_6t
Xbit_r1_c130 bl_130 br_130 wl_1 vdd gnd cell_6t
Xbit_r2_c130 bl_130 br_130 wl_2 vdd gnd cell_6t
Xbit_r3_c130 bl_130 br_130 wl_3 vdd gnd cell_6t
Xbit_r4_c130 bl_130 br_130 wl_4 vdd gnd cell_6t
Xbit_r5_c130 bl_130 br_130 wl_5 vdd gnd cell_6t
Xbit_r6_c130 bl_130 br_130 wl_6 vdd gnd cell_6t
Xbit_r7_c130 bl_130 br_130 wl_7 vdd gnd cell_6t
Xbit_r8_c130 bl_130 br_130 wl_8 vdd gnd cell_6t
Xbit_r9_c130 bl_130 br_130 wl_9 vdd gnd cell_6t
Xbit_r10_c130 bl_130 br_130 wl_10 vdd gnd cell_6t
Xbit_r11_c130 bl_130 br_130 wl_11 vdd gnd cell_6t
Xbit_r12_c130 bl_130 br_130 wl_12 vdd gnd cell_6t
Xbit_r13_c130 bl_130 br_130 wl_13 vdd gnd cell_6t
Xbit_r14_c130 bl_130 br_130 wl_14 vdd gnd cell_6t
Xbit_r15_c130 bl_130 br_130 wl_15 vdd gnd cell_6t
Xbit_r16_c130 bl_130 br_130 wl_16 vdd gnd cell_6t
Xbit_r17_c130 bl_130 br_130 wl_17 vdd gnd cell_6t
Xbit_r18_c130 bl_130 br_130 wl_18 vdd gnd cell_6t
Xbit_r19_c130 bl_130 br_130 wl_19 vdd gnd cell_6t
Xbit_r20_c130 bl_130 br_130 wl_20 vdd gnd cell_6t
Xbit_r21_c130 bl_130 br_130 wl_21 vdd gnd cell_6t
Xbit_r22_c130 bl_130 br_130 wl_22 vdd gnd cell_6t
Xbit_r23_c130 bl_130 br_130 wl_23 vdd gnd cell_6t
Xbit_r24_c130 bl_130 br_130 wl_24 vdd gnd cell_6t
Xbit_r25_c130 bl_130 br_130 wl_25 vdd gnd cell_6t
Xbit_r26_c130 bl_130 br_130 wl_26 vdd gnd cell_6t
Xbit_r27_c130 bl_130 br_130 wl_27 vdd gnd cell_6t
Xbit_r28_c130 bl_130 br_130 wl_28 vdd gnd cell_6t
Xbit_r29_c130 bl_130 br_130 wl_29 vdd gnd cell_6t
Xbit_r30_c130 bl_130 br_130 wl_30 vdd gnd cell_6t
Xbit_r31_c130 bl_130 br_130 wl_31 vdd gnd cell_6t
Xbit_r32_c130 bl_130 br_130 wl_32 vdd gnd cell_6t
Xbit_r33_c130 bl_130 br_130 wl_33 vdd gnd cell_6t
Xbit_r34_c130 bl_130 br_130 wl_34 vdd gnd cell_6t
Xbit_r35_c130 bl_130 br_130 wl_35 vdd gnd cell_6t
Xbit_r36_c130 bl_130 br_130 wl_36 vdd gnd cell_6t
Xbit_r37_c130 bl_130 br_130 wl_37 vdd gnd cell_6t
Xbit_r38_c130 bl_130 br_130 wl_38 vdd gnd cell_6t
Xbit_r39_c130 bl_130 br_130 wl_39 vdd gnd cell_6t
Xbit_r40_c130 bl_130 br_130 wl_40 vdd gnd cell_6t
Xbit_r41_c130 bl_130 br_130 wl_41 vdd gnd cell_6t
Xbit_r42_c130 bl_130 br_130 wl_42 vdd gnd cell_6t
Xbit_r43_c130 bl_130 br_130 wl_43 vdd gnd cell_6t
Xbit_r44_c130 bl_130 br_130 wl_44 vdd gnd cell_6t
Xbit_r45_c130 bl_130 br_130 wl_45 vdd gnd cell_6t
Xbit_r46_c130 bl_130 br_130 wl_46 vdd gnd cell_6t
Xbit_r47_c130 bl_130 br_130 wl_47 vdd gnd cell_6t
Xbit_r48_c130 bl_130 br_130 wl_48 vdd gnd cell_6t
Xbit_r49_c130 bl_130 br_130 wl_49 vdd gnd cell_6t
Xbit_r50_c130 bl_130 br_130 wl_50 vdd gnd cell_6t
Xbit_r51_c130 bl_130 br_130 wl_51 vdd gnd cell_6t
Xbit_r52_c130 bl_130 br_130 wl_52 vdd gnd cell_6t
Xbit_r53_c130 bl_130 br_130 wl_53 vdd gnd cell_6t
Xbit_r54_c130 bl_130 br_130 wl_54 vdd gnd cell_6t
Xbit_r55_c130 bl_130 br_130 wl_55 vdd gnd cell_6t
Xbit_r56_c130 bl_130 br_130 wl_56 vdd gnd cell_6t
Xbit_r57_c130 bl_130 br_130 wl_57 vdd gnd cell_6t
Xbit_r58_c130 bl_130 br_130 wl_58 vdd gnd cell_6t
Xbit_r59_c130 bl_130 br_130 wl_59 vdd gnd cell_6t
Xbit_r60_c130 bl_130 br_130 wl_60 vdd gnd cell_6t
Xbit_r61_c130 bl_130 br_130 wl_61 vdd gnd cell_6t
Xbit_r62_c130 bl_130 br_130 wl_62 vdd gnd cell_6t
Xbit_r63_c130 bl_130 br_130 wl_63 vdd gnd cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd cell_6t
Xbit_r1_c131 bl_131 br_131 wl_1 vdd gnd cell_6t
Xbit_r2_c131 bl_131 br_131 wl_2 vdd gnd cell_6t
Xbit_r3_c131 bl_131 br_131 wl_3 vdd gnd cell_6t
Xbit_r4_c131 bl_131 br_131 wl_4 vdd gnd cell_6t
Xbit_r5_c131 bl_131 br_131 wl_5 vdd gnd cell_6t
Xbit_r6_c131 bl_131 br_131 wl_6 vdd gnd cell_6t
Xbit_r7_c131 bl_131 br_131 wl_7 vdd gnd cell_6t
Xbit_r8_c131 bl_131 br_131 wl_8 vdd gnd cell_6t
Xbit_r9_c131 bl_131 br_131 wl_9 vdd gnd cell_6t
Xbit_r10_c131 bl_131 br_131 wl_10 vdd gnd cell_6t
Xbit_r11_c131 bl_131 br_131 wl_11 vdd gnd cell_6t
Xbit_r12_c131 bl_131 br_131 wl_12 vdd gnd cell_6t
Xbit_r13_c131 bl_131 br_131 wl_13 vdd gnd cell_6t
Xbit_r14_c131 bl_131 br_131 wl_14 vdd gnd cell_6t
Xbit_r15_c131 bl_131 br_131 wl_15 vdd gnd cell_6t
Xbit_r16_c131 bl_131 br_131 wl_16 vdd gnd cell_6t
Xbit_r17_c131 bl_131 br_131 wl_17 vdd gnd cell_6t
Xbit_r18_c131 bl_131 br_131 wl_18 vdd gnd cell_6t
Xbit_r19_c131 bl_131 br_131 wl_19 vdd gnd cell_6t
Xbit_r20_c131 bl_131 br_131 wl_20 vdd gnd cell_6t
Xbit_r21_c131 bl_131 br_131 wl_21 vdd gnd cell_6t
Xbit_r22_c131 bl_131 br_131 wl_22 vdd gnd cell_6t
Xbit_r23_c131 bl_131 br_131 wl_23 vdd gnd cell_6t
Xbit_r24_c131 bl_131 br_131 wl_24 vdd gnd cell_6t
Xbit_r25_c131 bl_131 br_131 wl_25 vdd gnd cell_6t
Xbit_r26_c131 bl_131 br_131 wl_26 vdd gnd cell_6t
Xbit_r27_c131 bl_131 br_131 wl_27 vdd gnd cell_6t
Xbit_r28_c131 bl_131 br_131 wl_28 vdd gnd cell_6t
Xbit_r29_c131 bl_131 br_131 wl_29 vdd gnd cell_6t
Xbit_r30_c131 bl_131 br_131 wl_30 vdd gnd cell_6t
Xbit_r31_c131 bl_131 br_131 wl_31 vdd gnd cell_6t
Xbit_r32_c131 bl_131 br_131 wl_32 vdd gnd cell_6t
Xbit_r33_c131 bl_131 br_131 wl_33 vdd gnd cell_6t
Xbit_r34_c131 bl_131 br_131 wl_34 vdd gnd cell_6t
Xbit_r35_c131 bl_131 br_131 wl_35 vdd gnd cell_6t
Xbit_r36_c131 bl_131 br_131 wl_36 vdd gnd cell_6t
Xbit_r37_c131 bl_131 br_131 wl_37 vdd gnd cell_6t
Xbit_r38_c131 bl_131 br_131 wl_38 vdd gnd cell_6t
Xbit_r39_c131 bl_131 br_131 wl_39 vdd gnd cell_6t
Xbit_r40_c131 bl_131 br_131 wl_40 vdd gnd cell_6t
Xbit_r41_c131 bl_131 br_131 wl_41 vdd gnd cell_6t
Xbit_r42_c131 bl_131 br_131 wl_42 vdd gnd cell_6t
Xbit_r43_c131 bl_131 br_131 wl_43 vdd gnd cell_6t
Xbit_r44_c131 bl_131 br_131 wl_44 vdd gnd cell_6t
Xbit_r45_c131 bl_131 br_131 wl_45 vdd gnd cell_6t
Xbit_r46_c131 bl_131 br_131 wl_46 vdd gnd cell_6t
Xbit_r47_c131 bl_131 br_131 wl_47 vdd gnd cell_6t
Xbit_r48_c131 bl_131 br_131 wl_48 vdd gnd cell_6t
Xbit_r49_c131 bl_131 br_131 wl_49 vdd gnd cell_6t
Xbit_r50_c131 bl_131 br_131 wl_50 vdd gnd cell_6t
Xbit_r51_c131 bl_131 br_131 wl_51 vdd gnd cell_6t
Xbit_r52_c131 bl_131 br_131 wl_52 vdd gnd cell_6t
Xbit_r53_c131 bl_131 br_131 wl_53 vdd gnd cell_6t
Xbit_r54_c131 bl_131 br_131 wl_54 vdd gnd cell_6t
Xbit_r55_c131 bl_131 br_131 wl_55 vdd gnd cell_6t
Xbit_r56_c131 bl_131 br_131 wl_56 vdd gnd cell_6t
Xbit_r57_c131 bl_131 br_131 wl_57 vdd gnd cell_6t
Xbit_r58_c131 bl_131 br_131 wl_58 vdd gnd cell_6t
Xbit_r59_c131 bl_131 br_131 wl_59 vdd gnd cell_6t
Xbit_r60_c131 bl_131 br_131 wl_60 vdd gnd cell_6t
Xbit_r61_c131 bl_131 br_131 wl_61 vdd gnd cell_6t
Xbit_r62_c131 bl_131 br_131 wl_62 vdd gnd cell_6t
Xbit_r63_c131 bl_131 br_131 wl_63 vdd gnd cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd cell_6t
Xbit_r1_c132 bl_132 br_132 wl_1 vdd gnd cell_6t
Xbit_r2_c132 bl_132 br_132 wl_2 vdd gnd cell_6t
Xbit_r3_c132 bl_132 br_132 wl_3 vdd gnd cell_6t
Xbit_r4_c132 bl_132 br_132 wl_4 vdd gnd cell_6t
Xbit_r5_c132 bl_132 br_132 wl_5 vdd gnd cell_6t
Xbit_r6_c132 bl_132 br_132 wl_6 vdd gnd cell_6t
Xbit_r7_c132 bl_132 br_132 wl_7 vdd gnd cell_6t
Xbit_r8_c132 bl_132 br_132 wl_8 vdd gnd cell_6t
Xbit_r9_c132 bl_132 br_132 wl_9 vdd gnd cell_6t
Xbit_r10_c132 bl_132 br_132 wl_10 vdd gnd cell_6t
Xbit_r11_c132 bl_132 br_132 wl_11 vdd gnd cell_6t
Xbit_r12_c132 bl_132 br_132 wl_12 vdd gnd cell_6t
Xbit_r13_c132 bl_132 br_132 wl_13 vdd gnd cell_6t
Xbit_r14_c132 bl_132 br_132 wl_14 vdd gnd cell_6t
Xbit_r15_c132 bl_132 br_132 wl_15 vdd gnd cell_6t
Xbit_r16_c132 bl_132 br_132 wl_16 vdd gnd cell_6t
Xbit_r17_c132 bl_132 br_132 wl_17 vdd gnd cell_6t
Xbit_r18_c132 bl_132 br_132 wl_18 vdd gnd cell_6t
Xbit_r19_c132 bl_132 br_132 wl_19 vdd gnd cell_6t
Xbit_r20_c132 bl_132 br_132 wl_20 vdd gnd cell_6t
Xbit_r21_c132 bl_132 br_132 wl_21 vdd gnd cell_6t
Xbit_r22_c132 bl_132 br_132 wl_22 vdd gnd cell_6t
Xbit_r23_c132 bl_132 br_132 wl_23 vdd gnd cell_6t
Xbit_r24_c132 bl_132 br_132 wl_24 vdd gnd cell_6t
Xbit_r25_c132 bl_132 br_132 wl_25 vdd gnd cell_6t
Xbit_r26_c132 bl_132 br_132 wl_26 vdd gnd cell_6t
Xbit_r27_c132 bl_132 br_132 wl_27 vdd gnd cell_6t
Xbit_r28_c132 bl_132 br_132 wl_28 vdd gnd cell_6t
Xbit_r29_c132 bl_132 br_132 wl_29 vdd gnd cell_6t
Xbit_r30_c132 bl_132 br_132 wl_30 vdd gnd cell_6t
Xbit_r31_c132 bl_132 br_132 wl_31 vdd gnd cell_6t
Xbit_r32_c132 bl_132 br_132 wl_32 vdd gnd cell_6t
Xbit_r33_c132 bl_132 br_132 wl_33 vdd gnd cell_6t
Xbit_r34_c132 bl_132 br_132 wl_34 vdd gnd cell_6t
Xbit_r35_c132 bl_132 br_132 wl_35 vdd gnd cell_6t
Xbit_r36_c132 bl_132 br_132 wl_36 vdd gnd cell_6t
Xbit_r37_c132 bl_132 br_132 wl_37 vdd gnd cell_6t
Xbit_r38_c132 bl_132 br_132 wl_38 vdd gnd cell_6t
Xbit_r39_c132 bl_132 br_132 wl_39 vdd gnd cell_6t
Xbit_r40_c132 bl_132 br_132 wl_40 vdd gnd cell_6t
Xbit_r41_c132 bl_132 br_132 wl_41 vdd gnd cell_6t
Xbit_r42_c132 bl_132 br_132 wl_42 vdd gnd cell_6t
Xbit_r43_c132 bl_132 br_132 wl_43 vdd gnd cell_6t
Xbit_r44_c132 bl_132 br_132 wl_44 vdd gnd cell_6t
Xbit_r45_c132 bl_132 br_132 wl_45 vdd gnd cell_6t
Xbit_r46_c132 bl_132 br_132 wl_46 vdd gnd cell_6t
Xbit_r47_c132 bl_132 br_132 wl_47 vdd gnd cell_6t
Xbit_r48_c132 bl_132 br_132 wl_48 vdd gnd cell_6t
Xbit_r49_c132 bl_132 br_132 wl_49 vdd gnd cell_6t
Xbit_r50_c132 bl_132 br_132 wl_50 vdd gnd cell_6t
Xbit_r51_c132 bl_132 br_132 wl_51 vdd gnd cell_6t
Xbit_r52_c132 bl_132 br_132 wl_52 vdd gnd cell_6t
Xbit_r53_c132 bl_132 br_132 wl_53 vdd gnd cell_6t
Xbit_r54_c132 bl_132 br_132 wl_54 vdd gnd cell_6t
Xbit_r55_c132 bl_132 br_132 wl_55 vdd gnd cell_6t
Xbit_r56_c132 bl_132 br_132 wl_56 vdd gnd cell_6t
Xbit_r57_c132 bl_132 br_132 wl_57 vdd gnd cell_6t
Xbit_r58_c132 bl_132 br_132 wl_58 vdd gnd cell_6t
Xbit_r59_c132 bl_132 br_132 wl_59 vdd gnd cell_6t
Xbit_r60_c132 bl_132 br_132 wl_60 vdd gnd cell_6t
Xbit_r61_c132 bl_132 br_132 wl_61 vdd gnd cell_6t
Xbit_r62_c132 bl_132 br_132 wl_62 vdd gnd cell_6t
Xbit_r63_c132 bl_132 br_132 wl_63 vdd gnd cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd cell_6t
Xbit_r1_c133 bl_133 br_133 wl_1 vdd gnd cell_6t
Xbit_r2_c133 bl_133 br_133 wl_2 vdd gnd cell_6t
Xbit_r3_c133 bl_133 br_133 wl_3 vdd gnd cell_6t
Xbit_r4_c133 bl_133 br_133 wl_4 vdd gnd cell_6t
Xbit_r5_c133 bl_133 br_133 wl_5 vdd gnd cell_6t
Xbit_r6_c133 bl_133 br_133 wl_6 vdd gnd cell_6t
Xbit_r7_c133 bl_133 br_133 wl_7 vdd gnd cell_6t
Xbit_r8_c133 bl_133 br_133 wl_8 vdd gnd cell_6t
Xbit_r9_c133 bl_133 br_133 wl_9 vdd gnd cell_6t
Xbit_r10_c133 bl_133 br_133 wl_10 vdd gnd cell_6t
Xbit_r11_c133 bl_133 br_133 wl_11 vdd gnd cell_6t
Xbit_r12_c133 bl_133 br_133 wl_12 vdd gnd cell_6t
Xbit_r13_c133 bl_133 br_133 wl_13 vdd gnd cell_6t
Xbit_r14_c133 bl_133 br_133 wl_14 vdd gnd cell_6t
Xbit_r15_c133 bl_133 br_133 wl_15 vdd gnd cell_6t
Xbit_r16_c133 bl_133 br_133 wl_16 vdd gnd cell_6t
Xbit_r17_c133 bl_133 br_133 wl_17 vdd gnd cell_6t
Xbit_r18_c133 bl_133 br_133 wl_18 vdd gnd cell_6t
Xbit_r19_c133 bl_133 br_133 wl_19 vdd gnd cell_6t
Xbit_r20_c133 bl_133 br_133 wl_20 vdd gnd cell_6t
Xbit_r21_c133 bl_133 br_133 wl_21 vdd gnd cell_6t
Xbit_r22_c133 bl_133 br_133 wl_22 vdd gnd cell_6t
Xbit_r23_c133 bl_133 br_133 wl_23 vdd gnd cell_6t
Xbit_r24_c133 bl_133 br_133 wl_24 vdd gnd cell_6t
Xbit_r25_c133 bl_133 br_133 wl_25 vdd gnd cell_6t
Xbit_r26_c133 bl_133 br_133 wl_26 vdd gnd cell_6t
Xbit_r27_c133 bl_133 br_133 wl_27 vdd gnd cell_6t
Xbit_r28_c133 bl_133 br_133 wl_28 vdd gnd cell_6t
Xbit_r29_c133 bl_133 br_133 wl_29 vdd gnd cell_6t
Xbit_r30_c133 bl_133 br_133 wl_30 vdd gnd cell_6t
Xbit_r31_c133 bl_133 br_133 wl_31 vdd gnd cell_6t
Xbit_r32_c133 bl_133 br_133 wl_32 vdd gnd cell_6t
Xbit_r33_c133 bl_133 br_133 wl_33 vdd gnd cell_6t
Xbit_r34_c133 bl_133 br_133 wl_34 vdd gnd cell_6t
Xbit_r35_c133 bl_133 br_133 wl_35 vdd gnd cell_6t
Xbit_r36_c133 bl_133 br_133 wl_36 vdd gnd cell_6t
Xbit_r37_c133 bl_133 br_133 wl_37 vdd gnd cell_6t
Xbit_r38_c133 bl_133 br_133 wl_38 vdd gnd cell_6t
Xbit_r39_c133 bl_133 br_133 wl_39 vdd gnd cell_6t
Xbit_r40_c133 bl_133 br_133 wl_40 vdd gnd cell_6t
Xbit_r41_c133 bl_133 br_133 wl_41 vdd gnd cell_6t
Xbit_r42_c133 bl_133 br_133 wl_42 vdd gnd cell_6t
Xbit_r43_c133 bl_133 br_133 wl_43 vdd gnd cell_6t
Xbit_r44_c133 bl_133 br_133 wl_44 vdd gnd cell_6t
Xbit_r45_c133 bl_133 br_133 wl_45 vdd gnd cell_6t
Xbit_r46_c133 bl_133 br_133 wl_46 vdd gnd cell_6t
Xbit_r47_c133 bl_133 br_133 wl_47 vdd gnd cell_6t
Xbit_r48_c133 bl_133 br_133 wl_48 vdd gnd cell_6t
Xbit_r49_c133 bl_133 br_133 wl_49 vdd gnd cell_6t
Xbit_r50_c133 bl_133 br_133 wl_50 vdd gnd cell_6t
Xbit_r51_c133 bl_133 br_133 wl_51 vdd gnd cell_6t
Xbit_r52_c133 bl_133 br_133 wl_52 vdd gnd cell_6t
Xbit_r53_c133 bl_133 br_133 wl_53 vdd gnd cell_6t
Xbit_r54_c133 bl_133 br_133 wl_54 vdd gnd cell_6t
Xbit_r55_c133 bl_133 br_133 wl_55 vdd gnd cell_6t
Xbit_r56_c133 bl_133 br_133 wl_56 vdd gnd cell_6t
Xbit_r57_c133 bl_133 br_133 wl_57 vdd gnd cell_6t
Xbit_r58_c133 bl_133 br_133 wl_58 vdd gnd cell_6t
Xbit_r59_c133 bl_133 br_133 wl_59 vdd gnd cell_6t
Xbit_r60_c133 bl_133 br_133 wl_60 vdd gnd cell_6t
Xbit_r61_c133 bl_133 br_133 wl_61 vdd gnd cell_6t
Xbit_r62_c133 bl_133 br_133 wl_62 vdd gnd cell_6t
Xbit_r63_c133 bl_133 br_133 wl_63 vdd gnd cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd cell_6t
Xbit_r1_c134 bl_134 br_134 wl_1 vdd gnd cell_6t
Xbit_r2_c134 bl_134 br_134 wl_2 vdd gnd cell_6t
Xbit_r3_c134 bl_134 br_134 wl_3 vdd gnd cell_6t
Xbit_r4_c134 bl_134 br_134 wl_4 vdd gnd cell_6t
Xbit_r5_c134 bl_134 br_134 wl_5 vdd gnd cell_6t
Xbit_r6_c134 bl_134 br_134 wl_6 vdd gnd cell_6t
Xbit_r7_c134 bl_134 br_134 wl_7 vdd gnd cell_6t
Xbit_r8_c134 bl_134 br_134 wl_8 vdd gnd cell_6t
Xbit_r9_c134 bl_134 br_134 wl_9 vdd gnd cell_6t
Xbit_r10_c134 bl_134 br_134 wl_10 vdd gnd cell_6t
Xbit_r11_c134 bl_134 br_134 wl_11 vdd gnd cell_6t
Xbit_r12_c134 bl_134 br_134 wl_12 vdd gnd cell_6t
Xbit_r13_c134 bl_134 br_134 wl_13 vdd gnd cell_6t
Xbit_r14_c134 bl_134 br_134 wl_14 vdd gnd cell_6t
Xbit_r15_c134 bl_134 br_134 wl_15 vdd gnd cell_6t
Xbit_r16_c134 bl_134 br_134 wl_16 vdd gnd cell_6t
Xbit_r17_c134 bl_134 br_134 wl_17 vdd gnd cell_6t
Xbit_r18_c134 bl_134 br_134 wl_18 vdd gnd cell_6t
Xbit_r19_c134 bl_134 br_134 wl_19 vdd gnd cell_6t
Xbit_r20_c134 bl_134 br_134 wl_20 vdd gnd cell_6t
Xbit_r21_c134 bl_134 br_134 wl_21 vdd gnd cell_6t
Xbit_r22_c134 bl_134 br_134 wl_22 vdd gnd cell_6t
Xbit_r23_c134 bl_134 br_134 wl_23 vdd gnd cell_6t
Xbit_r24_c134 bl_134 br_134 wl_24 vdd gnd cell_6t
Xbit_r25_c134 bl_134 br_134 wl_25 vdd gnd cell_6t
Xbit_r26_c134 bl_134 br_134 wl_26 vdd gnd cell_6t
Xbit_r27_c134 bl_134 br_134 wl_27 vdd gnd cell_6t
Xbit_r28_c134 bl_134 br_134 wl_28 vdd gnd cell_6t
Xbit_r29_c134 bl_134 br_134 wl_29 vdd gnd cell_6t
Xbit_r30_c134 bl_134 br_134 wl_30 vdd gnd cell_6t
Xbit_r31_c134 bl_134 br_134 wl_31 vdd gnd cell_6t
Xbit_r32_c134 bl_134 br_134 wl_32 vdd gnd cell_6t
Xbit_r33_c134 bl_134 br_134 wl_33 vdd gnd cell_6t
Xbit_r34_c134 bl_134 br_134 wl_34 vdd gnd cell_6t
Xbit_r35_c134 bl_134 br_134 wl_35 vdd gnd cell_6t
Xbit_r36_c134 bl_134 br_134 wl_36 vdd gnd cell_6t
Xbit_r37_c134 bl_134 br_134 wl_37 vdd gnd cell_6t
Xbit_r38_c134 bl_134 br_134 wl_38 vdd gnd cell_6t
Xbit_r39_c134 bl_134 br_134 wl_39 vdd gnd cell_6t
Xbit_r40_c134 bl_134 br_134 wl_40 vdd gnd cell_6t
Xbit_r41_c134 bl_134 br_134 wl_41 vdd gnd cell_6t
Xbit_r42_c134 bl_134 br_134 wl_42 vdd gnd cell_6t
Xbit_r43_c134 bl_134 br_134 wl_43 vdd gnd cell_6t
Xbit_r44_c134 bl_134 br_134 wl_44 vdd gnd cell_6t
Xbit_r45_c134 bl_134 br_134 wl_45 vdd gnd cell_6t
Xbit_r46_c134 bl_134 br_134 wl_46 vdd gnd cell_6t
Xbit_r47_c134 bl_134 br_134 wl_47 vdd gnd cell_6t
Xbit_r48_c134 bl_134 br_134 wl_48 vdd gnd cell_6t
Xbit_r49_c134 bl_134 br_134 wl_49 vdd gnd cell_6t
Xbit_r50_c134 bl_134 br_134 wl_50 vdd gnd cell_6t
Xbit_r51_c134 bl_134 br_134 wl_51 vdd gnd cell_6t
Xbit_r52_c134 bl_134 br_134 wl_52 vdd gnd cell_6t
Xbit_r53_c134 bl_134 br_134 wl_53 vdd gnd cell_6t
Xbit_r54_c134 bl_134 br_134 wl_54 vdd gnd cell_6t
Xbit_r55_c134 bl_134 br_134 wl_55 vdd gnd cell_6t
Xbit_r56_c134 bl_134 br_134 wl_56 vdd gnd cell_6t
Xbit_r57_c134 bl_134 br_134 wl_57 vdd gnd cell_6t
Xbit_r58_c134 bl_134 br_134 wl_58 vdd gnd cell_6t
Xbit_r59_c134 bl_134 br_134 wl_59 vdd gnd cell_6t
Xbit_r60_c134 bl_134 br_134 wl_60 vdd gnd cell_6t
Xbit_r61_c134 bl_134 br_134 wl_61 vdd gnd cell_6t
Xbit_r62_c134 bl_134 br_134 wl_62 vdd gnd cell_6t
Xbit_r63_c134 bl_134 br_134 wl_63 vdd gnd cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd cell_6t
Xbit_r1_c135 bl_135 br_135 wl_1 vdd gnd cell_6t
Xbit_r2_c135 bl_135 br_135 wl_2 vdd gnd cell_6t
Xbit_r3_c135 bl_135 br_135 wl_3 vdd gnd cell_6t
Xbit_r4_c135 bl_135 br_135 wl_4 vdd gnd cell_6t
Xbit_r5_c135 bl_135 br_135 wl_5 vdd gnd cell_6t
Xbit_r6_c135 bl_135 br_135 wl_6 vdd gnd cell_6t
Xbit_r7_c135 bl_135 br_135 wl_7 vdd gnd cell_6t
Xbit_r8_c135 bl_135 br_135 wl_8 vdd gnd cell_6t
Xbit_r9_c135 bl_135 br_135 wl_9 vdd gnd cell_6t
Xbit_r10_c135 bl_135 br_135 wl_10 vdd gnd cell_6t
Xbit_r11_c135 bl_135 br_135 wl_11 vdd gnd cell_6t
Xbit_r12_c135 bl_135 br_135 wl_12 vdd gnd cell_6t
Xbit_r13_c135 bl_135 br_135 wl_13 vdd gnd cell_6t
Xbit_r14_c135 bl_135 br_135 wl_14 vdd gnd cell_6t
Xbit_r15_c135 bl_135 br_135 wl_15 vdd gnd cell_6t
Xbit_r16_c135 bl_135 br_135 wl_16 vdd gnd cell_6t
Xbit_r17_c135 bl_135 br_135 wl_17 vdd gnd cell_6t
Xbit_r18_c135 bl_135 br_135 wl_18 vdd gnd cell_6t
Xbit_r19_c135 bl_135 br_135 wl_19 vdd gnd cell_6t
Xbit_r20_c135 bl_135 br_135 wl_20 vdd gnd cell_6t
Xbit_r21_c135 bl_135 br_135 wl_21 vdd gnd cell_6t
Xbit_r22_c135 bl_135 br_135 wl_22 vdd gnd cell_6t
Xbit_r23_c135 bl_135 br_135 wl_23 vdd gnd cell_6t
Xbit_r24_c135 bl_135 br_135 wl_24 vdd gnd cell_6t
Xbit_r25_c135 bl_135 br_135 wl_25 vdd gnd cell_6t
Xbit_r26_c135 bl_135 br_135 wl_26 vdd gnd cell_6t
Xbit_r27_c135 bl_135 br_135 wl_27 vdd gnd cell_6t
Xbit_r28_c135 bl_135 br_135 wl_28 vdd gnd cell_6t
Xbit_r29_c135 bl_135 br_135 wl_29 vdd gnd cell_6t
Xbit_r30_c135 bl_135 br_135 wl_30 vdd gnd cell_6t
Xbit_r31_c135 bl_135 br_135 wl_31 vdd gnd cell_6t
Xbit_r32_c135 bl_135 br_135 wl_32 vdd gnd cell_6t
Xbit_r33_c135 bl_135 br_135 wl_33 vdd gnd cell_6t
Xbit_r34_c135 bl_135 br_135 wl_34 vdd gnd cell_6t
Xbit_r35_c135 bl_135 br_135 wl_35 vdd gnd cell_6t
Xbit_r36_c135 bl_135 br_135 wl_36 vdd gnd cell_6t
Xbit_r37_c135 bl_135 br_135 wl_37 vdd gnd cell_6t
Xbit_r38_c135 bl_135 br_135 wl_38 vdd gnd cell_6t
Xbit_r39_c135 bl_135 br_135 wl_39 vdd gnd cell_6t
Xbit_r40_c135 bl_135 br_135 wl_40 vdd gnd cell_6t
Xbit_r41_c135 bl_135 br_135 wl_41 vdd gnd cell_6t
Xbit_r42_c135 bl_135 br_135 wl_42 vdd gnd cell_6t
Xbit_r43_c135 bl_135 br_135 wl_43 vdd gnd cell_6t
Xbit_r44_c135 bl_135 br_135 wl_44 vdd gnd cell_6t
Xbit_r45_c135 bl_135 br_135 wl_45 vdd gnd cell_6t
Xbit_r46_c135 bl_135 br_135 wl_46 vdd gnd cell_6t
Xbit_r47_c135 bl_135 br_135 wl_47 vdd gnd cell_6t
Xbit_r48_c135 bl_135 br_135 wl_48 vdd gnd cell_6t
Xbit_r49_c135 bl_135 br_135 wl_49 vdd gnd cell_6t
Xbit_r50_c135 bl_135 br_135 wl_50 vdd gnd cell_6t
Xbit_r51_c135 bl_135 br_135 wl_51 vdd gnd cell_6t
Xbit_r52_c135 bl_135 br_135 wl_52 vdd gnd cell_6t
Xbit_r53_c135 bl_135 br_135 wl_53 vdd gnd cell_6t
Xbit_r54_c135 bl_135 br_135 wl_54 vdd gnd cell_6t
Xbit_r55_c135 bl_135 br_135 wl_55 vdd gnd cell_6t
Xbit_r56_c135 bl_135 br_135 wl_56 vdd gnd cell_6t
Xbit_r57_c135 bl_135 br_135 wl_57 vdd gnd cell_6t
Xbit_r58_c135 bl_135 br_135 wl_58 vdd gnd cell_6t
Xbit_r59_c135 bl_135 br_135 wl_59 vdd gnd cell_6t
Xbit_r60_c135 bl_135 br_135 wl_60 vdd gnd cell_6t
Xbit_r61_c135 bl_135 br_135 wl_61 vdd gnd cell_6t
Xbit_r62_c135 bl_135 br_135 wl_62 vdd gnd cell_6t
Xbit_r63_c135 bl_135 br_135 wl_63 vdd gnd cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd cell_6t
Xbit_r1_c136 bl_136 br_136 wl_1 vdd gnd cell_6t
Xbit_r2_c136 bl_136 br_136 wl_2 vdd gnd cell_6t
Xbit_r3_c136 bl_136 br_136 wl_3 vdd gnd cell_6t
Xbit_r4_c136 bl_136 br_136 wl_4 vdd gnd cell_6t
Xbit_r5_c136 bl_136 br_136 wl_5 vdd gnd cell_6t
Xbit_r6_c136 bl_136 br_136 wl_6 vdd gnd cell_6t
Xbit_r7_c136 bl_136 br_136 wl_7 vdd gnd cell_6t
Xbit_r8_c136 bl_136 br_136 wl_8 vdd gnd cell_6t
Xbit_r9_c136 bl_136 br_136 wl_9 vdd gnd cell_6t
Xbit_r10_c136 bl_136 br_136 wl_10 vdd gnd cell_6t
Xbit_r11_c136 bl_136 br_136 wl_11 vdd gnd cell_6t
Xbit_r12_c136 bl_136 br_136 wl_12 vdd gnd cell_6t
Xbit_r13_c136 bl_136 br_136 wl_13 vdd gnd cell_6t
Xbit_r14_c136 bl_136 br_136 wl_14 vdd gnd cell_6t
Xbit_r15_c136 bl_136 br_136 wl_15 vdd gnd cell_6t
Xbit_r16_c136 bl_136 br_136 wl_16 vdd gnd cell_6t
Xbit_r17_c136 bl_136 br_136 wl_17 vdd gnd cell_6t
Xbit_r18_c136 bl_136 br_136 wl_18 vdd gnd cell_6t
Xbit_r19_c136 bl_136 br_136 wl_19 vdd gnd cell_6t
Xbit_r20_c136 bl_136 br_136 wl_20 vdd gnd cell_6t
Xbit_r21_c136 bl_136 br_136 wl_21 vdd gnd cell_6t
Xbit_r22_c136 bl_136 br_136 wl_22 vdd gnd cell_6t
Xbit_r23_c136 bl_136 br_136 wl_23 vdd gnd cell_6t
Xbit_r24_c136 bl_136 br_136 wl_24 vdd gnd cell_6t
Xbit_r25_c136 bl_136 br_136 wl_25 vdd gnd cell_6t
Xbit_r26_c136 bl_136 br_136 wl_26 vdd gnd cell_6t
Xbit_r27_c136 bl_136 br_136 wl_27 vdd gnd cell_6t
Xbit_r28_c136 bl_136 br_136 wl_28 vdd gnd cell_6t
Xbit_r29_c136 bl_136 br_136 wl_29 vdd gnd cell_6t
Xbit_r30_c136 bl_136 br_136 wl_30 vdd gnd cell_6t
Xbit_r31_c136 bl_136 br_136 wl_31 vdd gnd cell_6t
Xbit_r32_c136 bl_136 br_136 wl_32 vdd gnd cell_6t
Xbit_r33_c136 bl_136 br_136 wl_33 vdd gnd cell_6t
Xbit_r34_c136 bl_136 br_136 wl_34 vdd gnd cell_6t
Xbit_r35_c136 bl_136 br_136 wl_35 vdd gnd cell_6t
Xbit_r36_c136 bl_136 br_136 wl_36 vdd gnd cell_6t
Xbit_r37_c136 bl_136 br_136 wl_37 vdd gnd cell_6t
Xbit_r38_c136 bl_136 br_136 wl_38 vdd gnd cell_6t
Xbit_r39_c136 bl_136 br_136 wl_39 vdd gnd cell_6t
Xbit_r40_c136 bl_136 br_136 wl_40 vdd gnd cell_6t
Xbit_r41_c136 bl_136 br_136 wl_41 vdd gnd cell_6t
Xbit_r42_c136 bl_136 br_136 wl_42 vdd gnd cell_6t
Xbit_r43_c136 bl_136 br_136 wl_43 vdd gnd cell_6t
Xbit_r44_c136 bl_136 br_136 wl_44 vdd gnd cell_6t
Xbit_r45_c136 bl_136 br_136 wl_45 vdd gnd cell_6t
Xbit_r46_c136 bl_136 br_136 wl_46 vdd gnd cell_6t
Xbit_r47_c136 bl_136 br_136 wl_47 vdd gnd cell_6t
Xbit_r48_c136 bl_136 br_136 wl_48 vdd gnd cell_6t
Xbit_r49_c136 bl_136 br_136 wl_49 vdd gnd cell_6t
Xbit_r50_c136 bl_136 br_136 wl_50 vdd gnd cell_6t
Xbit_r51_c136 bl_136 br_136 wl_51 vdd gnd cell_6t
Xbit_r52_c136 bl_136 br_136 wl_52 vdd gnd cell_6t
Xbit_r53_c136 bl_136 br_136 wl_53 vdd gnd cell_6t
Xbit_r54_c136 bl_136 br_136 wl_54 vdd gnd cell_6t
Xbit_r55_c136 bl_136 br_136 wl_55 vdd gnd cell_6t
Xbit_r56_c136 bl_136 br_136 wl_56 vdd gnd cell_6t
Xbit_r57_c136 bl_136 br_136 wl_57 vdd gnd cell_6t
Xbit_r58_c136 bl_136 br_136 wl_58 vdd gnd cell_6t
Xbit_r59_c136 bl_136 br_136 wl_59 vdd gnd cell_6t
Xbit_r60_c136 bl_136 br_136 wl_60 vdd gnd cell_6t
Xbit_r61_c136 bl_136 br_136 wl_61 vdd gnd cell_6t
Xbit_r62_c136 bl_136 br_136 wl_62 vdd gnd cell_6t
Xbit_r63_c136 bl_136 br_136 wl_63 vdd gnd cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd cell_6t
Xbit_r1_c137 bl_137 br_137 wl_1 vdd gnd cell_6t
Xbit_r2_c137 bl_137 br_137 wl_2 vdd gnd cell_6t
Xbit_r3_c137 bl_137 br_137 wl_3 vdd gnd cell_6t
Xbit_r4_c137 bl_137 br_137 wl_4 vdd gnd cell_6t
Xbit_r5_c137 bl_137 br_137 wl_5 vdd gnd cell_6t
Xbit_r6_c137 bl_137 br_137 wl_6 vdd gnd cell_6t
Xbit_r7_c137 bl_137 br_137 wl_7 vdd gnd cell_6t
Xbit_r8_c137 bl_137 br_137 wl_8 vdd gnd cell_6t
Xbit_r9_c137 bl_137 br_137 wl_9 vdd gnd cell_6t
Xbit_r10_c137 bl_137 br_137 wl_10 vdd gnd cell_6t
Xbit_r11_c137 bl_137 br_137 wl_11 vdd gnd cell_6t
Xbit_r12_c137 bl_137 br_137 wl_12 vdd gnd cell_6t
Xbit_r13_c137 bl_137 br_137 wl_13 vdd gnd cell_6t
Xbit_r14_c137 bl_137 br_137 wl_14 vdd gnd cell_6t
Xbit_r15_c137 bl_137 br_137 wl_15 vdd gnd cell_6t
Xbit_r16_c137 bl_137 br_137 wl_16 vdd gnd cell_6t
Xbit_r17_c137 bl_137 br_137 wl_17 vdd gnd cell_6t
Xbit_r18_c137 bl_137 br_137 wl_18 vdd gnd cell_6t
Xbit_r19_c137 bl_137 br_137 wl_19 vdd gnd cell_6t
Xbit_r20_c137 bl_137 br_137 wl_20 vdd gnd cell_6t
Xbit_r21_c137 bl_137 br_137 wl_21 vdd gnd cell_6t
Xbit_r22_c137 bl_137 br_137 wl_22 vdd gnd cell_6t
Xbit_r23_c137 bl_137 br_137 wl_23 vdd gnd cell_6t
Xbit_r24_c137 bl_137 br_137 wl_24 vdd gnd cell_6t
Xbit_r25_c137 bl_137 br_137 wl_25 vdd gnd cell_6t
Xbit_r26_c137 bl_137 br_137 wl_26 vdd gnd cell_6t
Xbit_r27_c137 bl_137 br_137 wl_27 vdd gnd cell_6t
Xbit_r28_c137 bl_137 br_137 wl_28 vdd gnd cell_6t
Xbit_r29_c137 bl_137 br_137 wl_29 vdd gnd cell_6t
Xbit_r30_c137 bl_137 br_137 wl_30 vdd gnd cell_6t
Xbit_r31_c137 bl_137 br_137 wl_31 vdd gnd cell_6t
Xbit_r32_c137 bl_137 br_137 wl_32 vdd gnd cell_6t
Xbit_r33_c137 bl_137 br_137 wl_33 vdd gnd cell_6t
Xbit_r34_c137 bl_137 br_137 wl_34 vdd gnd cell_6t
Xbit_r35_c137 bl_137 br_137 wl_35 vdd gnd cell_6t
Xbit_r36_c137 bl_137 br_137 wl_36 vdd gnd cell_6t
Xbit_r37_c137 bl_137 br_137 wl_37 vdd gnd cell_6t
Xbit_r38_c137 bl_137 br_137 wl_38 vdd gnd cell_6t
Xbit_r39_c137 bl_137 br_137 wl_39 vdd gnd cell_6t
Xbit_r40_c137 bl_137 br_137 wl_40 vdd gnd cell_6t
Xbit_r41_c137 bl_137 br_137 wl_41 vdd gnd cell_6t
Xbit_r42_c137 bl_137 br_137 wl_42 vdd gnd cell_6t
Xbit_r43_c137 bl_137 br_137 wl_43 vdd gnd cell_6t
Xbit_r44_c137 bl_137 br_137 wl_44 vdd gnd cell_6t
Xbit_r45_c137 bl_137 br_137 wl_45 vdd gnd cell_6t
Xbit_r46_c137 bl_137 br_137 wl_46 vdd gnd cell_6t
Xbit_r47_c137 bl_137 br_137 wl_47 vdd gnd cell_6t
Xbit_r48_c137 bl_137 br_137 wl_48 vdd gnd cell_6t
Xbit_r49_c137 bl_137 br_137 wl_49 vdd gnd cell_6t
Xbit_r50_c137 bl_137 br_137 wl_50 vdd gnd cell_6t
Xbit_r51_c137 bl_137 br_137 wl_51 vdd gnd cell_6t
Xbit_r52_c137 bl_137 br_137 wl_52 vdd gnd cell_6t
Xbit_r53_c137 bl_137 br_137 wl_53 vdd gnd cell_6t
Xbit_r54_c137 bl_137 br_137 wl_54 vdd gnd cell_6t
Xbit_r55_c137 bl_137 br_137 wl_55 vdd gnd cell_6t
Xbit_r56_c137 bl_137 br_137 wl_56 vdd gnd cell_6t
Xbit_r57_c137 bl_137 br_137 wl_57 vdd gnd cell_6t
Xbit_r58_c137 bl_137 br_137 wl_58 vdd gnd cell_6t
Xbit_r59_c137 bl_137 br_137 wl_59 vdd gnd cell_6t
Xbit_r60_c137 bl_137 br_137 wl_60 vdd gnd cell_6t
Xbit_r61_c137 bl_137 br_137 wl_61 vdd gnd cell_6t
Xbit_r62_c137 bl_137 br_137 wl_62 vdd gnd cell_6t
Xbit_r63_c137 bl_137 br_137 wl_63 vdd gnd cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd cell_6t
Xbit_r1_c138 bl_138 br_138 wl_1 vdd gnd cell_6t
Xbit_r2_c138 bl_138 br_138 wl_2 vdd gnd cell_6t
Xbit_r3_c138 bl_138 br_138 wl_3 vdd gnd cell_6t
Xbit_r4_c138 bl_138 br_138 wl_4 vdd gnd cell_6t
Xbit_r5_c138 bl_138 br_138 wl_5 vdd gnd cell_6t
Xbit_r6_c138 bl_138 br_138 wl_6 vdd gnd cell_6t
Xbit_r7_c138 bl_138 br_138 wl_7 vdd gnd cell_6t
Xbit_r8_c138 bl_138 br_138 wl_8 vdd gnd cell_6t
Xbit_r9_c138 bl_138 br_138 wl_9 vdd gnd cell_6t
Xbit_r10_c138 bl_138 br_138 wl_10 vdd gnd cell_6t
Xbit_r11_c138 bl_138 br_138 wl_11 vdd gnd cell_6t
Xbit_r12_c138 bl_138 br_138 wl_12 vdd gnd cell_6t
Xbit_r13_c138 bl_138 br_138 wl_13 vdd gnd cell_6t
Xbit_r14_c138 bl_138 br_138 wl_14 vdd gnd cell_6t
Xbit_r15_c138 bl_138 br_138 wl_15 vdd gnd cell_6t
Xbit_r16_c138 bl_138 br_138 wl_16 vdd gnd cell_6t
Xbit_r17_c138 bl_138 br_138 wl_17 vdd gnd cell_6t
Xbit_r18_c138 bl_138 br_138 wl_18 vdd gnd cell_6t
Xbit_r19_c138 bl_138 br_138 wl_19 vdd gnd cell_6t
Xbit_r20_c138 bl_138 br_138 wl_20 vdd gnd cell_6t
Xbit_r21_c138 bl_138 br_138 wl_21 vdd gnd cell_6t
Xbit_r22_c138 bl_138 br_138 wl_22 vdd gnd cell_6t
Xbit_r23_c138 bl_138 br_138 wl_23 vdd gnd cell_6t
Xbit_r24_c138 bl_138 br_138 wl_24 vdd gnd cell_6t
Xbit_r25_c138 bl_138 br_138 wl_25 vdd gnd cell_6t
Xbit_r26_c138 bl_138 br_138 wl_26 vdd gnd cell_6t
Xbit_r27_c138 bl_138 br_138 wl_27 vdd gnd cell_6t
Xbit_r28_c138 bl_138 br_138 wl_28 vdd gnd cell_6t
Xbit_r29_c138 bl_138 br_138 wl_29 vdd gnd cell_6t
Xbit_r30_c138 bl_138 br_138 wl_30 vdd gnd cell_6t
Xbit_r31_c138 bl_138 br_138 wl_31 vdd gnd cell_6t
Xbit_r32_c138 bl_138 br_138 wl_32 vdd gnd cell_6t
Xbit_r33_c138 bl_138 br_138 wl_33 vdd gnd cell_6t
Xbit_r34_c138 bl_138 br_138 wl_34 vdd gnd cell_6t
Xbit_r35_c138 bl_138 br_138 wl_35 vdd gnd cell_6t
Xbit_r36_c138 bl_138 br_138 wl_36 vdd gnd cell_6t
Xbit_r37_c138 bl_138 br_138 wl_37 vdd gnd cell_6t
Xbit_r38_c138 bl_138 br_138 wl_38 vdd gnd cell_6t
Xbit_r39_c138 bl_138 br_138 wl_39 vdd gnd cell_6t
Xbit_r40_c138 bl_138 br_138 wl_40 vdd gnd cell_6t
Xbit_r41_c138 bl_138 br_138 wl_41 vdd gnd cell_6t
Xbit_r42_c138 bl_138 br_138 wl_42 vdd gnd cell_6t
Xbit_r43_c138 bl_138 br_138 wl_43 vdd gnd cell_6t
Xbit_r44_c138 bl_138 br_138 wl_44 vdd gnd cell_6t
Xbit_r45_c138 bl_138 br_138 wl_45 vdd gnd cell_6t
Xbit_r46_c138 bl_138 br_138 wl_46 vdd gnd cell_6t
Xbit_r47_c138 bl_138 br_138 wl_47 vdd gnd cell_6t
Xbit_r48_c138 bl_138 br_138 wl_48 vdd gnd cell_6t
Xbit_r49_c138 bl_138 br_138 wl_49 vdd gnd cell_6t
Xbit_r50_c138 bl_138 br_138 wl_50 vdd gnd cell_6t
Xbit_r51_c138 bl_138 br_138 wl_51 vdd gnd cell_6t
Xbit_r52_c138 bl_138 br_138 wl_52 vdd gnd cell_6t
Xbit_r53_c138 bl_138 br_138 wl_53 vdd gnd cell_6t
Xbit_r54_c138 bl_138 br_138 wl_54 vdd gnd cell_6t
Xbit_r55_c138 bl_138 br_138 wl_55 vdd gnd cell_6t
Xbit_r56_c138 bl_138 br_138 wl_56 vdd gnd cell_6t
Xbit_r57_c138 bl_138 br_138 wl_57 vdd gnd cell_6t
Xbit_r58_c138 bl_138 br_138 wl_58 vdd gnd cell_6t
Xbit_r59_c138 bl_138 br_138 wl_59 vdd gnd cell_6t
Xbit_r60_c138 bl_138 br_138 wl_60 vdd gnd cell_6t
Xbit_r61_c138 bl_138 br_138 wl_61 vdd gnd cell_6t
Xbit_r62_c138 bl_138 br_138 wl_62 vdd gnd cell_6t
Xbit_r63_c138 bl_138 br_138 wl_63 vdd gnd cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd cell_6t
Xbit_r1_c139 bl_139 br_139 wl_1 vdd gnd cell_6t
Xbit_r2_c139 bl_139 br_139 wl_2 vdd gnd cell_6t
Xbit_r3_c139 bl_139 br_139 wl_3 vdd gnd cell_6t
Xbit_r4_c139 bl_139 br_139 wl_4 vdd gnd cell_6t
Xbit_r5_c139 bl_139 br_139 wl_5 vdd gnd cell_6t
Xbit_r6_c139 bl_139 br_139 wl_6 vdd gnd cell_6t
Xbit_r7_c139 bl_139 br_139 wl_7 vdd gnd cell_6t
Xbit_r8_c139 bl_139 br_139 wl_8 vdd gnd cell_6t
Xbit_r9_c139 bl_139 br_139 wl_9 vdd gnd cell_6t
Xbit_r10_c139 bl_139 br_139 wl_10 vdd gnd cell_6t
Xbit_r11_c139 bl_139 br_139 wl_11 vdd gnd cell_6t
Xbit_r12_c139 bl_139 br_139 wl_12 vdd gnd cell_6t
Xbit_r13_c139 bl_139 br_139 wl_13 vdd gnd cell_6t
Xbit_r14_c139 bl_139 br_139 wl_14 vdd gnd cell_6t
Xbit_r15_c139 bl_139 br_139 wl_15 vdd gnd cell_6t
Xbit_r16_c139 bl_139 br_139 wl_16 vdd gnd cell_6t
Xbit_r17_c139 bl_139 br_139 wl_17 vdd gnd cell_6t
Xbit_r18_c139 bl_139 br_139 wl_18 vdd gnd cell_6t
Xbit_r19_c139 bl_139 br_139 wl_19 vdd gnd cell_6t
Xbit_r20_c139 bl_139 br_139 wl_20 vdd gnd cell_6t
Xbit_r21_c139 bl_139 br_139 wl_21 vdd gnd cell_6t
Xbit_r22_c139 bl_139 br_139 wl_22 vdd gnd cell_6t
Xbit_r23_c139 bl_139 br_139 wl_23 vdd gnd cell_6t
Xbit_r24_c139 bl_139 br_139 wl_24 vdd gnd cell_6t
Xbit_r25_c139 bl_139 br_139 wl_25 vdd gnd cell_6t
Xbit_r26_c139 bl_139 br_139 wl_26 vdd gnd cell_6t
Xbit_r27_c139 bl_139 br_139 wl_27 vdd gnd cell_6t
Xbit_r28_c139 bl_139 br_139 wl_28 vdd gnd cell_6t
Xbit_r29_c139 bl_139 br_139 wl_29 vdd gnd cell_6t
Xbit_r30_c139 bl_139 br_139 wl_30 vdd gnd cell_6t
Xbit_r31_c139 bl_139 br_139 wl_31 vdd gnd cell_6t
Xbit_r32_c139 bl_139 br_139 wl_32 vdd gnd cell_6t
Xbit_r33_c139 bl_139 br_139 wl_33 vdd gnd cell_6t
Xbit_r34_c139 bl_139 br_139 wl_34 vdd gnd cell_6t
Xbit_r35_c139 bl_139 br_139 wl_35 vdd gnd cell_6t
Xbit_r36_c139 bl_139 br_139 wl_36 vdd gnd cell_6t
Xbit_r37_c139 bl_139 br_139 wl_37 vdd gnd cell_6t
Xbit_r38_c139 bl_139 br_139 wl_38 vdd gnd cell_6t
Xbit_r39_c139 bl_139 br_139 wl_39 vdd gnd cell_6t
Xbit_r40_c139 bl_139 br_139 wl_40 vdd gnd cell_6t
Xbit_r41_c139 bl_139 br_139 wl_41 vdd gnd cell_6t
Xbit_r42_c139 bl_139 br_139 wl_42 vdd gnd cell_6t
Xbit_r43_c139 bl_139 br_139 wl_43 vdd gnd cell_6t
Xbit_r44_c139 bl_139 br_139 wl_44 vdd gnd cell_6t
Xbit_r45_c139 bl_139 br_139 wl_45 vdd gnd cell_6t
Xbit_r46_c139 bl_139 br_139 wl_46 vdd gnd cell_6t
Xbit_r47_c139 bl_139 br_139 wl_47 vdd gnd cell_6t
Xbit_r48_c139 bl_139 br_139 wl_48 vdd gnd cell_6t
Xbit_r49_c139 bl_139 br_139 wl_49 vdd gnd cell_6t
Xbit_r50_c139 bl_139 br_139 wl_50 vdd gnd cell_6t
Xbit_r51_c139 bl_139 br_139 wl_51 vdd gnd cell_6t
Xbit_r52_c139 bl_139 br_139 wl_52 vdd gnd cell_6t
Xbit_r53_c139 bl_139 br_139 wl_53 vdd gnd cell_6t
Xbit_r54_c139 bl_139 br_139 wl_54 vdd gnd cell_6t
Xbit_r55_c139 bl_139 br_139 wl_55 vdd gnd cell_6t
Xbit_r56_c139 bl_139 br_139 wl_56 vdd gnd cell_6t
Xbit_r57_c139 bl_139 br_139 wl_57 vdd gnd cell_6t
Xbit_r58_c139 bl_139 br_139 wl_58 vdd gnd cell_6t
Xbit_r59_c139 bl_139 br_139 wl_59 vdd gnd cell_6t
Xbit_r60_c139 bl_139 br_139 wl_60 vdd gnd cell_6t
Xbit_r61_c139 bl_139 br_139 wl_61 vdd gnd cell_6t
Xbit_r62_c139 bl_139 br_139 wl_62 vdd gnd cell_6t
Xbit_r63_c139 bl_139 br_139 wl_63 vdd gnd cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd cell_6t
Xbit_r1_c140 bl_140 br_140 wl_1 vdd gnd cell_6t
Xbit_r2_c140 bl_140 br_140 wl_2 vdd gnd cell_6t
Xbit_r3_c140 bl_140 br_140 wl_3 vdd gnd cell_6t
Xbit_r4_c140 bl_140 br_140 wl_4 vdd gnd cell_6t
Xbit_r5_c140 bl_140 br_140 wl_5 vdd gnd cell_6t
Xbit_r6_c140 bl_140 br_140 wl_6 vdd gnd cell_6t
Xbit_r7_c140 bl_140 br_140 wl_7 vdd gnd cell_6t
Xbit_r8_c140 bl_140 br_140 wl_8 vdd gnd cell_6t
Xbit_r9_c140 bl_140 br_140 wl_9 vdd gnd cell_6t
Xbit_r10_c140 bl_140 br_140 wl_10 vdd gnd cell_6t
Xbit_r11_c140 bl_140 br_140 wl_11 vdd gnd cell_6t
Xbit_r12_c140 bl_140 br_140 wl_12 vdd gnd cell_6t
Xbit_r13_c140 bl_140 br_140 wl_13 vdd gnd cell_6t
Xbit_r14_c140 bl_140 br_140 wl_14 vdd gnd cell_6t
Xbit_r15_c140 bl_140 br_140 wl_15 vdd gnd cell_6t
Xbit_r16_c140 bl_140 br_140 wl_16 vdd gnd cell_6t
Xbit_r17_c140 bl_140 br_140 wl_17 vdd gnd cell_6t
Xbit_r18_c140 bl_140 br_140 wl_18 vdd gnd cell_6t
Xbit_r19_c140 bl_140 br_140 wl_19 vdd gnd cell_6t
Xbit_r20_c140 bl_140 br_140 wl_20 vdd gnd cell_6t
Xbit_r21_c140 bl_140 br_140 wl_21 vdd gnd cell_6t
Xbit_r22_c140 bl_140 br_140 wl_22 vdd gnd cell_6t
Xbit_r23_c140 bl_140 br_140 wl_23 vdd gnd cell_6t
Xbit_r24_c140 bl_140 br_140 wl_24 vdd gnd cell_6t
Xbit_r25_c140 bl_140 br_140 wl_25 vdd gnd cell_6t
Xbit_r26_c140 bl_140 br_140 wl_26 vdd gnd cell_6t
Xbit_r27_c140 bl_140 br_140 wl_27 vdd gnd cell_6t
Xbit_r28_c140 bl_140 br_140 wl_28 vdd gnd cell_6t
Xbit_r29_c140 bl_140 br_140 wl_29 vdd gnd cell_6t
Xbit_r30_c140 bl_140 br_140 wl_30 vdd gnd cell_6t
Xbit_r31_c140 bl_140 br_140 wl_31 vdd gnd cell_6t
Xbit_r32_c140 bl_140 br_140 wl_32 vdd gnd cell_6t
Xbit_r33_c140 bl_140 br_140 wl_33 vdd gnd cell_6t
Xbit_r34_c140 bl_140 br_140 wl_34 vdd gnd cell_6t
Xbit_r35_c140 bl_140 br_140 wl_35 vdd gnd cell_6t
Xbit_r36_c140 bl_140 br_140 wl_36 vdd gnd cell_6t
Xbit_r37_c140 bl_140 br_140 wl_37 vdd gnd cell_6t
Xbit_r38_c140 bl_140 br_140 wl_38 vdd gnd cell_6t
Xbit_r39_c140 bl_140 br_140 wl_39 vdd gnd cell_6t
Xbit_r40_c140 bl_140 br_140 wl_40 vdd gnd cell_6t
Xbit_r41_c140 bl_140 br_140 wl_41 vdd gnd cell_6t
Xbit_r42_c140 bl_140 br_140 wl_42 vdd gnd cell_6t
Xbit_r43_c140 bl_140 br_140 wl_43 vdd gnd cell_6t
Xbit_r44_c140 bl_140 br_140 wl_44 vdd gnd cell_6t
Xbit_r45_c140 bl_140 br_140 wl_45 vdd gnd cell_6t
Xbit_r46_c140 bl_140 br_140 wl_46 vdd gnd cell_6t
Xbit_r47_c140 bl_140 br_140 wl_47 vdd gnd cell_6t
Xbit_r48_c140 bl_140 br_140 wl_48 vdd gnd cell_6t
Xbit_r49_c140 bl_140 br_140 wl_49 vdd gnd cell_6t
Xbit_r50_c140 bl_140 br_140 wl_50 vdd gnd cell_6t
Xbit_r51_c140 bl_140 br_140 wl_51 vdd gnd cell_6t
Xbit_r52_c140 bl_140 br_140 wl_52 vdd gnd cell_6t
Xbit_r53_c140 bl_140 br_140 wl_53 vdd gnd cell_6t
Xbit_r54_c140 bl_140 br_140 wl_54 vdd gnd cell_6t
Xbit_r55_c140 bl_140 br_140 wl_55 vdd gnd cell_6t
Xbit_r56_c140 bl_140 br_140 wl_56 vdd gnd cell_6t
Xbit_r57_c140 bl_140 br_140 wl_57 vdd gnd cell_6t
Xbit_r58_c140 bl_140 br_140 wl_58 vdd gnd cell_6t
Xbit_r59_c140 bl_140 br_140 wl_59 vdd gnd cell_6t
Xbit_r60_c140 bl_140 br_140 wl_60 vdd gnd cell_6t
Xbit_r61_c140 bl_140 br_140 wl_61 vdd gnd cell_6t
Xbit_r62_c140 bl_140 br_140 wl_62 vdd gnd cell_6t
Xbit_r63_c140 bl_140 br_140 wl_63 vdd gnd cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd cell_6t
Xbit_r1_c141 bl_141 br_141 wl_1 vdd gnd cell_6t
Xbit_r2_c141 bl_141 br_141 wl_2 vdd gnd cell_6t
Xbit_r3_c141 bl_141 br_141 wl_3 vdd gnd cell_6t
Xbit_r4_c141 bl_141 br_141 wl_4 vdd gnd cell_6t
Xbit_r5_c141 bl_141 br_141 wl_5 vdd gnd cell_6t
Xbit_r6_c141 bl_141 br_141 wl_6 vdd gnd cell_6t
Xbit_r7_c141 bl_141 br_141 wl_7 vdd gnd cell_6t
Xbit_r8_c141 bl_141 br_141 wl_8 vdd gnd cell_6t
Xbit_r9_c141 bl_141 br_141 wl_9 vdd gnd cell_6t
Xbit_r10_c141 bl_141 br_141 wl_10 vdd gnd cell_6t
Xbit_r11_c141 bl_141 br_141 wl_11 vdd gnd cell_6t
Xbit_r12_c141 bl_141 br_141 wl_12 vdd gnd cell_6t
Xbit_r13_c141 bl_141 br_141 wl_13 vdd gnd cell_6t
Xbit_r14_c141 bl_141 br_141 wl_14 vdd gnd cell_6t
Xbit_r15_c141 bl_141 br_141 wl_15 vdd gnd cell_6t
Xbit_r16_c141 bl_141 br_141 wl_16 vdd gnd cell_6t
Xbit_r17_c141 bl_141 br_141 wl_17 vdd gnd cell_6t
Xbit_r18_c141 bl_141 br_141 wl_18 vdd gnd cell_6t
Xbit_r19_c141 bl_141 br_141 wl_19 vdd gnd cell_6t
Xbit_r20_c141 bl_141 br_141 wl_20 vdd gnd cell_6t
Xbit_r21_c141 bl_141 br_141 wl_21 vdd gnd cell_6t
Xbit_r22_c141 bl_141 br_141 wl_22 vdd gnd cell_6t
Xbit_r23_c141 bl_141 br_141 wl_23 vdd gnd cell_6t
Xbit_r24_c141 bl_141 br_141 wl_24 vdd gnd cell_6t
Xbit_r25_c141 bl_141 br_141 wl_25 vdd gnd cell_6t
Xbit_r26_c141 bl_141 br_141 wl_26 vdd gnd cell_6t
Xbit_r27_c141 bl_141 br_141 wl_27 vdd gnd cell_6t
Xbit_r28_c141 bl_141 br_141 wl_28 vdd gnd cell_6t
Xbit_r29_c141 bl_141 br_141 wl_29 vdd gnd cell_6t
Xbit_r30_c141 bl_141 br_141 wl_30 vdd gnd cell_6t
Xbit_r31_c141 bl_141 br_141 wl_31 vdd gnd cell_6t
Xbit_r32_c141 bl_141 br_141 wl_32 vdd gnd cell_6t
Xbit_r33_c141 bl_141 br_141 wl_33 vdd gnd cell_6t
Xbit_r34_c141 bl_141 br_141 wl_34 vdd gnd cell_6t
Xbit_r35_c141 bl_141 br_141 wl_35 vdd gnd cell_6t
Xbit_r36_c141 bl_141 br_141 wl_36 vdd gnd cell_6t
Xbit_r37_c141 bl_141 br_141 wl_37 vdd gnd cell_6t
Xbit_r38_c141 bl_141 br_141 wl_38 vdd gnd cell_6t
Xbit_r39_c141 bl_141 br_141 wl_39 vdd gnd cell_6t
Xbit_r40_c141 bl_141 br_141 wl_40 vdd gnd cell_6t
Xbit_r41_c141 bl_141 br_141 wl_41 vdd gnd cell_6t
Xbit_r42_c141 bl_141 br_141 wl_42 vdd gnd cell_6t
Xbit_r43_c141 bl_141 br_141 wl_43 vdd gnd cell_6t
Xbit_r44_c141 bl_141 br_141 wl_44 vdd gnd cell_6t
Xbit_r45_c141 bl_141 br_141 wl_45 vdd gnd cell_6t
Xbit_r46_c141 bl_141 br_141 wl_46 vdd gnd cell_6t
Xbit_r47_c141 bl_141 br_141 wl_47 vdd gnd cell_6t
Xbit_r48_c141 bl_141 br_141 wl_48 vdd gnd cell_6t
Xbit_r49_c141 bl_141 br_141 wl_49 vdd gnd cell_6t
Xbit_r50_c141 bl_141 br_141 wl_50 vdd gnd cell_6t
Xbit_r51_c141 bl_141 br_141 wl_51 vdd gnd cell_6t
Xbit_r52_c141 bl_141 br_141 wl_52 vdd gnd cell_6t
Xbit_r53_c141 bl_141 br_141 wl_53 vdd gnd cell_6t
Xbit_r54_c141 bl_141 br_141 wl_54 vdd gnd cell_6t
Xbit_r55_c141 bl_141 br_141 wl_55 vdd gnd cell_6t
Xbit_r56_c141 bl_141 br_141 wl_56 vdd gnd cell_6t
Xbit_r57_c141 bl_141 br_141 wl_57 vdd gnd cell_6t
Xbit_r58_c141 bl_141 br_141 wl_58 vdd gnd cell_6t
Xbit_r59_c141 bl_141 br_141 wl_59 vdd gnd cell_6t
Xbit_r60_c141 bl_141 br_141 wl_60 vdd gnd cell_6t
Xbit_r61_c141 bl_141 br_141 wl_61 vdd gnd cell_6t
Xbit_r62_c141 bl_141 br_141 wl_62 vdd gnd cell_6t
Xbit_r63_c141 bl_141 br_141 wl_63 vdd gnd cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd cell_6t
Xbit_r1_c142 bl_142 br_142 wl_1 vdd gnd cell_6t
Xbit_r2_c142 bl_142 br_142 wl_2 vdd gnd cell_6t
Xbit_r3_c142 bl_142 br_142 wl_3 vdd gnd cell_6t
Xbit_r4_c142 bl_142 br_142 wl_4 vdd gnd cell_6t
Xbit_r5_c142 bl_142 br_142 wl_5 vdd gnd cell_6t
Xbit_r6_c142 bl_142 br_142 wl_6 vdd gnd cell_6t
Xbit_r7_c142 bl_142 br_142 wl_7 vdd gnd cell_6t
Xbit_r8_c142 bl_142 br_142 wl_8 vdd gnd cell_6t
Xbit_r9_c142 bl_142 br_142 wl_9 vdd gnd cell_6t
Xbit_r10_c142 bl_142 br_142 wl_10 vdd gnd cell_6t
Xbit_r11_c142 bl_142 br_142 wl_11 vdd gnd cell_6t
Xbit_r12_c142 bl_142 br_142 wl_12 vdd gnd cell_6t
Xbit_r13_c142 bl_142 br_142 wl_13 vdd gnd cell_6t
Xbit_r14_c142 bl_142 br_142 wl_14 vdd gnd cell_6t
Xbit_r15_c142 bl_142 br_142 wl_15 vdd gnd cell_6t
Xbit_r16_c142 bl_142 br_142 wl_16 vdd gnd cell_6t
Xbit_r17_c142 bl_142 br_142 wl_17 vdd gnd cell_6t
Xbit_r18_c142 bl_142 br_142 wl_18 vdd gnd cell_6t
Xbit_r19_c142 bl_142 br_142 wl_19 vdd gnd cell_6t
Xbit_r20_c142 bl_142 br_142 wl_20 vdd gnd cell_6t
Xbit_r21_c142 bl_142 br_142 wl_21 vdd gnd cell_6t
Xbit_r22_c142 bl_142 br_142 wl_22 vdd gnd cell_6t
Xbit_r23_c142 bl_142 br_142 wl_23 vdd gnd cell_6t
Xbit_r24_c142 bl_142 br_142 wl_24 vdd gnd cell_6t
Xbit_r25_c142 bl_142 br_142 wl_25 vdd gnd cell_6t
Xbit_r26_c142 bl_142 br_142 wl_26 vdd gnd cell_6t
Xbit_r27_c142 bl_142 br_142 wl_27 vdd gnd cell_6t
Xbit_r28_c142 bl_142 br_142 wl_28 vdd gnd cell_6t
Xbit_r29_c142 bl_142 br_142 wl_29 vdd gnd cell_6t
Xbit_r30_c142 bl_142 br_142 wl_30 vdd gnd cell_6t
Xbit_r31_c142 bl_142 br_142 wl_31 vdd gnd cell_6t
Xbit_r32_c142 bl_142 br_142 wl_32 vdd gnd cell_6t
Xbit_r33_c142 bl_142 br_142 wl_33 vdd gnd cell_6t
Xbit_r34_c142 bl_142 br_142 wl_34 vdd gnd cell_6t
Xbit_r35_c142 bl_142 br_142 wl_35 vdd gnd cell_6t
Xbit_r36_c142 bl_142 br_142 wl_36 vdd gnd cell_6t
Xbit_r37_c142 bl_142 br_142 wl_37 vdd gnd cell_6t
Xbit_r38_c142 bl_142 br_142 wl_38 vdd gnd cell_6t
Xbit_r39_c142 bl_142 br_142 wl_39 vdd gnd cell_6t
Xbit_r40_c142 bl_142 br_142 wl_40 vdd gnd cell_6t
Xbit_r41_c142 bl_142 br_142 wl_41 vdd gnd cell_6t
Xbit_r42_c142 bl_142 br_142 wl_42 vdd gnd cell_6t
Xbit_r43_c142 bl_142 br_142 wl_43 vdd gnd cell_6t
Xbit_r44_c142 bl_142 br_142 wl_44 vdd gnd cell_6t
Xbit_r45_c142 bl_142 br_142 wl_45 vdd gnd cell_6t
Xbit_r46_c142 bl_142 br_142 wl_46 vdd gnd cell_6t
Xbit_r47_c142 bl_142 br_142 wl_47 vdd gnd cell_6t
Xbit_r48_c142 bl_142 br_142 wl_48 vdd gnd cell_6t
Xbit_r49_c142 bl_142 br_142 wl_49 vdd gnd cell_6t
Xbit_r50_c142 bl_142 br_142 wl_50 vdd gnd cell_6t
Xbit_r51_c142 bl_142 br_142 wl_51 vdd gnd cell_6t
Xbit_r52_c142 bl_142 br_142 wl_52 vdd gnd cell_6t
Xbit_r53_c142 bl_142 br_142 wl_53 vdd gnd cell_6t
Xbit_r54_c142 bl_142 br_142 wl_54 vdd gnd cell_6t
Xbit_r55_c142 bl_142 br_142 wl_55 vdd gnd cell_6t
Xbit_r56_c142 bl_142 br_142 wl_56 vdd gnd cell_6t
Xbit_r57_c142 bl_142 br_142 wl_57 vdd gnd cell_6t
Xbit_r58_c142 bl_142 br_142 wl_58 vdd gnd cell_6t
Xbit_r59_c142 bl_142 br_142 wl_59 vdd gnd cell_6t
Xbit_r60_c142 bl_142 br_142 wl_60 vdd gnd cell_6t
Xbit_r61_c142 bl_142 br_142 wl_61 vdd gnd cell_6t
Xbit_r62_c142 bl_142 br_142 wl_62 vdd gnd cell_6t
Xbit_r63_c142 bl_142 br_142 wl_63 vdd gnd cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd cell_6t
Xbit_r1_c143 bl_143 br_143 wl_1 vdd gnd cell_6t
Xbit_r2_c143 bl_143 br_143 wl_2 vdd gnd cell_6t
Xbit_r3_c143 bl_143 br_143 wl_3 vdd gnd cell_6t
Xbit_r4_c143 bl_143 br_143 wl_4 vdd gnd cell_6t
Xbit_r5_c143 bl_143 br_143 wl_5 vdd gnd cell_6t
Xbit_r6_c143 bl_143 br_143 wl_6 vdd gnd cell_6t
Xbit_r7_c143 bl_143 br_143 wl_7 vdd gnd cell_6t
Xbit_r8_c143 bl_143 br_143 wl_8 vdd gnd cell_6t
Xbit_r9_c143 bl_143 br_143 wl_9 vdd gnd cell_6t
Xbit_r10_c143 bl_143 br_143 wl_10 vdd gnd cell_6t
Xbit_r11_c143 bl_143 br_143 wl_11 vdd gnd cell_6t
Xbit_r12_c143 bl_143 br_143 wl_12 vdd gnd cell_6t
Xbit_r13_c143 bl_143 br_143 wl_13 vdd gnd cell_6t
Xbit_r14_c143 bl_143 br_143 wl_14 vdd gnd cell_6t
Xbit_r15_c143 bl_143 br_143 wl_15 vdd gnd cell_6t
Xbit_r16_c143 bl_143 br_143 wl_16 vdd gnd cell_6t
Xbit_r17_c143 bl_143 br_143 wl_17 vdd gnd cell_6t
Xbit_r18_c143 bl_143 br_143 wl_18 vdd gnd cell_6t
Xbit_r19_c143 bl_143 br_143 wl_19 vdd gnd cell_6t
Xbit_r20_c143 bl_143 br_143 wl_20 vdd gnd cell_6t
Xbit_r21_c143 bl_143 br_143 wl_21 vdd gnd cell_6t
Xbit_r22_c143 bl_143 br_143 wl_22 vdd gnd cell_6t
Xbit_r23_c143 bl_143 br_143 wl_23 vdd gnd cell_6t
Xbit_r24_c143 bl_143 br_143 wl_24 vdd gnd cell_6t
Xbit_r25_c143 bl_143 br_143 wl_25 vdd gnd cell_6t
Xbit_r26_c143 bl_143 br_143 wl_26 vdd gnd cell_6t
Xbit_r27_c143 bl_143 br_143 wl_27 vdd gnd cell_6t
Xbit_r28_c143 bl_143 br_143 wl_28 vdd gnd cell_6t
Xbit_r29_c143 bl_143 br_143 wl_29 vdd gnd cell_6t
Xbit_r30_c143 bl_143 br_143 wl_30 vdd gnd cell_6t
Xbit_r31_c143 bl_143 br_143 wl_31 vdd gnd cell_6t
Xbit_r32_c143 bl_143 br_143 wl_32 vdd gnd cell_6t
Xbit_r33_c143 bl_143 br_143 wl_33 vdd gnd cell_6t
Xbit_r34_c143 bl_143 br_143 wl_34 vdd gnd cell_6t
Xbit_r35_c143 bl_143 br_143 wl_35 vdd gnd cell_6t
Xbit_r36_c143 bl_143 br_143 wl_36 vdd gnd cell_6t
Xbit_r37_c143 bl_143 br_143 wl_37 vdd gnd cell_6t
Xbit_r38_c143 bl_143 br_143 wl_38 vdd gnd cell_6t
Xbit_r39_c143 bl_143 br_143 wl_39 vdd gnd cell_6t
Xbit_r40_c143 bl_143 br_143 wl_40 vdd gnd cell_6t
Xbit_r41_c143 bl_143 br_143 wl_41 vdd gnd cell_6t
Xbit_r42_c143 bl_143 br_143 wl_42 vdd gnd cell_6t
Xbit_r43_c143 bl_143 br_143 wl_43 vdd gnd cell_6t
Xbit_r44_c143 bl_143 br_143 wl_44 vdd gnd cell_6t
Xbit_r45_c143 bl_143 br_143 wl_45 vdd gnd cell_6t
Xbit_r46_c143 bl_143 br_143 wl_46 vdd gnd cell_6t
Xbit_r47_c143 bl_143 br_143 wl_47 vdd gnd cell_6t
Xbit_r48_c143 bl_143 br_143 wl_48 vdd gnd cell_6t
Xbit_r49_c143 bl_143 br_143 wl_49 vdd gnd cell_6t
Xbit_r50_c143 bl_143 br_143 wl_50 vdd gnd cell_6t
Xbit_r51_c143 bl_143 br_143 wl_51 vdd gnd cell_6t
Xbit_r52_c143 bl_143 br_143 wl_52 vdd gnd cell_6t
Xbit_r53_c143 bl_143 br_143 wl_53 vdd gnd cell_6t
Xbit_r54_c143 bl_143 br_143 wl_54 vdd gnd cell_6t
Xbit_r55_c143 bl_143 br_143 wl_55 vdd gnd cell_6t
Xbit_r56_c143 bl_143 br_143 wl_56 vdd gnd cell_6t
Xbit_r57_c143 bl_143 br_143 wl_57 vdd gnd cell_6t
Xbit_r58_c143 bl_143 br_143 wl_58 vdd gnd cell_6t
Xbit_r59_c143 bl_143 br_143 wl_59 vdd gnd cell_6t
Xbit_r60_c143 bl_143 br_143 wl_60 vdd gnd cell_6t
Xbit_r61_c143 bl_143 br_143 wl_61 vdd gnd cell_6t
Xbit_r62_c143 bl_143 br_143 wl_62 vdd gnd cell_6t
Xbit_r63_c143 bl_143 br_143 wl_63 vdd gnd cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd cell_6t
Xbit_r1_c144 bl_144 br_144 wl_1 vdd gnd cell_6t
Xbit_r2_c144 bl_144 br_144 wl_2 vdd gnd cell_6t
Xbit_r3_c144 bl_144 br_144 wl_3 vdd gnd cell_6t
Xbit_r4_c144 bl_144 br_144 wl_4 vdd gnd cell_6t
Xbit_r5_c144 bl_144 br_144 wl_5 vdd gnd cell_6t
Xbit_r6_c144 bl_144 br_144 wl_6 vdd gnd cell_6t
Xbit_r7_c144 bl_144 br_144 wl_7 vdd gnd cell_6t
Xbit_r8_c144 bl_144 br_144 wl_8 vdd gnd cell_6t
Xbit_r9_c144 bl_144 br_144 wl_9 vdd gnd cell_6t
Xbit_r10_c144 bl_144 br_144 wl_10 vdd gnd cell_6t
Xbit_r11_c144 bl_144 br_144 wl_11 vdd gnd cell_6t
Xbit_r12_c144 bl_144 br_144 wl_12 vdd gnd cell_6t
Xbit_r13_c144 bl_144 br_144 wl_13 vdd gnd cell_6t
Xbit_r14_c144 bl_144 br_144 wl_14 vdd gnd cell_6t
Xbit_r15_c144 bl_144 br_144 wl_15 vdd gnd cell_6t
Xbit_r16_c144 bl_144 br_144 wl_16 vdd gnd cell_6t
Xbit_r17_c144 bl_144 br_144 wl_17 vdd gnd cell_6t
Xbit_r18_c144 bl_144 br_144 wl_18 vdd gnd cell_6t
Xbit_r19_c144 bl_144 br_144 wl_19 vdd gnd cell_6t
Xbit_r20_c144 bl_144 br_144 wl_20 vdd gnd cell_6t
Xbit_r21_c144 bl_144 br_144 wl_21 vdd gnd cell_6t
Xbit_r22_c144 bl_144 br_144 wl_22 vdd gnd cell_6t
Xbit_r23_c144 bl_144 br_144 wl_23 vdd gnd cell_6t
Xbit_r24_c144 bl_144 br_144 wl_24 vdd gnd cell_6t
Xbit_r25_c144 bl_144 br_144 wl_25 vdd gnd cell_6t
Xbit_r26_c144 bl_144 br_144 wl_26 vdd gnd cell_6t
Xbit_r27_c144 bl_144 br_144 wl_27 vdd gnd cell_6t
Xbit_r28_c144 bl_144 br_144 wl_28 vdd gnd cell_6t
Xbit_r29_c144 bl_144 br_144 wl_29 vdd gnd cell_6t
Xbit_r30_c144 bl_144 br_144 wl_30 vdd gnd cell_6t
Xbit_r31_c144 bl_144 br_144 wl_31 vdd gnd cell_6t
Xbit_r32_c144 bl_144 br_144 wl_32 vdd gnd cell_6t
Xbit_r33_c144 bl_144 br_144 wl_33 vdd gnd cell_6t
Xbit_r34_c144 bl_144 br_144 wl_34 vdd gnd cell_6t
Xbit_r35_c144 bl_144 br_144 wl_35 vdd gnd cell_6t
Xbit_r36_c144 bl_144 br_144 wl_36 vdd gnd cell_6t
Xbit_r37_c144 bl_144 br_144 wl_37 vdd gnd cell_6t
Xbit_r38_c144 bl_144 br_144 wl_38 vdd gnd cell_6t
Xbit_r39_c144 bl_144 br_144 wl_39 vdd gnd cell_6t
Xbit_r40_c144 bl_144 br_144 wl_40 vdd gnd cell_6t
Xbit_r41_c144 bl_144 br_144 wl_41 vdd gnd cell_6t
Xbit_r42_c144 bl_144 br_144 wl_42 vdd gnd cell_6t
Xbit_r43_c144 bl_144 br_144 wl_43 vdd gnd cell_6t
Xbit_r44_c144 bl_144 br_144 wl_44 vdd gnd cell_6t
Xbit_r45_c144 bl_144 br_144 wl_45 vdd gnd cell_6t
Xbit_r46_c144 bl_144 br_144 wl_46 vdd gnd cell_6t
Xbit_r47_c144 bl_144 br_144 wl_47 vdd gnd cell_6t
Xbit_r48_c144 bl_144 br_144 wl_48 vdd gnd cell_6t
Xbit_r49_c144 bl_144 br_144 wl_49 vdd gnd cell_6t
Xbit_r50_c144 bl_144 br_144 wl_50 vdd gnd cell_6t
Xbit_r51_c144 bl_144 br_144 wl_51 vdd gnd cell_6t
Xbit_r52_c144 bl_144 br_144 wl_52 vdd gnd cell_6t
Xbit_r53_c144 bl_144 br_144 wl_53 vdd gnd cell_6t
Xbit_r54_c144 bl_144 br_144 wl_54 vdd gnd cell_6t
Xbit_r55_c144 bl_144 br_144 wl_55 vdd gnd cell_6t
Xbit_r56_c144 bl_144 br_144 wl_56 vdd gnd cell_6t
Xbit_r57_c144 bl_144 br_144 wl_57 vdd gnd cell_6t
Xbit_r58_c144 bl_144 br_144 wl_58 vdd gnd cell_6t
Xbit_r59_c144 bl_144 br_144 wl_59 vdd gnd cell_6t
Xbit_r60_c144 bl_144 br_144 wl_60 vdd gnd cell_6t
Xbit_r61_c144 bl_144 br_144 wl_61 vdd gnd cell_6t
Xbit_r62_c144 bl_144 br_144 wl_62 vdd gnd cell_6t
Xbit_r63_c144 bl_144 br_144 wl_63 vdd gnd cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd cell_6t
Xbit_r1_c145 bl_145 br_145 wl_1 vdd gnd cell_6t
Xbit_r2_c145 bl_145 br_145 wl_2 vdd gnd cell_6t
Xbit_r3_c145 bl_145 br_145 wl_3 vdd gnd cell_6t
Xbit_r4_c145 bl_145 br_145 wl_4 vdd gnd cell_6t
Xbit_r5_c145 bl_145 br_145 wl_5 vdd gnd cell_6t
Xbit_r6_c145 bl_145 br_145 wl_6 vdd gnd cell_6t
Xbit_r7_c145 bl_145 br_145 wl_7 vdd gnd cell_6t
Xbit_r8_c145 bl_145 br_145 wl_8 vdd gnd cell_6t
Xbit_r9_c145 bl_145 br_145 wl_9 vdd gnd cell_6t
Xbit_r10_c145 bl_145 br_145 wl_10 vdd gnd cell_6t
Xbit_r11_c145 bl_145 br_145 wl_11 vdd gnd cell_6t
Xbit_r12_c145 bl_145 br_145 wl_12 vdd gnd cell_6t
Xbit_r13_c145 bl_145 br_145 wl_13 vdd gnd cell_6t
Xbit_r14_c145 bl_145 br_145 wl_14 vdd gnd cell_6t
Xbit_r15_c145 bl_145 br_145 wl_15 vdd gnd cell_6t
Xbit_r16_c145 bl_145 br_145 wl_16 vdd gnd cell_6t
Xbit_r17_c145 bl_145 br_145 wl_17 vdd gnd cell_6t
Xbit_r18_c145 bl_145 br_145 wl_18 vdd gnd cell_6t
Xbit_r19_c145 bl_145 br_145 wl_19 vdd gnd cell_6t
Xbit_r20_c145 bl_145 br_145 wl_20 vdd gnd cell_6t
Xbit_r21_c145 bl_145 br_145 wl_21 vdd gnd cell_6t
Xbit_r22_c145 bl_145 br_145 wl_22 vdd gnd cell_6t
Xbit_r23_c145 bl_145 br_145 wl_23 vdd gnd cell_6t
Xbit_r24_c145 bl_145 br_145 wl_24 vdd gnd cell_6t
Xbit_r25_c145 bl_145 br_145 wl_25 vdd gnd cell_6t
Xbit_r26_c145 bl_145 br_145 wl_26 vdd gnd cell_6t
Xbit_r27_c145 bl_145 br_145 wl_27 vdd gnd cell_6t
Xbit_r28_c145 bl_145 br_145 wl_28 vdd gnd cell_6t
Xbit_r29_c145 bl_145 br_145 wl_29 vdd gnd cell_6t
Xbit_r30_c145 bl_145 br_145 wl_30 vdd gnd cell_6t
Xbit_r31_c145 bl_145 br_145 wl_31 vdd gnd cell_6t
Xbit_r32_c145 bl_145 br_145 wl_32 vdd gnd cell_6t
Xbit_r33_c145 bl_145 br_145 wl_33 vdd gnd cell_6t
Xbit_r34_c145 bl_145 br_145 wl_34 vdd gnd cell_6t
Xbit_r35_c145 bl_145 br_145 wl_35 vdd gnd cell_6t
Xbit_r36_c145 bl_145 br_145 wl_36 vdd gnd cell_6t
Xbit_r37_c145 bl_145 br_145 wl_37 vdd gnd cell_6t
Xbit_r38_c145 bl_145 br_145 wl_38 vdd gnd cell_6t
Xbit_r39_c145 bl_145 br_145 wl_39 vdd gnd cell_6t
Xbit_r40_c145 bl_145 br_145 wl_40 vdd gnd cell_6t
Xbit_r41_c145 bl_145 br_145 wl_41 vdd gnd cell_6t
Xbit_r42_c145 bl_145 br_145 wl_42 vdd gnd cell_6t
Xbit_r43_c145 bl_145 br_145 wl_43 vdd gnd cell_6t
Xbit_r44_c145 bl_145 br_145 wl_44 vdd gnd cell_6t
Xbit_r45_c145 bl_145 br_145 wl_45 vdd gnd cell_6t
Xbit_r46_c145 bl_145 br_145 wl_46 vdd gnd cell_6t
Xbit_r47_c145 bl_145 br_145 wl_47 vdd gnd cell_6t
Xbit_r48_c145 bl_145 br_145 wl_48 vdd gnd cell_6t
Xbit_r49_c145 bl_145 br_145 wl_49 vdd gnd cell_6t
Xbit_r50_c145 bl_145 br_145 wl_50 vdd gnd cell_6t
Xbit_r51_c145 bl_145 br_145 wl_51 vdd gnd cell_6t
Xbit_r52_c145 bl_145 br_145 wl_52 vdd gnd cell_6t
Xbit_r53_c145 bl_145 br_145 wl_53 vdd gnd cell_6t
Xbit_r54_c145 bl_145 br_145 wl_54 vdd gnd cell_6t
Xbit_r55_c145 bl_145 br_145 wl_55 vdd gnd cell_6t
Xbit_r56_c145 bl_145 br_145 wl_56 vdd gnd cell_6t
Xbit_r57_c145 bl_145 br_145 wl_57 vdd gnd cell_6t
Xbit_r58_c145 bl_145 br_145 wl_58 vdd gnd cell_6t
Xbit_r59_c145 bl_145 br_145 wl_59 vdd gnd cell_6t
Xbit_r60_c145 bl_145 br_145 wl_60 vdd gnd cell_6t
Xbit_r61_c145 bl_145 br_145 wl_61 vdd gnd cell_6t
Xbit_r62_c145 bl_145 br_145 wl_62 vdd gnd cell_6t
Xbit_r63_c145 bl_145 br_145 wl_63 vdd gnd cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd cell_6t
Xbit_r1_c146 bl_146 br_146 wl_1 vdd gnd cell_6t
Xbit_r2_c146 bl_146 br_146 wl_2 vdd gnd cell_6t
Xbit_r3_c146 bl_146 br_146 wl_3 vdd gnd cell_6t
Xbit_r4_c146 bl_146 br_146 wl_4 vdd gnd cell_6t
Xbit_r5_c146 bl_146 br_146 wl_5 vdd gnd cell_6t
Xbit_r6_c146 bl_146 br_146 wl_6 vdd gnd cell_6t
Xbit_r7_c146 bl_146 br_146 wl_7 vdd gnd cell_6t
Xbit_r8_c146 bl_146 br_146 wl_8 vdd gnd cell_6t
Xbit_r9_c146 bl_146 br_146 wl_9 vdd gnd cell_6t
Xbit_r10_c146 bl_146 br_146 wl_10 vdd gnd cell_6t
Xbit_r11_c146 bl_146 br_146 wl_11 vdd gnd cell_6t
Xbit_r12_c146 bl_146 br_146 wl_12 vdd gnd cell_6t
Xbit_r13_c146 bl_146 br_146 wl_13 vdd gnd cell_6t
Xbit_r14_c146 bl_146 br_146 wl_14 vdd gnd cell_6t
Xbit_r15_c146 bl_146 br_146 wl_15 vdd gnd cell_6t
Xbit_r16_c146 bl_146 br_146 wl_16 vdd gnd cell_6t
Xbit_r17_c146 bl_146 br_146 wl_17 vdd gnd cell_6t
Xbit_r18_c146 bl_146 br_146 wl_18 vdd gnd cell_6t
Xbit_r19_c146 bl_146 br_146 wl_19 vdd gnd cell_6t
Xbit_r20_c146 bl_146 br_146 wl_20 vdd gnd cell_6t
Xbit_r21_c146 bl_146 br_146 wl_21 vdd gnd cell_6t
Xbit_r22_c146 bl_146 br_146 wl_22 vdd gnd cell_6t
Xbit_r23_c146 bl_146 br_146 wl_23 vdd gnd cell_6t
Xbit_r24_c146 bl_146 br_146 wl_24 vdd gnd cell_6t
Xbit_r25_c146 bl_146 br_146 wl_25 vdd gnd cell_6t
Xbit_r26_c146 bl_146 br_146 wl_26 vdd gnd cell_6t
Xbit_r27_c146 bl_146 br_146 wl_27 vdd gnd cell_6t
Xbit_r28_c146 bl_146 br_146 wl_28 vdd gnd cell_6t
Xbit_r29_c146 bl_146 br_146 wl_29 vdd gnd cell_6t
Xbit_r30_c146 bl_146 br_146 wl_30 vdd gnd cell_6t
Xbit_r31_c146 bl_146 br_146 wl_31 vdd gnd cell_6t
Xbit_r32_c146 bl_146 br_146 wl_32 vdd gnd cell_6t
Xbit_r33_c146 bl_146 br_146 wl_33 vdd gnd cell_6t
Xbit_r34_c146 bl_146 br_146 wl_34 vdd gnd cell_6t
Xbit_r35_c146 bl_146 br_146 wl_35 vdd gnd cell_6t
Xbit_r36_c146 bl_146 br_146 wl_36 vdd gnd cell_6t
Xbit_r37_c146 bl_146 br_146 wl_37 vdd gnd cell_6t
Xbit_r38_c146 bl_146 br_146 wl_38 vdd gnd cell_6t
Xbit_r39_c146 bl_146 br_146 wl_39 vdd gnd cell_6t
Xbit_r40_c146 bl_146 br_146 wl_40 vdd gnd cell_6t
Xbit_r41_c146 bl_146 br_146 wl_41 vdd gnd cell_6t
Xbit_r42_c146 bl_146 br_146 wl_42 vdd gnd cell_6t
Xbit_r43_c146 bl_146 br_146 wl_43 vdd gnd cell_6t
Xbit_r44_c146 bl_146 br_146 wl_44 vdd gnd cell_6t
Xbit_r45_c146 bl_146 br_146 wl_45 vdd gnd cell_6t
Xbit_r46_c146 bl_146 br_146 wl_46 vdd gnd cell_6t
Xbit_r47_c146 bl_146 br_146 wl_47 vdd gnd cell_6t
Xbit_r48_c146 bl_146 br_146 wl_48 vdd gnd cell_6t
Xbit_r49_c146 bl_146 br_146 wl_49 vdd gnd cell_6t
Xbit_r50_c146 bl_146 br_146 wl_50 vdd gnd cell_6t
Xbit_r51_c146 bl_146 br_146 wl_51 vdd gnd cell_6t
Xbit_r52_c146 bl_146 br_146 wl_52 vdd gnd cell_6t
Xbit_r53_c146 bl_146 br_146 wl_53 vdd gnd cell_6t
Xbit_r54_c146 bl_146 br_146 wl_54 vdd gnd cell_6t
Xbit_r55_c146 bl_146 br_146 wl_55 vdd gnd cell_6t
Xbit_r56_c146 bl_146 br_146 wl_56 vdd gnd cell_6t
Xbit_r57_c146 bl_146 br_146 wl_57 vdd gnd cell_6t
Xbit_r58_c146 bl_146 br_146 wl_58 vdd gnd cell_6t
Xbit_r59_c146 bl_146 br_146 wl_59 vdd gnd cell_6t
Xbit_r60_c146 bl_146 br_146 wl_60 vdd gnd cell_6t
Xbit_r61_c146 bl_146 br_146 wl_61 vdd gnd cell_6t
Xbit_r62_c146 bl_146 br_146 wl_62 vdd gnd cell_6t
Xbit_r63_c146 bl_146 br_146 wl_63 vdd gnd cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd cell_6t
Xbit_r1_c147 bl_147 br_147 wl_1 vdd gnd cell_6t
Xbit_r2_c147 bl_147 br_147 wl_2 vdd gnd cell_6t
Xbit_r3_c147 bl_147 br_147 wl_3 vdd gnd cell_6t
Xbit_r4_c147 bl_147 br_147 wl_4 vdd gnd cell_6t
Xbit_r5_c147 bl_147 br_147 wl_5 vdd gnd cell_6t
Xbit_r6_c147 bl_147 br_147 wl_6 vdd gnd cell_6t
Xbit_r7_c147 bl_147 br_147 wl_7 vdd gnd cell_6t
Xbit_r8_c147 bl_147 br_147 wl_8 vdd gnd cell_6t
Xbit_r9_c147 bl_147 br_147 wl_9 vdd gnd cell_6t
Xbit_r10_c147 bl_147 br_147 wl_10 vdd gnd cell_6t
Xbit_r11_c147 bl_147 br_147 wl_11 vdd gnd cell_6t
Xbit_r12_c147 bl_147 br_147 wl_12 vdd gnd cell_6t
Xbit_r13_c147 bl_147 br_147 wl_13 vdd gnd cell_6t
Xbit_r14_c147 bl_147 br_147 wl_14 vdd gnd cell_6t
Xbit_r15_c147 bl_147 br_147 wl_15 vdd gnd cell_6t
Xbit_r16_c147 bl_147 br_147 wl_16 vdd gnd cell_6t
Xbit_r17_c147 bl_147 br_147 wl_17 vdd gnd cell_6t
Xbit_r18_c147 bl_147 br_147 wl_18 vdd gnd cell_6t
Xbit_r19_c147 bl_147 br_147 wl_19 vdd gnd cell_6t
Xbit_r20_c147 bl_147 br_147 wl_20 vdd gnd cell_6t
Xbit_r21_c147 bl_147 br_147 wl_21 vdd gnd cell_6t
Xbit_r22_c147 bl_147 br_147 wl_22 vdd gnd cell_6t
Xbit_r23_c147 bl_147 br_147 wl_23 vdd gnd cell_6t
Xbit_r24_c147 bl_147 br_147 wl_24 vdd gnd cell_6t
Xbit_r25_c147 bl_147 br_147 wl_25 vdd gnd cell_6t
Xbit_r26_c147 bl_147 br_147 wl_26 vdd gnd cell_6t
Xbit_r27_c147 bl_147 br_147 wl_27 vdd gnd cell_6t
Xbit_r28_c147 bl_147 br_147 wl_28 vdd gnd cell_6t
Xbit_r29_c147 bl_147 br_147 wl_29 vdd gnd cell_6t
Xbit_r30_c147 bl_147 br_147 wl_30 vdd gnd cell_6t
Xbit_r31_c147 bl_147 br_147 wl_31 vdd gnd cell_6t
Xbit_r32_c147 bl_147 br_147 wl_32 vdd gnd cell_6t
Xbit_r33_c147 bl_147 br_147 wl_33 vdd gnd cell_6t
Xbit_r34_c147 bl_147 br_147 wl_34 vdd gnd cell_6t
Xbit_r35_c147 bl_147 br_147 wl_35 vdd gnd cell_6t
Xbit_r36_c147 bl_147 br_147 wl_36 vdd gnd cell_6t
Xbit_r37_c147 bl_147 br_147 wl_37 vdd gnd cell_6t
Xbit_r38_c147 bl_147 br_147 wl_38 vdd gnd cell_6t
Xbit_r39_c147 bl_147 br_147 wl_39 vdd gnd cell_6t
Xbit_r40_c147 bl_147 br_147 wl_40 vdd gnd cell_6t
Xbit_r41_c147 bl_147 br_147 wl_41 vdd gnd cell_6t
Xbit_r42_c147 bl_147 br_147 wl_42 vdd gnd cell_6t
Xbit_r43_c147 bl_147 br_147 wl_43 vdd gnd cell_6t
Xbit_r44_c147 bl_147 br_147 wl_44 vdd gnd cell_6t
Xbit_r45_c147 bl_147 br_147 wl_45 vdd gnd cell_6t
Xbit_r46_c147 bl_147 br_147 wl_46 vdd gnd cell_6t
Xbit_r47_c147 bl_147 br_147 wl_47 vdd gnd cell_6t
Xbit_r48_c147 bl_147 br_147 wl_48 vdd gnd cell_6t
Xbit_r49_c147 bl_147 br_147 wl_49 vdd gnd cell_6t
Xbit_r50_c147 bl_147 br_147 wl_50 vdd gnd cell_6t
Xbit_r51_c147 bl_147 br_147 wl_51 vdd gnd cell_6t
Xbit_r52_c147 bl_147 br_147 wl_52 vdd gnd cell_6t
Xbit_r53_c147 bl_147 br_147 wl_53 vdd gnd cell_6t
Xbit_r54_c147 bl_147 br_147 wl_54 vdd gnd cell_6t
Xbit_r55_c147 bl_147 br_147 wl_55 vdd gnd cell_6t
Xbit_r56_c147 bl_147 br_147 wl_56 vdd gnd cell_6t
Xbit_r57_c147 bl_147 br_147 wl_57 vdd gnd cell_6t
Xbit_r58_c147 bl_147 br_147 wl_58 vdd gnd cell_6t
Xbit_r59_c147 bl_147 br_147 wl_59 vdd gnd cell_6t
Xbit_r60_c147 bl_147 br_147 wl_60 vdd gnd cell_6t
Xbit_r61_c147 bl_147 br_147 wl_61 vdd gnd cell_6t
Xbit_r62_c147 bl_147 br_147 wl_62 vdd gnd cell_6t
Xbit_r63_c147 bl_147 br_147 wl_63 vdd gnd cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd cell_6t
Xbit_r1_c148 bl_148 br_148 wl_1 vdd gnd cell_6t
Xbit_r2_c148 bl_148 br_148 wl_2 vdd gnd cell_6t
Xbit_r3_c148 bl_148 br_148 wl_3 vdd gnd cell_6t
Xbit_r4_c148 bl_148 br_148 wl_4 vdd gnd cell_6t
Xbit_r5_c148 bl_148 br_148 wl_5 vdd gnd cell_6t
Xbit_r6_c148 bl_148 br_148 wl_6 vdd gnd cell_6t
Xbit_r7_c148 bl_148 br_148 wl_7 vdd gnd cell_6t
Xbit_r8_c148 bl_148 br_148 wl_8 vdd gnd cell_6t
Xbit_r9_c148 bl_148 br_148 wl_9 vdd gnd cell_6t
Xbit_r10_c148 bl_148 br_148 wl_10 vdd gnd cell_6t
Xbit_r11_c148 bl_148 br_148 wl_11 vdd gnd cell_6t
Xbit_r12_c148 bl_148 br_148 wl_12 vdd gnd cell_6t
Xbit_r13_c148 bl_148 br_148 wl_13 vdd gnd cell_6t
Xbit_r14_c148 bl_148 br_148 wl_14 vdd gnd cell_6t
Xbit_r15_c148 bl_148 br_148 wl_15 vdd gnd cell_6t
Xbit_r16_c148 bl_148 br_148 wl_16 vdd gnd cell_6t
Xbit_r17_c148 bl_148 br_148 wl_17 vdd gnd cell_6t
Xbit_r18_c148 bl_148 br_148 wl_18 vdd gnd cell_6t
Xbit_r19_c148 bl_148 br_148 wl_19 vdd gnd cell_6t
Xbit_r20_c148 bl_148 br_148 wl_20 vdd gnd cell_6t
Xbit_r21_c148 bl_148 br_148 wl_21 vdd gnd cell_6t
Xbit_r22_c148 bl_148 br_148 wl_22 vdd gnd cell_6t
Xbit_r23_c148 bl_148 br_148 wl_23 vdd gnd cell_6t
Xbit_r24_c148 bl_148 br_148 wl_24 vdd gnd cell_6t
Xbit_r25_c148 bl_148 br_148 wl_25 vdd gnd cell_6t
Xbit_r26_c148 bl_148 br_148 wl_26 vdd gnd cell_6t
Xbit_r27_c148 bl_148 br_148 wl_27 vdd gnd cell_6t
Xbit_r28_c148 bl_148 br_148 wl_28 vdd gnd cell_6t
Xbit_r29_c148 bl_148 br_148 wl_29 vdd gnd cell_6t
Xbit_r30_c148 bl_148 br_148 wl_30 vdd gnd cell_6t
Xbit_r31_c148 bl_148 br_148 wl_31 vdd gnd cell_6t
Xbit_r32_c148 bl_148 br_148 wl_32 vdd gnd cell_6t
Xbit_r33_c148 bl_148 br_148 wl_33 vdd gnd cell_6t
Xbit_r34_c148 bl_148 br_148 wl_34 vdd gnd cell_6t
Xbit_r35_c148 bl_148 br_148 wl_35 vdd gnd cell_6t
Xbit_r36_c148 bl_148 br_148 wl_36 vdd gnd cell_6t
Xbit_r37_c148 bl_148 br_148 wl_37 vdd gnd cell_6t
Xbit_r38_c148 bl_148 br_148 wl_38 vdd gnd cell_6t
Xbit_r39_c148 bl_148 br_148 wl_39 vdd gnd cell_6t
Xbit_r40_c148 bl_148 br_148 wl_40 vdd gnd cell_6t
Xbit_r41_c148 bl_148 br_148 wl_41 vdd gnd cell_6t
Xbit_r42_c148 bl_148 br_148 wl_42 vdd gnd cell_6t
Xbit_r43_c148 bl_148 br_148 wl_43 vdd gnd cell_6t
Xbit_r44_c148 bl_148 br_148 wl_44 vdd gnd cell_6t
Xbit_r45_c148 bl_148 br_148 wl_45 vdd gnd cell_6t
Xbit_r46_c148 bl_148 br_148 wl_46 vdd gnd cell_6t
Xbit_r47_c148 bl_148 br_148 wl_47 vdd gnd cell_6t
Xbit_r48_c148 bl_148 br_148 wl_48 vdd gnd cell_6t
Xbit_r49_c148 bl_148 br_148 wl_49 vdd gnd cell_6t
Xbit_r50_c148 bl_148 br_148 wl_50 vdd gnd cell_6t
Xbit_r51_c148 bl_148 br_148 wl_51 vdd gnd cell_6t
Xbit_r52_c148 bl_148 br_148 wl_52 vdd gnd cell_6t
Xbit_r53_c148 bl_148 br_148 wl_53 vdd gnd cell_6t
Xbit_r54_c148 bl_148 br_148 wl_54 vdd gnd cell_6t
Xbit_r55_c148 bl_148 br_148 wl_55 vdd gnd cell_6t
Xbit_r56_c148 bl_148 br_148 wl_56 vdd gnd cell_6t
Xbit_r57_c148 bl_148 br_148 wl_57 vdd gnd cell_6t
Xbit_r58_c148 bl_148 br_148 wl_58 vdd gnd cell_6t
Xbit_r59_c148 bl_148 br_148 wl_59 vdd gnd cell_6t
Xbit_r60_c148 bl_148 br_148 wl_60 vdd gnd cell_6t
Xbit_r61_c148 bl_148 br_148 wl_61 vdd gnd cell_6t
Xbit_r62_c148 bl_148 br_148 wl_62 vdd gnd cell_6t
Xbit_r63_c148 bl_148 br_148 wl_63 vdd gnd cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd cell_6t
Xbit_r1_c149 bl_149 br_149 wl_1 vdd gnd cell_6t
Xbit_r2_c149 bl_149 br_149 wl_2 vdd gnd cell_6t
Xbit_r3_c149 bl_149 br_149 wl_3 vdd gnd cell_6t
Xbit_r4_c149 bl_149 br_149 wl_4 vdd gnd cell_6t
Xbit_r5_c149 bl_149 br_149 wl_5 vdd gnd cell_6t
Xbit_r6_c149 bl_149 br_149 wl_6 vdd gnd cell_6t
Xbit_r7_c149 bl_149 br_149 wl_7 vdd gnd cell_6t
Xbit_r8_c149 bl_149 br_149 wl_8 vdd gnd cell_6t
Xbit_r9_c149 bl_149 br_149 wl_9 vdd gnd cell_6t
Xbit_r10_c149 bl_149 br_149 wl_10 vdd gnd cell_6t
Xbit_r11_c149 bl_149 br_149 wl_11 vdd gnd cell_6t
Xbit_r12_c149 bl_149 br_149 wl_12 vdd gnd cell_6t
Xbit_r13_c149 bl_149 br_149 wl_13 vdd gnd cell_6t
Xbit_r14_c149 bl_149 br_149 wl_14 vdd gnd cell_6t
Xbit_r15_c149 bl_149 br_149 wl_15 vdd gnd cell_6t
Xbit_r16_c149 bl_149 br_149 wl_16 vdd gnd cell_6t
Xbit_r17_c149 bl_149 br_149 wl_17 vdd gnd cell_6t
Xbit_r18_c149 bl_149 br_149 wl_18 vdd gnd cell_6t
Xbit_r19_c149 bl_149 br_149 wl_19 vdd gnd cell_6t
Xbit_r20_c149 bl_149 br_149 wl_20 vdd gnd cell_6t
Xbit_r21_c149 bl_149 br_149 wl_21 vdd gnd cell_6t
Xbit_r22_c149 bl_149 br_149 wl_22 vdd gnd cell_6t
Xbit_r23_c149 bl_149 br_149 wl_23 vdd gnd cell_6t
Xbit_r24_c149 bl_149 br_149 wl_24 vdd gnd cell_6t
Xbit_r25_c149 bl_149 br_149 wl_25 vdd gnd cell_6t
Xbit_r26_c149 bl_149 br_149 wl_26 vdd gnd cell_6t
Xbit_r27_c149 bl_149 br_149 wl_27 vdd gnd cell_6t
Xbit_r28_c149 bl_149 br_149 wl_28 vdd gnd cell_6t
Xbit_r29_c149 bl_149 br_149 wl_29 vdd gnd cell_6t
Xbit_r30_c149 bl_149 br_149 wl_30 vdd gnd cell_6t
Xbit_r31_c149 bl_149 br_149 wl_31 vdd gnd cell_6t
Xbit_r32_c149 bl_149 br_149 wl_32 vdd gnd cell_6t
Xbit_r33_c149 bl_149 br_149 wl_33 vdd gnd cell_6t
Xbit_r34_c149 bl_149 br_149 wl_34 vdd gnd cell_6t
Xbit_r35_c149 bl_149 br_149 wl_35 vdd gnd cell_6t
Xbit_r36_c149 bl_149 br_149 wl_36 vdd gnd cell_6t
Xbit_r37_c149 bl_149 br_149 wl_37 vdd gnd cell_6t
Xbit_r38_c149 bl_149 br_149 wl_38 vdd gnd cell_6t
Xbit_r39_c149 bl_149 br_149 wl_39 vdd gnd cell_6t
Xbit_r40_c149 bl_149 br_149 wl_40 vdd gnd cell_6t
Xbit_r41_c149 bl_149 br_149 wl_41 vdd gnd cell_6t
Xbit_r42_c149 bl_149 br_149 wl_42 vdd gnd cell_6t
Xbit_r43_c149 bl_149 br_149 wl_43 vdd gnd cell_6t
Xbit_r44_c149 bl_149 br_149 wl_44 vdd gnd cell_6t
Xbit_r45_c149 bl_149 br_149 wl_45 vdd gnd cell_6t
Xbit_r46_c149 bl_149 br_149 wl_46 vdd gnd cell_6t
Xbit_r47_c149 bl_149 br_149 wl_47 vdd gnd cell_6t
Xbit_r48_c149 bl_149 br_149 wl_48 vdd gnd cell_6t
Xbit_r49_c149 bl_149 br_149 wl_49 vdd gnd cell_6t
Xbit_r50_c149 bl_149 br_149 wl_50 vdd gnd cell_6t
Xbit_r51_c149 bl_149 br_149 wl_51 vdd gnd cell_6t
Xbit_r52_c149 bl_149 br_149 wl_52 vdd gnd cell_6t
Xbit_r53_c149 bl_149 br_149 wl_53 vdd gnd cell_6t
Xbit_r54_c149 bl_149 br_149 wl_54 vdd gnd cell_6t
Xbit_r55_c149 bl_149 br_149 wl_55 vdd gnd cell_6t
Xbit_r56_c149 bl_149 br_149 wl_56 vdd gnd cell_6t
Xbit_r57_c149 bl_149 br_149 wl_57 vdd gnd cell_6t
Xbit_r58_c149 bl_149 br_149 wl_58 vdd gnd cell_6t
Xbit_r59_c149 bl_149 br_149 wl_59 vdd gnd cell_6t
Xbit_r60_c149 bl_149 br_149 wl_60 vdd gnd cell_6t
Xbit_r61_c149 bl_149 br_149 wl_61 vdd gnd cell_6t
Xbit_r62_c149 bl_149 br_149 wl_62 vdd gnd cell_6t
Xbit_r63_c149 bl_149 br_149 wl_63 vdd gnd cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd cell_6t
Xbit_r1_c150 bl_150 br_150 wl_1 vdd gnd cell_6t
Xbit_r2_c150 bl_150 br_150 wl_2 vdd gnd cell_6t
Xbit_r3_c150 bl_150 br_150 wl_3 vdd gnd cell_6t
Xbit_r4_c150 bl_150 br_150 wl_4 vdd gnd cell_6t
Xbit_r5_c150 bl_150 br_150 wl_5 vdd gnd cell_6t
Xbit_r6_c150 bl_150 br_150 wl_6 vdd gnd cell_6t
Xbit_r7_c150 bl_150 br_150 wl_7 vdd gnd cell_6t
Xbit_r8_c150 bl_150 br_150 wl_8 vdd gnd cell_6t
Xbit_r9_c150 bl_150 br_150 wl_9 vdd gnd cell_6t
Xbit_r10_c150 bl_150 br_150 wl_10 vdd gnd cell_6t
Xbit_r11_c150 bl_150 br_150 wl_11 vdd gnd cell_6t
Xbit_r12_c150 bl_150 br_150 wl_12 vdd gnd cell_6t
Xbit_r13_c150 bl_150 br_150 wl_13 vdd gnd cell_6t
Xbit_r14_c150 bl_150 br_150 wl_14 vdd gnd cell_6t
Xbit_r15_c150 bl_150 br_150 wl_15 vdd gnd cell_6t
Xbit_r16_c150 bl_150 br_150 wl_16 vdd gnd cell_6t
Xbit_r17_c150 bl_150 br_150 wl_17 vdd gnd cell_6t
Xbit_r18_c150 bl_150 br_150 wl_18 vdd gnd cell_6t
Xbit_r19_c150 bl_150 br_150 wl_19 vdd gnd cell_6t
Xbit_r20_c150 bl_150 br_150 wl_20 vdd gnd cell_6t
Xbit_r21_c150 bl_150 br_150 wl_21 vdd gnd cell_6t
Xbit_r22_c150 bl_150 br_150 wl_22 vdd gnd cell_6t
Xbit_r23_c150 bl_150 br_150 wl_23 vdd gnd cell_6t
Xbit_r24_c150 bl_150 br_150 wl_24 vdd gnd cell_6t
Xbit_r25_c150 bl_150 br_150 wl_25 vdd gnd cell_6t
Xbit_r26_c150 bl_150 br_150 wl_26 vdd gnd cell_6t
Xbit_r27_c150 bl_150 br_150 wl_27 vdd gnd cell_6t
Xbit_r28_c150 bl_150 br_150 wl_28 vdd gnd cell_6t
Xbit_r29_c150 bl_150 br_150 wl_29 vdd gnd cell_6t
Xbit_r30_c150 bl_150 br_150 wl_30 vdd gnd cell_6t
Xbit_r31_c150 bl_150 br_150 wl_31 vdd gnd cell_6t
Xbit_r32_c150 bl_150 br_150 wl_32 vdd gnd cell_6t
Xbit_r33_c150 bl_150 br_150 wl_33 vdd gnd cell_6t
Xbit_r34_c150 bl_150 br_150 wl_34 vdd gnd cell_6t
Xbit_r35_c150 bl_150 br_150 wl_35 vdd gnd cell_6t
Xbit_r36_c150 bl_150 br_150 wl_36 vdd gnd cell_6t
Xbit_r37_c150 bl_150 br_150 wl_37 vdd gnd cell_6t
Xbit_r38_c150 bl_150 br_150 wl_38 vdd gnd cell_6t
Xbit_r39_c150 bl_150 br_150 wl_39 vdd gnd cell_6t
Xbit_r40_c150 bl_150 br_150 wl_40 vdd gnd cell_6t
Xbit_r41_c150 bl_150 br_150 wl_41 vdd gnd cell_6t
Xbit_r42_c150 bl_150 br_150 wl_42 vdd gnd cell_6t
Xbit_r43_c150 bl_150 br_150 wl_43 vdd gnd cell_6t
Xbit_r44_c150 bl_150 br_150 wl_44 vdd gnd cell_6t
Xbit_r45_c150 bl_150 br_150 wl_45 vdd gnd cell_6t
Xbit_r46_c150 bl_150 br_150 wl_46 vdd gnd cell_6t
Xbit_r47_c150 bl_150 br_150 wl_47 vdd gnd cell_6t
Xbit_r48_c150 bl_150 br_150 wl_48 vdd gnd cell_6t
Xbit_r49_c150 bl_150 br_150 wl_49 vdd gnd cell_6t
Xbit_r50_c150 bl_150 br_150 wl_50 vdd gnd cell_6t
Xbit_r51_c150 bl_150 br_150 wl_51 vdd gnd cell_6t
Xbit_r52_c150 bl_150 br_150 wl_52 vdd gnd cell_6t
Xbit_r53_c150 bl_150 br_150 wl_53 vdd gnd cell_6t
Xbit_r54_c150 bl_150 br_150 wl_54 vdd gnd cell_6t
Xbit_r55_c150 bl_150 br_150 wl_55 vdd gnd cell_6t
Xbit_r56_c150 bl_150 br_150 wl_56 vdd gnd cell_6t
Xbit_r57_c150 bl_150 br_150 wl_57 vdd gnd cell_6t
Xbit_r58_c150 bl_150 br_150 wl_58 vdd gnd cell_6t
Xbit_r59_c150 bl_150 br_150 wl_59 vdd gnd cell_6t
Xbit_r60_c150 bl_150 br_150 wl_60 vdd gnd cell_6t
Xbit_r61_c150 bl_150 br_150 wl_61 vdd gnd cell_6t
Xbit_r62_c150 bl_150 br_150 wl_62 vdd gnd cell_6t
Xbit_r63_c150 bl_150 br_150 wl_63 vdd gnd cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd cell_6t
Xbit_r1_c151 bl_151 br_151 wl_1 vdd gnd cell_6t
Xbit_r2_c151 bl_151 br_151 wl_2 vdd gnd cell_6t
Xbit_r3_c151 bl_151 br_151 wl_3 vdd gnd cell_6t
Xbit_r4_c151 bl_151 br_151 wl_4 vdd gnd cell_6t
Xbit_r5_c151 bl_151 br_151 wl_5 vdd gnd cell_6t
Xbit_r6_c151 bl_151 br_151 wl_6 vdd gnd cell_6t
Xbit_r7_c151 bl_151 br_151 wl_7 vdd gnd cell_6t
Xbit_r8_c151 bl_151 br_151 wl_8 vdd gnd cell_6t
Xbit_r9_c151 bl_151 br_151 wl_9 vdd gnd cell_6t
Xbit_r10_c151 bl_151 br_151 wl_10 vdd gnd cell_6t
Xbit_r11_c151 bl_151 br_151 wl_11 vdd gnd cell_6t
Xbit_r12_c151 bl_151 br_151 wl_12 vdd gnd cell_6t
Xbit_r13_c151 bl_151 br_151 wl_13 vdd gnd cell_6t
Xbit_r14_c151 bl_151 br_151 wl_14 vdd gnd cell_6t
Xbit_r15_c151 bl_151 br_151 wl_15 vdd gnd cell_6t
Xbit_r16_c151 bl_151 br_151 wl_16 vdd gnd cell_6t
Xbit_r17_c151 bl_151 br_151 wl_17 vdd gnd cell_6t
Xbit_r18_c151 bl_151 br_151 wl_18 vdd gnd cell_6t
Xbit_r19_c151 bl_151 br_151 wl_19 vdd gnd cell_6t
Xbit_r20_c151 bl_151 br_151 wl_20 vdd gnd cell_6t
Xbit_r21_c151 bl_151 br_151 wl_21 vdd gnd cell_6t
Xbit_r22_c151 bl_151 br_151 wl_22 vdd gnd cell_6t
Xbit_r23_c151 bl_151 br_151 wl_23 vdd gnd cell_6t
Xbit_r24_c151 bl_151 br_151 wl_24 vdd gnd cell_6t
Xbit_r25_c151 bl_151 br_151 wl_25 vdd gnd cell_6t
Xbit_r26_c151 bl_151 br_151 wl_26 vdd gnd cell_6t
Xbit_r27_c151 bl_151 br_151 wl_27 vdd gnd cell_6t
Xbit_r28_c151 bl_151 br_151 wl_28 vdd gnd cell_6t
Xbit_r29_c151 bl_151 br_151 wl_29 vdd gnd cell_6t
Xbit_r30_c151 bl_151 br_151 wl_30 vdd gnd cell_6t
Xbit_r31_c151 bl_151 br_151 wl_31 vdd gnd cell_6t
Xbit_r32_c151 bl_151 br_151 wl_32 vdd gnd cell_6t
Xbit_r33_c151 bl_151 br_151 wl_33 vdd gnd cell_6t
Xbit_r34_c151 bl_151 br_151 wl_34 vdd gnd cell_6t
Xbit_r35_c151 bl_151 br_151 wl_35 vdd gnd cell_6t
Xbit_r36_c151 bl_151 br_151 wl_36 vdd gnd cell_6t
Xbit_r37_c151 bl_151 br_151 wl_37 vdd gnd cell_6t
Xbit_r38_c151 bl_151 br_151 wl_38 vdd gnd cell_6t
Xbit_r39_c151 bl_151 br_151 wl_39 vdd gnd cell_6t
Xbit_r40_c151 bl_151 br_151 wl_40 vdd gnd cell_6t
Xbit_r41_c151 bl_151 br_151 wl_41 vdd gnd cell_6t
Xbit_r42_c151 bl_151 br_151 wl_42 vdd gnd cell_6t
Xbit_r43_c151 bl_151 br_151 wl_43 vdd gnd cell_6t
Xbit_r44_c151 bl_151 br_151 wl_44 vdd gnd cell_6t
Xbit_r45_c151 bl_151 br_151 wl_45 vdd gnd cell_6t
Xbit_r46_c151 bl_151 br_151 wl_46 vdd gnd cell_6t
Xbit_r47_c151 bl_151 br_151 wl_47 vdd gnd cell_6t
Xbit_r48_c151 bl_151 br_151 wl_48 vdd gnd cell_6t
Xbit_r49_c151 bl_151 br_151 wl_49 vdd gnd cell_6t
Xbit_r50_c151 bl_151 br_151 wl_50 vdd gnd cell_6t
Xbit_r51_c151 bl_151 br_151 wl_51 vdd gnd cell_6t
Xbit_r52_c151 bl_151 br_151 wl_52 vdd gnd cell_6t
Xbit_r53_c151 bl_151 br_151 wl_53 vdd gnd cell_6t
Xbit_r54_c151 bl_151 br_151 wl_54 vdd gnd cell_6t
Xbit_r55_c151 bl_151 br_151 wl_55 vdd gnd cell_6t
Xbit_r56_c151 bl_151 br_151 wl_56 vdd gnd cell_6t
Xbit_r57_c151 bl_151 br_151 wl_57 vdd gnd cell_6t
Xbit_r58_c151 bl_151 br_151 wl_58 vdd gnd cell_6t
Xbit_r59_c151 bl_151 br_151 wl_59 vdd gnd cell_6t
Xbit_r60_c151 bl_151 br_151 wl_60 vdd gnd cell_6t
Xbit_r61_c151 bl_151 br_151 wl_61 vdd gnd cell_6t
Xbit_r62_c151 bl_151 br_151 wl_62 vdd gnd cell_6t
Xbit_r63_c151 bl_151 br_151 wl_63 vdd gnd cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd cell_6t
Xbit_r1_c152 bl_152 br_152 wl_1 vdd gnd cell_6t
Xbit_r2_c152 bl_152 br_152 wl_2 vdd gnd cell_6t
Xbit_r3_c152 bl_152 br_152 wl_3 vdd gnd cell_6t
Xbit_r4_c152 bl_152 br_152 wl_4 vdd gnd cell_6t
Xbit_r5_c152 bl_152 br_152 wl_5 vdd gnd cell_6t
Xbit_r6_c152 bl_152 br_152 wl_6 vdd gnd cell_6t
Xbit_r7_c152 bl_152 br_152 wl_7 vdd gnd cell_6t
Xbit_r8_c152 bl_152 br_152 wl_8 vdd gnd cell_6t
Xbit_r9_c152 bl_152 br_152 wl_9 vdd gnd cell_6t
Xbit_r10_c152 bl_152 br_152 wl_10 vdd gnd cell_6t
Xbit_r11_c152 bl_152 br_152 wl_11 vdd gnd cell_6t
Xbit_r12_c152 bl_152 br_152 wl_12 vdd gnd cell_6t
Xbit_r13_c152 bl_152 br_152 wl_13 vdd gnd cell_6t
Xbit_r14_c152 bl_152 br_152 wl_14 vdd gnd cell_6t
Xbit_r15_c152 bl_152 br_152 wl_15 vdd gnd cell_6t
Xbit_r16_c152 bl_152 br_152 wl_16 vdd gnd cell_6t
Xbit_r17_c152 bl_152 br_152 wl_17 vdd gnd cell_6t
Xbit_r18_c152 bl_152 br_152 wl_18 vdd gnd cell_6t
Xbit_r19_c152 bl_152 br_152 wl_19 vdd gnd cell_6t
Xbit_r20_c152 bl_152 br_152 wl_20 vdd gnd cell_6t
Xbit_r21_c152 bl_152 br_152 wl_21 vdd gnd cell_6t
Xbit_r22_c152 bl_152 br_152 wl_22 vdd gnd cell_6t
Xbit_r23_c152 bl_152 br_152 wl_23 vdd gnd cell_6t
Xbit_r24_c152 bl_152 br_152 wl_24 vdd gnd cell_6t
Xbit_r25_c152 bl_152 br_152 wl_25 vdd gnd cell_6t
Xbit_r26_c152 bl_152 br_152 wl_26 vdd gnd cell_6t
Xbit_r27_c152 bl_152 br_152 wl_27 vdd gnd cell_6t
Xbit_r28_c152 bl_152 br_152 wl_28 vdd gnd cell_6t
Xbit_r29_c152 bl_152 br_152 wl_29 vdd gnd cell_6t
Xbit_r30_c152 bl_152 br_152 wl_30 vdd gnd cell_6t
Xbit_r31_c152 bl_152 br_152 wl_31 vdd gnd cell_6t
Xbit_r32_c152 bl_152 br_152 wl_32 vdd gnd cell_6t
Xbit_r33_c152 bl_152 br_152 wl_33 vdd gnd cell_6t
Xbit_r34_c152 bl_152 br_152 wl_34 vdd gnd cell_6t
Xbit_r35_c152 bl_152 br_152 wl_35 vdd gnd cell_6t
Xbit_r36_c152 bl_152 br_152 wl_36 vdd gnd cell_6t
Xbit_r37_c152 bl_152 br_152 wl_37 vdd gnd cell_6t
Xbit_r38_c152 bl_152 br_152 wl_38 vdd gnd cell_6t
Xbit_r39_c152 bl_152 br_152 wl_39 vdd gnd cell_6t
Xbit_r40_c152 bl_152 br_152 wl_40 vdd gnd cell_6t
Xbit_r41_c152 bl_152 br_152 wl_41 vdd gnd cell_6t
Xbit_r42_c152 bl_152 br_152 wl_42 vdd gnd cell_6t
Xbit_r43_c152 bl_152 br_152 wl_43 vdd gnd cell_6t
Xbit_r44_c152 bl_152 br_152 wl_44 vdd gnd cell_6t
Xbit_r45_c152 bl_152 br_152 wl_45 vdd gnd cell_6t
Xbit_r46_c152 bl_152 br_152 wl_46 vdd gnd cell_6t
Xbit_r47_c152 bl_152 br_152 wl_47 vdd gnd cell_6t
Xbit_r48_c152 bl_152 br_152 wl_48 vdd gnd cell_6t
Xbit_r49_c152 bl_152 br_152 wl_49 vdd gnd cell_6t
Xbit_r50_c152 bl_152 br_152 wl_50 vdd gnd cell_6t
Xbit_r51_c152 bl_152 br_152 wl_51 vdd gnd cell_6t
Xbit_r52_c152 bl_152 br_152 wl_52 vdd gnd cell_6t
Xbit_r53_c152 bl_152 br_152 wl_53 vdd gnd cell_6t
Xbit_r54_c152 bl_152 br_152 wl_54 vdd gnd cell_6t
Xbit_r55_c152 bl_152 br_152 wl_55 vdd gnd cell_6t
Xbit_r56_c152 bl_152 br_152 wl_56 vdd gnd cell_6t
Xbit_r57_c152 bl_152 br_152 wl_57 vdd gnd cell_6t
Xbit_r58_c152 bl_152 br_152 wl_58 vdd gnd cell_6t
Xbit_r59_c152 bl_152 br_152 wl_59 vdd gnd cell_6t
Xbit_r60_c152 bl_152 br_152 wl_60 vdd gnd cell_6t
Xbit_r61_c152 bl_152 br_152 wl_61 vdd gnd cell_6t
Xbit_r62_c152 bl_152 br_152 wl_62 vdd gnd cell_6t
Xbit_r63_c152 bl_152 br_152 wl_63 vdd gnd cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd cell_6t
Xbit_r1_c153 bl_153 br_153 wl_1 vdd gnd cell_6t
Xbit_r2_c153 bl_153 br_153 wl_2 vdd gnd cell_6t
Xbit_r3_c153 bl_153 br_153 wl_3 vdd gnd cell_6t
Xbit_r4_c153 bl_153 br_153 wl_4 vdd gnd cell_6t
Xbit_r5_c153 bl_153 br_153 wl_5 vdd gnd cell_6t
Xbit_r6_c153 bl_153 br_153 wl_6 vdd gnd cell_6t
Xbit_r7_c153 bl_153 br_153 wl_7 vdd gnd cell_6t
Xbit_r8_c153 bl_153 br_153 wl_8 vdd gnd cell_6t
Xbit_r9_c153 bl_153 br_153 wl_9 vdd gnd cell_6t
Xbit_r10_c153 bl_153 br_153 wl_10 vdd gnd cell_6t
Xbit_r11_c153 bl_153 br_153 wl_11 vdd gnd cell_6t
Xbit_r12_c153 bl_153 br_153 wl_12 vdd gnd cell_6t
Xbit_r13_c153 bl_153 br_153 wl_13 vdd gnd cell_6t
Xbit_r14_c153 bl_153 br_153 wl_14 vdd gnd cell_6t
Xbit_r15_c153 bl_153 br_153 wl_15 vdd gnd cell_6t
Xbit_r16_c153 bl_153 br_153 wl_16 vdd gnd cell_6t
Xbit_r17_c153 bl_153 br_153 wl_17 vdd gnd cell_6t
Xbit_r18_c153 bl_153 br_153 wl_18 vdd gnd cell_6t
Xbit_r19_c153 bl_153 br_153 wl_19 vdd gnd cell_6t
Xbit_r20_c153 bl_153 br_153 wl_20 vdd gnd cell_6t
Xbit_r21_c153 bl_153 br_153 wl_21 vdd gnd cell_6t
Xbit_r22_c153 bl_153 br_153 wl_22 vdd gnd cell_6t
Xbit_r23_c153 bl_153 br_153 wl_23 vdd gnd cell_6t
Xbit_r24_c153 bl_153 br_153 wl_24 vdd gnd cell_6t
Xbit_r25_c153 bl_153 br_153 wl_25 vdd gnd cell_6t
Xbit_r26_c153 bl_153 br_153 wl_26 vdd gnd cell_6t
Xbit_r27_c153 bl_153 br_153 wl_27 vdd gnd cell_6t
Xbit_r28_c153 bl_153 br_153 wl_28 vdd gnd cell_6t
Xbit_r29_c153 bl_153 br_153 wl_29 vdd gnd cell_6t
Xbit_r30_c153 bl_153 br_153 wl_30 vdd gnd cell_6t
Xbit_r31_c153 bl_153 br_153 wl_31 vdd gnd cell_6t
Xbit_r32_c153 bl_153 br_153 wl_32 vdd gnd cell_6t
Xbit_r33_c153 bl_153 br_153 wl_33 vdd gnd cell_6t
Xbit_r34_c153 bl_153 br_153 wl_34 vdd gnd cell_6t
Xbit_r35_c153 bl_153 br_153 wl_35 vdd gnd cell_6t
Xbit_r36_c153 bl_153 br_153 wl_36 vdd gnd cell_6t
Xbit_r37_c153 bl_153 br_153 wl_37 vdd gnd cell_6t
Xbit_r38_c153 bl_153 br_153 wl_38 vdd gnd cell_6t
Xbit_r39_c153 bl_153 br_153 wl_39 vdd gnd cell_6t
Xbit_r40_c153 bl_153 br_153 wl_40 vdd gnd cell_6t
Xbit_r41_c153 bl_153 br_153 wl_41 vdd gnd cell_6t
Xbit_r42_c153 bl_153 br_153 wl_42 vdd gnd cell_6t
Xbit_r43_c153 bl_153 br_153 wl_43 vdd gnd cell_6t
Xbit_r44_c153 bl_153 br_153 wl_44 vdd gnd cell_6t
Xbit_r45_c153 bl_153 br_153 wl_45 vdd gnd cell_6t
Xbit_r46_c153 bl_153 br_153 wl_46 vdd gnd cell_6t
Xbit_r47_c153 bl_153 br_153 wl_47 vdd gnd cell_6t
Xbit_r48_c153 bl_153 br_153 wl_48 vdd gnd cell_6t
Xbit_r49_c153 bl_153 br_153 wl_49 vdd gnd cell_6t
Xbit_r50_c153 bl_153 br_153 wl_50 vdd gnd cell_6t
Xbit_r51_c153 bl_153 br_153 wl_51 vdd gnd cell_6t
Xbit_r52_c153 bl_153 br_153 wl_52 vdd gnd cell_6t
Xbit_r53_c153 bl_153 br_153 wl_53 vdd gnd cell_6t
Xbit_r54_c153 bl_153 br_153 wl_54 vdd gnd cell_6t
Xbit_r55_c153 bl_153 br_153 wl_55 vdd gnd cell_6t
Xbit_r56_c153 bl_153 br_153 wl_56 vdd gnd cell_6t
Xbit_r57_c153 bl_153 br_153 wl_57 vdd gnd cell_6t
Xbit_r58_c153 bl_153 br_153 wl_58 vdd gnd cell_6t
Xbit_r59_c153 bl_153 br_153 wl_59 vdd gnd cell_6t
Xbit_r60_c153 bl_153 br_153 wl_60 vdd gnd cell_6t
Xbit_r61_c153 bl_153 br_153 wl_61 vdd gnd cell_6t
Xbit_r62_c153 bl_153 br_153 wl_62 vdd gnd cell_6t
Xbit_r63_c153 bl_153 br_153 wl_63 vdd gnd cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd cell_6t
Xbit_r1_c154 bl_154 br_154 wl_1 vdd gnd cell_6t
Xbit_r2_c154 bl_154 br_154 wl_2 vdd gnd cell_6t
Xbit_r3_c154 bl_154 br_154 wl_3 vdd gnd cell_6t
Xbit_r4_c154 bl_154 br_154 wl_4 vdd gnd cell_6t
Xbit_r5_c154 bl_154 br_154 wl_5 vdd gnd cell_6t
Xbit_r6_c154 bl_154 br_154 wl_6 vdd gnd cell_6t
Xbit_r7_c154 bl_154 br_154 wl_7 vdd gnd cell_6t
Xbit_r8_c154 bl_154 br_154 wl_8 vdd gnd cell_6t
Xbit_r9_c154 bl_154 br_154 wl_9 vdd gnd cell_6t
Xbit_r10_c154 bl_154 br_154 wl_10 vdd gnd cell_6t
Xbit_r11_c154 bl_154 br_154 wl_11 vdd gnd cell_6t
Xbit_r12_c154 bl_154 br_154 wl_12 vdd gnd cell_6t
Xbit_r13_c154 bl_154 br_154 wl_13 vdd gnd cell_6t
Xbit_r14_c154 bl_154 br_154 wl_14 vdd gnd cell_6t
Xbit_r15_c154 bl_154 br_154 wl_15 vdd gnd cell_6t
Xbit_r16_c154 bl_154 br_154 wl_16 vdd gnd cell_6t
Xbit_r17_c154 bl_154 br_154 wl_17 vdd gnd cell_6t
Xbit_r18_c154 bl_154 br_154 wl_18 vdd gnd cell_6t
Xbit_r19_c154 bl_154 br_154 wl_19 vdd gnd cell_6t
Xbit_r20_c154 bl_154 br_154 wl_20 vdd gnd cell_6t
Xbit_r21_c154 bl_154 br_154 wl_21 vdd gnd cell_6t
Xbit_r22_c154 bl_154 br_154 wl_22 vdd gnd cell_6t
Xbit_r23_c154 bl_154 br_154 wl_23 vdd gnd cell_6t
Xbit_r24_c154 bl_154 br_154 wl_24 vdd gnd cell_6t
Xbit_r25_c154 bl_154 br_154 wl_25 vdd gnd cell_6t
Xbit_r26_c154 bl_154 br_154 wl_26 vdd gnd cell_6t
Xbit_r27_c154 bl_154 br_154 wl_27 vdd gnd cell_6t
Xbit_r28_c154 bl_154 br_154 wl_28 vdd gnd cell_6t
Xbit_r29_c154 bl_154 br_154 wl_29 vdd gnd cell_6t
Xbit_r30_c154 bl_154 br_154 wl_30 vdd gnd cell_6t
Xbit_r31_c154 bl_154 br_154 wl_31 vdd gnd cell_6t
Xbit_r32_c154 bl_154 br_154 wl_32 vdd gnd cell_6t
Xbit_r33_c154 bl_154 br_154 wl_33 vdd gnd cell_6t
Xbit_r34_c154 bl_154 br_154 wl_34 vdd gnd cell_6t
Xbit_r35_c154 bl_154 br_154 wl_35 vdd gnd cell_6t
Xbit_r36_c154 bl_154 br_154 wl_36 vdd gnd cell_6t
Xbit_r37_c154 bl_154 br_154 wl_37 vdd gnd cell_6t
Xbit_r38_c154 bl_154 br_154 wl_38 vdd gnd cell_6t
Xbit_r39_c154 bl_154 br_154 wl_39 vdd gnd cell_6t
Xbit_r40_c154 bl_154 br_154 wl_40 vdd gnd cell_6t
Xbit_r41_c154 bl_154 br_154 wl_41 vdd gnd cell_6t
Xbit_r42_c154 bl_154 br_154 wl_42 vdd gnd cell_6t
Xbit_r43_c154 bl_154 br_154 wl_43 vdd gnd cell_6t
Xbit_r44_c154 bl_154 br_154 wl_44 vdd gnd cell_6t
Xbit_r45_c154 bl_154 br_154 wl_45 vdd gnd cell_6t
Xbit_r46_c154 bl_154 br_154 wl_46 vdd gnd cell_6t
Xbit_r47_c154 bl_154 br_154 wl_47 vdd gnd cell_6t
Xbit_r48_c154 bl_154 br_154 wl_48 vdd gnd cell_6t
Xbit_r49_c154 bl_154 br_154 wl_49 vdd gnd cell_6t
Xbit_r50_c154 bl_154 br_154 wl_50 vdd gnd cell_6t
Xbit_r51_c154 bl_154 br_154 wl_51 vdd gnd cell_6t
Xbit_r52_c154 bl_154 br_154 wl_52 vdd gnd cell_6t
Xbit_r53_c154 bl_154 br_154 wl_53 vdd gnd cell_6t
Xbit_r54_c154 bl_154 br_154 wl_54 vdd gnd cell_6t
Xbit_r55_c154 bl_154 br_154 wl_55 vdd gnd cell_6t
Xbit_r56_c154 bl_154 br_154 wl_56 vdd gnd cell_6t
Xbit_r57_c154 bl_154 br_154 wl_57 vdd gnd cell_6t
Xbit_r58_c154 bl_154 br_154 wl_58 vdd gnd cell_6t
Xbit_r59_c154 bl_154 br_154 wl_59 vdd gnd cell_6t
Xbit_r60_c154 bl_154 br_154 wl_60 vdd gnd cell_6t
Xbit_r61_c154 bl_154 br_154 wl_61 vdd gnd cell_6t
Xbit_r62_c154 bl_154 br_154 wl_62 vdd gnd cell_6t
Xbit_r63_c154 bl_154 br_154 wl_63 vdd gnd cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd cell_6t
Xbit_r1_c155 bl_155 br_155 wl_1 vdd gnd cell_6t
Xbit_r2_c155 bl_155 br_155 wl_2 vdd gnd cell_6t
Xbit_r3_c155 bl_155 br_155 wl_3 vdd gnd cell_6t
Xbit_r4_c155 bl_155 br_155 wl_4 vdd gnd cell_6t
Xbit_r5_c155 bl_155 br_155 wl_5 vdd gnd cell_6t
Xbit_r6_c155 bl_155 br_155 wl_6 vdd gnd cell_6t
Xbit_r7_c155 bl_155 br_155 wl_7 vdd gnd cell_6t
Xbit_r8_c155 bl_155 br_155 wl_8 vdd gnd cell_6t
Xbit_r9_c155 bl_155 br_155 wl_9 vdd gnd cell_6t
Xbit_r10_c155 bl_155 br_155 wl_10 vdd gnd cell_6t
Xbit_r11_c155 bl_155 br_155 wl_11 vdd gnd cell_6t
Xbit_r12_c155 bl_155 br_155 wl_12 vdd gnd cell_6t
Xbit_r13_c155 bl_155 br_155 wl_13 vdd gnd cell_6t
Xbit_r14_c155 bl_155 br_155 wl_14 vdd gnd cell_6t
Xbit_r15_c155 bl_155 br_155 wl_15 vdd gnd cell_6t
Xbit_r16_c155 bl_155 br_155 wl_16 vdd gnd cell_6t
Xbit_r17_c155 bl_155 br_155 wl_17 vdd gnd cell_6t
Xbit_r18_c155 bl_155 br_155 wl_18 vdd gnd cell_6t
Xbit_r19_c155 bl_155 br_155 wl_19 vdd gnd cell_6t
Xbit_r20_c155 bl_155 br_155 wl_20 vdd gnd cell_6t
Xbit_r21_c155 bl_155 br_155 wl_21 vdd gnd cell_6t
Xbit_r22_c155 bl_155 br_155 wl_22 vdd gnd cell_6t
Xbit_r23_c155 bl_155 br_155 wl_23 vdd gnd cell_6t
Xbit_r24_c155 bl_155 br_155 wl_24 vdd gnd cell_6t
Xbit_r25_c155 bl_155 br_155 wl_25 vdd gnd cell_6t
Xbit_r26_c155 bl_155 br_155 wl_26 vdd gnd cell_6t
Xbit_r27_c155 bl_155 br_155 wl_27 vdd gnd cell_6t
Xbit_r28_c155 bl_155 br_155 wl_28 vdd gnd cell_6t
Xbit_r29_c155 bl_155 br_155 wl_29 vdd gnd cell_6t
Xbit_r30_c155 bl_155 br_155 wl_30 vdd gnd cell_6t
Xbit_r31_c155 bl_155 br_155 wl_31 vdd gnd cell_6t
Xbit_r32_c155 bl_155 br_155 wl_32 vdd gnd cell_6t
Xbit_r33_c155 bl_155 br_155 wl_33 vdd gnd cell_6t
Xbit_r34_c155 bl_155 br_155 wl_34 vdd gnd cell_6t
Xbit_r35_c155 bl_155 br_155 wl_35 vdd gnd cell_6t
Xbit_r36_c155 bl_155 br_155 wl_36 vdd gnd cell_6t
Xbit_r37_c155 bl_155 br_155 wl_37 vdd gnd cell_6t
Xbit_r38_c155 bl_155 br_155 wl_38 vdd gnd cell_6t
Xbit_r39_c155 bl_155 br_155 wl_39 vdd gnd cell_6t
Xbit_r40_c155 bl_155 br_155 wl_40 vdd gnd cell_6t
Xbit_r41_c155 bl_155 br_155 wl_41 vdd gnd cell_6t
Xbit_r42_c155 bl_155 br_155 wl_42 vdd gnd cell_6t
Xbit_r43_c155 bl_155 br_155 wl_43 vdd gnd cell_6t
Xbit_r44_c155 bl_155 br_155 wl_44 vdd gnd cell_6t
Xbit_r45_c155 bl_155 br_155 wl_45 vdd gnd cell_6t
Xbit_r46_c155 bl_155 br_155 wl_46 vdd gnd cell_6t
Xbit_r47_c155 bl_155 br_155 wl_47 vdd gnd cell_6t
Xbit_r48_c155 bl_155 br_155 wl_48 vdd gnd cell_6t
Xbit_r49_c155 bl_155 br_155 wl_49 vdd gnd cell_6t
Xbit_r50_c155 bl_155 br_155 wl_50 vdd gnd cell_6t
Xbit_r51_c155 bl_155 br_155 wl_51 vdd gnd cell_6t
Xbit_r52_c155 bl_155 br_155 wl_52 vdd gnd cell_6t
Xbit_r53_c155 bl_155 br_155 wl_53 vdd gnd cell_6t
Xbit_r54_c155 bl_155 br_155 wl_54 vdd gnd cell_6t
Xbit_r55_c155 bl_155 br_155 wl_55 vdd gnd cell_6t
Xbit_r56_c155 bl_155 br_155 wl_56 vdd gnd cell_6t
Xbit_r57_c155 bl_155 br_155 wl_57 vdd gnd cell_6t
Xbit_r58_c155 bl_155 br_155 wl_58 vdd gnd cell_6t
Xbit_r59_c155 bl_155 br_155 wl_59 vdd gnd cell_6t
Xbit_r60_c155 bl_155 br_155 wl_60 vdd gnd cell_6t
Xbit_r61_c155 bl_155 br_155 wl_61 vdd gnd cell_6t
Xbit_r62_c155 bl_155 br_155 wl_62 vdd gnd cell_6t
Xbit_r63_c155 bl_155 br_155 wl_63 vdd gnd cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd cell_6t
Xbit_r1_c156 bl_156 br_156 wl_1 vdd gnd cell_6t
Xbit_r2_c156 bl_156 br_156 wl_2 vdd gnd cell_6t
Xbit_r3_c156 bl_156 br_156 wl_3 vdd gnd cell_6t
Xbit_r4_c156 bl_156 br_156 wl_4 vdd gnd cell_6t
Xbit_r5_c156 bl_156 br_156 wl_5 vdd gnd cell_6t
Xbit_r6_c156 bl_156 br_156 wl_6 vdd gnd cell_6t
Xbit_r7_c156 bl_156 br_156 wl_7 vdd gnd cell_6t
Xbit_r8_c156 bl_156 br_156 wl_8 vdd gnd cell_6t
Xbit_r9_c156 bl_156 br_156 wl_9 vdd gnd cell_6t
Xbit_r10_c156 bl_156 br_156 wl_10 vdd gnd cell_6t
Xbit_r11_c156 bl_156 br_156 wl_11 vdd gnd cell_6t
Xbit_r12_c156 bl_156 br_156 wl_12 vdd gnd cell_6t
Xbit_r13_c156 bl_156 br_156 wl_13 vdd gnd cell_6t
Xbit_r14_c156 bl_156 br_156 wl_14 vdd gnd cell_6t
Xbit_r15_c156 bl_156 br_156 wl_15 vdd gnd cell_6t
Xbit_r16_c156 bl_156 br_156 wl_16 vdd gnd cell_6t
Xbit_r17_c156 bl_156 br_156 wl_17 vdd gnd cell_6t
Xbit_r18_c156 bl_156 br_156 wl_18 vdd gnd cell_6t
Xbit_r19_c156 bl_156 br_156 wl_19 vdd gnd cell_6t
Xbit_r20_c156 bl_156 br_156 wl_20 vdd gnd cell_6t
Xbit_r21_c156 bl_156 br_156 wl_21 vdd gnd cell_6t
Xbit_r22_c156 bl_156 br_156 wl_22 vdd gnd cell_6t
Xbit_r23_c156 bl_156 br_156 wl_23 vdd gnd cell_6t
Xbit_r24_c156 bl_156 br_156 wl_24 vdd gnd cell_6t
Xbit_r25_c156 bl_156 br_156 wl_25 vdd gnd cell_6t
Xbit_r26_c156 bl_156 br_156 wl_26 vdd gnd cell_6t
Xbit_r27_c156 bl_156 br_156 wl_27 vdd gnd cell_6t
Xbit_r28_c156 bl_156 br_156 wl_28 vdd gnd cell_6t
Xbit_r29_c156 bl_156 br_156 wl_29 vdd gnd cell_6t
Xbit_r30_c156 bl_156 br_156 wl_30 vdd gnd cell_6t
Xbit_r31_c156 bl_156 br_156 wl_31 vdd gnd cell_6t
Xbit_r32_c156 bl_156 br_156 wl_32 vdd gnd cell_6t
Xbit_r33_c156 bl_156 br_156 wl_33 vdd gnd cell_6t
Xbit_r34_c156 bl_156 br_156 wl_34 vdd gnd cell_6t
Xbit_r35_c156 bl_156 br_156 wl_35 vdd gnd cell_6t
Xbit_r36_c156 bl_156 br_156 wl_36 vdd gnd cell_6t
Xbit_r37_c156 bl_156 br_156 wl_37 vdd gnd cell_6t
Xbit_r38_c156 bl_156 br_156 wl_38 vdd gnd cell_6t
Xbit_r39_c156 bl_156 br_156 wl_39 vdd gnd cell_6t
Xbit_r40_c156 bl_156 br_156 wl_40 vdd gnd cell_6t
Xbit_r41_c156 bl_156 br_156 wl_41 vdd gnd cell_6t
Xbit_r42_c156 bl_156 br_156 wl_42 vdd gnd cell_6t
Xbit_r43_c156 bl_156 br_156 wl_43 vdd gnd cell_6t
Xbit_r44_c156 bl_156 br_156 wl_44 vdd gnd cell_6t
Xbit_r45_c156 bl_156 br_156 wl_45 vdd gnd cell_6t
Xbit_r46_c156 bl_156 br_156 wl_46 vdd gnd cell_6t
Xbit_r47_c156 bl_156 br_156 wl_47 vdd gnd cell_6t
Xbit_r48_c156 bl_156 br_156 wl_48 vdd gnd cell_6t
Xbit_r49_c156 bl_156 br_156 wl_49 vdd gnd cell_6t
Xbit_r50_c156 bl_156 br_156 wl_50 vdd gnd cell_6t
Xbit_r51_c156 bl_156 br_156 wl_51 vdd gnd cell_6t
Xbit_r52_c156 bl_156 br_156 wl_52 vdd gnd cell_6t
Xbit_r53_c156 bl_156 br_156 wl_53 vdd gnd cell_6t
Xbit_r54_c156 bl_156 br_156 wl_54 vdd gnd cell_6t
Xbit_r55_c156 bl_156 br_156 wl_55 vdd gnd cell_6t
Xbit_r56_c156 bl_156 br_156 wl_56 vdd gnd cell_6t
Xbit_r57_c156 bl_156 br_156 wl_57 vdd gnd cell_6t
Xbit_r58_c156 bl_156 br_156 wl_58 vdd gnd cell_6t
Xbit_r59_c156 bl_156 br_156 wl_59 vdd gnd cell_6t
Xbit_r60_c156 bl_156 br_156 wl_60 vdd gnd cell_6t
Xbit_r61_c156 bl_156 br_156 wl_61 vdd gnd cell_6t
Xbit_r62_c156 bl_156 br_156 wl_62 vdd gnd cell_6t
Xbit_r63_c156 bl_156 br_156 wl_63 vdd gnd cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd cell_6t
Xbit_r1_c157 bl_157 br_157 wl_1 vdd gnd cell_6t
Xbit_r2_c157 bl_157 br_157 wl_2 vdd gnd cell_6t
Xbit_r3_c157 bl_157 br_157 wl_3 vdd gnd cell_6t
Xbit_r4_c157 bl_157 br_157 wl_4 vdd gnd cell_6t
Xbit_r5_c157 bl_157 br_157 wl_5 vdd gnd cell_6t
Xbit_r6_c157 bl_157 br_157 wl_6 vdd gnd cell_6t
Xbit_r7_c157 bl_157 br_157 wl_7 vdd gnd cell_6t
Xbit_r8_c157 bl_157 br_157 wl_8 vdd gnd cell_6t
Xbit_r9_c157 bl_157 br_157 wl_9 vdd gnd cell_6t
Xbit_r10_c157 bl_157 br_157 wl_10 vdd gnd cell_6t
Xbit_r11_c157 bl_157 br_157 wl_11 vdd gnd cell_6t
Xbit_r12_c157 bl_157 br_157 wl_12 vdd gnd cell_6t
Xbit_r13_c157 bl_157 br_157 wl_13 vdd gnd cell_6t
Xbit_r14_c157 bl_157 br_157 wl_14 vdd gnd cell_6t
Xbit_r15_c157 bl_157 br_157 wl_15 vdd gnd cell_6t
Xbit_r16_c157 bl_157 br_157 wl_16 vdd gnd cell_6t
Xbit_r17_c157 bl_157 br_157 wl_17 vdd gnd cell_6t
Xbit_r18_c157 bl_157 br_157 wl_18 vdd gnd cell_6t
Xbit_r19_c157 bl_157 br_157 wl_19 vdd gnd cell_6t
Xbit_r20_c157 bl_157 br_157 wl_20 vdd gnd cell_6t
Xbit_r21_c157 bl_157 br_157 wl_21 vdd gnd cell_6t
Xbit_r22_c157 bl_157 br_157 wl_22 vdd gnd cell_6t
Xbit_r23_c157 bl_157 br_157 wl_23 vdd gnd cell_6t
Xbit_r24_c157 bl_157 br_157 wl_24 vdd gnd cell_6t
Xbit_r25_c157 bl_157 br_157 wl_25 vdd gnd cell_6t
Xbit_r26_c157 bl_157 br_157 wl_26 vdd gnd cell_6t
Xbit_r27_c157 bl_157 br_157 wl_27 vdd gnd cell_6t
Xbit_r28_c157 bl_157 br_157 wl_28 vdd gnd cell_6t
Xbit_r29_c157 bl_157 br_157 wl_29 vdd gnd cell_6t
Xbit_r30_c157 bl_157 br_157 wl_30 vdd gnd cell_6t
Xbit_r31_c157 bl_157 br_157 wl_31 vdd gnd cell_6t
Xbit_r32_c157 bl_157 br_157 wl_32 vdd gnd cell_6t
Xbit_r33_c157 bl_157 br_157 wl_33 vdd gnd cell_6t
Xbit_r34_c157 bl_157 br_157 wl_34 vdd gnd cell_6t
Xbit_r35_c157 bl_157 br_157 wl_35 vdd gnd cell_6t
Xbit_r36_c157 bl_157 br_157 wl_36 vdd gnd cell_6t
Xbit_r37_c157 bl_157 br_157 wl_37 vdd gnd cell_6t
Xbit_r38_c157 bl_157 br_157 wl_38 vdd gnd cell_6t
Xbit_r39_c157 bl_157 br_157 wl_39 vdd gnd cell_6t
Xbit_r40_c157 bl_157 br_157 wl_40 vdd gnd cell_6t
Xbit_r41_c157 bl_157 br_157 wl_41 vdd gnd cell_6t
Xbit_r42_c157 bl_157 br_157 wl_42 vdd gnd cell_6t
Xbit_r43_c157 bl_157 br_157 wl_43 vdd gnd cell_6t
Xbit_r44_c157 bl_157 br_157 wl_44 vdd gnd cell_6t
Xbit_r45_c157 bl_157 br_157 wl_45 vdd gnd cell_6t
Xbit_r46_c157 bl_157 br_157 wl_46 vdd gnd cell_6t
Xbit_r47_c157 bl_157 br_157 wl_47 vdd gnd cell_6t
Xbit_r48_c157 bl_157 br_157 wl_48 vdd gnd cell_6t
Xbit_r49_c157 bl_157 br_157 wl_49 vdd gnd cell_6t
Xbit_r50_c157 bl_157 br_157 wl_50 vdd gnd cell_6t
Xbit_r51_c157 bl_157 br_157 wl_51 vdd gnd cell_6t
Xbit_r52_c157 bl_157 br_157 wl_52 vdd gnd cell_6t
Xbit_r53_c157 bl_157 br_157 wl_53 vdd gnd cell_6t
Xbit_r54_c157 bl_157 br_157 wl_54 vdd gnd cell_6t
Xbit_r55_c157 bl_157 br_157 wl_55 vdd gnd cell_6t
Xbit_r56_c157 bl_157 br_157 wl_56 vdd gnd cell_6t
Xbit_r57_c157 bl_157 br_157 wl_57 vdd gnd cell_6t
Xbit_r58_c157 bl_157 br_157 wl_58 vdd gnd cell_6t
Xbit_r59_c157 bl_157 br_157 wl_59 vdd gnd cell_6t
Xbit_r60_c157 bl_157 br_157 wl_60 vdd gnd cell_6t
Xbit_r61_c157 bl_157 br_157 wl_61 vdd gnd cell_6t
Xbit_r62_c157 bl_157 br_157 wl_62 vdd gnd cell_6t
Xbit_r63_c157 bl_157 br_157 wl_63 vdd gnd cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd cell_6t
Xbit_r1_c158 bl_158 br_158 wl_1 vdd gnd cell_6t
Xbit_r2_c158 bl_158 br_158 wl_2 vdd gnd cell_6t
Xbit_r3_c158 bl_158 br_158 wl_3 vdd gnd cell_6t
Xbit_r4_c158 bl_158 br_158 wl_4 vdd gnd cell_6t
Xbit_r5_c158 bl_158 br_158 wl_5 vdd gnd cell_6t
Xbit_r6_c158 bl_158 br_158 wl_6 vdd gnd cell_6t
Xbit_r7_c158 bl_158 br_158 wl_7 vdd gnd cell_6t
Xbit_r8_c158 bl_158 br_158 wl_8 vdd gnd cell_6t
Xbit_r9_c158 bl_158 br_158 wl_9 vdd gnd cell_6t
Xbit_r10_c158 bl_158 br_158 wl_10 vdd gnd cell_6t
Xbit_r11_c158 bl_158 br_158 wl_11 vdd gnd cell_6t
Xbit_r12_c158 bl_158 br_158 wl_12 vdd gnd cell_6t
Xbit_r13_c158 bl_158 br_158 wl_13 vdd gnd cell_6t
Xbit_r14_c158 bl_158 br_158 wl_14 vdd gnd cell_6t
Xbit_r15_c158 bl_158 br_158 wl_15 vdd gnd cell_6t
Xbit_r16_c158 bl_158 br_158 wl_16 vdd gnd cell_6t
Xbit_r17_c158 bl_158 br_158 wl_17 vdd gnd cell_6t
Xbit_r18_c158 bl_158 br_158 wl_18 vdd gnd cell_6t
Xbit_r19_c158 bl_158 br_158 wl_19 vdd gnd cell_6t
Xbit_r20_c158 bl_158 br_158 wl_20 vdd gnd cell_6t
Xbit_r21_c158 bl_158 br_158 wl_21 vdd gnd cell_6t
Xbit_r22_c158 bl_158 br_158 wl_22 vdd gnd cell_6t
Xbit_r23_c158 bl_158 br_158 wl_23 vdd gnd cell_6t
Xbit_r24_c158 bl_158 br_158 wl_24 vdd gnd cell_6t
Xbit_r25_c158 bl_158 br_158 wl_25 vdd gnd cell_6t
Xbit_r26_c158 bl_158 br_158 wl_26 vdd gnd cell_6t
Xbit_r27_c158 bl_158 br_158 wl_27 vdd gnd cell_6t
Xbit_r28_c158 bl_158 br_158 wl_28 vdd gnd cell_6t
Xbit_r29_c158 bl_158 br_158 wl_29 vdd gnd cell_6t
Xbit_r30_c158 bl_158 br_158 wl_30 vdd gnd cell_6t
Xbit_r31_c158 bl_158 br_158 wl_31 vdd gnd cell_6t
Xbit_r32_c158 bl_158 br_158 wl_32 vdd gnd cell_6t
Xbit_r33_c158 bl_158 br_158 wl_33 vdd gnd cell_6t
Xbit_r34_c158 bl_158 br_158 wl_34 vdd gnd cell_6t
Xbit_r35_c158 bl_158 br_158 wl_35 vdd gnd cell_6t
Xbit_r36_c158 bl_158 br_158 wl_36 vdd gnd cell_6t
Xbit_r37_c158 bl_158 br_158 wl_37 vdd gnd cell_6t
Xbit_r38_c158 bl_158 br_158 wl_38 vdd gnd cell_6t
Xbit_r39_c158 bl_158 br_158 wl_39 vdd gnd cell_6t
Xbit_r40_c158 bl_158 br_158 wl_40 vdd gnd cell_6t
Xbit_r41_c158 bl_158 br_158 wl_41 vdd gnd cell_6t
Xbit_r42_c158 bl_158 br_158 wl_42 vdd gnd cell_6t
Xbit_r43_c158 bl_158 br_158 wl_43 vdd gnd cell_6t
Xbit_r44_c158 bl_158 br_158 wl_44 vdd gnd cell_6t
Xbit_r45_c158 bl_158 br_158 wl_45 vdd gnd cell_6t
Xbit_r46_c158 bl_158 br_158 wl_46 vdd gnd cell_6t
Xbit_r47_c158 bl_158 br_158 wl_47 vdd gnd cell_6t
Xbit_r48_c158 bl_158 br_158 wl_48 vdd gnd cell_6t
Xbit_r49_c158 bl_158 br_158 wl_49 vdd gnd cell_6t
Xbit_r50_c158 bl_158 br_158 wl_50 vdd gnd cell_6t
Xbit_r51_c158 bl_158 br_158 wl_51 vdd gnd cell_6t
Xbit_r52_c158 bl_158 br_158 wl_52 vdd gnd cell_6t
Xbit_r53_c158 bl_158 br_158 wl_53 vdd gnd cell_6t
Xbit_r54_c158 bl_158 br_158 wl_54 vdd gnd cell_6t
Xbit_r55_c158 bl_158 br_158 wl_55 vdd gnd cell_6t
Xbit_r56_c158 bl_158 br_158 wl_56 vdd gnd cell_6t
Xbit_r57_c158 bl_158 br_158 wl_57 vdd gnd cell_6t
Xbit_r58_c158 bl_158 br_158 wl_58 vdd gnd cell_6t
Xbit_r59_c158 bl_158 br_158 wl_59 vdd gnd cell_6t
Xbit_r60_c158 bl_158 br_158 wl_60 vdd gnd cell_6t
Xbit_r61_c158 bl_158 br_158 wl_61 vdd gnd cell_6t
Xbit_r62_c158 bl_158 br_158 wl_62 vdd gnd cell_6t
Xbit_r63_c158 bl_158 br_158 wl_63 vdd gnd cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd cell_6t
Xbit_r1_c159 bl_159 br_159 wl_1 vdd gnd cell_6t
Xbit_r2_c159 bl_159 br_159 wl_2 vdd gnd cell_6t
Xbit_r3_c159 bl_159 br_159 wl_3 vdd gnd cell_6t
Xbit_r4_c159 bl_159 br_159 wl_4 vdd gnd cell_6t
Xbit_r5_c159 bl_159 br_159 wl_5 vdd gnd cell_6t
Xbit_r6_c159 bl_159 br_159 wl_6 vdd gnd cell_6t
Xbit_r7_c159 bl_159 br_159 wl_7 vdd gnd cell_6t
Xbit_r8_c159 bl_159 br_159 wl_8 vdd gnd cell_6t
Xbit_r9_c159 bl_159 br_159 wl_9 vdd gnd cell_6t
Xbit_r10_c159 bl_159 br_159 wl_10 vdd gnd cell_6t
Xbit_r11_c159 bl_159 br_159 wl_11 vdd gnd cell_6t
Xbit_r12_c159 bl_159 br_159 wl_12 vdd gnd cell_6t
Xbit_r13_c159 bl_159 br_159 wl_13 vdd gnd cell_6t
Xbit_r14_c159 bl_159 br_159 wl_14 vdd gnd cell_6t
Xbit_r15_c159 bl_159 br_159 wl_15 vdd gnd cell_6t
Xbit_r16_c159 bl_159 br_159 wl_16 vdd gnd cell_6t
Xbit_r17_c159 bl_159 br_159 wl_17 vdd gnd cell_6t
Xbit_r18_c159 bl_159 br_159 wl_18 vdd gnd cell_6t
Xbit_r19_c159 bl_159 br_159 wl_19 vdd gnd cell_6t
Xbit_r20_c159 bl_159 br_159 wl_20 vdd gnd cell_6t
Xbit_r21_c159 bl_159 br_159 wl_21 vdd gnd cell_6t
Xbit_r22_c159 bl_159 br_159 wl_22 vdd gnd cell_6t
Xbit_r23_c159 bl_159 br_159 wl_23 vdd gnd cell_6t
Xbit_r24_c159 bl_159 br_159 wl_24 vdd gnd cell_6t
Xbit_r25_c159 bl_159 br_159 wl_25 vdd gnd cell_6t
Xbit_r26_c159 bl_159 br_159 wl_26 vdd gnd cell_6t
Xbit_r27_c159 bl_159 br_159 wl_27 vdd gnd cell_6t
Xbit_r28_c159 bl_159 br_159 wl_28 vdd gnd cell_6t
Xbit_r29_c159 bl_159 br_159 wl_29 vdd gnd cell_6t
Xbit_r30_c159 bl_159 br_159 wl_30 vdd gnd cell_6t
Xbit_r31_c159 bl_159 br_159 wl_31 vdd gnd cell_6t
Xbit_r32_c159 bl_159 br_159 wl_32 vdd gnd cell_6t
Xbit_r33_c159 bl_159 br_159 wl_33 vdd gnd cell_6t
Xbit_r34_c159 bl_159 br_159 wl_34 vdd gnd cell_6t
Xbit_r35_c159 bl_159 br_159 wl_35 vdd gnd cell_6t
Xbit_r36_c159 bl_159 br_159 wl_36 vdd gnd cell_6t
Xbit_r37_c159 bl_159 br_159 wl_37 vdd gnd cell_6t
Xbit_r38_c159 bl_159 br_159 wl_38 vdd gnd cell_6t
Xbit_r39_c159 bl_159 br_159 wl_39 vdd gnd cell_6t
Xbit_r40_c159 bl_159 br_159 wl_40 vdd gnd cell_6t
Xbit_r41_c159 bl_159 br_159 wl_41 vdd gnd cell_6t
Xbit_r42_c159 bl_159 br_159 wl_42 vdd gnd cell_6t
Xbit_r43_c159 bl_159 br_159 wl_43 vdd gnd cell_6t
Xbit_r44_c159 bl_159 br_159 wl_44 vdd gnd cell_6t
Xbit_r45_c159 bl_159 br_159 wl_45 vdd gnd cell_6t
Xbit_r46_c159 bl_159 br_159 wl_46 vdd gnd cell_6t
Xbit_r47_c159 bl_159 br_159 wl_47 vdd gnd cell_6t
Xbit_r48_c159 bl_159 br_159 wl_48 vdd gnd cell_6t
Xbit_r49_c159 bl_159 br_159 wl_49 vdd gnd cell_6t
Xbit_r50_c159 bl_159 br_159 wl_50 vdd gnd cell_6t
Xbit_r51_c159 bl_159 br_159 wl_51 vdd gnd cell_6t
Xbit_r52_c159 bl_159 br_159 wl_52 vdd gnd cell_6t
Xbit_r53_c159 bl_159 br_159 wl_53 vdd gnd cell_6t
Xbit_r54_c159 bl_159 br_159 wl_54 vdd gnd cell_6t
Xbit_r55_c159 bl_159 br_159 wl_55 vdd gnd cell_6t
Xbit_r56_c159 bl_159 br_159 wl_56 vdd gnd cell_6t
Xbit_r57_c159 bl_159 br_159 wl_57 vdd gnd cell_6t
Xbit_r58_c159 bl_159 br_159 wl_58 vdd gnd cell_6t
Xbit_r59_c159 bl_159 br_159 wl_59 vdd gnd cell_6t
Xbit_r60_c159 bl_159 br_159 wl_60 vdd gnd cell_6t
Xbit_r61_c159 bl_159 br_159 wl_61 vdd gnd cell_6t
Xbit_r62_c159 bl_159 br_159 wl_62 vdd gnd cell_6t
Xbit_r63_c159 bl_159 br_159 wl_63 vdd gnd cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd cell_6t
Xbit_r1_c160 bl_160 br_160 wl_1 vdd gnd cell_6t
Xbit_r2_c160 bl_160 br_160 wl_2 vdd gnd cell_6t
Xbit_r3_c160 bl_160 br_160 wl_3 vdd gnd cell_6t
Xbit_r4_c160 bl_160 br_160 wl_4 vdd gnd cell_6t
Xbit_r5_c160 bl_160 br_160 wl_5 vdd gnd cell_6t
Xbit_r6_c160 bl_160 br_160 wl_6 vdd gnd cell_6t
Xbit_r7_c160 bl_160 br_160 wl_7 vdd gnd cell_6t
Xbit_r8_c160 bl_160 br_160 wl_8 vdd gnd cell_6t
Xbit_r9_c160 bl_160 br_160 wl_9 vdd gnd cell_6t
Xbit_r10_c160 bl_160 br_160 wl_10 vdd gnd cell_6t
Xbit_r11_c160 bl_160 br_160 wl_11 vdd gnd cell_6t
Xbit_r12_c160 bl_160 br_160 wl_12 vdd gnd cell_6t
Xbit_r13_c160 bl_160 br_160 wl_13 vdd gnd cell_6t
Xbit_r14_c160 bl_160 br_160 wl_14 vdd gnd cell_6t
Xbit_r15_c160 bl_160 br_160 wl_15 vdd gnd cell_6t
Xbit_r16_c160 bl_160 br_160 wl_16 vdd gnd cell_6t
Xbit_r17_c160 bl_160 br_160 wl_17 vdd gnd cell_6t
Xbit_r18_c160 bl_160 br_160 wl_18 vdd gnd cell_6t
Xbit_r19_c160 bl_160 br_160 wl_19 vdd gnd cell_6t
Xbit_r20_c160 bl_160 br_160 wl_20 vdd gnd cell_6t
Xbit_r21_c160 bl_160 br_160 wl_21 vdd gnd cell_6t
Xbit_r22_c160 bl_160 br_160 wl_22 vdd gnd cell_6t
Xbit_r23_c160 bl_160 br_160 wl_23 vdd gnd cell_6t
Xbit_r24_c160 bl_160 br_160 wl_24 vdd gnd cell_6t
Xbit_r25_c160 bl_160 br_160 wl_25 vdd gnd cell_6t
Xbit_r26_c160 bl_160 br_160 wl_26 vdd gnd cell_6t
Xbit_r27_c160 bl_160 br_160 wl_27 vdd gnd cell_6t
Xbit_r28_c160 bl_160 br_160 wl_28 vdd gnd cell_6t
Xbit_r29_c160 bl_160 br_160 wl_29 vdd gnd cell_6t
Xbit_r30_c160 bl_160 br_160 wl_30 vdd gnd cell_6t
Xbit_r31_c160 bl_160 br_160 wl_31 vdd gnd cell_6t
Xbit_r32_c160 bl_160 br_160 wl_32 vdd gnd cell_6t
Xbit_r33_c160 bl_160 br_160 wl_33 vdd gnd cell_6t
Xbit_r34_c160 bl_160 br_160 wl_34 vdd gnd cell_6t
Xbit_r35_c160 bl_160 br_160 wl_35 vdd gnd cell_6t
Xbit_r36_c160 bl_160 br_160 wl_36 vdd gnd cell_6t
Xbit_r37_c160 bl_160 br_160 wl_37 vdd gnd cell_6t
Xbit_r38_c160 bl_160 br_160 wl_38 vdd gnd cell_6t
Xbit_r39_c160 bl_160 br_160 wl_39 vdd gnd cell_6t
Xbit_r40_c160 bl_160 br_160 wl_40 vdd gnd cell_6t
Xbit_r41_c160 bl_160 br_160 wl_41 vdd gnd cell_6t
Xbit_r42_c160 bl_160 br_160 wl_42 vdd gnd cell_6t
Xbit_r43_c160 bl_160 br_160 wl_43 vdd gnd cell_6t
Xbit_r44_c160 bl_160 br_160 wl_44 vdd gnd cell_6t
Xbit_r45_c160 bl_160 br_160 wl_45 vdd gnd cell_6t
Xbit_r46_c160 bl_160 br_160 wl_46 vdd gnd cell_6t
Xbit_r47_c160 bl_160 br_160 wl_47 vdd gnd cell_6t
Xbit_r48_c160 bl_160 br_160 wl_48 vdd gnd cell_6t
Xbit_r49_c160 bl_160 br_160 wl_49 vdd gnd cell_6t
Xbit_r50_c160 bl_160 br_160 wl_50 vdd gnd cell_6t
Xbit_r51_c160 bl_160 br_160 wl_51 vdd gnd cell_6t
Xbit_r52_c160 bl_160 br_160 wl_52 vdd gnd cell_6t
Xbit_r53_c160 bl_160 br_160 wl_53 vdd gnd cell_6t
Xbit_r54_c160 bl_160 br_160 wl_54 vdd gnd cell_6t
Xbit_r55_c160 bl_160 br_160 wl_55 vdd gnd cell_6t
Xbit_r56_c160 bl_160 br_160 wl_56 vdd gnd cell_6t
Xbit_r57_c160 bl_160 br_160 wl_57 vdd gnd cell_6t
Xbit_r58_c160 bl_160 br_160 wl_58 vdd gnd cell_6t
Xbit_r59_c160 bl_160 br_160 wl_59 vdd gnd cell_6t
Xbit_r60_c160 bl_160 br_160 wl_60 vdd gnd cell_6t
Xbit_r61_c160 bl_160 br_160 wl_61 vdd gnd cell_6t
Xbit_r62_c160 bl_160 br_160 wl_62 vdd gnd cell_6t
Xbit_r63_c160 bl_160 br_160 wl_63 vdd gnd cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd cell_6t
Xbit_r1_c161 bl_161 br_161 wl_1 vdd gnd cell_6t
Xbit_r2_c161 bl_161 br_161 wl_2 vdd gnd cell_6t
Xbit_r3_c161 bl_161 br_161 wl_3 vdd gnd cell_6t
Xbit_r4_c161 bl_161 br_161 wl_4 vdd gnd cell_6t
Xbit_r5_c161 bl_161 br_161 wl_5 vdd gnd cell_6t
Xbit_r6_c161 bl_161 br_161 wl_6 vdd gnd cell_6t
Xbit_r7_c161 bl_161 br_161 wl_7 vdd gnd cell_6t
Xbit_r8_c161 bl_161 br_161 wl_8 vdd gnd cell_6t
Xbit_r9_c161 bl_161 br_161 wl_9 vdd gnd cell_6t
Xbit_r10_c161 bl_161 br_161 wl_10 vdd gnd cell_6t
Xbit_r11_c161 bl_161 br_161 wl_11 vdd gnd cell_6t
Xbit_r12_c161 bl_161 br_161 wl_12 vdd gnd cell_6t
Xbit_r13_c161 bl_161 br_161 wl_13 vdd gnd cell_6t
Xbit_r14_c161 bl_161 br_161 wl_14 vdd gnd cell_6t
Xbit_r15_c161 bl_161 br_161 wl_15 vdd gnd cell_6t
Xbit_r16_c161 bl_161 br_161 wl_16 vdd gnd cell_6t
Xbit_r17_c161 bl_161 br_161 wl_17 vdd gnd cell_6t
Xbit_r18_c161 bl_161 br_161 wl_18 vdd gnd cell_6t
Xbit_r19_c161 bl_161 br_161 wl_19 vdd gnd cell_6t
Xbit_r20_c161 bl_161 br_161 wl_20 vdd gnd cell_6t
Xbit_r21_c161 bl_161 br_161 wl_21 vdd gnd cell_6t
Xbit_r22_c161 bl_161 br_161 wl_22 vdd gnd cell_6t
Xbit_r23_c161 bl_161 br_161 wl_23 vdd gnd cell_6t
Xbit_r24_c161 bl_161 br_161 wl_24 vdd gnd cell_6t
Xbit_r25_c161 bl_161 br_161 wl_25 vdd gnd cell_6t
Xbit_r26_c161 bl_161 br_161 wl_26 vdd gnd cell_6t
Xbit_r27_c161 bl_161 br_161 wl_27 vdd gnd cell_6t
Xbit_r28_c161 bl_161 br_161 wl_28 vdd gnd cell_6t
Xbit_r29_c161 bl_161 br_161 wl_29 vdd gnd cell_6t
Xbit_r30_c161 bl_161 br_161 wl_30 vdd gnd cell_6t
Xbit_r31_c161 bl_161 br_161 wl_31 vdd gnd cell_6t
Xbit_r32_c161 bl_161 br_161 wl_32 vdd gnd cell_6t
Xbit_r33_c161 bl_161 br_161 wl_33 vdd gnd cell_6t
Xbit_r34_c161 bl_161 br_161 wl_34 vdd gnd cell_6t
Xbit_r35_c161 bl_161 br_161 wl_35 vdd gnd cell_6t
Xbit_r36_c161 bl_161 br_161 wl_36 vdd gnd cell_6t
Xbit_r37_c161 bl_161 br_161 wl_37 vdd gnd cell_6t
Xbit_r38_c161 bl_161 br_161 wl_38 vdd gnd cell_6t
Xbit_r39_c161 bl_161 br_161 wl_39 vdd gnd cell_6t
Xbit_r40_c161 bl_161 br_161 wl_40 vdd gnd cell_6t
Xbit_r41_c161 bl_161 br_161 wl_41 vdd gnd cell_6t
Xbit_r42_c161 bl_161 br_161 wl_42 vdd gnd cell_6t
Xbit_r43_c161 bl_161 br_161 wl_43 vdd gnd cell_6t
Xbit_r44_c161 bl_161 br_161 wl_44 vdd gnd cell_6t
Xbit_r45_c161 bl_161 br_161 wl_45 vdd gnd cell_6t
Xbit_r46_c161 bl_161 br_161 wl_46 vdd gnd cell_6t
Xbit_r47_c161 bl_161 br_161 wl_47 vdd gnd cell_6t
Xbit_r48_c161 bl_161 br_161 wl_48 vdd gnd cell_6t
Xbit_r49_c161 bl_161 br_161 wl_49 vdd gnd cell_6t
Xbit_r50_c161 bl_161 br_161 wl_50 vdd gnd cell_6t
Xbit_r51_c161 bl_161 br_161 wl_51 vdd gnd cell_6t
Xbit_r52_c161 bl_161 br_161 wl_52 vdd gnd cell_6t
Xbit_r53_c161 bl_161 br_161 wl_53 vdd gnd cell_6t
Xbit_r54_c161 bl_161 br_161 wl_54 vdd gnd cell_6t
Xbit_r55_c161 bl_161 br_161 wl_55 vdd gnd cell_6t
Xbit_r56_c161 bl_161 br_161 wl_56 vdd gnd cell_6t
Xbit_r57_c161 bl_161 br_161 wl_57 vdd gnd cell_6t
Xbit_r58_c161 bl_161 br_161 wl_58 vdd gnd cell_6t
Xbit_r59_c161 bl_161 br_161 wl_59 vdd gnd cell_6t
Xbit_r60_c161 bl_161 br_161 wl_60 vdd gnd cell_6t
Xbit_r61_c161 bl_161 br_161 wl_61 vdd gnd cell_6t
Xbit_r62_c161 bl_161 br_161 wl_62 vdd gnd cell_6t
Xbit_r63_c161 bl_161 br_161 wl_63 vdd gnd cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd cell_6t
Xbit_r1_c162 bl_162 br_162 wl_1 vdd gnd cell_6t
Xbit_r2_c162 bl_162 br_162 wl_2 vdd gnd cell_6t
Xbit_r3_c162 bl_162 br_162 wl_3 vdd gnd cell_6t
Xbit_r4_c162 bl_162 br_162 wl_4 vdd gnd cell_6t
Xbit_r5_c162 bl_162 br_162 wl_5 vdd gnd cell_6t
Xbit_r6_c162 bl_162 br_162 wl_6 vdd gnd cell_6t
Xbit_r7_c162 bl_162 br_162 wl_7 vdd gnd cell_6t
Xbit_r8_c162 bl_162 br_162 wl_8 vdd gnd cell_6t
Xbit_r9_c162 bl_162 br_162 wl_9 vdd gnd cell_6t
Xbit_r10_c162 bl_162 br_162 wl_10 vdd gnd cell_6t
Xbit_r11_c162 bl_162 br_162 wl_11 vdd gnd cell_6t
Xbit_r12_c162 bl_162 br_162 wl_12 vdd gnd cell_6t
Xbit_r13_c162 bl_162 br_162 wl_13 vdd gnd cell_6t
Xbit_r14_c162 bl_162 br_162 wl_14 vdd gnd cell_6t
Xbit_r15_c162 bl_162 br_162 wl_15 vdd gnd cell_6t
Xbit_r16_c162 bl_162 br_162 wl_16 vdd gnd cell_6t
Xbit_r17_c162 bl_162 br_162 wl_17 vdd gnd cell_6t
Xbit_r18_c162 bl_162 br_162 wl_18 vdd gnd cell_6t
Xbit_r19_c162 bl_162 br_162 wl_19 vdd gnd cell_6t
Xbit_r20_c162 bl_162 br_162 wl_20 vdd gnd cell_6t
Xbit_r21_c162 bl_162 br_162 wl_21 vdd gnd cell_6t
Xbit_r22_c162 bl_162 br_162 wl_22 vdd gnd cell_6t
Xbit_r23_c162 bl_162 br_162 wl_23 vdd gnd cell_6t
Xbit_r24_c162 bl_162 br_162 wl_24 vdd gnd cell_6t
Xbit_r25_c162 bl_162 br_162 wl_25 vdd gnd cell_6t
Xbit_r26_c162 bl_162 br_162 wl_26 vdd gnd cell_6t
Xbit_r27_c162 bl_162 br_162 wl_27 vdd gnd cell_6t
Xbit_r28_c162 bl_162 br_162 wl_28 vdd gnd cell_6t
Xbit_r29_c162 bl_162 br_162 wl_29 vdd gnd cell_6t
Xbit_r30_c162 bl_162 br_162 wl_30 vdd gnd cell_6t
Xbit_r31_c162 bl_162 br_162 wl_31 vdd gnd cell_6t
Xbit_r32_c162 bl_162 br_162 wl_32 vdd gnd cell_6t
Xbit_r33_c162 bl_162 br_162 wl_33 vdd gnd cell_6t
Xbit_r34_c162 bl_162 br_162 wl_34 vdd gnd cell_6t
Xbit_r35_c162 bl_162 br_162 wl_35 vdd gnd cell_6t
Xbit_r36_c162 bl_162 br_162 wl_36 vdd gnd cell_6t
Xbit_r37_c162 bl_162 br_162 wl_37 vdd gnd cell_6t
Xbit_r38_c162 bl_162 br_162 wl_38 vdd gnd cell_6t
Xbit_r39_c162 bl_162 br_162 wl_39 vdd gnd cell_6t
Xbit_r40_c162 bl_162 br_162 wl_40 vdd gnd cell_6t
Xbit_r41_c162 bl_162 br_162 wl_41 vdd gnd cell_6t
Xbit_r42_c162 bl_162 br_162 wl_42 vdd gnd cell_6t
Xbit_r43_c162 bl_162 br_162 wl_43 vdd gnd cell_6t
Xbit_r44_c162 bl_162 br_162 wl_44 vdd gnd cell_6t
Xbit_r45_c162 bl_162 br_162 wl_45 vdd gnd cell_6t
Xbit_r46_c162 bl_162 br_162 wl_46 vdd gnd cell_6t
Xbit_r47_c162 bl_162 br_162 wl_47 vdd gnd cell_6t
Xbit_r48_c162 bl_162 br_162 wl_48 vdd gnd cell_6t
Xbit_r49_c162 bl_162 br_162 wl_49 vdd gnd cell_6t
Xbit_r50_c162 bl_162 br_162 wl_50 vdd gnd cell_6t
Xbit_r51_c162 bl_162 br_162 wl_51 vdd gnd cell_6t
Xbit_r52_c162 bl_162 br_162 wl_52 vdd gnd cell_6t
Xbit_r53_c162 bl_162 br_162 wl_53 vdd gnd cell_6t
Xbit_r54_c162 bl_162 br_162 wl_54 vdd gnd cell_6t
Xbit_r55_c162 bl_162 br_162 wl_55 vdd gnd cell_6t
Xbit_r56_c162 bl_162 br_162 wl_56 vdd gnd cell_6t
Xbit_r57_c162 bl_162 br_162 wl_57 vdd gnd cell_6t
Xbit_r58_c162 bl_162 br_162 wl_58 vdd gnd cell_6t
Xbit_r59_c162 bl_162 br_162 wl_59 vdd gnd cell_6t
Xbit_r60_c162 bl_162 br_162 wl_60 vdd gnd cell_6t
Xbit_r61_c162 bl_162 br_162 wl_61 vdd gnd cell_6t
Xbit_r62_c162 bl_162 br_162 wl_62 vdd gnd cell_6t
Xbit_r63_c162 bl_162 br_162 wl_63 vdd gnd cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd cell_6t
Xbit_r1_c163 bl_163 br_163 wl_1 vdd gnd cell_6t
Xbit_r2_c163 bl_163 br_163 wl_2 vdd gnd cell_6t
Xbit_r3_c163 bl_163 br_163 wl_3 vdd gnd cell_6t
Xbit_r4_c163 bl_163 br_163 wl_4 vdd gnd cell_6t
Xbit_r5_c163 bl_163 br_163 wl_5 vdd gnd cell_6t
Xbit_r6_c163 bl_163 br_163 wl_6 vdd gnd cell_6t
Xbit_r7_c163 bl_163 br_163 wl_7 vdd gnd cell_6t
Xbit_r8_c163 bl_163 br_163 wl_8 vdd gnd cell_6t
Xbit_r9_c163 bl_163 br_163 wl_9 vdd gnd cell_6t
Xbit_r10_c163 bl_163 br_163 wl_10 vdd gnd cell_6t
Xbit_r11_c163 bl_163 br_163 wl_11 vdd gnd cell_6t
Xbit_r12_c163 bl_163 br_163 wl_12 vdd gnd cell_6t
Xbit_r13_c163 bl_163 br_163 wl_13 vdd gnd cell_6t
Xbit_r14_c163 bl_163 br_163 wl_14 vdd gnd cell_6t
Xbit_r15_c163 bl_163 br_163 wl_15 vdd gnd cell_6t
Xbit_r16_c163 bl_163 br_163 wl_16 vdd gnd cell_6t
Xbit_r17_c163 bl_163 br_163 wl_17 vdd gnd cell_6t
Xbit_r18_c163 bl_163 br_163 wl_18 vdd gnd cell_6t
Xbit_r19_c163 bl_163 br_163 wl_19 vdd gnd cell_6t
Xbit_r20_c163 bl_163 br_163 wl_20 vdd gnd cell_6t
Xbit_r21_c163 bl_163 br_163 wl_21 vdd gnd cell_6t
Xbit_r22_c163 bl_163 br_163 wl_22 vdd gnd cell_6t
Xbit_r23_c163 bl_163 br_163 wl_23 vdd gnd cell_6t
Xbit_r24_c163 bl_163 br_163 wl_24 vdd gnd cell_6t
Xbit_r25_c163 bl_163 br_163 wl_25 vdd gnd cell_6t
Xbit_r26_c163 bl_163 br_163 wl_26 vdd gnd cell_6t
Xbit_r27_c163 bl_163 br_163 wl_27 vdd gnd cell_6t
Xbit_r28_c163 bl_163 br_163 wl_28 vdd gnd cell_6t
Xbit_r29_c163 bl_163 br_163 wl_29 vdd gnd cell_6t
Xbit_r30_c163 bl_163 br_163 wl_30 vdd gnd cell_6t
Xbit_r31_c163 bl_163 br_163 wl_31 vdd gnd cell_6t
Xbit_r32_c163 bl_163 br_163 wl_32 vdd gnd cell_6t
Xbit_r33_c163 bl_163 br_163 wl_33 vdd gnd cell_6t
Xbit_r34_c163 bl_163 br_163 wl_34 vdd gnd cell_6t
Xbit_r35_c163 bl_163 br_163 wl_35 vdd gnd cell_6t
Xbit_r36_c163 bl_163 br_163 wl_36 vdd gnd cell_6t
Xbit_r37_c163 bl_163 br_163 wl_37 vdd gnd cell_6t
Xbit_r38_c163 bl_163 br_163 wl_38 vdd gnd cell_6t
Xbit_r39_c163 bl_163 br_163 wl_39 vdd gnd cell_6t
Xbit_r40_c163 bl_163 br_163 wl_40 vdd gnd cell_6t
Xbit_r41_c163 bl_163 br_163 wl_41 vdd gnd cell_6t
Xbit_r42_c163 bl_163 br_163 wl_42 vdd gnd cell_6t
Xbit_r43_c163 bl_163 br_163 wl_43 vdd gnd cell_6t
Xbit_r44_c163 bl_163 br_163 wl_44 vdd gnd cell_6t
Xbit_r45_c163 bl_163 br_163 wl_45 vdd gnd cell_6t
Xbit_r46_c163 bl_163 br_163 wl_46 vdd gnd cell_6t
Xbit_r47_c163 bl_163 br_163 wl_47 vdd gnd cell_6t
Xbit_r48_c163 bl_163 br_163 wl_48 vdd gnd cell_6t
Xbit_r49_c163 bl_163 br_163 wl_49 vdd gnd cell_6t
Xbit_r50_c163 bl_163 br_163 wl_50 vdd gnd cell_6t
Xbit_r51_c163 bl_163 br_163 wl_51 vdd gnd cell_6t
Xbit_r52_c163 bl_163 br_163 wl_52 vdd gnd cell_6t
Xbit_r53_c163 bl_163 br_163 wl_53 vdd gnd cell_6t
Xbit_r54_c163 bl_163 br_163 wl_54 vdd gnd cell_6t
Xbit_r55_c163 bl_163 br_163 wl_55 vdd gnd cell_6t
Xbit_r56_c163 bl_163 br_163 wl_56 vdd gnd cell_6t
Xbit_r57_c163 bl_163 br_163 wl_57 vdd gnd cell_6t
Xbit_r58_c163 bl_163 br_163 wl_58 vdd gnd cell_6t
Xbit_r59_c163 bl_163 br_163 wl_59 vdd gnd cell_6t
Xbit_r60_c163 bl_163 br_163 wl_60 vdd gnd cell_6t
Xbit_r61_c163 bl_163 br_163 wl_61 vdd gnd cell_6t
Xbit_r62_c163 bl_163 br_163 wl_62 vdd gnd cell_6t
Xbit_r63_c163 bl_163 br_163 wl_63 vdd gnd cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd cell_6t
Xbit_r1_c164 bl_164 br_164 wl_1 vdd gnd cell_6t
Xbit_r2_c164 bl_164 br_164 wl_2 vdd gnd cell_6t
Xbit_r3_c164 bl_164 br_164 wl_3 vdd gnd cell_6t
Xbit_r4_c164 bl_164 br_164 wl_4 vdd gnd cell_6t
Xbit_r5_c164 bl_164 br_164 wl_5 vdd gnd cell_6t
Xbit_r6_c164 bl_164 br_164 wl_6 vdd gnd cell_6t
Xbit_r7_c164 bl_164 br_164 wl_7 vdd gnd cell_6t
Xbit_r8_c164 bl_164 br_164 wl_8 vdd gnd cell_6t
Xbit_r9_c164 bl_164 br_164 wl_9 vdd gnd cell_6t
Xbit_r10_c164 bl_164 br_164 wl_10 vdd gnd cell_6t
Xbit_r11_c164 bl_164 br_164 wl_11 vdd gnd cell_6t
Xbit_r12_c164 bl_164 br_164 wl_12 vdd gnd cell_6t
Xbit_r13_c164 bl_164 br_164 wl_13 vdd gnd cell_6t
Xbit_r14_c164 bl_164 br_164 wl_14 vdd gnd cell_6t
Xbit_r15_c164 bl_164 br_164 wl_15 vdd gnd cell_6t
Xbit_r16_c164 bl_164 br_164 wl_16 vdd gnd cell_6t
Xbit_r17_c164 bl_164 br_164 wl_17 vdd gnd cell_6t
Xbit_r18_c164 bl_164 br_164 wl_18 vdd gnd cell_6t
Xbit_r19_c164 bl_164 br_164 wl_19 vdd gnd cell_6t
Xbit_r20_c164 bl_164 br_164 wl_20 vdd gnd cell_6t
Xbit_r21_c164 bl_164 br_164 wl_21 vdd gnd cell_6t
Xbit_r22_c164 bl_164 br_164 wl_22 vdd gnd cell_6t
Xbit_r23_c164 bl_164 br_164 wl_23 vdd gnd cell_6t
Xbit_r24_c164 bl_164 br_164 wl_24 vdd gnd cell_6t
Xbit_r25_c164 bl_164 br_164 wl_25 vdd gnd cell_6t
Xbit_r26_c164 bl_164 br_164 wl_26 vdd gnd cell_6t
Xbit_r27_c164 bl_164 br_164 wl_27 vdd gnd cell_6t
Xbit_r28_c164 bl_164 br_164 wl_28 vdd gnd cell_6t
Xbit_r29_c164 bl_164 br_164 wl_29 vdd gnd cell_6t
Xbit_r30_c164 bl_164 br_164 wl_30 vdd gnd cell_6t
Xbit_r31_c164 bl_164 br_164 wl_31 vdd gnd cell_6t
Xbit_r32_c164 bl_164 br_164 wl_32 vdd gnd cell_6t
Xbit_r33_c164 bl_164 br_164 wl_33 vdd gnd cell_6t
Xbit_r34_c164 bl_164 br_164 wl_34 vdd gnd cell_6t
Xbit_r35_c164 bl_164 br_164 wl_35 vdd gnd cell_6t
Xbit_r36_c164 bl_164 br_164 wl_36 vdd gnd cell_6t
Xbit_r37_c164 bl_164 br_164 wl_37 vdd gnd cell_6t
Xbit_r38_c164 bl_164 br_164 wl_38 vdd gnd cell_6t
Xbit_r39_c164 bl_164 br_164 wl_39 vdd gnd cell_6t
Xbit_r40_c164 bl_164 br_164 wl_40 vdd gnd cell_6t
Xbit_r41_c164 bl_164 br_164 wl_41 vdd gnd cell_6t
Xbit_r42_c164 bl_164 br_164 wl_42 vdd gnd cell_6t
Xbit_r43_c164 bl_164 br_164 wl_43 vdd gnd cell_6t
Xbit_r44_c164 bl_164 br_164 wl_44 vdd gnd cell_6t
Xbit_r45_c164 bl_164 br_164 wl_45 vdd gnd cell_6t
Xbit_r46_c164 bl_164 br_164 wl_46 vdd gnd cell_6t
Xbit_r47_c164 bl_164 br_164 wl_47 vdd gnd cell_6t
Xbit_r48_c164 bl_164 br_164 wl_48 vdd gnd cell_6t
Xbit_r49_c164 bl_164 br_164 wl_49 vdd gnd cell_6t
Xbit_r50_c164 bl_164 br_164 wl_50 vdd gnd cell_6t
Xbit_r51_c164 bl_164 br_164 wl_51 vdd gnd cell_6t
Xbit_r52_c164 bl_164 br_164 wl_52 vdd gnd cell_6t
Xbit_r53_c164 bl_164 br_164 wl_53 vdd gnd cell_6t
Xbit_r54_c164 bl_164 br_164 wl_54 vdd gnd cell_6t
Xbit_r55_c164 bl_164 br_164 wl_55 vdd gnd cell_6t
Xbit_r56_c164 bl_164 br_164 wl_56 vdd gnd cell_6t
Xbit_r57_c164 bl_164 br_164 wl_57 vdd gnd cell_6t
Xbit_r58_c164 bl_164 br_164 wl_58 vdd gnd cell_6t
Xbit_r59_c164 bl_164 br_164 wl_59 vdd gnd cell_6t
Xbit_r60_c164 bl_164 br_164 wl_60 vdd gnd cell_6t
Xbit_r61_c164 bl_164 br_164 wl_61 vdd gnd cell_6t
Xbit_r62_c164 bl_164 br_164 wl_62 vdd gnd cell_6t
Xbit_r63_c164 bl_164 br_164 wl_63 vdd gnd cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd cell_6t
Xbit_r1_c165 bl_165 br_165 wl_1 vdd gnd cell_6t
Xbit_r2_c165 bl_165 br_165 wl_2 vdd gnd cell_6t
Xbit_r3_c165 bl_165 br_165 wl_3 vdd gnd cell_6t
Xbit_r4_c165 bl_165 br_165 wl_4 vdd gnd cell_6t
Xbit_r5_c165 bl_165 br_165 wl_5 vdd gnd cell_6t
Xbit_r6_c165 bl_165 br_165 wl_6 vdd gnd cell_6t
Xbit_r7_c165 bl_165 br_165 wl_7 vdd gnd cell_6t
Xbit_r8_c165 bl_165 br_165 wl_8 vdd gnd cell_6t
Xbit_r9_c165 bl_165 br_165 wl_9 vdd gnd cell_6t
Xbit_r10_c165 bl_165 br_165 wl_10 vdd gnd cell_6t
Xbit_r11_c165 bl_165 br_165 wl_11 vdd gnd cell_6t
Xbit_r12_c165 bl_165 br_165 wl_12 vdd gnd cell_6t
Xbit_r13_c165 bl_165 br_165 wl_13 vdd gnd cell_6t
Xbit_r14_c165 bl_165 br_165 wl_14 vdd gnd cell_6t
Xbit_r15_c165 bl_165 br_165 wl_15 vdd gnd cell_6t
Xbit_r16_c165 bl_165 br_165 wl_16 vdd gnd cell_6t
Xbit_r17_c165 bl_165 br_165 wl_17 vdd gnd cell_6t
Xbit_r18_c165 bl_165 br_165 wl_18 vdd gnd cell_6t
Xbit_r19_c165 bl_165 br_165 wl_19 vdd gnd cell_6t
Xbit_r20_c165 bl_165 br_165 wl_20 vdd gnd cell_6t
Xbit_r21_c165 bl_165 br_165 wl_21 vdd gnd cell_6t
Xbit_r22_c165 bl_165 br_165 wl_22 vdd gnd cell_6t
Xbit_r23_c165 bl_165 br_165 wl_23 vdd gnd cell_6t
Xbit_r24_c165 bl_165 br_165 wl_24 vdd gnd cell_6t
Xbit_r25_c165 bl_165 br_165 wl_25 vdd gnd cell_6t
Xbit_r26_c165 bl_165 br_165 wl_26 vdd gnd cell_6t
Xbit_r27_c165 bl_165 br_165 wl_27 vdd gnd cell_6t
Xbit_r28_c165 bl_165 br_165 wl_28 vdd gnd cell_6t
Xbit_r29_c165 bl_165 br_165 wl_29 vdd gnd cell_6t
Xbit_r30_c165 bl_165 br_165 wl_30 vdd gnd cell_6t
Xbit_r31_c165 bl_165 br_165 wl_31 vdd gnd cell_6t
Xbit_r32_c165 bl_165 br_165 wl_32 vdd gnd cell_6t
Xbit_r33_c165 bl_165 br_165 wl_33 vdd gnd cell_6t
Xbit_r34_c165 bl_165 br_165 wl_34 vdd gnd cell_6t
Xbit_r35_c165 bl_165 br_165 wl_35 vdd gnd cell_6t
Xbit_r36_c165 bl_165 br_165 wl_36 vdd gnd cell_6t
Xbit_r37_c165 bl_165 br_165 wl_37 vdd gnd cell_6t
Xbit_r38_c165 bl_165 br_165 wl_38 vdd gnd cell_6t
Xbit_r39_c165 bl_165 br_165 wl_39 vdd gnd cell_6t
Xbit_r40_c165 bl_165 br_165 wl_40 vdd gnd cell_6t
Xbit_r41_c165 bl_165 br_165 wl_41 vdd gnd cell_6t
Xbit_r42_c165 bl_165 br_165 wl_42 vdd gnd cell_6t
Xbit_r43_c165 bl_165 br_165 wl_43 vdd gnd cell_6t
Xbit_r44_c165 bl_165 br_165 wl_44 vdd gnd cell_6t
Xbit_r45_c165 bl_165 br_165 wl_45 vdd gnd cell_6t
Xbit_r46_c165 bl_165 br_165 wl_46 vdd gnd cell_6t
Xbit_r47_c165 bl_165 br_165 wl_47 vdd gnd cell_6t
Xbit_r48_c165 bl_165 br_165 wl_48 vdd gnd cell_6t
Xbit_r49_c165 bl_165 br_165 wl_49 vdd gnd cell_6t
Xbit_r50_c165 bl_165 br_165 wl_50 vdd gnd cell_6t
Xbit_r51_c165 bl_165 br_165 wl_51 vdd gnd cell_6t
Xbit_r52_c165 bl_165 br_165 wl_52 vdd gnd cell_6t
Xbit_r53_c165 bl_165 br_165 wl_53 vdd gnd cell_6t
Xbit_r54_c165 bl_165 br_165 wl_54 vdd gnd cell_6t
Xbit_r55_c165 bl_165 br_165 wl_55 vdd gnd cell_6t
Xbit_r56_c165 bl_165 br_165 wl_56 vdd gnd cell_6t
Xbit_r57_c165 bl_165 br_165 wl_57 vdd gnd cell_6t
Xbit_r58_c165 bl_165 br_165 wl_58 vdd gnd cell_6t
Xbit_r59_c165 bl_165 br_165 wl_59 vdd gnd cell_6t
Xbit_r60_c165 bl_165 br_165 wl_60 vdd gnd cell_6t
Xbit_r61_c165 bl_165 br_165 wl_61 vdd gnd cell_6t
Xbit_r62_c165 bl_165 br_165 wl_62 vdd gnd cell_6t
Xbit_r63_c165 bl_165 br_165 wl_63 vdd gnd cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd cell_6t
Xbit_r1_c166 bl_166 br_166 wl_1 vdd gnd cell_6t
Xbit_r2_c166 bl_166 br_166 wl_2 vdd gnd cell_6t
Xbit_r3_c166 bl_166 br_166 wl_3 vdd gnd cell_6t
Xbit_r4_c166 bl_166 br_166 wl_4 vdd gnd cell_6t
Xbit_r5_c166 bl_166 br_166 wl_5 vdd gnd cell_6t
Xbit_r6_c166 bl_166 br_166 wl_6 vdd gnd cell_6t
Xbit_r7_c166 bl_166 br_166 wl_7 vdd gnd cell_6t
Xbit_r8_c166 bl_166 br_166 wl_8 vdd gnd cell_6t
Xbit_r9_c166 bl_166 br_166 wl_9 vdd gnd cell_6t
Xbit_r10_c166 bl_166 br_166 wl_10 vdd gnd cell_6t
Xbit_r11_c166 bl_166 br_166 wl_11 vdd gnd cell_6t
Xbit_r12_c166 bl_166 br_166 wl_12 vdd gnd cell_6t
Xbit_r13_c166 bl_166 br_166 wl_13 vdd gnd cell_6t
Xbit_r14_c166 bl_166 br_166 wl_14 vdd gnd cell_6t
Xbit_r15_c166 bl_166 br_166 wl_15 vdd gnd cell_6t
Xbit_r16_c166 bl_166 br_166 wl_16 vdd gnd cell_6t
Xbit_r17_c166 bl_166 br_166 wl_17 vdd gnd cell_6t
Xbit_r18_c166 bl_166 br_166 wl_18 vdd gnd cell_6t
Xbit_r19_c166 bl_166 br_166 wl_19 vdd gnd cell_6t
Xbit_r20_c166 bl_166 br_166 wl_20 vdd gnd cell_6t
Xbit_r21_c166 bl_166 br_166 wl_21 vdd gnd cell_6t
Xbit_r22_c166 bl_166 br_166 wl_22 vdd gnd cell_6t
Xbit_r23_c166 bl_166 br_166 wl_23 vdd gnd cell_6t
Xbit_r24_c166 bl_166 br_166 wl_24 vdd gnd cell_6t
Xbit_r25_c166 bl_166 br_166 wl_25 vdd gnd cell_6t
Xbit_r26_c166 bl_166 br_166 wl_26 vdd gnd cell_6t
Xbit_r27_c166 bl_166 br_166 wl_27 vdd gnd cell_6t
Xbit_r28_c166 bl_166 br_166 wl_28 vdd gnd cell_6t
Xbit_r29_c166 bl_166 br_166 wl_29 vdd gnd cell_6t
Xbit_r30_c166 bl_166 br_166 wl_30 vdd gnd cell_6t
Xbit_r31_c166 bl_166 br_166 wl_31 vdd gnd cell_6t
Xbit_r32_c166 bl_166 br_166 wl_32 vdd gnd cell_6t
Xbit_r33_c166 bl_166 br_166 wl_33 vdd gnd cell_6t
Xbit_r34_c166 bl_166 br_166 wl_34 vdd gnd cell_6t
Xbit_r35_c166 bl_166 br_166 wl_35 vdd gnd cell_6t
Xbit_r36_c166 bl_166 br_166 wl_36 vdd gnd cell_6t
Xbit_r37_c166 bl_166 br_166 wl_37 vdd gnd cell_6t
Xbit_r38_c166 bl_166 br_166 wl_38 vdd gnd cell_6t
Xbit_r39_c166 bl_166 br_166 wl_39 vdd gnd cell_6t
Xbit_r40_c166 bl_166 br_166 wl_40 vdd gnd cell_6t
Xbit_r41_c166 bl_166 br_166 wl_41 vdd gnd cell_6t
Xbit_r42_c166 bl_166 br_166 wl_42 vdd gnd cell_6t
Xbit_r43_c166 bl_166 br_166 wl_43 vdd gnd cell_6t
Xbit_r44_c166 bl_166 br_166 wl_44 vdd gnd cell_6t
Xbit_r45_c166 bl_166 br_166 wl_45 vdd gnd cell_6t
Xbit_r46_c166 bl_166 br_166 wl_46 vdd gnd cell_6t
Xbit_r47_c166 bl_166 br_166 wl_47 vdd gnd cell_6t
Xbit_r48_c166 bl_166 br_166 wl_48 vdd gnd cell_6t
Xbit_r49_c166 bl_166 br_166 wl_49 vdd gnd cell_6t
Xbit_r50_c166 bl_166 br_166 wl_50 vdd gnd cell_6t
Xbit_r51_c166 bl_166 br_166 wl_51 vdd gnd cell_6t
Xbit_r52_c166 bl_166 br_166 wl_52 vdd gnd cell_6t
Xbit_r53_c166 bl_166 br_166 wl_53 vdd gnd cell_6t
Xbit_r54_c166 bl_166 br_166 wl_54 vdd gnd cell_6t
Xbit_r55_c166 bl_166 br_166 wl_55 vdd gnd cell_6t
Xbit_r56_c166 bl_166 br_166 wl_56 vdd gnd cell_6t
Xbit_r57_c166 bl_166 br_166 wl_57 vdd gnd cell_6t
Xbit_r58_c166 bl_166 br_166 wl_58 vdd gnd cell_6t
Xbit_r59_c166 bl_166 br_166 wl_59 vdd gnd cell_6t
Xbit_r60_c166 bl_166 br_166 wl_60 vdd gnd cell_6t
Xbit_r61_c166 bl_166 br_166 wl_61 vdd gnd cell_6t
Xbit_r62_c166 bl_166 br_166 wl_62 vdd gnd cell_6t
Xbit_r63_c166 bl_166 br_166 wl_63 vdd gnd cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd cell_6t
Xbit_r1_c167 bl_167 br_167 wl_1 vdd gnd cell_6t
Xbit_r2_c167 bl_167 br_167 wl_2 vdd gnd cell_6t
Xbit_r3_c167 bl_167 br_167 wl_3 vdd gnd cell_6t
Xbit_r4_c167 bl_167 br_167 wl_4 vdd gnd cell_6t
Xbit_r5_c167 bl_167 br_167 wl_5 vdd gnd cell_6t
Xbit_r6_c167 bl_167 br_167 wl_6 vdd gnd cell_6t
Xbit_r7_c167 bl_167 br_167 wl_7 vdd gnd cell_6t
Xbit_r8_c167 bl_167 br_167 wl_8 vdd gnd cell_6t
Xbit_r9_c167 bl_167 br_167 wl_9 vdd gnd cell_6t
Xbit_r10_c167 bl_167 br_167 wl_10 vdd gnd cell_6t
Xbit_r11_c167 bl_167 br_167 wl_11 vdd gnd cell_6t
Xbit_r12_c167 bl_167 br_167 wl_12 vdd gnd cell_6t
Xbit_r13_c167 bl_167 br_167 wl_13 vdd gnd cell_6t
Xbit_r14_c167 bl_167 br_167 wl_14 vdd gnd cell_6t
Xbit_r15_c167 bl_167 br_167 wl_15 vdd gnd cell_6t
Xbit_r16_c167 bl_167 br_167 wl_16 vdd gnd cell_6t
Xbit_r17_c167 bl_167 br_167 wl_17 vdd gnd cell_6t
Xbit_r18_c167 bl_167 br_167 wl_18 vdd gnd cell_6t
Xbit_r19_c167 bl_167 br_167 wl_19 vdd gnd cell_6t
Xbit_r20_c167 bl_167 br_167 wl_20 vdd gnd cell_6t
Xbit_r21_c167 bl_167 br_167 wl_21 vdd gnd cell_6t
Xbit_r22_c167 bl_167 br_167 wl_22 vdd gnd cell_6t
Xbit_r23_c167 bl_167 br_167 wl_23 vdd gnd cell_6t
Xbit_r24_c167 bl_167 br_167 wl_24 vdd gnd cell_6t
Xbit_r25_c167 bl_167 br_167 wl_25 vdd gnd cell_6t
Xbit_r26_c167 bl_167 br_167 wl_26 vdd gnd cell_6t
Xbit_r27_c167 bl_167 br_167 wl_27 vdd gnd cell_6t
Xbit_r28_c167 bl_167 br_167 wl_28 vdd gnd cell_6t
Xbit_r29_c167 bl_167 br_167 wl_29 vdd gnd cell_6t
Xbit_r30_c167 bl_167 br_167 wl_30 vdd gnd cell_6t
Xbit_r31_c167 bl_167 br_167 wl_31 vdd gnd cell_6t
Xbit_r32_c167 bl_167 br_167 wl_32 vdd gnd cell_6t
Xbit_r33_c167 bl_167 br_167 wl_33 vdd gnd cell_6t
Xbit_r34_c167 bl_167 br_167 wl_34 vdd gnd cell_6t
Xbit_r35_c167 bl_167 br_167 wl_35 vdd gnd cell_6t
Xbit_r36_c167 bl_167 br_167 wl_36 vdd gnd cell_6t
Xbit_r37_c167 bl_167 br_167 wl_37 vdd gnd cell_6t
Xbit_r38_c167 bl_167 br_167 wl_38 vdd gnd cell_6t
Xbit_r39_c167 bl_167 br_167 wl_39 vdd gnd cell_6t
Xbit_r40_c167 bl_167 br_167 wl_40 vdd gnd cell_6t
Xbit_r41_c167 bl_167 br_167 wl_41 vdd gnd cell_6t
Xbit_r42_c167 bl_167 br_167 wl_42 vdd gnd cell_6t
Xbit_r43_c167 bl_167 br_167 wl_43 vdd gnd cell_6t
Xbit_r44_c167 bl_167 br_167 wl_44 vdd gnd cell_6t
Xbit_r45_c167 bl_167 br_167 wl_45 vdd gnd cell_6t
Xbit_r46_c167 bl_167 br_167 wl_46 vdd gnd cell_6t
Xbit_r47_c167 bl_167 br_167 wl_47 vdd gnd cell_6t
Xbit_r48_c167 bl_167 br_167 wl_48 vdd gnd cell_6t
Xbit_r49_c167 bl_167 br_167 wl_49 vdd gnd cell_6t
Xbit_r50_c167 bl_167 br_167 wl_50 vdd gnd cell_6t
Xbit_r51_c167 bl_167 br_167 wl_51 vdd gnd cell_6t
Xbit_r52_c167 bl_167 br_167 wl_52 vdd gnd cell_6t
Xbit_r53_c167 bl_167 br_167 wl_53 vdd gnd cell_6t
Xbit_r54_c167 bl_167 br_167 wl_54 vdd gnd cell_6t
Xbit_r55_c167 bl_167 br_167 wl_55 vdd gnd cell_6t
Xbit_r56_c167 bl_167 br_167 wl_56 vdd gnd cell_6t
Xbit_r57_c167 bl_167 br_167 wl_57 vdd gnd cell_6t
Xbit_r58_c167 bl_167 br_167 wl_58 vdd gnd cell_6t
Xbit_r59_c167 bl_167 br_167 wl_59 vdd gnd cell_6t
Xbit_r60_c167 bl_167 br_167 wl_60 vdd gnd cell_6t
Xbit_r61_c167 bl_167 br_167 wl_61 vdd gnd cell_6t
Xbit_r62_c167 bl_167 br_167 wl_62 vdd gnd cell_6t
Xbit_r63_c167 bl_167 br_167 wl_63 vdd gnd cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd cell_6t
Xbit_r1_c168 bl_168 br_168 wl_1 vdd gnd cell_6t
Xbit_r2_c168 bl_168 br_168 wl_2 vdd gnd cell_6t
Xbit_r3_c168 bl_168 br_168 wl_3 vdd gnd cell_6t
Xbit_r4_c168 bl_168 br_168 wl_4 vdd gnd cell_6t
Xbit_r5_c168 bl_168 br_168 wl_5 vdd gnd cell_6t
Xbit_r6_c168 bl_168 br_168 wl_6 vdd gnd cell_6t
Xbit_r7_c168 bl_168 br_168 wl_7 vdd gnd cell_6t
Xbit_r8_c168 bl_168 br_168 wl_8 vdd gnd cell_6t
Xbit_r9_c168 bl_168 br_168 wl_9 vdd gnd cell_6t
Xbit_r10_c168 bl_168 br_168 wl_10 vdd gnd cell_6t
Xbit_r11_c168 bl_168 br_168 wl_11 vdd gnd cell_6t
Xbit_r12_c168 bl_168 br_168 wl_12 vdd gnd cell_6t
Xbit_r13_c168 bl_168 br_168 wl_13 vdd gnd cell_6t
Xbit_r14_c168 bl_168 br_168 wl_14 vdd gnd cell_6t
Xbit_r15_c168 bl_168 br_168 wl_15 vdd gnd cell_6t
Xbit_r16_c168 bl_168 br_168 wl_16 vdd gnd cell_6t
Xbit_r17_c168 bl_168 br_168 wl_17 vdd gnd cell_6t
Xbit_r18_c168 bl_168 br_168 wl_18 vdd gnd cell_6t
Xbit_r19_c168 bl_168 br_168 wl_19 vdd gnd cell_6t
Xbit_r20_c168 bl_168 br_168 wl_20 vdd gnd cell_6t
Xbit_r21_c168 bl_168 br_168 wl_21 vdd gnd cell_6t
Xbit_r22_c168 bl_168 br_168 wl_22 vdd gnd cell_6t
Xbit_r23_c168 bl_168 br_168 wl_23 vdd gnd cell_6t
Xbit_r24_c168 bl_168 br_168 wl_24 vdd gnd cell_6t
Xbit_r25_c168 bl_168 br_168 wl_25 vdd gnd cell_6t
Xbit_r26_c168 bl_168 br_168 wl_26 vdd gnd cell_6t
Xbit_r27_c168 bl_168 br_168 wl_27 vdd gnd cell_6t
Xbit_r28_c168 bl_168 br_168 wl_28 vdd gnd cell_6t
Xbit_r29_c168 bl_168 br_168 wl_29 vdd gnd cell_6t
Xbit_r30_c168 bl_168 br_168 wl_30 vdd gnd cell_6t
Xbit_r31_c168 bl_168 br_168 wl_31 vdd gnd cell_6t
Xbit_r32_c168 bl_168 br_168 wl_32 vdd gnd cell_6t
Xbit_r33_c168 bl_168 br_168 wl_33 vdd gnd cell_6t
Xbit_r34_c168 bl_168 br_168 wl_34 vdd gnd cell_6t
Xbit_r35_c168 bl_168 br_168 wl_35 vdd gnd cell_6t
Xbit_r36_c168 bl_168 br_168 wl_36 vdd gnd cell_6t
Xbit_r37_c168 bl_168 br_168 wl_37 vdd gnd cell_6t
Xbit_r38_c168 bl_168 br_168 wl_38 vdd gnd cell_6t
Xbit_r39_c168 bl_168 br_168 wl_39 vdd gnd cell_6t
Xbit_r40_c168 bl_168 br_168 wl_40 vdd gnd cell_6t
Xbit_r41_c168 bl_168 br_168 wl_41 vdd gnd cell_6t
Xbit_r42_c168 bl_168 br_168 wl_42 vdd gnd cell_6t
Xbit_r43_c168 bl_168 br_168 wl_43 vdd gnd cell_6t
Xbit_r44_c168 bl_168 br_168 wl_44 vdd gnd cell_6t
Xbit_r45_c168 bl_168 br_168 wl_45 vdd gnd cell_6t
Xbit_r46_c168 bl_168 br_168 wl_46 vdd gnd cell_6t
Xbit_r47_c168 bl_168 br_168 wl_47 vdd gnd cell_6t
Xbit_r48_c168 bl_168 br_168 wl_48 vdd gnd cell_6t
Xbit_r49_c168 bl_168 br_168 wl_49 vdd gnd cell_6t
Xbit_r50_c168 bl_168 br_168 wl_50 vdd gnd cell_6t
Xbit_r51_c168 bl_168 br_168 wl_51 vdd gnd cell_6t
Xbit_r52_c168 bl_168 br_168 wl_52 vdd gnd cell_6t
Xbit_r53_c168 bl_168 br_168 wl_53 vdd gnd cell_6t
Xbit_r54_c168 bl_168 br_168 wl_54 vdd gnd cell_6t
Xbit_r55_c168 bl_168 br_168 wl_55 vdd gnd cell_6t
Xbit_r56_c168 bl_168 br_168 wl_56 vdd gnd cell_6t
Xbit_r57_c168 bl_168 br_168 wl_57 vdd gnd cell_6t
Xbit_r58_c168 bl_168 br_168 wl_58 vdd gnd cell_6t
Xbit_r59_c168 bl_168 br_168 wl_59 vdd gnd cell_6t
Xbit_r60_c168 bl_168 br_168 wl_60 vdd gnd cell_6t
Xbit_r61_c168 bl_168 br_168 wl_61 vdd gnd cell_6t
Xbit_r62_c168 bl_168 br_168 wl_62 vdd gnd cell_6t
Xbit_r63_c168 bl_168 br_168 wl_63 vdd gnd cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd cell_6t
Xbit_r1_c169 bl_169 br_169 wl_1 vdd gnd cell_6t
Xbit_r2_c169 bl_169 br_169 wl_2 vdd gnd cell_6t
Xbit_r3_c169 bl_169 br_169 wl_3 vdd gnd cell_6t
Xbit_r4_c169 bl_169 br_169 wl_4 vdd gnd cell_6t
Xbit_r5_c169 bl_169 br_169 wl_5 vdd gnd cell_6t
Xbit_r6_c169 bl_169 br_169 wl_6 vdd gnd cell_6t
Xbit_r7_c169 bl_169 br_169 wl_7 vdd gnd cell_6t
Xbit_r8_c169 bl_169 br_169 wl_8 vdd gnd cell_6t
Xbit_r9_c169 bl_169 br_169 wl_9 vdd gnd cell_6t
Xbit_r10_c169 bl_169 br_169 wl_10 vdd gnd cell_6t
Xbit_r11_c169 bl_169 br_169 wl_11 vdd gnd cell_6t
Xbit_r12_c169 bl_169 br_169 wl_12 vdd gnd cell_6t
Xbit_r13_c169 bl_169 br_169 wl_13 vdd gnd cell_6t
Xbit_r14_c169 bl_169 br_169 wl_14 vdd gnd cell_6t
Xbit_r15_c169 bl_169 br_169 wl_15 vdd gnd cell_6t
Xbit_r16_c169 bl_169 br_169 wl_16 vdd gnd cell_6t
Xbit_r17_c169 bl_169 br_169 wl_17 vdd gnd cell_6t
Xbit_r18_c169 bl_169 br_169 wl_18 vdd gnd cell_6t
Xbit_r19_c169 bl_169 br_169 wl_19 vdd gnd cell_6t
Xbit_r20_c169 bl_169 br_169 wl_20 vdd gnd cell_6t
Xbit_r21_c169 bl_169 br_169 wl_21 vdd gnd cell_6t
Xbit_r22_c169 bl_169 br_169 wl_22 vdd gnd cell_6t
Xbit_r23_c169 bl_169 br_169 wl_23 vdd gnd cell_6t
Xbit_r24_c169 bl_169 br_169 wl_24 vdd gnd cell_6t
Xbit_r25_c169 bl_169 br_169 wl_25 vdd gnd cell_6t
Xbit_r26_c169 bl_169 br_169 wl_26 vdd gnd cell_6t
Xbit_r27_c169 bl_169 br_169 wl_27 vdd gnd cell_6t
Xbit_r28_c169 bl_169 br_169 wl_28 vdd gnd cell_6t
Xbit_r29_c169 bl_169 br_169 wl_29 vdd gnd cell_6t
Xbit_r30_c169 bl_169 br_169 wl_30 vdd gnd cell_6t
Xbit_r31_c169 bl_169 br_169 wl_31 vdd gnd cell_6t
Xbit_r32_c169 bl_169 br_169 wl_32 vdd gnd cell_6t
Xbit_r33_c169 bl_169 br_169 wl_33 vdd gnd cell_6t
Xbit_r34_c169 bl_169 br_169 wl_34 vdd gnd cell_6t
Xbit_r35_c169 bl_169 br_169 wl_35 vdd gnd cell_6t
Xbit_r36_c169 bl_169 br_169 wl_36 vdd gnd cell_6t
Xbit_r37_c169 bl_169 br_169 wl_37 vdd gnd cell_6t
Xbit_r38_c169 bl_169 br_169 wl_38 vdd gnd cell_6t
Xbit_r39_c169 bl_169 br_169 wl_39 vdd gnd cell_6t
Xbit_r40_c169 bl_169 br_169 wl_40 vdd gnd cell_6t
Xbit_r41_c169 bl_169 br_169 wl_41 vdd gnd cell_6t
Xbit_r42_c169 bl_169 br_169 wl_42 vdd gnd cell_6t
Xbit_r43_c169 bl_169 br_169 wl_43 vdd gnd cell_6t
Xbit_r44_c169 bl_169 br_169 wl_44 vdd gnd cell_6t
Xbit_r45_c169 bl_169 br_169 wl_45 vdd gnd cell_6t
Xbit_r46_c169 bl_169 br_169 wl_46 vdd gnd cell_6t
Xbit_r47_c169 bl_169 br_169 wl_47 vdd gnd cell_6t
Xbit_r48_c169 bl_169 br_169 wl_48 vdd gnd cell_6t
Xbit_r49_c169 bl_169 br_169 wl_49 vdd gnd cell_6t
Xbit_r50_c169 bl_169 br_169 wl_50 vdd gnd cell_6t
Xbit_r51_c169 bl_169 br_169 wl_51 vdd gnd cell_6t
Xbit_r52_c169 bl_169 br_169 wl_52 vdd gnd cell_6t
Xbit_r53_c169 bl_169 br_169 wl_53 vdd gnd cell_6t
Xbit_r54_c169 bl_169 br_169 wl_54 vdd gnd cell_6t
Xbit_r55_c169 bl_169 br_169 wl_55 vdd gnd cell_6t
Xbit_r56_c169 bl_169 br_169 wl_56 vdd gnd cell_6t
Xbit_r57_c169 bl_169 br_169 wl_57 vdd gnd cell_6t
Xbit_r58_c169 bl_169 br_169 wl_58 vdd gnd cell_6t
Xbit_r59_c169 bl_169 br_169 wl_59 vdd gnd cell_6t
Xbit_r60_c169 bl_169 br_169 wl_60 vdd gnd cell_6t
Xbit_r61_c169 bl_169 br_169 wl_61 vdd gnd cell_6t
Xbit_r62_c169 bl_169 br_169 wl_62 vdd gnd cell_6t
Xbit_r63_c169 bl_169 br_169 wl_63 vdd gnd cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd cell_6t
Xbit_r1_c170 bl_170 br_170 wl_1 vdd gnd cell_6t
Xbit_r2_c170 bl_170 br_170 wl_2 vdd gnd cell_6t
Xbit_r3_c170 bl_170 br_170 wl_3 vdd gnd cell_6t
Xbit_r4_c170 bl_170 br_170 wl_4 vdd gnd cell_6t
Xbit_r5_c170 bl_170 br_170 wl_5 vdd gnd cell_6t
Xbit_r6_c170 bl_170 br_170 wl_6 vdd gnd cell_6t
Xbit_r7_c170 bl_170 br_170 wl_7 vdd gnd cell_6t
Xbit_r8_c170 bl_170 br_170 wl_8 vdd gnd cell_6t
Xbit_r9_c170 bl_170 br_170 wl_9 vdd gnd cell_6t
Xbit_r10_c170 bl_170 br_170 wl_10 vdd gnd cell_6t
Xbit_r11_c170 bl_170 br_170 wl_11 vdd gnd cell_6t
Xbit_r12_c170 bl_170 br_170 wl_12 vdd gnd cell_6t
Xbit_r13_c170 bl_170 br_170 wl_13 vdd gnd cell_6t
Xbit_r14_c170 bl_170 br_170 wl_14 vdd gnd cell_6t
Xbit_r15_c170 bl_170 br_170 wl_15 vdd gnd cell_6t
Xbit_r16_c170 bl_170 br_170 wl_16 vdd gnd cell_6t
Xbit_r17_c170 bl_170 br_170 wl_17 vdd gnd cell_6t
Xbit_r18_c170 bl_170 br_170 wl_18 vdd gnd cell_6t
Xbit_r19_c170 bl_170 br_170 wl_19 vdd gnd cell_6t
Xbit_r20_c170 bl_170 br_170 wl_20 vdd gnd cell_6t
Xbit_r21_c170 bl_170 br_170 wl_21 vdd gnd cell_6t
Xbit_r22_c170 bl_170 br_170 wl_22 vdd gnd cell_6t
Xbit_r23_c170 bl_170 br_170 wl_23 vdd gnd cell_6t
Xbit_r24_c170 bl_170 br_170 wl_24 vdd gnd cell_6t
Xbit_r25_c170 bl_170 br_170 wl_25 vdd gnd cell_6t
Xbit_r26_c170 bl_170 br_170 wl_26 vdd gnd cell_6t
Xbit_r27_c170 bl_170 br_170 wl_27 vdd gnd cell_6t
Xbit_r28_c170 bl_170 br_170 wl_28 vdd gnd cell_6t
Xbit_r29_c170 bl_170 br_170 wl_29 vdd gnd cell_6t
Xbit_r30_c170 bl_170 br_170 wl_30 vdd gnd cell_6t
Xbit_r31_c170 bl_170 br_170 wl_31 vdd gnd cell_6t
Xbit_r32_c170 bl_170 br_170 wl_32 vdd gnd cell_6t
Xbit_r33_c170 bl_170 br_170 wl_33 vdd gnd cell_6t
Xbit_r34_c170 bl_170 br_170 wl_34 vdd gnd cell_6t
Xbit_r35_c170 bl_170 br_170 wl_35 vdd gnd cell_6t
Xbit_r36_c170 bl_170 br_170 wl_36 vdd gnd cell_6t
Xbit_r37_c170 bl_170 br_170 wl_37 vdd gnd cell_6t
Xbit_r38_c170 bl_170 br_170 wl_38 vdd gnd cell_6t
Xbit_r39_c170 bl_170 br_170 wl_39 vdd gnd cell_6t
Xbit_r40_c170 bl_170 br_170 wl_40 vdd gnd cell_6t
Xbit_r41_c170 bl_170 br_170 wl_41 vdd gnd cell_6t
Xbit_r42_c170 bl_170 br_170 wl_42 vdd gnd cell_6t
Xbit_r43_c170 bl_170 br_170 wl_43 vdd gnd cell_6t
Xbit_r44_c170 bl_170 br_170 wl_44 vdd gnd cell_6t
Xbit_r45_c170 bl_170 br_170 wl_45 vdd gnd cell_6t
Xbit_r46_c170 bl_170 br_170 wl_46 vdd gnd cell_6t
Xbit_r47_c170 bl_170 br_170 wl_47 vdd gnd cell_6t
Xbit_r48_c170 bl_170 br_170 wl_48 vdd gnd cell_6t
Xbit_r49_c170 bl_170 br_170 wl_49 vdd gnd cell_6t
Xbit_r50_c170 bl_170 br_170 wl_50 vdd gnd cell_6t
Xbit_r51_c170 bl_170 br_170 wl_51 vdd gnd cell_6t
Xbit_r52_c170 bl_170 br_170 wl_52 vdd gnd cell_6t
Xbit_r53_c170 bl_170 br_170 wl_53 vdd gnd cell_6t
Xbit_r54_c170 bl_170 br_170 wl_54 vdd gnd cell_6t
Xbit_r55_c170 bl_170 br_170 wl_55 vdd gnd cell_6t
Xbit_r56_c170 bl_170 br_170 wl_56 vdd gnd cell_6t
Xbit_r57_c170 bl_170 br_170 wl_57 vdd gnd cell_6t
Xbit_r58_c170 bl_170 br_170 wl_58 vdd gnd cell_6t
Xbit_r59_c170 bl_170 br_170 wl_59 vdd gnd cell_6t
Xbit_r60_c170 bl_170 br_170 wl_60 vdd gnd cell_6t
Xbit_r61_c170 bl_170 br_170 wl_61 vdd gnd cell_6t
Xbit_r62_c170 bl_170 br_170 wl_62 vdd gnd cell_6t
Xbit_r63_c170 bl_170 br_170 wl_63 vdd gnd cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd cell_6t
Xbit_r1_c171 bl_171 br_171 wl_1 vdd gnd cell_6t
Xbit_r2_c171 bl_171 br_171 wl_2 vdd gnd cell_6t
Xbit_r3_c171 bl_171 br_171 wl_3 vdd gnd cell_6t
Xbit_r4_c171 bl_171 br_171 wl_4 vdd gnd cell_6t
Xbit_r5_c171 bl_171 br_171 wl_5 vdd gnd cell_6t
Xbit_r6_c171 bl_171 br_171 wl_6 vdd gnd cell_6t
Xbit_r7_c171 bl_171 br_171 wl_7 vdd gnd cell_6t
Xbit_r8_c171 bl_171 br_171 wl_8 vdd gnd cell_6t
Xbit_r9_c171 bl_171 br_171 wl_9 vdd gnd cell_6t
Xbit_r10_c171 bl_171 br_171 wl_10 vdd gnd cell_6t
Xbit_r11_c171 bl_171 br_171 wl_11 vdd gnd cell_6t
Xbit_r12_c171 bl_171 br_171 wl_12 vdd gnd cell_6t
Xbit_r13_c171 bl_171 br_171 wl_13 vdd gnd cell_6t
Xbit_r14_c171 bl_171 br_171 wl_14 vdd gnd cell_6t
Xbit_r15_c171 bl_171 br_171 wl_15 vdd gnd cell_6t
Xbit_r16_c171 bl_171 br_171 wl_16 vdd gnd cell_6t
Xbit_r17_c171 bl_171 br_171 wl_17 vdd gnd cell_6t
Xbit_r18_c171 bl_171 br_171 wl_18 vdd gnd cell_6t
Xbit_r19_c171 bl_171 br_171 wl_19 vdd gnd cell_6t
Xbit_r20_c171 bl_171 br_171 wl_20 vdd gnd cell_6t
Xbit_r21_c171 bl_171 br_171 wl_21 vdd gnd cell_6t
Xbit_r22_c171 bl_171 br_171 wl_22 vdd gnd cell_6t
Xbit_r23_c171 bl_171 br_171 wl_23 vdd gnd cell_6t
Xbit_r24_c171 bl_171 br_171 wl_24 vdd gnd cell_6t
Xbit_r25_c171 bl_171 br_171 wl_25 vdd gnd cell_6t
Xbit_r26_c171 bl_171 br_171 wl_26 vdd gnd cell_6t
Xbit_r27_c171 bl_171 br_171 wl_27 vdd gnd cell_6t
Xbit_r28_c171 bl_171 br_171 wl_28 vdd gnd cell_6t
Xbit_r29_c171 bl_171 br_171 wl_29 vdd gnd cell_6t
Xbit_r30_c171 bl_171 br_171 wl_30 vdd gnd cell_6t
Xbit_r31_c171 bl_171 br_171 wl_31 vdd gnd cell_6t
Xbit_r32_c171 bl_171 br_171 wl_32 vdd gnd cell_6t
Xbit_r33_c171 bl_171 br_171 wl_33 vdd gnd cell_6t
Xbit_r34_c171 bl_171 br_171 wl_34 vdd gnd cell_6t
Xbit_r35_c171 bl_171 br_171 wl_35 vdd gnd cell_6t
Xbit_r36_c171 bl_171 br_171 wl_36 vdd gnd cell_6t
Xbit_r37_c171 bl_171 br_171 wl_37 vdd gnd cell_6t
Xbit_r38_c171 bl_171 br_171 wl_38 vdd gnd cell_6t
Xbit_r39_c171 bl_171 br_171 wl_39 vdd gnd cell_6t
Xbit_r40_c171 bl_171 br_171 wl_40 vdd gnd cell_6t
Xbit_r41_c171 bl_171 br_171 wl_41 vdd gnd cell_6t
Xbit_r42_c171 bl_171 br_171 wl_42 vdd gnd cell_6t
Xbit_r43_c171 bl_171 br_171 wl_43 vdd gnd cell_6t
Xbit_r44_c171 bl_171 br_171 wl_44 vdd gnd cell_6t
Xbit_r45_c171 bl_171 br_171 wl_45 vdd gnd cell_6t
Xbit_r46_c171 bl_171 br_171 wl_46 vdd gnd cell_6t
Xbit_r47_c171 bl_171 br_171 wl_47 vdd gnd cell_6t
Xbit_r48_c171 bl_171 br_171 wl_48 vdd gnd cell_6t
Xbit_r49_c171 bl_171 br_171 wl_49 vdd gnd cell_6t
Xbit_r50_c171 bl_171 br_171 wl_50 vdd gnd cell_6t
Xbit_r51_c171 bl_171 br_171 wl_51 vdd gnd cell_6t
Xbit_r52_c171 bl_171 br_171 wl_52 vdd gnd cell_6t
Xbit_r53_c171 bl_171 br_171 wl_53 vdd gnd cell_6t
Xbit_r54_c171 bl_171 br_171 wl_54 vdd gnd cell_6t
Xbit_r55_c171 bl_171 br_171 wl_55 vdd gnd cell_6t
Xbit_r56_c171 bl_171 br_171 wl_56 vdd gnd cell_6t
Xbit_r57_c171 bl_171 br_171 wl_57 vdd gnd cell_6t
Xbit_r58_c171 bl_171 br_171 wl_58 vdd gnd cell_6t
Xbit_r59_c171 bl_171 br_171 wl_59 vdd gnd cell_6t
Xbit_r60_c171 bl_171 br_171 wl_60 vdd gnd cell_6t
Xbit_r61_c171 bl_171 br_171 wl_61 vdd gnd cell_6t
Xbit_r62_c171 bl_171 br_171 wl_62 vdd gnd cell_6t
Xbit_r63_c171 bl_171 br_171 wl_63 vdd gnd cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd cell_6t
Xbit_r1_c172 bl_172 br_172 wl_1 vdd gnd cell_6t
Xbit_r2_c172 bl_172 br_172 wl_2 vdd gnd cell_6t
Xbit_r3_c172 bl_172 br_172 wl_3 vdd gnd cell_6t
Xbit_r4_c172 bl_172 br_172 wl_4 vdd gnd cell_6t
Xbit_r5_c172 bl_172 br_172 wl_5 vdd gnd cell_6t
Xbit_r6_c172 bl_172 br_172 wl_6 vdd gnd cell_6t
Xbit_r7_c172 bl_172 br_172 wl_7 vdd gnd cell_6t
Xbit_r8_c172 bl_172 br_172 wl_8 vdd gnd cell_6t
Xbit_r9_c172 bl_172 br_172 wl_9 vdd gnd cell_6t
Xbit_r10_c172 bl_172 br_172 wl_10 vdd gnd cell_6t
Xbit_r11_c172 bl_172 br_172 wl_11 vdd gnd cell_6t
Xbit_r12_c172 bl_172 br_172 wl_12 vdd gnd cell_6t
Xbit_r13_c172 bl_172 br_172 wl_13 vdd gnd cell_6t
Xbit_r14_c172 bl_172 br_172 wl_14 vdd gnd cell_6t
Xbit_r15_c172 bl_172 br_172 wl_15 vdd gnd cell_6t
Xbit_r16_c172 bl_172 br_172 wl_16 vdd gnd cell_6t
Xbit_r17_c172 bl_172 br_172 wl_17 vdd gnd cell_6t
Xbit_r18_c172 bl_172 br_172 wl_18 vdd gnd cell_6t
Xbit_r19_c172 bl_172 br_172 wl_19 vdd gnd cell_6t
Xbit_r20_c172 bl_172 br_172 wl_20 vdd gnd cell_6t
Xbit_r21_c172 bl_172 br_172 wl_21 vdd gnd cell_6t
Xbit_r22_c172 bl_172 br_172 wl_22 vdd gnd cell_6t
Xbit_r23_c172 bl_172 br_172 wl_23 vdd gnd cell_6t
Xbit_r24_c172 bl_172 br_172 wl_24 vdd gnd cell_6t
Xbit_r25_c172 bl_172 br_172 wl_25 vdd gnd cell_6t
Xbit_r26_c172 bl_172 br_172 wl_26 vdd gnd cell_6t
Xbit_r27_c172 bl_172 br_172 wl_27 vdd gnd cell_6t
Xbit_r28_c172 bl_172 br_172 wl_28 vdd gnd cell_6t
Xbit_r29_c172 bl_172 br_172 wl_29 vdd gnd cell_6t
Xbit_r30_c172 bl_172 br_172 wl_30 vdd gnd cell_6t
Xbit_r31_c172 bl_172 br_172 wl_31 vdd gnd cell_6t
Xbit_r32_c172 bl_172 br_172 wl_32 vdd gnd cell_6t
Xbit_r33_c172 bl_172 br_172 wl_33 vdd gnd cell_6t
Xbit_r34_c172 bl_172 br_172 wl_34 vdd gnd cell_6t
Xbit_r35_c172 bl_172 br_172 wl_35 vdd gnd cell_6t
Xbit_r36_c172 bl_172 br_172 wl_36 vdd gnd cell_6t
Xbit_r37_c172 bl_172 br_172 wl_37 vdd gnd cell_6t
Xbit_r38_c172 bl_172 br_172 wl_38 vdd gnd cell_6t
Xbit_r39_c172 bl_172 br_172 wl_39 vdd gnd cell_6t
Xbit_r40_c172 bl_172 br_172 wl_40 vdd gnd cell_6t
Xbit_r41_c172 bl_172 br_172 wl_41 vdd gnd cell_6t
Xbit_r42_c172 bl_172 br_172 wl_42 vdd gnd cell_6t
Xbit_r43_c172 bl_172 br_172 wl_43 vdd gnd cell_6t
Xbit_r44_c172 bl_172 br_172 wl_44 vdd gnd cell_6t
Xbit_r45_c172 bl_172 br_172 wl_45 vdd gnd cell_6t
Xbit_r46_c172 bl_172 br_172 wl_46 vdd gnd cell_6t
Xbit_r47_c172 bl_172 br_172 wl_47 vdd gnd cell_6t
Xbit_r48_c172 bl_172 br_172 wl_48 vdd gnd cell_6t
Xbit_r49_c172 bl_172 br_172 wl_49 vdd gnd cell_6t
Xbit_r50_c172 bl_172 br_172 wl_50 vdd gnd cell_6t
Xbit_r51_c172 bl_172 br_172 wl_51 vdd gnd cell_6t
Xbit_r52_c172 bl_172 br_172 wl_52 vdd gnd cell_6t
Xbit_r53_c172 bl_172 br_172 wl_53 vdd gnd cell_6t
Xbit_r54_c172 bl_172 br_172 wl_54 vdd gnd cell_6t
Xbit_r55_c172 bl_172 br_172 wl_55 vdd gnd cell_6t
Xbit_r56_c172 bl_172 br_172 wl_56 vdd gnd cell_6t
Xbit_r57_c172 bl_172 br_172 wl_57 vdd gnd cell_6t
Xbit_r58_c172 bl_172 br_172 wl_58 vdd gnd cell_6t
Xbit_r59_c172 bl_172 br_172 wl_59 vdd gnd cell_6t
Xbit_r60_c172 bl_172 br_172 wl_60 vdd gnd cell_6t
Xbit_r61_c172 bl_172 br_172 wl_61 vdd gnd cell_6t
Xbit_r62_c172 bl_172 br_172 wl_62 vdd gnd cell_6t
Xbit_r63_c172 bl_172 br_172 wl_63 vdd gnd cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd cell_6t
Xbit_r1_c173 bl_173 br_173 wl_1 vdd gnd cell_6t
Xbit_r2_c173 bl_173 br_173 wl_2 vdd gnd cell_6t
Xbit_r3_c173 bl_173 br_173 wl_3 vdd gnd cell_6t
Xbit_r4_c173 bl_173 br_173 wl_4 vdd gnd cell_6t
Xbit_r5_c173 bl_173 br_173 wl_5 vdd gnd cell_6t
Xbit_r6_c173 bl_173 br_173 wl_6 vdd gnd cell_6t
Xbit_r7_c173 bl_173 br_173 wl_7 vdd gnd cell_6t
Xbit_r8_c173 bl_173 br_173 wl_8 vdd gnd cell_6t
Xbit_r9_c173 bl_173 br_173 wl_9 vdd gnd cell_6t
Xbit_r10_c173 bl_173 br_173 wl_10 vdd gnd cell_6t
Xbit_r11_c173 bl_173 br_173 wl_11 vdd gnd cell_6t
Xbit_r12_c173 bl_173 br_173 wl_12 vdd gnd cell_6t
Xbit_r13_c173 bl_173 br_173 wl_13 vdd gnd cell_6t
Xbit_r14_c173 bl_173 br_173 wl_14 vdd gnd cell_6t
Xbit_r15_c173 bl_173 br_173 wl_15 vdd gnd cell_6t
Xbit_r16_c173 bl_173 br_173 wl_16 vdd gnd cell_6t
Xbit_r17_c173 bl_173 br_173 wl_17 vdd gnd cell_6t
Xbit_r18_c173 bl_173 br_173 wl_18 vdd gnd cell_6t
Xbit_r19_c173 bl_173 br_173 wl_19 vdd gnd cell_6t
Xbit_r20_c173 bl_173 br_173 wl_20 vdd gnd cell_6t
Xbit_r21_c173 bl_173 br_173 wl_21 vdd gnd cell_6t
Xbit_r22_c173 bl_173 br_173 wl_22 vdd gnd cell_6t
Xbit_r23_c173 bl_173 br_173 wl_23 vdd gnd cell_6t
Xbit_r24_c173 bl_173 br_173 wl_24 vdd gnd cell_6t
Xbit_r25_c173 bl_173 br_173 wl_25 vdd gnd cell_6t
Xbit_r26_c173 bl_173 br_173 wl_26 vdd gnd cell_6t
Xbit_r27_c173 bl_173 br_173 wl_27 vdd gnd cell_6t
Xbit_r28_c173 bl_173 br_173 wl_28 vdd gnd cell_6t
Xbit_r29_c173 bl_173 br_173 wl_29 vdd gnd cell_6t
Xbit_r30_c173 bl_173 br_173 wl_30 vdd gnd cell_6t
Xbit_r31_c173 bl_173 br_173 wl_31 vdd gnd cell_6t
Xbit_r32_c173 bl_173 br_173 wl_32 vdd gnd cell_6t
Xbit_r33_c173 bl_173 br_173 wl_33 vdd gnd cell_6t
Xbit_r34_c173 bl_173 br_173 wl_34 vdd gnd cell_6t
Xbit_r35_c173 bl_173 br_173 wl_35 vdd gnd cell_6t
Xbit_r36_c173 bl_173 br_173 wl_36 vdd gnd cell_6t
Xbit_r37_c173 bl_173 br_173 wl_37 vdd gnd cell_6t
Xbit_r38_c173 bl_173 br_173 wl_38 vdd gnd cell_6t
Xbit_r39_c173 bl_173 br_173 wl_39 vdd gnd cell_6t
Xbit_r40_c173 bl_173 br_173 wl_40 vdd gnd cell_6t
Xbit_r41_c173 bl_173 br_173 wl_41 vdd gnd cell_6t
Xbit_r42_c173 bl_173 br_173 wl_42 vdd gnd cell_6t
Xbit_r43_c173 bl_173 br_173 wl_43 vdd gnd cell_6t
Xbit_r44_c173 bl_173 br_173 wl_44 vdd gnd cell_6t
Xbit_r45_c173 bl_173 br_173 wl_45 vdd gnd cell_6t
Xbit_r46_c173 bl_173 br_173 wl_46 vdd gnd cell_6t
Xbit_r47_c173 bl_173 br_173 wl_47 vdd gnd cell_6t
Xbit_r48_c173 bl_173 br_173 wl_48 vdd gnd cell_6t
Xbit_r49_c173 bl_173 br_173 wl_49 vdd gnd cell_6t
Xbit_r50_c173 bl_173 br_173 wl_50 vdd gnd cell_6t
Xbit_r51_c173 bl_173 br_173 wl_51 vdd gnd cell_6t
Xbit_r52_c173 bl_173 br_173 wl_52 vdd gnd cell_6t
Xbit_r53_c173 bl_173 br_173 wl_53 vdd gnd cell_6t
Xbit_r54_c173 bl_173 br_173 wl_54 vdd gnd cell_6t
Xbit_r55_c173 bl_173 br_173 wl_55 vdd gnd cell_6t
Xbit_r56_c173 bl_173 br_173 wl_56 vdd gnd cell_6t
Xbit_r57_c173 bl_173 br_173 wl_57 vdd gnd cell_6t
Xbit_r58_c173 bl_173 br_173 wl_58 vdd gnd cell_6t
Xbit_r59_c173 bl_173 br_173 wl_59 vdd gnd cell_6t
Xbit_r60_c173 bl_173 br_173 wl_60 vdd gnd cell_6t
Xbit_r61_c173 bl_173 br_173 wl_61 vdd gnd cell_6t
Xbit_r62_c173 bl_173 br_173 wl_62 vdd gnd cell_6t
Xbit_r63_c173 bl_173 br_173 wl_63 vdd gnd cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd cell_6t
Xbit_r1_c174 bl_174 br_174 wl_1 vdd gnd cell_6t
Xbit_r2_c174 bl_174 br_174 wl_2 vdd gnd cell_6t
Xbit_r3_c174 bl_174 br_174 wl_3 vdd gnd cell_6t
Xbit_r4_c174 bl_174 br_174 wl_4 vdd gnd cell_6t
Xbit_r5_c174 bl_174 br_174 wl_5 vdd gnd cell_6t
Xbit_r6_c174 bl_174 br_174 wl_6 vdd gnd cell_6t
Xbit_r7_c174 bl_174 br_174 wl_7 vdd gnd cell_6t
Xbit_r8_c174 bl_174 br_174 wl_8 vdd gnd cell_6t
Xbit_r9_c174 bl_174 br_174 wl_9 vdd gnd cell_6t
Xbit_r10_c174 bl_174 br_174 wl_10 vdd gnd cell_6t
Xbit_r11_c174 bl_174 br_174 wl_11 vdd gnd cell_6t
Xbit_r12_c174 bl_174 br_174 wl_12 vdd gnd cell_6t
Xbit_r13_c174 bl_174 br_174 wl_13 vdd gnd cell_6t
Xbit_r14_c174 bl_174 br_174 wl_14 vdd gnd cell_6t
Xbit_r15_c174 bl_174 br_174 wl_15 vdd gnd cell_6t
Xbit_r16_c174 bl_174 br_174 wl_16 vdd gnd cell_6t
Xbit_r17_c174 bl_174 br_174 wl_17 vdd gnd cell_6t
Xbit_r18_c174 bl_174 br_174 wl_18 vdd gnd cell_6t
Xbit_r19_c174 bl_174 br_174 wl_19 vdd gnd cell_6t
Xbit_r20_c174 bl_174 br_174 wl_20 vdd gnd cell_6t
Xbit_r21_c174 bl_174 br_174 wl_21 vdd gnd cell_6t
Xbit_r22_c174 bl_174 br_174 wl_22 vdd gnd cell_6t
Xbit_r23_c174 bl_174 br_174 wl_23 vdd gnd cell_6t
Xbit_r24_c174 bl_174 br_174 wl_24 vdd gnd cell_6t
Xbit_r25_c174 bl_174 br_174 wl_25 vdd gnd cell_6t
Xbit_r26_c174 bl_174 br_174 wl_26 vdd gnd cell_6t
Xbit_r27_c174 bl_174 br_174 wl_27 vdd gnd cell_6t
Xbit_r28_c174 bl_174 br_174 wl_28 vdd gnd cell_6t
Xbit_r29_c174 bl_174 br_174 wl_29 vdd gnd cell_6t
Xbit_r30_c174 bl_174 br_174 wl_30 vdd gnd cell_6t
Xbit_r31_c174 bl_174 br_174 wl_31 vdd gnd cell_6t
Xbit_r32_c174 bl_174 br_174 wl_32 vdd gnd cell_6t
Xbit_r33_c174 bl_174 br_174 wl_33 vdd gnd cell_6t
Xbit_r34_c174 bl_174 br_174 wl_34 vdd gnd cell_6t
Xbit_r35_c174 bl_174 br_174 wl_35 vdd gnd cell_6t
Xbit_r36_c174 bl_174 br_174 wl_36 vdd gnd cell_6t
Xbit_r37_c174 bl_174 br_174 wl_37 vdd gnd cell_6t
Xbit_r38_c174 bl_174 br_174 wl_38 vdd gnd cell_6t
Xbit_r39_c174 bl_174 br_174 wl_39 vdd gnd cell_6t
Xbit_r40_c174 bl_174 br_174 wl_40 vdd gnd cell_6t
Xbit_r41_c174 bl_174 br_174 wl_41 vdd gnd cell_6t
Xbit_r42_c174 bl_174 br_174 wl_42 vdd gnd cell_6t
Xbit_r43_c174 bl_174 br_174 wl_43 vdd gnd cell_6t
Xbit_r44_c174 bl_174 br_174 wl_44 vdd gnd cell_6t
Xbit_r45_c174 bl_174 br_174 wl_45 vdd gnd cell_6t
Xbit_r46_c174 bl_174 br_174 wl_46 vdd gnd cell_6t
Xbit_r47_c174 bl_174 br_174 wl_47 vdd gnd cell_6t
Xbit_r48_c174 bl_174 br_174 wl_48 vdd gnd cell_6t
Xbit_r49_c174 bl_174 br_174 wl_49 vdd gnd cell_6t
Xbit_r50_c174 bl_174 br_174 wl_50 vdd gnd cell_6t
Xbit_r51_c174 bl_174 br_174 wl_51 vdd gnd cell_6t
Xbit_r52_c174 bl_174 br_174 wl_52 vdd gnd cell_6t
Xbit_r53_c174 bl_174 br_174 wl_53 vdd gnd cell_6t
Xbit_r54_c174 bl_174 br_174 wl_54 vdd gnd cell_6t
Xbit_r55_c174 bl_174 br_174 wl_55 vdd gnd cell_6t
Xbit_r56_c174 bl_174 br_174 wl_56 vdd gnd cell_6t
Xbit_r57_c174 bl_174 br_174 wl_57 vdd gnd cell_6t
Xbit_r58_c174 bl_174 br_174 wl_58 vdd gnd cell_6t
Xbit_r59_c174 bl_174 br_174 wl_59 vdd gnd cell_6t
Xbit_r60_c174 bl_174 br_174 wl_60 vdd gnd cell_6t
Xbit_r61_c174 bl_174 br_174 wl_61 vdd gnd cell_6t
Xbit_r62_c174 bl_174 br_174 wl_62 vdd gnd cell_6t
Xbit_r63_c174 bl_174 br_174 wl_63 vdd gnd cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd cell_6t
Xbit_r1_c175 bl_175 br_175 wl_1 vdd gnd cell_6t
Xbit_r2_c175 bl_175 br_175 wl_2 vdd gnd cell_6t
Xbit_r3_c175 bl_175 br_175 wl_3 vdd gnd cell_6t
Xbit_r4_c175 bl_175 br_175 wl_4 vdd gnd cell_6t
Xbit_r5_c175 bl_175 br_175 wl_5 vdd gnd cell_6t
Xbit_r6_c175 bl_175 br_175 wl_6 vdd gnd cell_6t
Xbit_r7_c175 bl_175 br_175 wl_7 vdd gnd cell_6t
Xbit_r8_c175 bl_175 br_175 wl_8 vdd gnd cell_6t
Xbit_r9_c175 bl_175 br_175 wl_9 vdd gnd cell_6t
Xbit_r10_c175 bl_175 br_175 wl_10 vdd gnd cell_6t
Xbit_r11_c175 bl_175 br_175 wl_11 vdd gnd cell_6t
Xbit_r12_c175 bl_175 br_175 wl_12 vdd gnd cell_6t
Xbit_r13_c175 bl_175 br_175 wl_13 vdd gnd cell_6t
Xbit_r14_c175 bl_175 br_175 wl_14 vdd gnd cell_6t
Xbit_r15_c175 bl_175 br_175 wl_15 vdd gnd cell_6t
Xbit_r16_c175 bl_175 br_175 wl_16 vdd gnd cell_6t
Xbit_r17_c175 bl_175 br_175 wl_17 vdd gnd cell_6t
Xbit_r18_c175 bl_175 br_175 wl_18 vdd gnd cell_6t
Xbit_r19_c175 bl_175 br_175 wl_19 vdd gnd cell_6t
Xbit_r20_c175 bl_175 br_175 wl_20 vdd gnd cell_6t
Xbit_r21_c175 bl_175 br_175 wl_21 vdd gnd cell_6t
Xbit_r22_c175 bl_175 br_175 wl_22 vdd gnd cell_6t
Xbit_r23_c175 bl_175 br_175 wl_23 vdd gnd cell_6t
Xbit_r24_c175 bl_175 br_175 wl_24 vdd gnd cell_6t
Xbit_r25_c175 bl_175 br_175 wl_25 vdd gnd cell_6t
Xbit_r26_c175 bl_175 br_175 wl_26 vdd gnd cell_6t
Xbit_r27_c175 bl_175 br_175 wl_27 vdd gnd cell_6t
Xbit_r28_c175 bl_175 br_175 wl_28 vdd gnd cell_6t
Xbit_r29_c175 bl_175 br_175 wl_29 vdd gnd cell_6t
Xbit_r30_c175 bl_175 br_175 wl_30 vdd gnd cell_6t
Xbit_r31_c175 bl_175 br_175 wl_31 vdd gnd cell_6t
Xbit_r32_c175 bl_175 br_175 wl_32 vdd gnd cell_6t
Xbit_r33_c175 bl_175 br_175 wl_33 vdd gnd cell_6t
Xbit_r34_c175 bl_175 br_175 wl_34 vdd gnd cell_6t
Xbit_r35_c175 bl_175 br_175 wl_35 vdd gnd cell_6t
Xbit_r36_c175 bl_175 br_175 wl_36 vdd gnd cell_6t
Xbit_r37_c175 bl_175 br_175 wl_37 vdd gnd cell_6t
Xbit_r38_c175 bl_175 br_175 wl_38 vdd gnd cell_6t
Xbit_r39_c175 bl_175 br_175 wl_39 vdd gnd cell_6t
Xbit_r40_c175 bl_175 br_175 wl_40 vdd gnd cell_6t
Xbit_r41_c175 bl_175 br_175 wl_41 vdd gnd cell_6t
Xbit_r42_c175 bl_175 br_175 wl_42 vdd gnd cell_6t
Xbit_r43_c175 bl_175 br_175 wl_43 vdd gnd cell_6t
Xbit_r44_c175 bl_175 br_175 wl_44 vdd gnd cell_6t
Xbit_r45_c175 bl_175 br_175 wl_45 vdd gnd cell_6t
Xbit_r46_c175 bl_175 br_175 wl_46 vdd gnd cell_6t
Xbit_r47_c175 bl_175 br_175 wl_47 vdd gnd cell_6t
Xbit_r48_c175 bl_175 br_175 wl_48 vdd gnd cell_6t
Xbit_r49_c175 bl_175 br_175 wl_49 vdd gnd cell_6t
Xbit_r50_c175 bl_175 br_175 wl_50 vdd gnd cell_6t
Xbit_r51_c175 bl_175 br_175 wl_51 vdd gnd cell_6t
Xbit_r52_c175 bl_175 br_175 wl_52 vdd gnd cell_6t
Xbit_r53_c175 bl_175 br_175 wl_53 vdd gnd cell_6t
Xbit_r54_c175 bl_175 br_175 wl_54 vdd gnd cell_6t
Xbit_r55_c175 bl_175 br_175 wl_55 vdd gnd cell_6t
Xbit_r56_c175 bl_175 br_175 wl_56 vdd gnd cell_6t
Xbit_r57_c175 bl_175 br_175 wl_57 vdd gnd cell_6t
Xbit_r58_c175 bl_175 br_175 wl_58 vdd gnd cell_6t
Xbit_r59_c175 bl_175 br_175 wl_59 vdd gnd cell_6t
Xbit_r60_c175 bl_175 br_175 wl_60 vdd gnd cell_6t
Xbit_r61_c175 bl_175 br_175 wl_61 vdd gnd cell_6t
Xbit_r62_c175 bl_175 br_175 wl_62 vdd gnd cell_6t
Xbit_r63_c175 bl_175 br_175 wl_63 vdd gnd cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd cell_6t
Xbit_r1_c176 bl_176 br_176 wl_1 vdd gnd cell_6t
Xbit_r2_c176 bl_176 br_176 wl_2 vdd gnd cell_6t
Xbit_r3_c176 bl_176 br_176 wl_3 vdd gnd cell_6t
Xbit_r4_c176 bl_176 br_176 wl_4 vdd gnd cell_6t
Xbit_r5_c176 bl_176 br_176 wl_5 vdd gnd cell_6t
Xbit_r6_c176 bl_176 br_176 wl_6 vdd gnd cell_6t
Xbit_r7_c176 bl_176 br_176 wl_7 vdd gnd cell_6t
Xbit_r8_c176 bl_176 br_176 wl_8 vdd gnd cell_6t
Xbit_r9_c176 bl_176 br_176 wl_9 vdd gnd cell_6t
Xbit_r10_c176 bl_176 br_176 wl_10 vdd gnd cell_6t
Xbit_r11_c176 bl_176 br_176 wl_11 vdd gnd cell_6t
Xbit_r12_c176 bl_176 br_176 wl_12 vdd gnd cell_6t
Xbit_r13_c176 bl_176 br_176 wl_13 vdd gnd cell_6t
Xbit_r14_c176 bl_176 br_176 wl_14 vdd gnd cell_6t
Xbit_r15_c176 bl_176 br_176 wl_15 vdd gnd cell_6t
Xbit_r16_c176 bl_176 br_176 wl_16 vdd gnd cell_6t
Xbit_r17_c176 bl_176 br_176 wl_17 vdd gnd cell_6t
Xbit_r18_c176 bl_176 br_176 wl_18 vdd gnd cell_6t
Xbit_r19_c176 bl_176 br_176 wl_19 vdd gnd cell_6t
Xbit_r20_c176 bl_176 br_176 wl_20 vdd gnd cell_6t
Xbit_r21_c176 bl_176 br_176 wl_21 vdd gnd cell_6t
Xbit_r22_c176 bl_176 br_176 wl_22 vdd gnd cell_6t
Xbit_r23_c176 bl_176 br_176 wl_23 vdd gnd cell_6t
Xbit_r24_c176 bl_176 br_176 wl_24 vdd gnd cell_6t
Xbit_r25_c176 bl_176 br_176 wl_25 vdd gnd cell_6t
Xbit_r26_c176 bl_176 br_176 wl_26 vdd gnd cell_6t
Xbit_r27_c176 bl_176 br_176 wl_27 vdd gnd cell_6t
Xbit_r28_c176 bl_176 br_176 wl_28 vdd gnd cell_6t
Xbit_r29_c176 bl_176 br_176 wl_29 vdd gnd cell_6t
Xbit_r30_c176 bl_176 br_176 wl_30 vdd gnd cell_6t
Xbit_r31_c176 bl_176 br_176 wl_31 vdd gnd cell_6t
Xbit_r32_c176 bl_176 br_176 wl_32 vdd gnd cell_6t
Xbit_r33_c176 bl_176 br_176 wl_33 vdd gnd cell_6t
Xbit_r34_c176 bl_176 br_176 wl_34 vdd gnd cell_6t
Xbit_r35_c176 bl_176 br_176 wl_35 vdd gnd cell_6t
Xbit_r36_c176 bl_176 br_176 wl_36 vdd gnd cell_6t
Xbit_r37_c176 bl_176 br_176 wl_37 vdd gnd cell_6t
Xbit_r38_c176 bl_176 br_176 wl_38 vdd gnd cell_6t
Xbit_r39_c176 bl_176 br_176 wl_39 vdd gnd cell_6t
Xbit_r40_c176 bl_176 br_176 wl_40 vdd gnd cell_6t
Xbit_r41_c176 bl_176 br_176 wl_41 vdd gnd cell_6t
Xbit_r42_c176 bl_176 br_176 wl_42 vdd gnd cell_6t
Xbit_r43_c176 bl_176 br_176 wl_43 vdd gnd cell_6t
Xbit_r44_c176 bl_176 br_176 wl_44 vdd gnd cell_6t
Xbit_r45_c176 bl_176 br_176 wl_45 vdd gnd cell_6t
Xbit_r46_c176 bl_176 br_176 wl_46 vdd gnd cell_6t
Xbit_r47_c176 bl_176 br_176 wl_47 vdd gnd cell_6t
Xbit_r48_c176 bl_176 br_176 wl_48 vdd gnd cell_6t
Xbit_r49_c176 bl_176 br_176 wl_49 vdd gnd cell_6t
Xbit_r50_c176 bl_176 br_176 wl_50 vdd gnd cell_6t
Xbit_r51_c176 bl_176 br_176 wl_51 vdd gnd cell_6t
Xbit_r52_c176 bl_176 br_176 wl_52 vdd gnd cell_6t
Xbit_r53_c176 bl_176 br_176 wl_53 vdd gnd cell_6t
Xbit_r54_c176 bl_176 br_176 wl_54 vdd gnd cell_6t
Xbit_r55_c176 bl_176 br_176 wl_55 vdd gnd cell_6t
Xbit_r56_c176 bl_176 br_176 wl_56 vdd gnd cell_6t
Xbit_r57_c176 bl_176 br_176 wl_57 vdd gnd cell_6t
Xbit_r58_c176 bl_176 br_176 wl_58 vdd gnd cell_6t
Xbit_r59_c176 bl_176 br_176 wl_59 vdd gnd cell_6t
Xbit_r60_c176 bl_176 br_176 wl_60 vdd gnd cell_6t
Xbit_r61_c176 bl_176 br_176 wl_61 vdd gnd cell_6t
Xbit_r62_c176 bl_176 br_176 wl_62 vdd gnd cell_6t
Xbit_r63_c176 bl_176 br_176 wl_63 vdd gnd cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd cell_6t
Xbit_r1_c177 bl_177 br_177 wl_1 vdd gnd cell_6t
Xbit_r2_c177 bl_177 br_177 wl_2 vdd gnd cell_6t
Xbit_r3_c177 bl_177 br_177 wl_3 vdd gnd cell_6t
Xbit_r4_c177 bl_177 br_177 wl_4 vdd gnd cell_6t
Xbit_r5_c177 bl_177 br_177 wl_5 vdd gnd cell_6t
Xbit_r6_c177 bl_177 br_177 wl_6 vdd gnd cell_6t
Xbit_r7_c177 bl_177 br_177 wl_7 vdd gnd cell_6t
Xbit_r8_c177 bl_177 br_177 wl_8 vdd gnd cell_6t
Xbit_r9_c177 bl_177 br_177 wl_9 vdd gnd cell_6t
Xbit_r10_c177 bl_177 br_177 wl_10 vdd gnd cell_6t
Xbit_r11_c177 bl_177 br_177 wl_11 vdd gnd cell_6t
Xbit_r12_c177 bl_177 br_177 wl_12 vdd gnd cell_6t
Xbit_r13_c177 bl_177 br_177 wl_13 vdd gnd cell_6t
Xbit_r14_c177 bl_177 br_177 wl_14 vdd gnd cell_6t
Xbit_r15_c177 bl_177 br_177 wl_15 vdd gnd cell_6t
Xbit_r16_c177 bl_177 br_177 wl_16 vdd gnd cell_6t
Xbit_r17_c177 bl_177 br_177 wl_17 vdd gnd cell_6t
Xbit_r18_c177 bl_177 br_177 wl_18 vdd gnd cell_6t
Xbit_r19_c177 bl_177 br_177 wl_19 vdd gnd cell_6t
Xbit_r20_c177 bl_177 br_177 wl_20 vdd gnd cell_6t
Xbit_r21_c177 bl_177 br_177 wl_21 vdd gnd cell_6t
Xbit_r22_c177 bl_177 br_177 wl_22 vdd gnd cell_6t
Xbit_r23_c177 bl_177 br_177 wl_23 vdd gnd cell_6t
Xbit_r24_c177 bl_177 br_177 wl_24 vdd gnd cell_6t
Xbit_r25_c177 bl_177 br_177 wl_25 vdd gnd cell_6t
Xbit_r26_c177 bl_177 br_177 wl_26 vdd gnd cell_6t
Xbit_r27_c177 bl_177 br_177 wl_27 vdd gnd cell_6t
Xbit_r28_c177 bl_177 br_177 wl_28 vdd gnd cell_6t
Xbit_r29_c177 bl_177 br_177 wl_29 vdd gnd cell_6t
Xbit_r30_c177 bl_177 br_177 wl_30 vdd gnd cell_6t
Xbit_r31_c177 bl_177 br_177 wl_31 vdd gnd cell_6t
Xbit_r32_c177 bl_177 br_177 wl_32 vdd gnd cell_6t
Xbit_r33_c177 bl_177 br_177 wl_33 vdd gnd cell_6t
Xbit_r34_c177 bl_177 br_177 wl_34 vdd gnd cell_6t
Xbit_r35_c177 bl_177 br_177 wl_35 vdd gnd cell_6t
Xbit_r36_c177 bl_177 br_177 wl_36 vdd gnd cell_6t
Xbit_r37_c177 bl_177 br_177 wl_37 vdd gnd cell_6t
Xbit_r38_c177 bl_177 br_177 wl_38 vdd gnd cell_6t
Xbit_r39_c177 bl_177 br_177 wl_39 vdd gnd cell_6t
Xbit_r40_c177 bl_177 br_177 wl_40 vdd gnd cell_6t
Xbit_r41_c177 bl_177 br_177 wl_41 vdd gnd cell_6t
Xbit_r42_c177 bl_177 br_177 wl_42 vdd gnd cell_6t
Xbit_r43_c177 bl_177 br_177 wl_43 vdd gnd cell_6t
Xbit_r44_c177 bl_177 br_177 wl_44 vdd gnd cell_6t
Xbit_r45_c177 bl_177 br_177 wl_45 vdd gnd cell_6t
Xbit_r46_c177 bl_177 br_177 wl_46 vdd gnd cell_6t
Xbit_r47_c177 bl_177 br_177 wl_47 vdd gnd cell_6t
Xbit_r48_c177 bl_177 br_177 wl_48 vdd gnd cell_6t
Xbit_r49_c177 bl_177 br_177 wl_49 vdd gnd cell_6t
Xbit_r50_c177 bl_177 br_177 wl_50 vdd gnd cell_6t
Xbit_r51_c177 bl_177 br_177 wl_51 vdd gnd cell_6t
Xbit_r52_c177 bl_177 br_177 wl_52 vdd gnd cell_6t
Xbit_r53_c177 bl_177 br_177 wl_53 vdd gnd cell_6t
Xbit_r54_c177 bl_177 br_177 wl_54 vdd gnd cell_6t
Xbit_r55_c177 bl_177 br_177 wl_55 vdd gnd cell_6t
Xbit_r56_c177 bl_177 br_177 wl_56 vdd gnd cell_6t
Xbit_r57_c177 bl_177 br_177 wl_57 vdd gnd cell_6t
Xbit_r58_c177 bl_177 br_177 wl_58 vdd gnd cell_6t
Xbit_r59_c177 bl_177 br_177 wl_59 vdd gnd cell_6t
Xbit_r60_c177 bl_177 br_177 wl_60 vdd gnd cell_6t
Xbit_r61_c177 bl_177 br_177 wl_61 vdd gnd cell_6t
Xbit_r62_c177 bl_177 br_177 wl_62 vdd gnd cell_6t
Xbit_r63_c177 bl_177 br_177 wl_63 vdd gnd cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd cell_6t
Xbit_r1_c178 bl_178 br_178 wl_1 vdd gnd cell_6t
Xbit_r2_c178 bl_178 br_178 wl_2 vdd gnd cell_6t
Xbit_r3_c178 bl_178 br_178 wl_3 vdd gnd cell_6t
Xbit_r4_c178 bl_178 br_178 wl_4 vdd gnd cell_6t
Xbit_r5_c178 bl_178 br_178 wl_5 vdd gnd cell_6t
Xbit_r6_c178 bl_178 br_178 wl_6 vdd gnd cell_6t
Xbit_r7_c178 bl_178 br_178 wl_7 vdd gnd cell_6t
Xbit_r8_c178 bl_178 br_178 wl_8 vdd gnd cell_6t
Xbit_r9_c178 bl_178 br_178 wl_9 vdd gnd cell_6t
Xbit_r10_c178 bl_178 br_178 wl_10 vdd gnd cell_6t
Xbit_r11_c178 bl_178 br_178 wl_11 vdd gnd cell_6t
Xbit_r12_c178 bl_178 br_178 wl_12 vdd gnd cell_6t
Xbit_r13_c178 bl_178 br_178 wl_13 vdd gnd cell_6t
Xbit_r14_c178 bl_178 br_178 wl_14 vdd gnd cell_6t
Xbit_r15_c178 bl_178 br_178 wl_15 vdd gnd cell_6t
Xbit_r16_c178 bl_178 br_178 wl_16 vdd gnd cell_6t
Xbit_r17_c178 bl_178 br_178 wl_17 vdd gnd cell_6t
Xbit_r18_c178 bl_178 br_178 wl_18 vdd gnd cell_6t
Xbit_r19_c178 bl_178 br_178 wl_19 vdd gnd cell_6t
Xbit_r20_c178 bl_178 br_178 wl_20 vdd gnd cell_6t
Xbit_r21_c178 bl_178 br_178 wl_21 vdd gnd cell_6t
Xbit_r22_c178 bl_178 br_178 wl_22 vdd gnd cell_6t
Xbit_r23_c178 bl_178 br_178 wl_23 vdd gnd cell_6t
Xbit_r24_c178 bl_178 br_178 wl_24 vdd gnd cell_6t
Xbit_r25_c178 bl_178 br_178 wl_25 vdd gnd cell_6t
Xbit_r26_c178 bl_178 br_178 wl_26 vdd gnd cell_6t
Xbit_r27_c178 bl_178 br_178 wl_27 vdd gnd cell_6t
Xbit_r28_c178 bl_178 br_178 wl_28 vdd gnd cell_6t
Xbit_r29_c178 bl_178 br_178 wl_29 vdd gnd cell_6t
Xbit_r30_c178 bl_178 br_178 wl_30 vdd gnd cell_6t
Xbit_r31_c178 bl_178 br_178 wl_31 vdd gnd cell_6t
Xbit_r32_c178 bl_178 br_178 wl_32 vdd gnd cell_6t
Xbit_r33_c178 bl_178 br_178 wl_33 vdd gnd cell_6t
Xbit_r34_c178 bl_178 br_178 wl_34 vdd gnd cell_6t
Xbit_r35_c178 bl_178 br_178 wl_35 vdd gnd cell_6t
Xbit_r36_c178 bl_178 br_178 wl_36 vdd gnd cell_6t
Xbit_r37_c178 bl_178 br_178 wl_37 vdd gnd cell_6t
Xbit_r38_c178 bl_178 br_178 wl_38 vdd gnd cell_6t
Xbit_r39_c178 bl_178 br_178 wl_39 vdd gnd cell_6t
Xbit_r40_c178 bl_178 br_178 wl_40 vdd gnd cell_6t
Xbit_r41_c178 bl_178 br_178 wl_41 vdd gnd cell_6t
Xbit_r42_c178 bl_178 br_178 wl_42 vdd gnd cell_6t
Xbit_r43_c178 bl_178 br_178 wl_43 vdd gnd cell_6t
Xbit_r44_c178 bl_178 br_178 wl_44 vdd gnd cell_6t
Xbit_r45_c178 bl_178 br_178 wl_45 vdd gnd cell_6t
Xbit_r46_c178 bl_178 br_178 wl_46 vdd gnd cell_6t
Xbit_r47_c178 bl_178 br_178 wl_47 vdd gnd cell_6t
Xbit_r48_c178 bl_178 br_178 wl_48 vdd gnd cell_6t
Xbit_r49_c178 bl_178 br_178 wl_49 vdd gnd cell_6t
Xbit_r50_c178 bl_178 br_178 wl_50 vdd gnd cell_6t
Xbit_r51_c178 bl_178 br_178 wl_51 vdd gnd cell_6t
Xbit_r52_c178 bl_178 br_178 wl_52 vdd gnd cell_6t
Xbit_r53_c178 bl_178 br_178 wl_53 vdd gnd cell_6t
Xbit_r54_c178 bl_178 br_178 wl_54 vdd gnd cell_6t
Xbit_r55_c178 bl_178 br_178 wl_55 vdd gnd cell_6t
Xbit_r56_c178 bl_178 br_178 wl_56 vdd gnd cell_6t
Xbit_r57_c178 bl_178 br_178 wl_57 vdd gnd cell_6t
Xbit_r58_c178 bl_178 br_178 wl_58 vdd gnd cell_6t
Xbit_r59_c178 bl_178 br_178 wl_59 vdd gnd cell_6t
Xbit_r60_c178 bl_178 br_178 wl_60 vdd gnd cell_6t
Xbit_r61_c178 bl_178 br_178 wl_61 vdd gnd cell_6t
Xbit_r62_c178 bl_178 br_178 wl_62 vdd gnd cell_6t
Xbit_r63_c178 bl_178 br_178 wl_63 vdd gnd cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd cell_6t
Xbit_r1_c179 bl_179 br_179 wl_1 vdd gnd cell_6t
Xbit_r2_c179 bl_179 br_179 wl_2 vdd gnd cell_6t
Xbit_r3_c179 bl_179 br_179 wl_3 vdd gnd cell_6t
Xbit_r4_c179 bl_179 br_179 wl_4 vdd gnd cell_6t
Xbit_r5_c179 bl_179 br_179 wl_5 vdd gnd cell_6t
Xbit_r6_c179 bl_179 br_179 wl_6 vdd gnd cell_6t
Xbit_r7_c179 bl_179 br_179 wl_7 vdd gnd cell_6t
Xbit_r8_c179 bl_179 br_179 wl_8 vdd gnd cell_6t
Xbit_r9_c179 bl_179 br_179 wl_9 vdd gnd cell_6t
Xbit_r10_c179 bl_179 br_179 wl_10 vdd gnd cell_6t
Xbit_r11_c179 bl_179 br_179 wl_11 vdd gnd cell_6t
Xbit_r12_c179 bl_179 br_179 wl_12 vdd gnd cell_6t
Xbit_r13_c179 bl_179 br_179 wl_13 vdd gnd cell_6t
Xbit_r14_c179 bl_179 br_179 wl_14 vdd gnd cell_6t
Xbit_r15_c179 bl_179 br_179 wl_15 vdd gnd cell_6t
Xbit_r16_c179 bl_179 br_179 wl_16 vdd gnd cell_6t
Xbit_r17_c179 bl_179 br_179 wl_17 vdd gnd cell_6t
Xbit_r18_c179 bl_179 br_179 wl_18 vdd gnd cell_6t
Xbit_r19_c179 bl_179 br_179 wl_19 vdd gnd cell_6t
Xbit_r20_c179 bl_179 br_179 wl_20 vdd gnd cell_6t
Xbit_r21_c179 bl_179 br_179 wl_21 vdd gnd cell_6t
Xbit_r22_c179 bl_179 br_179 wl_22 vdd gnd cell_6t
Xbit_r23_c179 bl_179 br_179 wl_23 vdd gnd cell_6t
Xbit_r24_c179 bl_179 br_179 wl_24 vdd gnd cell_6t
Xbit_r25_c179 bl_179 br_179 wl_25 vdd gnd cell_6t
Xbit_r26_c179 bl_179 br_179 wl_26 vdd gnd cell_6t
Xbit_r27_c179 bl_179 br_179 wl_27 vdd gnd cell_6t
Xbit_r28_c179 bl_179 br_179 wl_28 vdd gnd cell_6t
Xbit_r29_c179 bl_179 br_179 wl_29 vdd gnd cell_6t
Xbit_r30_c179 bl_179 br_179 wl_30 vdd gnd cell_6t
Xbit_r31_c179 bl_179 br_179 wl_31 vdd gnd cell_6t
Xbit_r32_c179 bl_179 br_179 wl_32 vdd gnd cell_6t
Xbit_r33_c179 bl_179 br_179 wl_33 vdd gnd cell_6t
Xbit_r34_c179 bl_179 br_179 wl_34 vdd gnd cell_6t
Xbit_r35_c179 bl_179 br_179 wl_35 vdd gnd cell_6t
Xbit_r36_c179 bl_179 br_179 wl_36 vdd gnd cell_6t
Xbit_r37_c179 bl_179 br_179 wl_37 vdd gnd cell_6t
Xbit_r38_c179 bl_179 br_179 wl_38 vdd gnd cell_6t
Xbit_r39_c179 bl_179 br_179 wl_39 vdd gnd cell_6t
Xbit_r40_c179 bl_179 br_179 wl_40 vdd gnd cell_6t
Xbit_r41_c179 bl_179 br_179 wl_41 vdd gnd cell_6t
Xbit_r42_c179 bl_179 br_179 wl_42 vdd gnd cell_6t
Xbit_r43_c179 bl_179 br_179 wl_43 vdd gnd cell_6t
Xbit_r44_c179 bl_179 br_179 wl_44 vdd gnd cell_6t
Xbit_r45_c179 bl_179 br_179 wl_45 vdd gnd cell_6t
Xbit_r46_c179 bl_179 br_179 wl_46 vdd gnd cell_6t
Xbit_r47_c179 bl_179 br_179 wl_47 vdd gnd cell_6t
Xbit_r48_c179 bl_179 br_179 wl_48 vdd gnd cell_6t
Xbit_r49_c179 bl_179 br_179 wl_49 vdd gnd cell_6t
Xbit_r50_c179 bl_179 br_179 wl_50 vdd gnd cell_6t
Xbit_r51_c179 bl_179 br_179 wl_51 vdd gnd cell_6t
Xbit_r52_c179 bl_179 br_179 wl_52 vdd gnd cell_6t
Xbit_r53_c179 bl_179 br_179 wl_53 vdd gnd cell_6t
Xbit_r54_c179 bl_179 br_179 wl_54 vdd gnd cell_6t
Xbit_r55_c179 bl_179 br_179 wl_55 vdd gnd cell_6t
Xbit_r56_c179 bl_179 br_179 wl_56 vdd gnd cell_6t
Xbit_r57_c179 bl_179 br_179 wl_57 vdd gnd cell_6t
Xbit_r58_c179 bl_179 br_179 wl_58 vdd gnd cell_6t
Xbit_r59_c179 bl_179 br_179 wl_59 vdd gnd cell_6t
Xbit_r60_c179 bl_179 br_179 wl_60 vdd gnd cell_6t
Xbit_r61_c179 bl_179 br_179 wl_61 vdd gnd cell_6t
Xbit_r62_c179 bl_179 br_179 wl_62 vdd gnd cell_6t
Xbit_r63_c179 bl_179 br_179 wl_63 vdd gnd cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd cell_6t
Xbit_r1_c180 bl_180 br_180 wl_1 vdd gnd cell_6t
Xbit_r2_c180 bl_180 br_180 wl_2 vdd gnd cell_6t
Xbit_r3_c180 bl_180 br_180 wl_3 vdd gnd cell_6t
Xbit_r4_c180 bl_180 br_180 wl_4 vdd gnd cell_6t
Xbit_r5_c180 bl_180 br_180 wl_5 vdd gnd cell_6t
Xbit_r6_c180 bl_180 br_180 wl_6 vdd gnd cell_6t
Xbit_r7_c180 bl_180 br_180 wl_7 vdd gnd cell_6t
Xbit_r8_c180 bl_180 br_180 wl_8 vdd gnd cell_6t
Xbit_r9_c180 bl_180 br_180 wl_9 vdd gnd cell_6t
Xbit_r10_c180 bl_180 br_180 wl_10 vdd gnd cell_6t
Xbit_r11_c180 bl_180 br_180 wl_11 vdd gnd cell_6t
Xbit_r12_c180 bl_180 br_180 wl_12 vdd gnd cell_6t
Xbit_r13_c180 bl_180 br_180 wl_13 vdd gnd cell_6t
Xbit_r14_c180 bl_180 br_180 wl_14 vdd gnd cell_6t
Xbit_r15_c180 bl_180 br_180 wl_15 vdd gnd cell_6t
Xbit_r16_c180 bl_180 br_180 wl_16 vdd gnd cell_6t
Xbit_r17_c180 bl_180 br_180 wl_17 vdd gnd cell_6t
Xbit_r18_c180 bl_180 br_180 wl_18 vdd gnd cell_6t
Xbit_r19_c180 bl_180 br_180 wl_19 vdd gnd cell_6t
Xbit_r20_c180 bl_180 br_180 wl_20 vdd gnd cell_6t
Xbit_r21_c180 bl_180 br_180 wl_21 vdd gnd cell_6t
Xbit_r22_c180 bl_180 br_180 wl_22 vdd gnd cell_6t
Xbit_r23_c180 bl_180 br_180 wl_23 vdd gnd cell_6t
Xbit_r24_c180 bl_180 br_180 wl_24 vdd gnd cell_6t
Xbit_r25_c180 bl_180 br_180 wl_25 vdd gnd cell_6t
Xbit_r26_c180 bl_180 br_180 wl_26 vdd gnd cell_6t
Xbit_r27_c180 bl_180 br_180 wl_27 vdd gnd cell_6t
Xbit_r28_c180 bl_180 br_180 wl_28 vdd gnd cell_6t
Xbit_r29_c180 bl_180 br_180 wl_29 vdd gnd cell_6t
Xbit_r30_c180 bl_180 br_180 wl_30 vdd gnd cell_6t
Xbit_r31_c180 bl_180 br_180 wl_31 vdd gnd cell_6t
Xbit_r32_c180 bl_180 br_180 wl_32 vdd gnd cell_6t
Xbit_r33_c180 bl_180 br_180 wl_33 vdd gnd cell_6t
Xbit_r34_c180 bl_180 br_180 wl_34 vdd gnd cell_6t
Xbit_r35_c180 bl_180 br_180 wl_35 vdd gnd cell_6t
Xbit_r36_c180 bl_180 br_180 wl_36 vdd gnd cell_6t
Xbit_r37_c180 bl_180 br_180 wl_37 vdd gnd cell_6t
Xbit_r38_c180 bl_180 br_180 wl_38 vdd gnd cell_6t
Xbit_r39_c180 bl_180 br_180 wl_39 vdd gnd cell_6t
Xbit_r40_c180 bl_180 br_180 wl_40 vdd gnd cell_6t
Xbit_r41_c180 bl_180 br_180 wl_41 vdd gnd cell_6t
Xbit_r42_c180 bl_180 br_180 wl_42 vdd gnd cell_6t
Xbit_r43_c180 bl_180 br_180 wl_43 vdd gnd cell_6t
Xbit_r44_c180 bl_180 br_180 wl_44 vdd gnd cell_6t
Xbit_r45_c180 bl_180 br_180 wl_45 vdd gnd cell_6t
Xbit_r46_c180 bl_180 br_180 wl_46 vdd gnd cell_6t
Xbit_r47_c180 bl_180 br_180 wl_47 vdd gnd cell_6t
Xbit_r48_c180 bl_180 br_180 wl_48 vdd gnd cell_6t
Xbit_r49_c180 bl_180 br_180 wl_49 vdd gnd cell_6t
Xbit_r50_c180 bl_180 br_180 wl_50 vdd gnd cell_6t
Xbit_r51_c180 bl_180 br_180 wl_51 vdd gnd cell_6t
Xbit_r52_c180 bl_180 br_180 wl_52 vdd gnd cell_6t
Xbit_r53_c180 bl_180 br_180 wl_53 vdd gnd cell_6t
Xbit_r54_c180 bl_180 br_180 wl_54 vdd gnd cell_6t
Xbit_r55_c180 bl_180 br_180 wl_55 vdd gnd cell_6t
Xbit_r56_c180 bl_180 br_180 wl_56 vdd gnd cell_6t
Xbit_r57_c180 bl_180 br_180 wl_57 vdd gnd cell_6t
Xbit_r58_c180 bl_180 br_180 wl_58 vdd gnd cell_6t
Xbit_r59_c180 bl_180 br_180 wl_59 vdd gnd cell_6t
Xbit_r60_c180 bl_180 br_180 wl_60 vdd gnd cell_6t
Xbit_r61_c180 bl_180 br_180 wl_61 vdd gnd cell_6t
Xbit_r62_c180 bl_180 br_180 wl_62 vdd gnd cell_6t
Xbit_r63_c180 bl_180 br_180 wl_63 vdd gnd cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd cell_6t
Xbit_r1_c181 bl_181 br_181 wl_1 vdd gnd cell_6t
Xbit_r2_c181 bl_181 br_181 wl_2 vdd gnd cell_6t
Xbit_r3_c181 bl_181 br_181 wl_3 vdd gnd cell_6t
Xbit_r4_c181 bl_181 br_181 wl_4 vdd gnd cell_6t
Xbit_r5_c181 bl_181 br_181 wl_5 vdd gnd cell_6t
Xbit_r6_c181 bl_181 br_181 wl_6 vdd gnd cell_6t
Xbit_r7_c181 bl_181 br_181 wl_7 vdd gnd cell_6t
Xbit_r8_c181 bl_181 br_181 wl_8 vdd gnd cell_6t
Xbit_r9_c181 bl_181 br_181 wl_9 vdd gnd cell_6t
Xbit_r10_c181 bl_181 br_181 wl_10 vdd gnd cell_6t
Xbit_r11_c181 bl_181 br_181 wl_11 vdd gnd cell_6t
Xbit_r12_c181 bl_181 br_181 wl_12 vdd gnd cell_6t
Xbit_r13_c181 bl_181 br_181 wl_13 vdd gnd cell_6t
Xbit_r14_c181 bl_181 br_181 wl_14 vdd gnd cell_6t
Xbit_r15_c181 bl_181 br_181 wl_15 vdd gnd cell_6t
Xbit_r16_c181 bl_181 br_181 wl_16 vdd gnd cell_6t
Xbit_r17_c181 bl_181 br_181 wl_17 vdd gnd cell_6t
Xbit_r18_c181 bl_181 br_181 wl_18 vdd gnd cell_6t
Xbit_r19_c181 bl_181 br_181 wl_19 vdd gnd cell_6t
Xbit_r20_c181 bl_181 br_181 wl_20 vdd gnd cell_6t
Xbit_r21_c181 bl_181 br_181 wl_21 vdd gnd cell_6t
Xbit_r22_c181 bl_181 br_181 wl_22 vdd gnd cell_6t
Xbit_r23_c181 bl_181 br_181 wl_23 vdd gnd cell_6t
Xbit_r24_c181 bl_181 br_181 wl_24 vdd gnd cell_6t
Xbit_r25_c181 bl_181 br_181 wl_25 vdd gnd cell_6t
Xbit_r26_c181 bl_181 br_181 wl_26 vdd gnd cell_6t
Xbit_r27_c181 bl_181 br_181 wl_27 vdd gnd cell_6t
Xbit_r28_c181 bl_181 br_181 wl_28 vdd gnd cell_6t
Xbit_r29_c181 bl_181 br_181 wl_29 vdd gnd cell_6t
Xbit_r30_c181 bl_181 br_181 wl_30 vdd gnd cell_6t
Xbit_r31_c181 bl_181 br_181 wl_31 vdd gnd cell_6t
Xbit_r32_c181 bl_181 br_181 wl_32 vdd gnd cell_6t
Xbit_r33_c181 bl_181 br_181 wl_33 vdd gnd cell_6t
Xbit_r34_c181 bl_181 br_181 wl_34 vdd gnd cell_6t
Xbit_r35_c181 bl_181 br_181 wl_35 vdd gnd cell_6t
Xbit_r36_c181 bl_181 br_181 wl_36 vdd gnd cell_6t
Xbit_r37_c181 bl_181 br_181 wl_37 vdd gnd cell_6t
Xbit_r38_c181 bl_181 br_181 wl_38 vdd gnd cell_6t
Xbit_r39_c181 bl_181 br_181 wl_39 vdd gnd cell_6t
Xbit_r40_c181 bl_181 br_181 wl_40 vdd gnd cell_6t
Xbit_r41_c181 bl_181 br_181 wl_41 vdd gnd cell_6t
Xbit_r42_c181 bl_181 br_181 wl_42 vdd gnd cell_6t
Xbit_r43_c181 bl_181 br_181 wl_43 vdd gnd cell_6t
Xbit_r44_c181 bl_181 br_181 wl_44 vdd gnd cell_6t
Xbit_r45_c181 bl_181 br_181 wl_45 vdd gnd cell_6t
Xbit_r46_c181 bl_181 br_181 wl_46 vdd gnd cell_6t
Xbit_r47_c181 bl_181 br_181 wl_47 vdd gnd cell_6t
Xbit_r48_c181 bl_181 br_181 wl_48 vdd gnd cell_6t
Xbit_r49_c181 bl_181 br_181 wl_49 vdd gnd cell_6t
Xbit_r50_c181 bl_181 br_181 wl_50 vdd gnd cell_6t
Xbit_r51_c181 bl_181 br_181 wl_51 vdd gnd cell_6t
Xbit_r52_c181 bl_181 br_181 wl_52 vdd gnd cell_6t
Xbit_r53_c181 bl_181 br_181 wl_53 vdd gnd cell_6t
Xbit_r54_c181 bl_181 br_181 wl_54 vdd gnd cell_6t
Xbit_r55_c181 bl_181 br_181 wl_55 vdd gnd cell_6t
Xbit_r56_c181 bl_181 br_181 wl_56 vdd gnd cell_6t
Xbit_r57_c181 bl_181 br_181 wl_57 vdd gnd cell_6t
Xbit_r58_c181 bl_181 br_181 wl_58 vdd gnd cell_6t
Xbit_r59_c181 bl_181 br_181 wl_59 vdd gnd cell_6t
Xbit_r60_c181 bl_181 br_181 wl_60 vdd gnd cell_6t
Xbit_r61_c181 bl_181 br_181 wl_61 vdd gnd cell_6t
Xbit_r62_c181 bl_181 br_181 wl_62 vdd gnd cell_6t
Xbit_r63_c181 bl_181 br_181 wl_63 vdd gnd cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd cell_6t
Xbit_r1_c182 bl_182 br_182 wl_1 vdd gnd cell_6t
Xbit_r2_c182 bl_182 br_182 wl_2 vdd gnd cell_6t
Xbit_r3_c182 bl_182 br_182 wl_3 vdd gnd cell_6t
Xbit_r4_c182 bl_182 br_182 wl_4 vdd gnd cell_6t
Xbit_r5_c182 bl_182 br_182 wl_5 vdd gnd cell_6t
Xbit_r6_c182 bl_182 br_182 wl_6 vdd gnd cell_6t
Xbit_r7_c182 bl_182 br_182 wl_7 vdd gnd cell_6t
Xbit_r8_c182 bl_182 br_182 wl_8 vdd gnd cell_6t
Xbit_r9_c182 bl_182 br_182 wl_9 vdd gnd cell_6t
Xbit_r10_c182 bl_182 br_182 wl_10 vdd gnd cell_6t
Xbit_r11_c182 bl_182 br_182 wl_11 vdd gnd cell_6t
Xbit_r12_c182 bl_182 br_182 wl_12 vdd gnd cell_6t
Xbit_r13_c182 bl_182 br_182 wl_13 vdd gnd cell_6t
Xbit_r14_c182 bl_182 br_182 wl_14 vdd gnd cell_6t
Xbit_r15_c182 bl_182 br_182 wl_15 vdd gnd cell_6t
Xbit_r16_c182 bl_182 br_182 wl_16 vdd gnd cell_6t
Xbit_r17_c182 bl_182 br_182 wl_17 vdd gnd cell_6t
Xbit_r18_c182 bl_182 br_182 wl_18 vdd gnd cell_6t
Xbit_r19_c182 bl_182 br_182 wl_19 vdd gnd cell_6t
Xbit_r20_c182 bl_182 br_182 wl_20 vdd gnd cell_6t
Xbit_r21_c182 bl_182 br_182 wl_21 vdd gnd cell_6t
Xbit_r22_c182 bl_182 br_182 wl_22 vdd gnd cell_6t
Xbit_r23_c182 bl_182 br_182 wl_23 vdd gnd cell_6t
Xbit_r24_c182 bl_182 br_182 wl_24 vdd gnd cell_6t
Xbit_r25_c182 bl_182 br_182 wl_25 vdd gnd cell_6t
Xbit_r26_c182 bl_182 br_182 wl_26 vdd gnd cell_6t
Xbit_r27_c182 bl_182 br_182 wl_27 vdd gnd cell_6t
Xbit_r28_c182 bl_182 br_182 wl_28 vdd gnd cell_6t
Xbit_r29_c182 bl_182 br_182 wl_29 vdd gnd cell_6t
Xbit_r30_c182 bl_182 br_182 wl_30 vdd gnd cell_6t
Xbit_r31_c182 bl_182 br_182 wl_31 vdd gnd cell_6t
Xbit_r32_c182 bl_182 br_182 wl_32 vdd gnd cell_6t
Xbit_r33_c182 bl_182 br_182 wl_33 vdd gnd cell_6t
Xbit_r34_c182 bl_182 br_182 wl_34 vdd gnd cell_6t
Xbit_r35_c182 bl_182 br_182 wl_35 vdd gnd cell_6t
Xbit_r36_c182 bl_182 br_182 wl_36 vdd gnd cell_6t
Xbit_r37_c182 bl_182 br_182 wl_37 vdd gnd cell_6t
Xbit_r38_c182 bl_182 br_182 wl_38 vdd gnd cell_6t
Xbit_r39_c182 bl_182 br_182 wl_39 vdd gnd cell_6t
Xbit_r40_c182 bl_182 br_182 wl_40 vdd gnd cell_6t
Xbit_r41_c182 bl_182 br_182 wl_41 vdd gnd cell_6t
Xbit_r42_c182 bl_182 br_182 wl_42 vdd gnd cell_6t
Xbit_r43_c182 bl_182 br_182 wl_43 vdd gnd cell_6t
Xbit_r44_c182 bl_182 br_182 wl_44 vdd gnd cell_6t
Xbit_r45_c182 bl_182 br_182 wl_45 vdd gnd cell_6t
Xbit_r46_c182 bl_182 br_182 wl_46 vdd gnd cell_6t
Xbit_r47_c182 bl_182 br_182 wl_47 vdd gnd cell_6t
Xbit_r48_c182 bl_182 br_182 wl_48 vdd gnd cell_6t
Xbit_r49_c182 bl_182 br_182 wl_49 vdd gnd cell_6t
Xbit_r50_c182 bl_182 br_182 wl_50 vdd gnd cell_6t
Xbit_r51_c182 bl_182 br_182 wl_51 vdd gnd cell_6t
Xbit_r52_c182 bl_182 br_182 wl_52 vdd gnd cell_6t
Xbit_r53_c182 bl_182 br_182 wl_53 vdd gnd cell_6t
Xbit_r54_c182 bl_182 br_182 wl_54 vdd gnd cell_6t
Xbit_r55_c182 bl_182 br_182 wl_55 vdd gnd cell_6t
Xbit_r56_c182 bl_182 br_182 wl_56 vdd gnd cell_6t
Xbit_r57_c182 bl_182 br_182 wl_57 vdd gnd cell_6t
Xbit_r58_c182 bl_182 br_182 wl_58 vdd gnd cell_6t
Xbit_r59_c182 bl_182 br_182 wl_59 vdd gnd cell_6t
Xbit_r60_c182 bl_182 br_182 wl_60 vdd gnd cell_6t
Xbit_r61_c182 bl_182 br_182 wl_61 vdd gnd cell_6t
Xbit_r62_c182 bl_182 br_182 wl_62 vdd gnd cell_6t
Xbit_r63_c182 bl_182 br_182 wl_63 vdd gnd cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd cell_6t
Xbit_r1_c183 bl_183 br_183 wl_1 vdd gnd cell_6t
Xbit_r2_c183 bl_183 br_183 wl_2 vdd gnd cell_6t
Xbit_r3_c183 bl_183 br_183 wl_3 vdd gnd cell_6t
Xbit_r4_c183 bl_183 br_183 wl_4 vdd gnd cell_6t
Xbit_r5_c183 bl_183 br_183 wl_5 vdd gnd cell_6t
Xbit_r6_c183 bl_183 br_183 wl_6 vdd gnd cell_6t
Xbit_r7_c183 bl_183 br_183 wl_7 vdd gnd cell_6t
Xbit_r8_c183 bl_183 br_183 wl_8 vdd gnd cell_6t
Xbit_r9_c183 bl_183 br_183 wl_9 vdd gnd cell_6t
Xbit_r10_c183 bl_183 br_183 wl_10 vdd gnd cell_6t
Xbit_r11_c183 bl_183 br_183 wl_11 vdd gnd cell_6t
Xbit_r12_c183 bl_183 br_183 wl_12 vdd gnd cell_6t
Xbit_r13_c183 bl_183 br_183 wl_13 vdd gnd cell_6t
Xbit_r14_c183 bl_183 br_183 wl_14 vdd gnd cell_6t
Xbit_r15_c183 bl_183 br_183 wl_15 vdd gnd cell_6t
Xbit_r16_c183 bl_183 br_183 wl_16 vdd gnd cell_6t
Xbit_r17_c183 bl_183 br_183 wl_17 vdd gnd cell_6t
Xbit_r18_c183 bl_183 br_183 wl_18 vdd gnd cell_6t
Xbit_r19_c183 bl_183 br_183 wl_19 vdd gnd cell_6t
Xbit_r20_c183 bl_183 br_183 wl_20 vdd gnd cell_6t
Xbit_r21_c183 bl_183 br_183 wl_21 vdd gnd cell_6t
Xbit_r22_c183 bl_183 br_183 wl_22 vdd gnd cell_6t
Xbit_r23_c183 bl_183 br_183 wl_23 vdd gnd cell_6t
Xbit_r24_c183 bl_183 br_183 wl_24 vdd gnd cell_6t
Xbit_r25_c183 bl_183 br_183 wl_25 vdd gnd cell_6t
Xbit_r26_c183 bl_183 br_183 wl_26 vdd gnd cell_6t
Xbit_r27_c183 bl_183 br_183 wl_27 vdd gnd cell_6t
Xbit_r28_c183 bl_183 br_183 wl_28 vdd gnd cell_6t
Xbit_r29_c183 bl_183 br_183 wl_29 vdd gnd cell_6t
Xbit_r30_c183 bl_183 br_183 wl_30 vdd gnd cell_6t
Xbit_r31_c183 bl_183 br_183 wl_31 vdd gnd cell_6t
Xbit_r32_c183 bl_183 br_183 wl_32 vdd gnd cell_6t
Xbit_r33_c183 bl_183 br_183 wl_33 vdd gnd cell_6t
Xbit_r34_c183 bl_183 br_183 wl_34 vdd gnd cell_6t
Xbit_r35_c183 bl_183 br_183 wl_35 vdd gnd cell_6t
Xbit_r36_c183 bl_183 br_183 wl_36 vdd gnd cell_6t
Xbit_r37_c183 bl_183 br_183 wl_37 vdd gnd cell_6t
Xbit_r38_c183 bl_183 br_183 wl_38 vdd gnd cell_6t
Xbit_r39_c183 bl_183 br_183 wl_39 vdd gnd cell_6t
Xbit_r40_c183 bl_183 br_183 wl_40 vdd gnd cell_6t
Xbit_r41_c183 bl_183 br_183 wl_41 vdd gnd cell_6t
Xbit_r42_c183 bl_183 br_183 wl_42 vdd gnd cell_6t
Xbit_r43_c183 bl_183 br_183 wl_43 vdd gnd cell_6t
Xbit_r44_c183 bl_183 br_183 wl_44 vdd gnd cell_6t
Xbit_r45_c183 bl_183 br_183 wl_45 vdd gnd cell_6t
Xbit_r46_c183 bl_183 br_183 wl_46 vdd gnd cell_6t
Xbit_r47_c183 bl_183 br_183 wl_47 vdd gnd cell_6t
Xbit_r48_c183 bl_183 br_183 wl_48 vdd gnd cell_6t
Xbit_r49_c183 bl_183 br_183 wl_49 vdd gnd cell_6t
Xbit_r50_c183 bl_183 br_183 wl_50 vdd gnd cell_6t
Xbit_r51_c183 bl_183 br_183 wl_51 vdd gnd cell_6t
Xbit_r52_c183 bl_183 br_183 wl_52 vdd gnd cell_6t
Xbit_r53_c183 bl_183 br_183 wl_53 vdd gnd cell_6t
Xbit_r54_c183 bl_183 br_183 wl_54 vdd gnd cell_6t
Xbit_r55_c183 bl_183 br_183 wl_55 vdd gnd cell_6t
Xbit_r56_c183 bl_183 br_183 wl_56 vdd gnd cell_6t
Xbit_r57_c183 bl_183 br_183 wl_57 vdd gnd cell_6t
Xbit_r58_c183 bl_183 br_183 wl_58 vdd gnd cell_6t
Xbit_r59_c183 bl_183 br_183 wl_59 vdd gnd cell_6t
Xbit_r60_c183 bl_183 br_183 wl_60 vdd gnd cell_6t
Xbit_r61_c183 bl_183 br_183 wl_61 vdd gnd cell_6t
Xbit_r62_c183 bl_183 br_183 wl_62 vdd gnd cell_6t
Xbit_r63_c183 bl_183 br_183 wl_63 vdd gnd cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd cell_6t
Xbit_r1_c184 bl_184 br_184 wl_1 vdd gnd cell_6t
Xbit_r2_c184 bl_184 br_184 wl_2 vdd gnd cell_6t
Xbit_r3_c184 bl_184 br_184 wl_3 vdd gnd cell_6t
Xbit_r4_c184 bl_184 br_184 wl_4 vdd gnd cell_6t
Xbit_r5_c184 bl_184 br_184 wl_5 vdd gnd cell_6t
Xbit_r6_c184 bl_184 br_184 wl_6 vdd gnd cell_6t
Xbit_r7_c184 bl_184 br_184 wl_7 vdd gnd cell_6t
Xbit_r8_c184 bl_184 br_184 wl_8 vdd gnd cell_6t
Xbit_r9_c184 bl_184 br_184 wl_9 vdd gnd cell_6t
Xbit_r10_c184 bl_184 br_184 wl_10 vdd gnd cell_6t
Xbit_r11_c184 bl_184 br_184 wl_11 vdd gnd cell_6t
Xbit_r12_c184 bl_184 br_184 wl_12 vdd gnd cell_6t
Xbit_r13_c184 bl_184 br_184 wl_13 vdd gnd cell_6t
Xbit_r14_c184 bl_184 br_184 wl_14 vdd gnd cell_6t
Xbit_r15_c184 bl_184 br_184 wl_15 vdd gnd cell_6t
Xbit_r16_c184 bl_184 br_184 wl_16 vdd gnd cell_6t
Xbit_r17_c184 bl_184 br_184 wl_17 vdd gnd cell_6t
Xbit_r18_c184 bl_184 br_184 wl_18 vdd gnd cell_6t
Xbit_r19_c184 bl_184 br_184 wl_19 vdd gnd cell_6t
Xbit_r20_c184 bl_184 br_184 wl_20 vdd gnd cell_6t
Xbit_r21_c184 bl_184 br_184 wl_21 vdd gnd cell_6t
Xbit_r22_c184 bl_184 br_184 wl_22 vdd gnd cell_6t
Xbit_r23_c184 bl_184 br_184 wl_23 vdd gnd cell_6t
Xbit_r24_c184 bl_184 br_184 wl_24 vdd gnd cell_6t
Xbit_r25_c184 bl_184 br_184 wl_25 vdd gnd cell_6t
Xbit_r26_c184 bl_184 br_184 wl_26 vdd gnd cell_6t
Xbit_r27_c184 bl_184 br_184 wl_27 vdd gnd cell_6t
Xbit_r28_c184 bl_184 br_184 wl_28 vdd gnd cell_6t
Xbit_r29_c184 bl_184 br_184 wl_29 vdd gnd cell_6t
Xbit_r30_c184 bl_184 br_184 wl_30 vdd gnd cell_6t
Xbit_r31_c184 bl_184 br_184 wl_31 vdd gnd cell_6t
Xbit_r32_c184 bl_184 br_184 wl_32 vdd gnd cell_6t
Xbit_r33_c184 bl_184 br_184 wl_33 vdd gnd cell_6t
Xbit_r34_c184 bl_184 br_184 wl_34 vdd gnd cell_6t
Xbit_r35_c184 bl_184 br_184 wl_35 vdd gnd cell_6t
Xbit_r36_c184 bl_184 br_184 wl_36 vdd gnd cell_6t
Xbit_r37_c184 bl_184 br_184 wl_37 vdd gnd cell_6t
Xbit_r38_c184 bl_184 br_184 wl_38 vdd gnd cell_6t
Xbit_r39_c184 bl_184 br_184 wl_39 vdd gnd cell_6t
Xbit_r40_c184 bl_184 br_184 wl_40 vdd gnd cell_6t
Xbit_r41_c184 bl_184 br_184 wl_41 vdd gnd cell_6t
Xbit_r42_c184 bl_184 br_184 wl_42 vdd gnd cell_6t
Xbit_r43_c184 bl_184 br_184 wl_43 vdd gnd cell_6t
Xbit_r44_c184 bl_184 br_184 wl_44 vdd gnd cell_6t
Xbit_r45_c184 bl_184 br_184 wl_45 vdd gnd cell_6t
Xbit_r46_c184 bl_184 br_184 wl_46 vdd gnd cell_6t
Xbit_r47_c184 bl_184 br_184 wl_47 vdd gnd cell_6t
Xbit_r48_c184 bl_184 br_184 wl_48 vdd gnd cell_6t
Xbit_r49_c184 bl_184 br_184 wl_49 vdd gnd cell_6t
Xbit_r50_c184 bl_184 br_184 wl_50 vdd gnd cell_6t
Xbit_r51_c184 bl_184 br_184 wl_51 vdd gnd cell_6t
Xbit_r52_c184 bl_184 br_184 wl_52 vdd gnd cell_6t
Xbit_r53_c184 bl_184 br_184 wl_53 vdd gnd cell_6t
Xbit_r54_c184 bl_184 br_184 wl_54 vdd gnd cell_6t
Xbit_r55_c184 bl_184 br_184 wl_55 vdd gnd cell_6t
Xbit_r56_c184 bl_184 br_184 wl_56 vdd gnd cell_6t
Xbit_r57_c184 bl_184 br_184 wl_57 vdd gnd cell_6t
Xbit_r58_c184 bl_184 br_184 wl_58 vdd gnd cell_6t
Xbit_r59_c184 bl_184 br_184 wl_59 vdd gnd cell_6t
Xbit_r60_c184 bl_184 br_184 wl_60 vdd gnd cell_6t
Xbit_r61_c184 bl_184 br_184 wl_61 vdd gnd cell_6t
Xbit_r62_c184 bl_184 br_184 wl_62 vdd gnd cell_6t
Xbit_r63_c184 bl_184 br_184 wl_63 vdd gnd cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd cell_6t
Xbit_r1_c185 bl_185 br_185 wl_1 vdd gnd cell_6t
Xbit_r2_c185 bl_185 br_185 wl_2 vdd gnd cell_6t
Xbit_r3_c185 bl_185 br_185 wl_3 vdd gnd cell_6t
Xbit_r4_c185 bl_185 br_185 wl_4 vdd gnd cell_6t
Xbit_r5_c185 bl_185 br_185 wl_5 vdd gnd cell_6t
Xbit_r6_c185 bl_185 br_185 wl_6 vdd gnd cell_6t
Xbit_r7_c185 bl_185 br_185 wl_7 vdd gnd cell_6t
Xbit_r8_c185 bl_185 br_185 wl_8 vdd gnd cell_6t
Xbit_r9_c185 bl_185 br_185 wl_9 vdd gnd cell_6t
Xbit_r10_c185 bl_185 br_185 wl_10 vdd gnd cell_6t
Xbit_r11_c185 bl_185 br_185 wl_11 vdd gnd cell_6t
Xbit_r12_c185 bl_185 br_185 wl_12 vdd gnd cell_6t
Xbit_r13_c185 bl_185 br_185 wl_13 vdd gnd cell_6t
Xbit_r14_c185 bl_185 br_185 wl_14 vdd gnd cell_6t
Xbit_r15_c185 bl_185 br_185 wl_15 vdd gnd cell_6t
Xbit_r16_c185 bl_185 br_185 wl_16 vdd gnd cell_6t
Xbit_r17_c185 bl_185 br_185 wl_17 vdd gnd cell_6t
Xbit_r18_c185 bl_185 br_185 wl_18 vdd gnd cell_6t
Xbit_r19_c185 bl_185 br_185 wl_19 vdd gnd cell_6t
Xbit_r20_c185 bl_185 br_185 wl_20 vdd gnd cell_6t
Xbit_r21_c185 bl_185 br_185 wl_21 vdd gnd cell_6t
Xbit_r22_c185 bl_185 br_185 wl_22 vdd gnd cell_6t
Xbit_r23_c185 bl_185 br_185 wl_23 vdd gnd cell_6t
Xbit_r24_c185 bl_185 br_185 wl_24 vdd gnd cell_6t
Xbit_r25_c185 bl_185 br_185 wl_25 vdd gnd cell_6t
Xbit_r26_c185 bl_185 br_185 wl_26 vdd gnd cell_6t
Xbit_r27_c185 bl_185 br_185 wl_27 vdd gnd cell_6t
Xbit_r28_c185 bl_185 br_185 wl_28 vdd gnd cell_6t
Xbit_r29_c185 bl_185 br_185 wl_29 vdd gnd cell_6t
Xbit_r30_c185 bl_185 br_185 wl_30 vdd gnd cell_6t
Xbit_r31_c185 bl_185 br_185 wl_31 vdd gnd cell_6t
Xbit_r32_c185 bl_185 br_185 wl_32 vdd gnd cell_6t
Xbit_r33_c185 bl_185 br_185 wl_33 vdd gnd cell_6t
Xbit_r34_c185 bl_185 br_185 wl_34 vdd gnd cell_6t
Xbit_r35_c185 bl_185 br_185 wl_35 vdd gnd cell_6t
Xbit_r36_c185 bl_185 br_185 wl_36 vdd gnd cell_6t
Xbit_r37_c185 bl_185 br_185 wl_37 vdd gnd cell_6t
Xbit_r38_c185 bl_185 br_185 wl_38 vdd gnd cell_6t
Xbit_r39_c185 bl_185 br_185 wl_39 vdd gnd cell_6t
Xbit_r40_c185 bl_185 br_185 wl_40 vdd gnd cell_6t
Xbit_r41_c185 bl_185 br_185 wl_41 vdd gnd cell_6t
Xbit_r42_c185 bl_185 br_185 wl_42 vdd gnd cell_6t
Xbit_r43_c185 bl_185 br_185 wl_43 vdd gnd cell_6t
Xbit_r44_c185 bl_185 br_185 wl_44 vdd gnd cell_6t
Xbit_r45_c185 bl_185 br_185 wl_45 vdd gnd cell_6t
Xbit_r46_c185 bl_185 br_185 wl_46 vdd gnd cell_6t
Xbit_r47_c185 bl_185 br_185 wl_47 vdd gnd cell_6t
Xbit_r48_c185 bl_185 br_185 wl_48 vdd gnd cell_6t
Xbit_r49_c185 bl_185 br_185 wl_49 vdd gnd cell_6t
Xbit_r50_c185 bl_185 br_185 wl_50 vdd gnd cell_6t
Xbit_r51_c185 bl_185 br_185 wl_51 vdd gnd cell_6t
Xbit_r52_c185 bl_185 br_185 wl_52 vdd gnd cell_6t
Xbit_r53_c185 bl_185 br_185 wl_53 vdd gnd cell_6t
Xbit_r54_c185 bl_185 br_185 wl_54 vdd gnd cell_6t
Xbit_r55_c185 bl_185 br_185 wl_55 vdd gnd cell_6t
Xbit_r56_c185 bl_185 br_185 wl_56 vdd gnd cell_6t
Xbit_r57_c185 bl_185 br_185 wl_57 vdd gnd cell_6t
Xbit_r58_c185 bl_185 br_185 wl_58 vdd gnd cell_6t
Xbit_r59_c185 bl_185 br_185 wl_59 vdd gnd cell_6t
Xbit_r60_c185 bl_185 br_185 wl_60 vdd gnd cell_6t
Xbit_r61_c185 bl_185 br_185 wl_61 vdd gnd cell_6t
Xbit_r62_c185 bl_185 br_185 wl_62 vdd gnd cell_6t
Xbit_r63_c185 bl_185 br_185 wl_63 vdd gnd cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd cell_6t
Xbit_r1_c186 bl_186 br_186 wl_1 vdd gnd cell_6t
Xbit_r2_c186 bl_186 br_186 wl_2 vdd gnd cell_6t
Xbit_r3_c186 bl_186 br_186 wl_3 vdd gnd cell_6t
Xbit_r4_c186 bl_186 br_186 wl_4 vdd gnd cell_6t
Xbit_r5_c186 bl_186 br_186 wl_5 vdd gnd cell_6t
Xbit_r6_c186 bl_186 br_186 wl_6 vdd gnd cell_6t
Xbit_r7_c186 bl_186 br_186 wl_7 vdd gnd cell_6t
Xbit_r8_c186 bl_186 br_186 wl_8 vdd gnd cell_6t
Xbit_r9_c186 bl_186 br_186 wl_9 vdd gnd cell_6t
Xbit_r10_c186 bl_186 br_186 wl_10 vdd gnd cell_6t
Xbit_r11_c186 bl_186 br_186 wl_11 vdd gnd cell_6t
Xbit_r12_c186 bl_186 br_186 wl_12 vdd gnd cell_6t
Xbit_r13_c186 bl_186 br_186 wl_13 vdd gnd cell_6t
Xbit_r14_c186 bl_186 br_186 wl_14 vdd gnd cell_6t
Xbit_r15_c186 bl_186 br_186 wl_15 vdd gnd cell_6t
Xbit_r16_c186 bl_186 br_186 wl_16 vdd gnd cell_6t
Xbit_r17_c186 bl_186 br_186 wl_17 vdd gnd cell_6t
Xbit_r18_c186 bl_186 br_186 wl_18 vdd gnd cell_6t
Xbit_r19_c186 bl_186 br_186 wl_19 vdd gnd cell_6t
Xbit_r20_c186 bl_186 br_186 wl_20 vdd gnd cell_6t
Xbit_r21_c186 bl_186 br_186 wl_21 vdd gnd cell_6t
Xbit_r22_c186 bl_186 br_186 wl_22 vdd gnd cell_6t
Xbit_r23_c186 bl_186 br_186 wl_23 vdd gnd cell_6t
Xbit_r24_c186 bl_186 br_186 wl_24 vdd gnd cell_6t
Xbit_r25_c186 bl_186 br_186 wl_25 vdd gnd cell_6t
Xbit_r26_c186 bl_186 br_186 wl_26 vdd gnd cell_6t
Xbit_r27_c186 bl_186 br_186 wl_27 vdd gnd cell_6t
Xbit_r28_c186 bl_186 br_186 wl_28 vdd gnd cell_6t
Xbit_r29_c186 bl_186 br_186 wl_29 vdd gnd cell_6t
Xbit_r30_c186 bl_186 br_186 wl_30 vdd gnd cell_6t
Xbit_r31_c186 bl_186 br_186 wl_31 vdd gnd cell_6t
Xbit_r32_c186 bl_186 br_186 wl_32 vdd gnd cell_6t
Xbit_r33_c186 bl_186 br_186 wl_33 vdd gnd cell_6t
Xbit_r34_c186 bl_186 br_186 wl_34 vdd gnd cell_6t
Xbit_r35_c186 bl_186 br_186 wl_35 vdd gnd cell_6t
Xbit_r36_c186 bl_186 br_186 wl_36 vdd gnd cell_6t
Xbit_r37_c186 bl_186 br_186 wl_37 vdd gnd cell_6t
Xbit_r38_c186 bl_186 br_186 wl_38 vdd gnd cell_6t
Xbit_r39_c186 bl_186 br_186 wl_39 vdd gnd cell_6t
Xbit_r40_c186 bl_186 br_186 wl_40 vdd gnd cell_6t
Xbit_r41_c186 bl_186 br_186 wl_41 vdd gnd cell_6t
Xbit_r42_c186 bl_186 br_186 wl_42 vdd gnd cell_6t
Xbit_r43_c186 bl_186 br_186 wl_43 vdd gnd cell_6t
Xbit_r44_c186 bl_186 br_186 wl_44 vdd gnd cell_6t
Xbit_r45_c186 bl_186 br_186 wl_45 vdd gnd cell_6t
Xbit_r46_c186 bl_186 br_186 wl_46 vdd gnd cell_6t
Xbit_r47_c186 bl_186 br_186 wl_47 vdd gnd cell_6t
Xbit_r48_c186 bl_186 br_186 wl_48 vdd gnd cell_6t
Xbit_r49_c186 bl_186 br_186 wl_49 vdd gnd cell_6t
Xbit_r50_c186 bl_186 br_186 wl_50 vdd gnd cell_6t
Xbit_r51_c186 bl_186 br_186 wl_51 vdd gnd cell_6t
Xbit_r52_c186 bl_186 br_186 wl_52 vdd gnd cell_6t
Xbit_r53_c186 bl_186 br_186 wl_53 vdd gnd cell_6t
Xbit_r54_c186 bl_186 br_186 wl_54 vdd gnd cell_6t
Xbit_r55_c186 bl_186 br_186 wl_55 vdd gnd cell_6t
Xbit_r56_c186 bl_186 br_186 wl_56 vdd gnd cell_6t
Xbit_r57_c186 bl_186 br_186 wl_57 vdd gnd cell_6t
Xbit_r58_c186 bl_186 br_186 wl_58 vdd gnd cell_6t
Xbit_r59_c186 bl_186 br_186 wl_59 vdd gnd cell_6t
Xbit_r60_c186 bl_186 br_186 wl_60 vdd gnd cell_6t
Xbit_r61_c186 bl_186 br_186 wl_61 vdd gnd cell_6t
Xbit_r62_c186 bl_186 br_186 wl_62 vdd gnd cell_6t
Xbit_r63_c186 bl_186 br_186 wl_63 vdd gnd cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd cell_6t
Xbit_r1_c187 bl_187 br_187 wl_1 vdd gnd cell_6t
Xbit_r2_c187 bl_187 br_187 wl_2 vdd gnd cell_6t
Xbit_r3_c187 bl_187 br_187 wl_3 vdd gnd cell_6t
Xbit_r4_c187 bl_187 br_187 wl_4 vdd gnd cell_6t
Xbit_r5_c187 bl_187 br_187 wl_5 vdd gnd cell_6t
Xbit_r6_c187 bl_187 br_187 wl_6 vdd gnd cell_6t
Xbit_r7_c187 bl_187 br_187 wl_7 vdd gnd cell_6t
Xbit_r8_c187 bl_187 br_187 wl_8 vdd gnd cell_6t
Xbit_r9_c187 bl_187 br_187 wl_9 vdd gnd cell_6t
Xbit_r10_c187 bl_187 br_187 wl_10 vdd gnd cell_6t
Xbit_r11_c187 bl_187 br_187 wl_11 vdd gnd cell_6t
Xbit_r12_c187 bl_187 br_187 wl_12 vdd gnd cell_6t
Xbit_r13_c187 bl_187 br_187 wl_13 vdd gnd cell_6t
Xbit_r14_c187 bl_187 br_187 wl_14 vdd gnd cell_6t
Xbit_r15_c187 bl_187 br_187 wl_15 vdd gnd cell_6t
Xbit_r16_c187 bl_187 br_187 wl_16 vdd gnd cell_6t
Xbit_r17_c187 bl_187 br_187 wl_17 vdd gnd cell_6t
Xbit_r18_c187 bl_187 br_187 wl_18 vdd gnd cell_6t
Xbit_r19_c187 bl_187 br_187 wl_19 vdd gnd cell_6t
Xbit_r20_c187 bl_187 br_187 wl_20 vdd gnd cell_6t
Xbit_r21_c187 bl_187 br_187 wl_21 vdd gnd cell_6t
Xbit_r22_c187 bl_187 br_187 wl_22 vdd gnd cell_6t
Xbit_r23_c187 bl_187 br_187 wl_23 vdd gnd cell_6t
Xbit_r24_c187 bl_187 br_187 wl_24 vdd gnd cell_6t
Xbit_r25_c187 bl_187 br_187 wl_25 vdd gnd cell_6t
Xbit_r26_c187 bl_187 br_187 wl_26 vdd gnd cell_6t
Xbit_r27_c187 bl_187 br_187 wl_27 vdd gnd cell_6t
Xbit_r28_c187 bl_187 br_187 wl_28 vdd gnd cell_6t
Xbit_r29_c187 bl_187 br_187 wl_29 vdd gnd cell_6t
Xbit_r30_c187 bl_187 br_187 wl_30 vdd gnd cell_6t
Xbit_r31_c187 bl_187 br_187 wl_31 vdd gnd cell_6t
Xbit_r32_c187 bl_187 br_187 wl_32 vdd gnd cell_6t
Xbit_r33_c187 bl_187 br_187 wl_33 vdd gnd cell_6t
Xbit_r34_c187 bl_187 br_187 wl_34 vdd gnd cell_6t
Xbit_r35_c187 bl_187 br_187 wl_35 vdd gnd cell_6t
Xbit_r36_c187 bl_187 br_187 wl_36 vdd gnd cell_6t
Xbit_r37_c187 bl_187 br_187 wl_37 vdd gnd cell_6t
Xbit_r38_c187 bl_187 br_187 wl_38 vdd gnd cell_6t
Xbit_r39_c187 bl_187 br_187 wl_39 vdd gnd cell_6t
Xbit_r40_c187 bl_187 br_187 wl_40 vdd gnd cell_6t
Xbit_r41_c187 bl_187 br_187 wl_41 vdd gnd cell_6t
Xbit_r42_c187 bl_187 br_187 wl_42 vdd gnd cell_6t
Xbit_r43_c187 bl_187 br_187 wl_43 vdd gnd cell_6t
Xbit_r44_c187 bl_187 br_187 wl_44 vdd gnd cell_6t
Xbit_r45_c187 bl_187 br_187 wl_45 vdd gnd cell_6t
Xbit_r46_c187 bl_187 br_187 wl_46 vdd gnd cell_6t
Xbit_r47_c187 bl_187 br_187 wl_47 vdd gnd cell_6t
Xbit_r48_c187 bl_187 br_187 wl_48 vdd gnd cell_6t
Xbit_r49_c187 bl_187 br_187 wl_49 vdd gnd cell_6t
Xbit_r50_c187 bl_187 br_187 wl_50 vdd gnd cell_6t
Xbit_r51_c187 bl_187 br_187 wl_51 vdd gnd cell_6t
Xbit_r52_c187 bl_187 br_187 wl_52 vdd gnd cell_6t
Xbit_r53_c187 bl_187 br_187 wl_53 vdd gnd cell_6t
Xbit_r54_c187 bl_187 br_187 wl_54 vdd gnd cell_6t
Xbit_r55_c187 bl_187 br_187 wl_55 vdd gnd cell_6t
Xbit_r56_c187 bl_187 br_187 wl_56 vdd gnd cell_6t
Xbit_r57_c187 bl_187 br_187 wl_57 vdd gnd cell_6t
Xbit_r58_c187 bl_187 br_187 wl_58 vdd gnd cell_6t
Xbit_r59_c187 bl_187 br_187 wl_59 vdd gnd cell_6t
Xbit_r60_c187 bl_187 br_187 wl_60 vdd gnd cell_6t
Xbit_r61_c187 bl_187 br_187 wl_61 vdd gnd cell_6t
Xbit_r62_c187 bl_187 br_187 wl_62 vdd gnd cell_6t
Xbit_r63_c187 bl_187 br_187 wl_63 vdd gnd cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd cell_6t
Xbit_r1_c188 bl_188 br_188 wl_1 vdd gnd cell_6t
Xbit_r2_c188 bl_188 br_188 wl_2 vdd gnd cell_6t
Xbit_r3_c188 bl_188 br_188 wl_3 vdd gnd cell_6t
Xbit_r4_c188 bl_188 br_188 wl_4 vdd gnd cell_6t
Xbit_r5_c188 bl_188 br_188 wl_5 vdd gnd cell_6t
Xbit_r6_c188 bl_188 br_188 wl_6 vdd gnd cell_6t
Xbit_r7_c188 bl_188 br_188 wl_7 vdd gnd cell_6t
Xbit_r8_c188 bl_188 br_188 wl_8 vdd gnd cell_6t
Xbit_r9_c188 bl_188 br_188 wl_9 vdd gnd cell_6t
Xbit_r10_c188 bl_188 br_188 wl_10 vdd gnd cell_6t
Xbit_r11_c188 bl_188 br_188 wl_11 vdd gnd cell_6t
Xbit_r12_c188 bl_188 br_188 wl_12 vdd gnd cell_6t
Xbit_r13_c188 bl_188 br_188 wl_13 vdd gnd cell_6t
Xbit_r14_c188 bl_188 br_188 wl_14 vdd gnd cell_6t
Xbit_r15_c188 bl_188 br_188 wl_15 vdd gnd cell_6t
Xbit_r16_c188 bl_188 br_188 wl_16 vdd gnd cell_6t
Xbit_r17_c188 bl_188 br_188 wl_17 vdd gnd cell_6t
Xbit_r18_c188 bl_188 br_188 wl_18 vdd gnd cell_6t
Xbit_r19_c188 bl_188 br_188 wl_19 vdd gnd cell_6t
Xbit_r20_c188 bl_188 br_188 wl_20 vdd gnd cell_6t
Xbit_r21_c188 bl_188 br_188 wl_21 vdd gnd cell_6t
Xbit_r22_c188 bl_188 br_188 wl_22 vdd gnd cell_6t
Xbit_r23_c188 bl_188 br_188 wl_23 vdd gnd cell_6t
Xbit_r24_c188 bl_188 br_188 wl_24 vdd gnd cell_6t
Xbit_r25_c188 bl_188 br_188 wl_25 vdd gnd cell_6t
Xbit_r26_c188 bl_188 br_188 wl_26 vdd gnd cell_6t
Xbit_r27_c188 bl_188 br_188 wl_27 vdd gnd cell_6t
Xbit_r28_c188 bl_188 br_188 wl_28 vdd gnd cell_6t
Xbit_r29_c188 bl_188 br_188 wl_29 vdd gnd cell_6t
Xbit_r30_c188 bl_188 br_188 wl_30 vdd gnd cell_6t
Xbit_r31_c188 bl_188 br_188 wl_31 vdd gnd cell_6t
Xbit_r32_c188 bl_188 br_188 wl_32 vdd gnd cell_6t
Xbit_r33_c188 bl_188 br_188 wl_33 vdd gnd cell_6t
Xbit_r34_c188 bl_188 br_188 wl_34 vdd gnd cell_6t
Xbit_r35_c188 bl_188 br_188 wl_35 vdd gnd cell_6t
Xbit_r36_c188 bl_188 br_188 wl_36 vdd gnd cell_6t
Xbit_r37_c188 bl_188 br_188 wl_37 vdd gnd cell_6t
Xbit_r38_c188 bl_188 br_188 wl_38 vdd gnd cell_6t
Xbit_r39_c188 bl_188 br_188 wl_39 vdd gnd cell_6t
Xbit_r40_c188 bl_188 br_188 wl_40 vdd gnd cell_6t
Xbit_r41_c188 bl_188 br_188 wl_41 vdd gnd cell_6t
Xbit_r42_c188 bl_188 br_188 wl_42 vdd gnd cell_6t
Xbit_r43_c188 bl_188 br_188 wl_43 vdd gnd cell_6t
Xbit_r44_c188 bl_188 br_188 wl_44 vdd gnd cell_6t
Xbit_r45_c188 bl_188 br_188 wl_45 vdd gnd cell_6t
Xbit_r46_c188 bl_188 br_188 wl_46 vdd gnd cell_6t
Xbit_r47_c188 bl_188 br_188 wl_47 vdd gnd cell_6t
Xbit_r48_c188 bl_188 br_188 wl_48 vdd gnd cell_6t
Xbit_r49_c188 bl_188 br_188 wl_49 vdd gnd cell_6t
Xbit_r50_c188 bl_188 br_188 wl_50 vdd gnd cell_6t
Xbit_r51_c188 bl_188 br_188 wl_51 vdd gnd cell_6t
Xbit_r52_c188 bl_188 br_188 wl_52 vdd gnd cell_6t
Xbit_r53_c188 bl_188 br_188 wl_53 vdd gnd cell_6t
Xbit_r54_c188 bl_188 br_188 wl_54 vdd gnd cell_6t
Xbit_r55_c188 bl_188 br_188 wl_55 vdd gnd cell_6t
Xbit_r56_c188 bl_188 br_188 wl_56 vdd gnd cell_6t
Xbit_r57_c188 bl_188 br_188 wl_57 vdd gnd cell_6t
Xbit_r58_c188 bl_188 br_188 wl_58 vdd gnd cell_6t
Xbit_r59_c188 bl_188 br_188 wl_59 vdd gnd cell_6t
Xbit_r60_c188 bl_188 br_188 wl_60 vdd gnd cell_6t
Xbit_r61_c188 bl_188 br_188 wl_61 vdd gnd cell_6t
Xbit_r62_c188 bl_188 br_188 wl_62 vdd gnd cell_6t
Xbit_r63_c188 bl_188 br_188 wl_63 vdd gnd cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd cell_6t
Xbit_r1_c189 bl_189 br_189 wl_1 vdd gnd cell_6t
Xbit_r2_c189 bl_189 br_189 wl_2 vdd gnd cell_6t
Xbit_r3_c189 bl_189 br_189 wl_3 vdd gnd cell_6t
Xbit_r4_c189 bl_189 br_189 wl_4 vdd gnd cell_6t
Xbit_r5_c189 bl_189 br_189 wl_5 vdd gnd cell_6t
Xbit_r6_c189 bl_189 br_189 wl_6 vdd gnd cell_6t
Xbit_r7_c189 bl_189 br_189 wl_7 vdd gnd cell_6t
Xbit_r8_c189 bl_189 br_189 wl_8 vdd gnd cell_6t
Xbit_r9_c189 bl_189 br_189 wl_9 vdd gnd cell_6t
Xbit_r10_c189 bl_189 br_189 wl_10 vdd gnd cell_6t
Xbit_r11_c189 bl_189 br_189 wl_11 vdd gnd cell_6t
Xbit_r12_c189 bl_189 br_189 wl_12 vdd gnd cell_6t
Xbit_r13_c189 bl_189 br_189 wl_13 vdd gnd cell_6t
Xbit_r14_c189 bl_189 br_189 wl_14 vdd gnd cell_6t
Xbit_r15_c189 bl_189 br_189 wl_15 vdd gnd cell_6t
Xbit_r16_c189 bl_189 br_189 wl_16 vdd gnd cell_6t
Xbit_r17_c189 bl_189 br_189 wl_17 vdd gnd cell_6t
Xbit_r18_c189 bl_189 br_189 wl_18 vdd gnd cell_6t
Xbit_r19_c189 bl_189 br_189 wl_19 vdd gnd cell_6t
Xbit_r20_c189 bl_189 br_189 wl_20 vdd gnd cell_6t
Xbit_r21_c189 bl_189 br_189 wl_21 vdd gnd cell_6t
Xbit_r22_c189 bl_189 br_189 wl_22 vdd gnd cell_6t
Xbit_r23_c189 bl_189 br_189 wl_23 vdd gnd cell_6t
Xbit_r24_c189 bl_189 br_189 wl_24 vdd gnd cell_6t
Xbit_r25_c189 bl_189 br_189 wl_25 vdd gnd cell_6t
Xbit_r26_c189 bl_189 br_189 wl_26 vdd gnd cell_6t
Xbit_r27_c189 bl_189 br_189 wl_27 vdd gnd cell_6t
Xbit_r28_c189 bl_189 br_189 wl_28 vdd gnd cell_6t
Xbit_r29_c189 bl_189 br_189 wl_29 vdd gnd cell_6t
Xbit_r30_c189 bl_189 br_189 wl_30 vdd gnd cell_6t
Xbit_r31_c189 bl_189 br_189 wl_31 vdd gnd cell_6t
Xbit_r32_c189 bl_189 br_189 wl_32 vdd gnd cell_6t
Xbit_r33_c189 bl_189 br_189 wl_33 vdd gnd cell_6t
Xbit_r34_c189 bl_189 br_189 wl_34 vdd gnd cell_6t
Xbit_r35_c189 bl_189 br_189 wl_35 vdd gnd cell_6t
Xbit_r36_c189 bl_189 br_189 wl_36 vdd gnd cell_6t
Xbit_r37_c189 bl_189 br_189 wl_37 vdd gnd cell_6t
Xbit_r38_c189 bl_189 br_189 wl_38 vdd gnd cell_6t
Xbit_r39_c189 bl_189 br_189 wl_39 vdd gnd cell_6t
Xbit_r40_c189 bl_189 br_189 wl_40 vdd gnd cell_6t
Xbit_r41_c189 bl_189 br_189 wl_41 vdd gnd cell_6t
Xbit_r42_c189 bl_189 br_189 wl_42 vdd gnd cell_6t
Xbit_r43_c189 bl_189 br_189 wl_43 vdd gnd cell_6t
Xbit_r44_c189 bl_189 br_189 wl_44 vdd gnd cell_6t
Xbit_r45_c189 bl_189 br_189 wl_45 vdd gnd cell_6t
Xbit_r46_c189 bl_189 br_189 wl_46 vdd gnd cell_6t
Xbit_r47_c189 bl_189 br_189 wl_47 vdd gnd cell_6t
Xbit_r48_c189 bl_189 br_189 wl_48 vdd gnd cell_6t
Xbit_r49_c189 bl_189 br_189 wl_49 vdd gnd cell_6t
Xbit_r50_c189 bl_189 br_189 wl_50 vdd gnd cell_6t
Xbit_r51_c189 bl_189 br_189 wl_51 vdd gnd cell_6t
Xbit_r52_c189 bl_189 br_189 wl_52 vdd gnd cell_6t
Xbit_r53_c189 bl_189 br_189 wl_53 vdd gnd cell_6t
Xbit_r54_c189 bl_189 br_189 wl_54 vdd gnd cell_6t
Xbit_r55_c189 bl_189 br_189 wl_55 vdd gnd cell_6t
Xbit_r56_c189 bl_189 br_189 wl_56 vdd gnd cell_6t
Xbit_r57_c189 bl_189 br_189 wl_57 vdd gnd cell_6t
Xbit_r58_c189 bl_189 br_189 wl_58 vdd gnd cell_6t
Xbit_r59_c189 bl_189 br_189 wl_59 vdd gnd cell_6t
Xbit_r60_c189 bl_189 br_189 wl_60 vdd gnd cell_6t
Xbit_r61_c189 bl_189 br_189 wl_61 vdd gnd cell_6t
Xbit_r62_c189 bl_189 br_189 wl_62 vdd gnd cell_6t
Xbit_r63_c189 bl_189 br_189 wl_63 vdd gnd cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd cell_6t
Xbit_r1_c190 bl_190 br_190 wl_1 vdd gnd cell_6t
Xbit_r2_c190 bl_190 br_190 wl_2 vdd gnd cell_6t
Xbit_r3_c190 bl_190 br_190 wl_3 vdd gnd cell_6t
Xbit_r4_c190 bl_190 br_190 wl_4 vdd gnd cell_6t
Xbit_r5_c190 bl_190 br_190 wl_5 vdd gnd cell_6t
Xbit_r6_c190 bl_190 br_190 wl_6 vdd gnd cell_6t
Xbit_r7_c190 bl_190 br_190 wl_7 vdd gnd cell_6t
Xbit_r8_c190 bl_190 br_190 wl_8 vdd gnd cell_6t
Xbit_r9_c190 bl_190 br_190 wl_9 vdd gnd cell_6t
Xbit_r10_c190 bl_190 br_190 wl_10 vdd gnd cell_6t
Xbit_r11_c190 bl_190 br_190 wl_11 vdd gnd cell_6t
Xbit_r12_c190 bl_190 br_190 wl_12 vdd gnd cell_6t
Xbit_r13_c190 bl_190 br_190 wl_13 vdd gnd cell_6t
Xbit_r14_c190 bl_190 br_190 wl_14 vdd gnd cell_6t
Xbit_r15_c190 bl_190 br_190 wl_15 vdd gnd cell_6t
Xbit_r16_c190 bl_190 br_190 wl_16 vdd gnd cell_6t
Xbit_r17_c190 bl_190 br_190 wl_17 vdd gnd cell_6t
Xbit_r18_c190 bl_190 br_190 wl_18 vdd gnd cell_6t
Xbit_r19_c190 bl_190 br_190 wl_19 vdd gnd cell_6t
Xbit_r20_c190 bl_190 br_190 wl_20 vdd gnd cell_6t
Xbit_r21_c190 bl_190 br_190 wl_21 vdd gnd cell_6t
Xbit_r22_c190 bl_190 br_190 wl_22 vdd gnd cell_6t
Xbit_r23_c190 bl_190 br_190 wl_23 vdd gnd cell_6t
Xbit_r24_c190 bl_190 br_190 wl_24 vdd gnd cell_6t
Xbit_r25_c190 bl_190 br_190 wl_25 vdd gnd cell_6t
Xbit_r26_c190 bl_190 br_190 wl_26 vdd gnd cell_6t
Xbit_r27_c190 bl_190 br_190 wl_27 vdd gnd cell_6t
Xbit_r28_c190 bl_190 br_190 wl_28 vdd gnd cell_6t
Xbit_r29_c190 bl_190 br_190 wl_29 vdd gnd cell_6t
Xbit_r30_c190 bl_190 br_190 wl_30 vdd gnd cell_6t
Xbit_r31_c190 bl_190 br_190 wl_31 vdd gnd cell_6t
Xbit_r32_c190 bl_190 br_190 wl_32 vdd gnd cell_6t
Xbit_r33_c190 bl_190 br_190 wl_33 vdd gnd cell_6t
Xbit_r34_c190 bl_190 br_190 wl_34 vdd gnd cell_6t
Xbit_r35_c190 bl_190 br_190 wl_35 vdd gnd cell_6t
Xbit_r36_c190 bl_190 br_190 wl_36 vdd gnd cell_6t
Xbit_r37_c190 bl_190 br_190 wl_37 vdd gnd cell_6t
Xbit_r38_c190 bl_190 br_190 wl_38 vdd gnd cell_6t
Xbit_r39_c190 bl_190 br_190 wl_39 vdd gnd cell_6t
Xbit_r40_c190 bl_190 br_190 wl_40 vdd gnd cell_6t
Xbit_r41_c190 bl_190 br_190 wl_41 vdd gnd cell_6t
Xbit_r42_c190 bl_190 br_190 wl_42 vdd gnd cell_6t
Xbit_r43_c190 bl_190 br_190 wl_43 vdd gnd cell_6t
Xbit_r44_c190 bl_190 br_190 wl_44 vdd gnd cell_6t
Xbit_r45_c190 bl_190 br_190 wl_45 vdd gnd cell_6t
Xbit_r46_c190 bl_190 br_190 wl_46 vdd gnd cell_6t
Xbit_r47_c190 bl_190 br_190 wl_47 vdd gnd cell_6t
Xbit_r48_c190 bl_190 br_190 wl_48 vdd gnd cell_6t
Xbit_r49_c190 bl_190 br_190 wl_49 vdd gnd cell_6t
Xbit_r50_c190 bl_190 br_190 wl_50 vdd gnd cell_6t
Xbit_r51_c190 bl_190 br_190 wl_51 vdd gnd cell_6t
Xbit_r52_c190 bl_190 br_190 wl_52 vdd gnd cell_6t
Xbit_r53_c190 bl_190 br_190 wl_53 vdd gnd cell_6t
Xbit_r54_c190 bl_190 br_190 wl_54 vdd gnd cell_6t
Xbit_r55_c190 bl_190 br_190 wl_55 vdd gnd cell_6t
Xbit_r56_c190 bl_190 br_190 wl_56 vdd gnd cell_6t
Xbit_r57_c190 bl_190 br_190 wl_57 vdd gnd cell_6t
Xbit_r58_c190 bl_190 br_190 wl_58 vdd gnd cell_6t
Xbit_r59_c190 bl_190 br_190 wl_59 vdd gnd cell_6t
Xbit_r60_c190 bl_190 br_190 wl_60 vdd gnd cell_6t
Xbit_r61_c190 bl_190 br_190 wl_61 vdd gnd cell_6t
Xbit_r62_c190 bl_190 br_190 wl_62 vdd gnd cell_6t
Xbit_r63_c190 bl_190 br_190 wl_63 vdd gnd cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd cell_6t
Xbit_r1_c191 bl_191 br_191 wl_1 vdd gnd cell_6t
Xbit_r2_c191 bl_191 br_191 wl_2 vdd gnd cell_6t
Xbit_r3_c191 bl_191 br_191 wl_3 vdd gnd cell_6t
Xbit_r4_c191 bl_191 br_191 wl_4 vdd gnd cell_6t
Xbit_r5_c191 bl_191 br_191 wl_5 vdd gnd cell_6t
Xbit_r6_c191 bl_191 br_191 wl_6 vdd gnd cell_6t
Xbit_r7_c191 bl_191 br_191 wl_7 vdd gnd cell_6t
Xbit_r8_c191 bl_191 br_191 wl_8 vdd gnd cell_6t
Xbit_r9_c191 bl_191 br_191 wl_9 vdd gnd cell_6t
Xbit_r10_c191 bl_191 br_191 wl_10 vdd gnd cell_6t
Xbit_r11_c191 bl_191 br_191 wl_11 vdd gnd cell_6t
Xbit_r12_c191 bl_191 br_191 wl_12 vdd gnd cell_6t
Xbit_r13_c191 bl_191 br_191 wl_13 vdd gnd cell_6t
Xbit_r14_c191 bl_191 br_191 wl_14 vdd gnd cell_6t
Xbit_r15_c191 bl_191 br_191 wl_15 vdd gnd cell_6t
Xbit_r16_c191 bl_191 br_191 wl_16 vdd gnd cell_6t
Xbit_r17_c191 bl_191 br_191 wl_17 vdd gnd cell_6t
Xbit_r18_c191 bl_191 br_191 wl_18 vdd gnd cell_6t
Xbit_r19_c191 bl_191 br_191 wl_19 vdd gnd cell_6t
Xbit_r20_c191 bl_191 br_191 wl_20 vdd gnd cell_6t
Xbit_r21_c191 bl_191 br_191 wl_21 vdd gnd cell_6t
Xbit_r22_c191 bl_191 br_191 wl_22 vdd gnd cell_6t
Xbit_r23_c191 bl_191 br_191 wl_23 vdd gnd cell_6t
Xbit_r24_c191 bl_191 br_191 wl_24 vdd gnd cell_6t
Xbit_r25_c191 bl_191 br_191 wl_25 vdd gnd cell_6t
Xbit_r26_c191 bl_191 br_191 wl_26 vdd gnd cell_6t
Xbit_r27_c191 bl_191 br_191 wl_27 vdd gnd cell_6t
Xbit_r28_c191 bl_191 br_191 wl_28 vdd gnd cell_6t
Xbit_r29_c191 bl_191 br_191 wl_29 vdd gnd cell_6t
Xbit_r30_c191 bl_191 br_191 wl_30 vdd gnd cell_6t
Xbit_r31_c191 bl_191 br_191 wl_31 vdd gnd cell_6t
Xbit_r32_c191 bl_191 br_191 wl_32 vdd gnd cell_6t
Xbit_r33_c191 bl_191 br_191 wl_33 vdd gnd cell_6t
Xbit_r34_c191 bl_191 br_191 wl_34 vdd gnd cell_6t
Xbit_r35_c191 bl_191 br_191 wl_35 vdd gnd cell_6t
Xbit_r36_c191 bl_191 br_191 wl_36 vdd gnd cell_6t
Xbit_r37_c191 bl_191 br_191 wl_37 vdd gnd cell_6t
Xbit_r38_c191 bl_191 br_191 wl_38 vdd gnd cell_6t
Xbit_r39_c191 bl_191 br_191 wl_39 vdd gnd cell_6t
Xbit_r40_c191 bl_191 br_191 wl_40 vdd gnd cell_6t
Xbit_r41_c191 bl_191 br_191 wl_41 vdd gnd cell_6t
Xbit_r42_c191 bl_191 br_191 wl_42 vdd gnd cell_6t
Xbit_r43_c191 bl_191 br_191 wl_43 vdd gnd cell_6t
Xbit_r44_c191 bl_191 br_191 wl_44 vdd gnd cell_6t
Xbit_r45_c191 bl_191 br_191 wl_45 vdd gnd cell_6t
Xbit_r46_c191 bl_191 br_191 wl_46 vdd gnd cell_6t
Xbit_r47_c191 bl_191 br_191 wl_47 vdd gnd cell_6t
Xbit_r48_c191 bl_191 br_191 wl_48 vdd gnd cell_6t
Xbit_r49_c191 bl_191 br_191 wl_49 vdd gnd cell_6t
Xbit_r50_c191 bl_191 br_191 wl_50 vdd gnd cell_6t
Xbit_r51_c191 bl_191 br_191 wl_51 vdd gnd cell_6t
Xbit_r52_c191 bl_191 br_191 wl_52 vdd gnd cell_6t
Xbit_r53_c191 bl_191 br_191 wl_53 vdd gnd cell_6t
Xbit_r54_c191 bl_191 br_191 wl_54 vdd gnd cell_6t
Xbit_r55_c191 bl_191 br_191 wl_55 vdd gnd cell_6t
Xbit_r56_c191 bl_191 br_191 wl_56 vdd gnd cell_6t
Xbit_r57_c191 bl_191 br_191 wl_57 vdd gnd cell_6t
Xbit_r58_c191 bl_191 br_191 wl_58 vdd gnd cell_6t
Xbit_r59_c191 bl_191 br_191 wl_59 vdd gnd cell_6t
Xbit_r60_c191 bl_191 br_191 wl_60 vdd gnd cell_6t
Xbit_r61_c191 bl_191 br_191 wl_61 vdd gnd cell_6t
Xbit_r62_c191 bl_191 br_191 wl_62 vdd gnd cell_6t
Xbit_r63_c191 bl_191 br_191 wl_63 vdd gnd cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd cell_6t
Xbit_r1_c192 bl_192 br_192 wl_1 vdd gnd cell_6t
Xbit_r2_c192 bl_192 br_192 wl_2 vdd gnd cell_6t
Xbit_r3_c192 bl_192 br_192 wl_3 vdd gnd cell_6t
Xbit_r4_c192 bl_192 br_192 wl_4 vdd gnd cell_6t
Xbit_r5_c192 bl_192 br_192 wl_5 vdd gnd cell_6t
Xbit_r6_c192 bl_192 br_192 wl_6 vdd gnd cell_6t
Xbit_r7_c192 bl_192 br_192 wl_7 vdd gnd cell_6t
Xbit_r8_c192 bl_192 br_192 wl_8 vdd gnd cell_6t
Xbit_r9_c192 bl_192 br_192 wl_9 vdd gnd cell_6t
Xbit_r10_c192 bl_192 br_192 wl_10 vdd gnd cell_6t
Xbit_r11_c192 bl_192 br_192 wl_11 vdd gnd cell_6t
Xbit_r12_c192 bl_192 br_192 wl_12 vdd gnd cell_6t
Xbit_r13_c192 bl_192 br_192 wl_13 vdd gnd cell_6t
Xbit_r14_c192 bl_192 br_192 wl_14 vdd gnd cell_6t
Xbit_r15_c192 bl_192 br_192 wl_15 vdd gnd cell_6t
Xbit_r16_c192 bl_192 br_192 wl_16 vdd gnd cell_6t
Xbit_r17_c192 bl_192 br_192 wl_17 vdd gnd cell_6t
Xbit_r18_c192 bl_192 br_192 wl_18 vdd gnd cell_6t
Xbit_r19_c192 bl_192 br_192 wl_19 vdd gnd cell_6t
Xbit_r20_c192 bl_192 br_192 wl_20 vdd gnd cell_6t
Xbit_r21_c192 bl_192 br_192 wl_21 vdd gnd cell_6t
Xbit_r22_c192 bl_192 br_192 wl_22 vdd gnd cell_6t
Xbit_r23_c192 bl_192 br_192 wl_23 vdd gnd cell_6t
Xbit_r24_c192 bl_192 br_192 wl_24 vdd gnd cell_6t
Xbit_r25_c192 bl_192 br_192 wl_25 vdd gnd cell_6t
Xbit_r26_c192 bl_192 br_192 wl_26 vdd gnd cell_6t
Xbit_r27_c192 bl_192 br_192 wl_27 vdd gnd cell_6t
Xbit_r28_c192 bl_192 br_192 wl_28 vdd gnd cell_6t
Xbit_r29_c192 bl_192 br_192 wl_29 vdd gnd cell_6t
Xbit_r30_c192 bl_192 br_192 wl_30 vdd gnd cell_6t
Xbit_r31_c192 bl_192 br_192 wl_31 vdd gnd cell_6t
Xbit_r32_c192 bl_192 br_192 wl_32 vdd gnd cell_6t
Xbit_r33_c192 bl_192 br_192 wl_33 vdd gnd cell_6t
Xbit_r34_c192 bl_192 br_192 wl_34 vdd gnd cell_6t
Xbit_r35_c192 bl_192 br_192 wl_35 vdd gnd cell_6t
Xbit_r36_c192 bl_192 br_192 wl_36 vdd gnd cell_6t
Xbit_r37_c192 bl_192 br_192 wl_37 vdd gnd cell_6t
Xbit_r38_c192 bl_192 br_192 wl_38 vdd gnd cell_6t
Xbit_r39_c192 bl_192 br_192 wl_39 vdd gnd cell_6t
Xbit_r40_c192 bl_192 br_192 wl_40 vdd gnd cell_6t
Xbit_r41_c192 bl_192 br_192 wl_41 vdd gnd cell_6t
Xbit_r42_c192 bl_192 br_192 wl_42 vdd gnd cell_6t
Xbit_r43_c192 bl_192 br_192 wl_43 vdd gnd cell_6t
Xbit_r44_c192 bl_192 br_192 wl_44 vdd gnd cell_6t
Xbit_r45_c192 bl_192 br_192 wl_45 vdd gnd cell_6t
Xbit_r46_c192 bl_192 br_192 wl_46 vdd gnd cell_6t
Xbit_r47_c192 bl_192 br_192 wl_47 vdd gnd cell_6t
Xbit_r48_c192 bl_192 br_192 wl_48 vdd gnd cell_6t
Xbit_r49_c192 bl_192 br_192 wl_49 vdd gnd cell_6t
Xbit_r50_c192 bl_192 br_192 wl_50 vdd gnd cell_6t
Xbit_r51_c192 bl_192 br_192 wl_51 vdd gnd cell_6t
Xbit_r52_c192 bl_192 br_192 wl_52 vdd gnd cell_6t
Xbit_r53_c192 bl_192 br_192 wl_53 vdd gnd cell_6t
Xbit_r54_c192 bl_192 br_192 wl_54 vdd gnd cell_6t
Xbit_r55_c192 bl_192 br_192 wl_55 vdd gnd cell_6t
Xbit_r56_c192 bl_192 br_192 wl_56 vdd gnd cell_6t
Xbit_r57_c192 bl_192 br_192 wl_57 vdd gnd cell_6t
Xbit_r58_c192 bl_192 br_192 wl_58 vdd gnd cell_6t
Xbit_r59_c192 bl_192 br_192 wl_59 vdd gnd cell_6t
Xbit_r60_c192 bl_192 br_192 wl_60 vdd gnd cell_6t
Xbit_r61_c192 bl_192 br_192 wl_61 vdd gnd cell_6t
Xbit_r62_c192 bl_192 br_192 wl_62 vdd gnd cell_6t
Xbit_r63_c192 bl_192 br_192 wl_63 vdd gnd cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd cell_6t
Xbit_r1_c193 bl_193 br_193 wl_1 vdd gnd cell_6t
Xbit_r2_c193 bl_193 br_193 wl_2 vdd gnd cell_6t
Xbit_r3_c193 bl_193 br_193 wl_3 vdd gnd cell_6t
Xbit_r4_c193 bl_193 br_193 wl_4 vdd gnd cell_6t
Xbit_r5_c193 bl_193 br_193 wl_5 vdd gnd cell_6t
Xbit_r6_c193 bl_193 br_193 wl_6 vdd gnd cell_6t
Xbit_r7_c193 bl_193 br_193 wl_7 vdd gnd cell_6t
Xbit_r8_c193 bl_193 br_193 wl_8 vdd gnd cell_6t
Xbit_r9_c193 bl_193 br_193 wl_9 vdd gnd cell_6t
Xbit_r10_c193 bl_193 br_193 wl_10 vdd gnd cell_6t
Xbit_r11_c193 bl_193 br_193 wl_11 vdd gnd cell_6t
Xbit_r12_c193 bl_193 br_193 wl_12 vdd gnd cell_6t
Xbit_r13_c193 bl_193 br_193 wl_13 vdd gnd cell_6t
Xbit_r14_c193 bl_193 br_193 wl_14 vdd gnd cell_6t
Xbit_r15_c193 bl_193 br_193 wl_15 vdd gnd cell_6t
Xbit_r16_c193 bl_193 br_193 wl_16 vdd gnd cell_6t
Xbit_r17_c193 bl_193 br_193 wl_17 vdd gnd cell_6t
Xbit_r18_c193 bl_193 br_193 wl_18 vdd gnd cell_6t
Xbit_r19_c193 bl_193 br_193 wl_19 vdd gnd cell_6t
Xbit_r20_c193 bl_193 br_193 wl_20 vdd gnd cell_6t
Xbit_r21_c193 bl_193 br_193 wl_21 vdd gnd cell_6t
Xbit_r22_c193 bl_193 br_193 wl_22 vdd gnd cell_6t
Xbit_r23_c193 bl_193 br_193 wl_23 vdd gnd cell_6t
Xbit_r24_c193 bl_193 br_193 wl_24 vdd gnd cell_6t
Xbit_r25_c193 bl_193 br_193 wl_25 vdd gnd cell_6t
Xbit_r26_c193 bl_193 br_193 wl_26 vdd gnd cell_6t
Xbit_r27_c193 bl_193 br_193 wl_27 vdd gnd cell_6t
Xbit_r28_c193 bl_193 br_193 wl_28 vdd gnd cell_6t
Xbit_r29_c193 bl_193 br_193 wl_29 vdd gnd cell_6t
Xbit_r30_c193 bl_193 br_193 wl_30 vdd gnd cell_6t
Xbit_r31_c193 bl_193 br_193 wl_31 vdd gnd cell_6t
Xbit_r32_c193 bl_193 br_193 wl_32 vdd gnd cell_6t
Xbit_r33_c193 bl_193 br_193 wl_33 vdd gnd cell_6t
Xbit_r34_c193 bl_193 br_193 wl_34 vdd gnd cell_6t
Xbit_r35_c193 bl_193 br_193 wl_35 vdd gnd cell_6t
Xbit_r36_c193 bl_193 br_193 wl_36 vdd gnd cell_6t
Xbit_r37_c193 bl_193 br_193 wl_37 vdd gnd cell_6t
Xbit_r38_c193 bl_193 br_193 wl_38 vdd gnd cell_6t
Xbit_r39_c193 bl_193 br_193 wl_39 vdd gnd cell_6t
Xbit_r40_c193 bl_193 br_193 wl_40 vdd gnd cell_6t
Xbit_r41_c193 bl_193 br_193 wl_41 vdd gnd cell_6t
Xbit_r42_c193 bl_193 br_193 wl_42 vdd gnd cell_6t
Xbit_r43_c193 bl_193 br_193 wl_43 vdd gnd cell_6t
Xbit_r44_c193 bl_193 br_193 wl_44 vdd gnd cell_6t
Xbit_r45_c193 bl_193 br_193 wl_45 vdd gnd cell_6t
Xbit_r46_c193 bl_193 br_193 wl_46 vdd gnd cell_6t
Xbit_r47_c193 bl_193 br_193 wl_47 vdd gnd cell_6t
Xbit_r48_c193 bl_193 br_193 wl_48 vdd gnd cell_6t
Xbit_r49_c193 bl_193 br_193 wl_49 vdd gnd cell_6t
Xbit_r50_c193 bl_193 br_193 wl_50 vdd gnd cell_6t
Xbit_r51_c193 bl_193 br_193 wl_51 vdd gnd cell_6t
Xbit_r52_c193 bl_193 br_193 wl_52 vdd gnd cell_6t
Xbit_r53_c193 bl_193 br_193 wl_53 vdd gnd cell_6t
Xbit_r54_c193 bl_193 br_193 wl_54 vdd gnd cell_6t
Xbit_r55_c193 bl_193 br_193 wl_55 vdd gnd cell_6t
Xbit_r56_c193 bl_193 br_193 wl_56 vdd gnd cell_6t
Xbit_r57_c193 bl_193 br_193 wl_57 vdd gnd cell_6t
Xbit_r58_c193 bl_193 br_193 wl_58 vdd gnd cell_6t
Xbit_r59_c193 bl_193 br_193 wl_59 vdd gnd cell_6t
Xbit_r60_c193 bl_193 br_193 wl_60 vdd gnd cell_6t
Xbit_r61_c193 bl_193 br_193 wl_61 vdd gnd cell_6t
Xbit_r62_c193 bl_193 br_193 wl_62 vdd gnd cell_6t
Xbit_r63_c193 bl_193 br_193 wl_63 vdd gnd cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd cell_6t
Xbit_r1_c194 bl_194 br_194 wl_1 vdd gnd cell_6t
Xbit_r2_c194 bl_194 br_194 wl_2 vdd gnd cell_6t
Xbit_r3_c194 bl_194 br_194 wl_3 vdd gnd cell_6t
Xbit_r4_c194 bl_194 br_194 wl_4 vdd gnd cell_6t
Xbit_r5_c194 bl_194 br_194 wl_5 vdd gnd cell_6t
Xbit_r6_c194 bl_194 br_194 wl_6 vdd gnd cell_6t
Xbit_r7_c194 bl_194 br_194 wl_7 vdd gnd cell_6t
Xbit_r8_c194 bl_194 br_194 wl_8 vdd gnd cell_6t
Xbit_r9_c194 bl_194 br_194 wl_9 vdd gnd cell_6t
Xbit_r10_c194 bl_194 br_194 wl_10 vdd gnd cell_6t
Xbit_r11_c194 bl_194 br_194 wl_11 vdd gnd cell_6t
Xbit_r12_c194 bl_194 br_194 wl_12 vdd gnd cell_6t
Xbit_r13_c194 bl_194 br_194 wl_13 vdd gnd cell_6t
Xbit_r14_c194 bl_194 br_194 wl_14 vdd gnd cell_6t
Xbit_r15_c194 bl_194 br_194 wl_15 vdd gnd cell_6t
Xbit_r16_c194 bl_194 br_194 wl_16 vdd gnd cell_6t
Xbit_r17_c194 bl_194 br_194 wl_17 vdd gnd cell_6t
Xbit_r18_c194 bl_194 br_194 wl_18 vdd gnd cell_6t
Xbit_r19_c194 bl_194 br_194 wl_19 vdd gnd cell_6t
Xbit_r20_c194 bl_194 br_194 wl_20 vdd gnd cell_6t
Xbit_r21_c194 bl_194 br_194 wl_21 vdd gnd cell_6t
Xbit_r22_c194 bl_194 br_194 wl_22 vdd gnd cell_6t
Xbit_r23_c194 bl_194 br_194 wl_23 vdd gnd cell_6t
Xbit_r24_c194 bl_194 br_194 wl_24 vdd gnd cell_6t
Xbit_r25_c194 bl_194 br_194 wl_25 vdd gnd cell_6t
Xbit_r26_c194 bl_194 br_194 wl_26 vdd gnd cell_6t
Xbit_r27_c194 bl_194 br_194 wl_27 vdd gnd cell_6t
Xbit_r28_c194 bl_194 br_194 wl_28 vdd gnd cell_6t
Xbit_r29_c194 bl_194 br_194 wl_29 vdd gnd cell_6t
Xbit_r30_c194 bl_194 br_194 wl_30 vdd gnd cell_6t
Xbit_r31_c194 bl_194 br_194 wl_31 vdd gnd cell_6t
Xbit_r32_c194 bl_194 br_194 wl_32 vdd gnd cell_6t
Xbit_r33_c194 bl_194 br_194 wl_33 vdd gnd cell_6t
Xbit_r34_c194 bl_194 br_194 wl_34 vdd gnd cell_6t
Xbit_r35_c194 bl_194 br_194 wl_35 vdd gnd cell_6t
Xbit_r36_c194 bl_194 br_194 wl_36 vdd gnd cell_6t
Xbit_r37_c194 bl_194 br_194 wl_37 vdd gnd cell_6t
Xbit_r38_c194 bl_194 br_194 wl_38 vdd gnd cell_6t
Xbit_r39_c194 bl_194 br_194 wl_39 vdd gnd cell_6t
Xbit_r40_c194 bl_194 br_194 wl_40 vdd gnd cell_6t
Xbit_r41_c194 bl_194 br_194 wl_41 vdd gnd cell_6t
Xbit_r42_c194 bl_194 br_194 wl_42 vdd gnd cell_6t
Xbit_r43_c194 bl_194 br_194 wl_43 vdd gnd cell_6t
Xbit_r44_c194 bl_194 br_194 wl_44 vdd gnd cell_6t
Xbit_r45_c194 bl_194 br_194 wl_45 vdd gnd cell_6t
Xbit_r46_c194 bl_194 br_194 wl_46 vdd gnd cell_6t
Xbit_r47_c194 bl_194 br_194 wl_47 vdd gnd cell_6t
Xbit_r48_c194 bl_194 br_194 wl_48 vdd gnd cell_6t
Xbit_r49_c194 bl_194 br_194 wl_49 vdd gnd cell_6t
Xbit_r50_c194 bl_194 br_194 wl_50 vdd gnd cell_6t
Xbit_r51_c194 bl_194 br_194 wl_51 vdd gnd cell_6t
Xbit_r52_c194 bl_194 br_194 wl_52 vdd gnd cell_6t
Xbit_r53_c194 bl_194 br_194 wl_53 vdd gnd cell_6t
Xbit_r54_c194 bl_194 br_194 wl_54 vdd gnd cell_6t
Xbit_r55_c194 bl_194 br_194 wl_55 vdd gnd cell_6t
Xbit_r56_c194 bl_194 br_194 wl_56 vdd gnd cell_6t
Xbit_r57_c194 bl_194 br_194 wl_57 vdd gnd cell_6t
Xbit_r58_c194 bl_194 br_194 wl_58 vdd gnd cell_6t
Xbit_r59_c194 bl_194 br_194 wl_59 vdd gnd cell_6t
Xbit_r60_c194 bl_194 br_194 wl_60 vdd gnd cell_6t
Xbit_r61_c194 bl_194 br_194 wl_61 vdd gnd cell_6t
Xbit_r62_c194 bl_194 br_194 wl_62 vdd gnd cell_6t
Xbit_r63_c194 bl_194 br_194 wl_63 vdd gnd cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd cell_6t
Xbit_r1_c195 bl_195 br_195 wl_1 vdd gnd cell_6t
Xbit_r2_c195 bl_195 br_195 wl_2 vdd gnd cell_6t
Xbit_r3_c195 bl_195 br_195 wl_3 vdd gnd cell_6t
Xbit_r4_c195 bl_195 br_195 wl_4 vdd gnd cell_6t
Xbit_r5_c195 bl_195 br_195 wl_5 vdd gnd cell_6t
Xbit_r6_c195 bl_195 br_195 wl_6 vdd gnd cell_6t
Xbit_r7_c195 bl_195 br_195 wl_7 vdd gnd cell_6t
Xbit_r8_c195 bl_195 br_195 wl_8 vdd gnd cell_6t
Xbit_r9_c195 bl_195 br_195 wl_9 vdd gnd cell_6t
Xbit_r10_c195 bl_195 br_195 wl_10 vdd gnd cell_6t
Xbit_r11_c195 bl_195 br_195 wl_11 vdd gnd cell_6t
Xbit_r12_c195 bl_195 br_195 wl_12 vdd gnd cell_6t
Xbit_r13_c195 bl_195 br_195 wl_13 vdd gnd cell_6t
Xbit_r14_c195 bl_195 br_195 wl_14 vdd gnd cell_6t
Xbit_r15_c195 bl_195 br_195 wl_15 vdd gnd cell_6t
Xbit_r16_c195 bl_195 br_195 wl_16 vdd gnd cell_6t
Xbit_r17_c195 bl_195 br_195 wl_17 vdd gnd cell_6t
Xbit_r18_c195 bl_195 br_195 wl_18 vdd gnd cell_6t
Xbit_r19_c195 bl_195 br_195 wl_19 vdd gnd cell_6t
Xbit_r20_c195 bl_195 br_195 wl_20 vdd gnd cell_6t
Xbit_r21_c195 bl_195 br_195 wl_21 vdd gnd cell_6t
Xbit_r22_c195 bl_195 br_195 wl_22 vdd gnd cell_6t
Xbit_r23_c195 bl_195 br_195 wl_23 vdd gnd cell_6t
Xbit_r24_c195 bl_195 br_195 wl_24 vdd gnd cell_6t
Xbit_r25_c195 bl_195 br_195 wl_25 vdd gnd cell_6t
Xbit_r26_c195 bl_195 br_195 wl_26 vdd gnd cell_6t
Xbit_r27_c195 bl_195 br_195 wl_27 vdd gnd cell_6t
Xbit_r28_c195 bl_195 br_195 wl_28 vdd gnd cell_6t
Xbit_r29_c195 bl_195 br_195 wl_29 vdd gnd cell_6t
Xbit_r30_c195 bl_195 br_195 wl_30 vdd gnd cell_6t
Xbit_r31_c195 bl_195 br_195 wl_31 vdd gnd cell_6t
Xbit_r32_c195 bl_195 br_195 wl_32 vdd gnd cell_6t
Xbit_r33_c195 bl_195 br_195 wl_33 vdd gnd cell_6t
Xbit_r34_c195 bl_195 br_195 wl_34 vdd gnd cell_6t
Xbit_r35_c195 bl_195 br_195 wl_35 vdd gnd cell_6t
Xbit_r36_c195 bl_195 br_195 wl_36 vdd gnd cell_6t
Xbit_r37_c195 bl_195 br_195 wl_37 vdd gnd cell_6t
Xbit_r38_c195 bl_195 br_195 wl_38 vdd gnd cell_6t
Xbit_r39_c195 bl_195 br_195 wl_39 vdd gnd cell_6t
Xbit_r40_c195 bl_195 br_195 wl_40 vdd gnd cell_6t
Xbit_r41_c195 bl_195 br_195 wl_41 vdd gnd cell_6t
Xbit_r42_c195 bl_195 br_195 wl_42 vdd gnd cell_6t
Xbit_r43_c195 bl_195 br_195 wl_43 vdd gnd cell_6t
Xbit_r44_c195 bl_195 br_195 wl_44 vdd gnd cell_6t
Xbit_r45_c195 bl_195 br_195 wl_45 vdd gnd cell_6t
Xbit_r46_c195 bl_195 br_195 wl_46 vdd gnd cell_6t
Xbit_r47_c195 bl_195 br_195 wl_47 vdd gnd cell_6t
Xbit_r48_c195 bl_195 br_195 wl_48 vdd gnd cell_6t
Xbit_r49_c195 bl_195 br_195 wl_49 vdd gnd cell_6t
Xbit_r50_c195 bl_195 br_195 wl_50 vdd gnd cell_6t
Xbit_r51_c195 bl_195 br_195 wl_51 vdd gnd cell_6t
Xbit_r52_c195 bl_195 br_195 wl_52 vdd gnd cell_6t
Xbit_r53_c195 bl_195 br_195 wl_53 vdd gnd cell_6t
Xbit_r54_c195 bl_195 br_195 wl_54 vdd gnd cell_6t
Xbit_r55_c195 bl_195 br_195 wl_55 vdd gnd cell_6t
Xbit_r56_c195 bl_195 br_195 wl_56 vdd gnd cell_6t
Xbit_r57_c195 bl_195 br_195 wl_57 vdd gnd cell_6t
Xbit_r58_c195 bl_195 br_195 wl_58 vdd gnd cell_6t
Xbit_r59_c195 bl_195 br_195 wl_59 vdd gnd cell_6t
Xbit_r60_c195 bl_195 br_195 wl_60 vdd gnd cell_6t
Xbit_r61_c195 bl_195 br_195 wl_61 vdd gnd cell_6t
Xbit_r62_c195 bl_195 br_195 wl_62 vdd gnd cell_6t
Xbit_r63_c195 bl_195 br_195 wl_63 vdd gnd cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd cell_6t
Xbit_r1_c196 bl_196 br_196 wl_1 vdd gnd cell_6t
Xbit_r2_c196 bl_196 br_196 wl_2 vdd gnd cell_6t
Xbit_r3_c196 bl_196 br_196 wl_3 vdd gnd cell_6t
Xbit_r4_c196 bl_196 br_196 wl_4 vdd gnd cell_6t
Xbit_r5_c196 bl_196 br_196 wl_5 vdd gnd cell_6t
Xbit_r6_c196 bl_196 br_196 wl_6 vdd gnd cell_6t
Xbit_r7_c196 bl_196 br_196 wl_7 vdd gnd cell_6t
Xbit_r8_c196 bl_196 br_196 wl_8 vdd gnd cell_6t
Xbit_r9_c196 bl_196 br_196 wl_9 vdd gnd cell_6t
Xbit_r10_c196 bl_196 br_196 wl_10 vdd gnd cell_6t
Xbit_r11_c196 bl_196 br_196 wl_11 vdd gnd cell_6t
Xbit_r12_c196 bl_196 br_196 wl_12 vdd gnd cell_6t
Xbit_r13_c196 bl_196 br_196 wl_13 vdd gnd cell_6t
Xbit_r14_c196 bl_196 br_196 wl_14 vdd gnd cell_6t
Xbit_r15_c196 bl_196 br_196 wl_15 vdd gnd cell_6t
Xbit_r16_c196 bl_196 br_196 wl_16 vdd gnd cell_6t
Xbit_r17_c196 bl_196 br_196 wl_17 vdd gnd cell_6t
Xbit_r18_c196 bl_196 br_196 wl_18 vdd gnd cell_6t
Xbit_r19_c196 bl_196 br_196 wl_19 vdd gnd cell_6t
Xbit_r20_c196 bl_196 br_196 wl_20 vdd gnd cell_6t
Xbit_r21_c196 bl_196 br_196 wl_21 vdd gnd cell_6t
Xbit_r22_c196 bl_196 br_196 wl_22 vdd gnd cell_6t
Xbit_r23_c196 bl_196 br_196 wl_23 vdd gnd cell_6t
Xbit_r24_c196 bl_196 br_196 wl_24 vdd gnd cell_6t
Xbit_r25_c196 bl_196 br_196 wl_25 vdd gnd cell_6t
Xbit_r26_c196 bl_196 br_196 wl_26 vdd gnd cell_6t
Xbit_r27_c196 bl_196 br_196 wl_27 vdd gnd cell_6t
Xbit_r28_c196 bl_196 br_196 wl_28 vdd gnd cell_6t
Xbit_r29_c196 bl_196 br_196 wl_29 vdd gnd cell_6t
Xbit_r30_c196 bl_196 br_196 wl_30 vdd gnd cell_6t
Xbit_r31_c196 bl_196 br_196 wl_31 vdd gnd cell_6t
Xbit_r32_c196 bl_196 br_196 wl_32 vdd gnd cell_6t
Xbit_r33_c196 bl_196 br_196 wl_33 vdd gnd cell_6t
Xbit_r34_c196 bl_196 br_196 wl_34 vdd gnd cell_6t
Xbit_r35_c196 bl_196 br_196 wl_35 vdd gnd cell_6t
Xbit_r36_c196 bl_196 br_196 wl_36 vdd gnd cell_6t
Xbit_r37_c196 bl_196 br_196 wl_37 vdd gnd cell_6t
Xbit_r38_c196 bl_196 br_196 wl_38 vdd gnd cell_6t
Xbit_r39_c196 bl_196 br_196 wl_39 vdd gnd cell_6t
Xbit_r40_c196 bl_196 br_196 wl_40 vdd gnd cell_6t
Xbit_r41_c196 bl_196 br_196 wl_41 vdd gnd cell_6t
Xbit_r42_c196 bl_196 br_196 wl_42 vdd gnd cell_6t
Xbit_r43_c196 bl_196 br_196 wl_43 vdd gnd cell_6t
Xbit_r44_c196 bl_196 br_196 wl_44 vdd gnd cell_6t
Xbit_r45_c196 bl_196 br_196 wl_45 vdd gnd cell_6t
Xbit_r46_c196 bl_196 br_196 wl_46 vdd gnd cell_6t
Xbit_r47_c196 bl_196 br_196 wl_47 vdd gnd cell_6t
Xbit_r48_c196 bl_196 br_196 wl_48 vdd gnd cell_6t
Xbit_r49_c196 bl_196 br_196 wl_49 vdd gnd cell_6t
Xbit_r50_c196 bl_196 br_196 wl_50 vdd gnd cell_6t
Xbit_r51_c196 bl_196 br_196 wl_51 vdd gnd cell_6t
Xbit_r52_c196 bl_196 br_196 wl_52 vdd gnd cell_6t
Xbit_r53_c196 bl_196 br_196 wl_53 vdd gnd cell_6t
Xbit_r54_c196 bl_196 br_196 wl_54 vdd gnd cell_6t
Xbit_r55_c196 bl_196 br_196 wl_55 vdd gnd cell_6t
Xbit_r56_c196 bl_196 br_196 wl_56 vdd gnd cell_6t
Xbit_r57_c196 bl_196 br_196 wl_57 vdd gnd cell_6t
Xbit_r58_c196 bl_196 br_196 wl_58 vdd gnd cell_6t
Xbit_r59_c196 bl_196 br_196 wl_59 vdd gnd cell_6t
Xbit_r60_c196 bl_196 br_196 wl_60 vdd gnd cell_6t
Xbit_r61_c196 bl_196 br_196 wl_61 vdd gnd cell_6t
Xbit_r62_c196 bl_196 br_196 wl_62 vdd gnd cell_6t
Xbit_r63_c196 bl_196 br_196 wl_63 vdd gnd cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd cell_6t
Xbit_r1_c197 bl_197 br_197 wl_1 vdd gnd cell_6t
Xbit_r2_c197 bl_197 br_197 wl_2 vdd gnd cell_6t
Xbit_r3_c197 bl_197 br_197 wl_3 vdd gnd cell_6t
Xbit_r4_c197 bl_197 br_197 wl_4 vdd gnd cell_6t
Xbit_r5_c197 bl_197 br_197 wl_5 vdd gnd cell_6t
Xbit_r6_c197 bl_197 br_197 wl_6 vdd gnd cell_6t
Xbit_r7_c197 bl_197 br_197 wl_7 vdd gnd cell_6t
Xbit_r8_c197 bl_197 br_197 wl_8 vdd gnd cell_6t
Xbit_r9_c197 bl_197 br_197 wl_9 vdd gnd cell_6t
Xbit_r10_c197 bl_197 br_197 wl_10 vdd gnd cell_6t
Xbit_r11_c197 bl_197 br_197 wl_11 vdd gnd cell_6t
Xbit_r12_c197 bl_197 br_197 wl_12 vdd gnd cell_6t
Xbit_r13_c197 bl_197 br_197 wl_13 vdd gnd cell_6t
Xbit_r14_c197 bl_197 br_197 wl_14 vdd gnd cell_6t
Xbit_r15_c197 bl_197 br_197 wl_15 vdd gnd cell_6t
Xbit_r16_c197 bl_197 br_197 wl_16 vdd gnd cell_6t
Xbit_r17_c197 bl_197 br_197 wl_17 vdd gnd cell_6t
Xbit_r18_c197 bl_197 br_197 wl_18 vdd gnd cell_6t
Xbit_r19_c197 bl_197 br_197 wl_19 vdd gnd cell_6t
Xbit_r20_c197 bl_197 br_197 wl_20 vdd gnd cell_6t
Xbit_r21_c197 bl_197 br_197 wl_21 vdd gnd cell_6t
Xbit_r22_c197 bl_197 br_197 wl_22 vdd gnd cell_6t
Xbit_r23_c197 bl_197 br_197 wl_23 vdd gnd cell_6t
Xbit_r24_c197 bl_197 br_197 wl_24 vdd gnd cell_6t
Xbit_r25_c197 bl_197 br_197 wl_25 vdd gnd cell_6t
Xbit_r26_c197 bl_197 br_197 wl_26 vdd gnd cell_6t
Xbit_r27_c197 bl_197 br_197 wl_27 vdd gnd cell_6t
Xbit_r28_c197 bl_197 br_197 wl_28 vdd gnd cell_6t
Xbit_r29_c197 bl_197 br_197 wl_29 vdd gnd cell_6t
Xbit_r30_c197 bl_197 br_197 wl_30 vdd gnd cell_6t
Xbit_r31_c197 bl_197 br_197 wl_31 vdd gnd cell_6t
Xbit_r32_c197 bl_197 br_197 wl_32 vdd gnd cell_6t
Xbit_r33_c197 bl_197 br_197 wl_33 vdd gnd cell_6t
Xbit_r34_c197 bl_197 br_197 wl_34 vdd gnd cell_6t
Xbit_r35_c197 bl_197 br_197 wl_35 vdd gnd cell_6t
Xbit_r36_c197 bl_197 br_197 wl_36 vdd gnd cell_6t
Xbit_r37_c197 bl_197 br_197 wl_37 vdd gnd cell_6t
Xbit_r38_c197 bl_197 br_197 wl_38 vdd gnd cell_6t
Xbit_r39_c197 bl_197 br_197 wl_39 vdd gnd cell_6t
Xbit_r40_c197 bl_197 br_197 wl_40 vdd gnd cell_6t
Xbit_r41_c197 bl_197 br_197 wl_41 vdd gnd cell_6t
Xbit_r42_c197 bl_197 br_197 wl_42 vdd gnd cell_6t
Xbit_r43_c197 bl_197 br_197 wl_43 vdd gnd cell_6t
Xbit_r44_c197 bl_197 br_197 wl_44 vdd gnd cell_6t
Xbit_r45_c197 bl_197 br_197 wl_45 vdd gnd cell_6t
Xbit_r46_c197 bl_197 br_197 wl_46 vdd gnd cell_6t
Xbit_r47_c197 bl_197 br_197 wl_47 vdd gnd cell_6t
Xbit_r48_c197 bl_197 br_197 wl_48 vdd gnd cell_6t
Xbit_r49_c197 bl_197 br_197 wl_49 vdd gnd cell_6t
Xbit_r50_c197 bl_197 br_197 wl_50 vdd gnd cell_6t
Xbit_r51_c197 bl_197 br_197 wl_51 vdd gnd cell_6t
Xbit_r52_c197 bl_197 br_197 wl_52 vdd gnd cell_6t
Xbit_r53_c197 bl_197 br_197 wl_53 vdd gnd cell_6t
Xbit_r54_c197 bl_197 br_197 wl_54 vdd gnd cell_6t
Xbit_r55_c197 bl_197 br_197 wl_55 vdd gnd cell_6t
Xbit_r56_c197 bl_197 br_197 wl_56 vdd gnd cell_6t
Xbit_r57_c197 bl_197 br_197 wl_57 vdd gnd cell_6t
Xbit_r58_c197 bl_197 br_197 wl_58 vdd gnd cell_6t
Xbit_r59_c197 bl_197 br_197 wl_59 vdd gnd cell_6t
Xbit_r60_c197 bl_197 br_197 wl_60 vdd gnd cell_6t
Xbit_r61_c197 bl_197 br_197 wl_61 vdd gnd cell_6t
Xbit_r62_c197 bl_197 br_197 wl_62 vdd gnd cell_6t
Xbit_r63_c197 bl_197 br_197 wl_63 vdd gnd cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd cell_6t
Xbit_r1_c198 bl_198 br_198 wl_1 vdd gnd cell_6t
Xbit_r2_c198 bl_198 br_198 wl_2 vdd gnd cell_6t
Xbit_r3_c198 bl_198 br_198 wl_3 vdd gnd cell_6t
Xbit_r4_c198 bl_198 br_198 wl_4 vdd gnd cell_6t
Xbit_r5_c198 bl_198 br_198 wl_5 vdd gnd cell_6t
Xbit_r6_c198 bl_198 br_198 wl_6 vdd gnd cell_6t
Xbit_r7_c198 bl_198 br_198 wl_7 vdd gnd cell_6t
Xbit_r8_c198 bl_198 br_198 wl_8 vdd gnd cell_6t
Xbit_r9_c198 bl_198 br_198 wl_9 vdd gnd cell_6t
Xbit_r10_c198 bl_198 br_198 wl_10 vdd gnd cell_6t
Xbit_r11_c198 bl_198 br_198 wl_11 vdd gnd cell_6t
Xbit_r12_c198 bl_198 br_198 wl_12 vdd gnd cell_6t
Xbit_r13_c198 bl_198 br_198 wl_13 vdd gnd cell_6t
Xbit_r14_c198 bl_198 br_198 wl_14 vdd gnd cell_6t
Xbit_r15_c198 bl_198 br_198 wl_15 vdd gnd cell_6t
Xbit_r16_c198 bl_198 br_198 wl_16 vdd gnd cell_6t
Xbit_r17_c198 bl_198 br_198 wl_17 vdd gnd cell_6t
Xbit_r18_c198 bl_198 br_198 wl_18 vdd gnd cell_6t
Xbit_r19_c198 bl_198 br_198 wl_19 vdd gnd cell_6t
Xbit_r20_c198 bl_198 br_198 wl_20 vdd gnd cell_6t
Xbit_r21_c198 bl_198 br_198 wl_21 vdd gnd cell_6t
Xbit_r22_c198 bl_198 br_198 wl_22 vdd gnd cell_6t
Xbit_r23_c198 bl_198 br_198 wl_23 vdd gnd cell_6t
Xbit_r24_c198 bl_198 br_198 wl_24 vdd gnd cell_6t
Xbit_r25_c198 bl_198 br_198 wl_25 vdd gnd cell_6t
Xbit_r26_c198 bl_198 br_198 wl_26 vdd gnd cell_6t
Xbit_r27_c198 bl_198 br_198 wl_27 vdd gnd cell_6t
Xbit_r28_c198 bl_198 br_198 wl_28 vdd gnd cell_6t
Xbit_r29_c198 bl_198 br_198 wl_29 vdd gnd cell_6t
Xbit_r30_c198 bl_198 br_198 wl_30 vdd gnd cell_6t
Xbit_r31_c198 bl_198 br_198 wl_31 vdd gnd cell_6t
Xbit_r32_c198 bl_198 br_198 wl_32 vdd gnd cell_6t
Xbit_r33_c198 bl_198 br_198 wl_33 vdd gnd cell_6t
Xbit_r34_c198 bl_198 br_198 wl_34 vdd gnd cell_6t
Xbit_r35_c198 bl_198 br_198 wl_35 vdd gnd cell_6t
Xbit_r36_c198 bl_198 br_198 wl_36 vdd gnd cell_6t
Xbit_r37_c198 bl_198 br_198 wl_37 vdd gnd cell_6t
Xbit_r38_c198 bl_198 br_198 wl_38 vdd gnd cell_6t
Xbit_r39_c198 bl_198 br_198 wl_39 vdd gnd cell_6t
Xbit_r40_c198 bl_198 br_198 wl_40 vdd gnd cell_6t
Xbit_r41_c198 bl_198 br_198 wl_41 vdd gnd cell_6t
Xbit_r42_c198 bl_198 br_198 wl_42 vdd gnd cell_6t
Xbit_r43_c198 bl_198 br_198 wl_43 vdd gnd cell_6t
Xbit_r44_c198 bl_198 br_198 wl_44 vdd gnd cell_6t
Xbit_r45_c198 bl_198 br_198 wl_45 vdd gnd cell_6t
Xbit_r46_c198 bl_198 br_198 wl_46 vdd gnd cell_6t
Xbit_r47_c198 bl_198 br_198 wl_47 vdd gnd cell_6t
Xbit_r48_c198 bl_198 br_198 wl_48 vdd gnd cell_6t
Xbit_r49_c198 bl_198 br_198 wl_49 vdd gnd cell_6t
Xbit_r50_c198 bl_198 br_198 wl_50 vdd gnd cell_6t
Xbit_r51_c198 bl_198 br_198 wl_51 vdd gnd cell_6t
Xbit_r52_c198 bl_198 br_198 wl_52 vdd gnd cell_6t
Xbit_r53_c198 bl_198 br_198 wl_53 vdd gnd cell_6t
Xbit_r54_c198 bl_198 br_198 wl_54 vdd gnd cell_6t
Xbit_r55_c198 bl_198 br_198 wl_55 vdd gnd cell_6t
Xbit_r56_c198 bl_198 br_198 wl_56 vdd gnd cell_6t
Xbit_r57_c198 bl_198 br_198 wl_57 vdd gnd cell_6t
Xbit_r58_c198 bl_198 br_198 wl_58 vdd gnd cell_6t
Xbit_r59_c198 bl_198 br_198 wl_59 vdd gnd cell_6t
Xbit_r60_c198 bl_198 br_198 wl_60 vdd gnd cell_6t
Xbit_r61_c198 bl_198 br_198 wl_61 vdd gnd cell_6t
Xbit_r62_c198 bl_198 br_198 wl_62 vdd gnd cell_6t
Xbit_r63_c198 bl_198 br_198 wl_63 vdd gnd cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd cell_6t
Xbit_r1_c199 bl_199 br_199 wl_1 vdd gnd cell_6t
Xbit_r2_c199 bl_199 br_199 wl_2 vdd gnd cell_6t
Xbit_r3_c199 bl_199 br_199 wl_3 vdd gnd cell_6t
Xbit_r4_c199 bl_199 br_199 wl_4 vdd gnd cell_6t
Xbit_r5_c199 bl_199 br_199 wl_5 vdd gnd cell_6t
Xbit_r6_c199 bl_199 br_199 wl_6 vdd gnd cell_6t
Xbit_r7_c199 bl_199 br_199 wl_7 vdd gnd cell_6t
Xbit_r8_c199 bl_199 br_199 wl_8 vdd gnd cell_6t
Xbit_r9_c199 bl_199 br_199 wl_9 vdd gnd cell_6t
Xbit_r10_c199 bl_199 br_199 wl_10 vdd gnd cell_6t
Xbit_r11_c199 bl_199 br_199 wl_11 vdd gnd cell_6t
Xbit_r12_c199 bl_199 br_199 wl_12 vdd gnd cell_6t
Xbit_r13_c199 bl_199 br_199 wl_13 vdd gnd cell_6t
Xbit_r14_c199 bl_199 br_199 wl_14 vdd gnd cell_6t
Xbit_r15_c199 bl_199 br_199 wl_15 vdd gnd cell_6t
Xbit_r16_c199 bl_199 br_199 wl_16 vdd gnd cell_6t
Xbit_r17_c199 bl_199 br_199 wl_17 vdd gnd cell_6t
Xbit_r18_c199 bl_199 br_199 wl_18 vdd gnd cell_6t
Xbit_r19_c199 bl_199 br_199 wl_19 vdd gnd cell_6t
Xbit_r20_c199 bl_199 br_199 wl_20 vdd gnd cell_6t
Xbit_r21_c199 bl_199 br_199 wl_21 vdd gnd cell_6t
Xbit_r22_c199 bl_199 br_199 wl_22 vdd gnd cell_6t
Xbit_r23_c199 bl_199 br_199 wl_23 vdd gnd cell_6t
Xbit_r24_c199 bl_199 br_199 wl_24 vdd gnd cell_6t
Xbit_r25_c199 bl_199 br_199 wl_25 vdd gnd cell_6t
Xbit_r26_c199 bl_199 br_199 wl_26 vdd gnd cell_6t
Xbit_r27_c199 bl_199 br_199 wl_27 vdd gnd cell_6t
Xbit_r28_c199 bl_199 br_199 wl_28 vdd gnd cell_6t
Xbit_r29_c199 bl_199 br_199 wl_29 vdd gnd cell_6t
Xbit_r30_c199 bl_199 br_199 wl_30 vdd gnd cell_6t
Xbit_r31_c199 bl_199 br_199 wl_31 vdd gnd cell_6t
Xbit_r32_c199 bl_199 br_199 wl_32 vdd gnd cell_6t
Xbit_r33_c199 bl_199 br_199 wl_33 vdd gnd cell_6t
Xbit_r34_c199 bl_199 br_199 wl_34 vdd gnd cell_6t
Xbit_r35_c199 bl_199 br_199 wl_35 vdd gnd cell_6t
Xbit_r36_c199 bl_199 br_199 wl_36 vdd gnd cell_6t
Xbit_r37_c199 bl_199 br_199 wl_37 vdd gnd cell_6t
Xbit_r38_c199 bl_199 br_199 wl_38 vdd gnd cell_6t
Xbit_r39_c199 bl_199 br_199 wl_39 vdd gnd cell_6t
Xbit_r40_c199 bl_199 br_199 wl_40 vdd gnd cell_6t
Xbit_r41_c199 bl_199 br_199 wl_41 vdd gnd cell_6t
Xbit_r42_c199 bl_199 br_199 wl_42 vdd gnd cell_6t
Xbit_r43_c199 bl_199 br_199 wl_43 vdd gnd cell_6t
Xbit_r44_c199 bl_199 br_199 wl_44 vdd gnd cell_6t
Xbit_r45_c199 bl_199 br_199 wl_45 vdd gnd cell_6t
Xbit_r46_c199 bl_199 br_199 wl_46 vdd gnd cell_6t
Xbit_r47_c199 bl_199 br_199 wl_47 vdd gnd cell_6t
Xbit_r48_c199 bl_199 br_199 wl_48 vdd gnd cell_6t
Xbit_r49_c199 bl_199 br_199 wl_49 vdd gnd cell_6t
Xbit_r50_c199 bl_199 br_199 wl_50 vdd gnd cell_6t
Xbit_r51_c199 bl_199 br_199 wl_51 vdd gnd cell_6t
Xbit_r52_c199 bl_199 br_199 wl_52 vdd gnd cell_6t
Xbit_r53_c199 bl_199 br_199 wl_53 vdd gnd cell_6t
Xbit_r54_c199 bl_199 br_199 wl_54 vdd gnd cell_6t
Xbit_r55_c199 bl_199 br_199 wl_55 vdd gnd cell_6t
Xbit_r56_c199 bl_199 br_199 wl_56 vdd gnd cell_6t
Xbit_r57_c199 bl_199 br_199 wl_57 vdd gnd cell_6t
Xbit_r58_c199 bl_199 br_199 wl_58 vdd gnd cell_6t
Xbit_r59_c199 bl_199 br_199 wl_59 vdd gnd cell_6t
Xbit_r60_c199 bl_199 br_199 wl_60 vdd gnd cell_6t
Xbit_r61_c199 bl_199 br_199 wl_61 vdd gnd cell_6t
Xbit_r62_c199 bl_199 br_199 wl_62 vdd gnd cell_6t
Xbit_r63_c199 bl_199 br_199 wl_63 vdd gnd cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd cell_6t
Xbit_r1_c200 bl_200 br_200 wl_1 vdd gnd cell_6t
Xbit_r2_c200 bl_200 br_200 wl_2 vdd gnd cell_6t
Xbit_r3_c200 bl_200 br_200 wl_3 vdd gnd cell_6t
Xbit_r4_c200 bl_200 br_200 wl_4 vdd gnd cell_6t
Xbit_r5_c200 bl_200 br_200 wl_5 vdd gnd cell_6t
Xbit_r6_c200 bl_200 br_200 wl_6 vdd gnd cell_6t
Xbit_r7_c200 bl_200 br_200 wl_7 vdd gnd cell_6t
Xbit_r8_c200 bl_200 br_200 wl_8 vdd gnd cell_6t
Xbit_r9_c200 bl_200 br_200 wl_9 vdd gnd cell_6t
Xbit_r10_c200 bl_200 br_200 wl_10 vdd gnd cell_6t
Xbit_r11_c200 bl_200 br_200 wl_11 vdd gnd cell_6t
Xbit_r12_c200 bl_200 br_200 wl_12 vdd gnd cell_6t
Xbit_r13_c200 bl_200 br_200 wl_13 vdd gnd cell_6t
Xbit_r14_c200 bl_200 br_200 wl_14 vdd gnd cell_6t
Xbit_r15_c200 bl_200 br_200 wl_15 vdd gnd cell_6t
Xbit_r16_c200 bl_200 br_200 wl_16 vdd gnd cell_6t
Xbit_r17_c200 bl_200 br_200 wl_17 vdd gnd cell_6t
Xbit_r18_c200 bl_200 br_200 wl_18 vdd gnd cell_6t
Xbit_r19_c200 bl_200 br_200 wl_19 vdd gnd cell_6t
Xbit_r20_c200 bl_200 br_200 wl_20 vdd gnd cell_6t
Xbit_r21_c200 bl_200 br_200 wl_21 vdd gnd cell_6t
Xbit_r22_c200 bl_200 br_200 wl_22 vdd gnd cell_6t
Xbit_r23_c200 bl_200 br_200 wl_23 vdd gnd cell_6t
Xbit_r24_c200 bl_200 br_200 wl_24 vdd gnd cell_6t
Xbit_r25_c200 bl_200 br_200 wl_25 vdd gnd cell_6t
Xbit_r26_c200 bl_200 br_200 wl_26 vdd gnd cell_6t
Xbit_r27_c200 bl_200 br_200 wl_27 vdd gnd cell_6t
Xbit_r28_c200 bl_200 br_200 wl_28 vdd gnd cell_6t
Xbit_r29_c200 bl_200 br_200 wl_29 vdd gnd cell_6t
Xbit_r30_c200 bl_200 br_200 wl_30 vdd gnd cell_6t
Xbit_r31_c200 bl_200 br_200 wl_31 vdd gnd cell_6t
Xbit_r32_c200 bl_200 br_200 wl_32 vdd gnd cell_6t
Xbit_r33_c200 bl_200 br_200 wl_33 vdd gnd cell_6t
Xbit_r34_c200 bl_200 br_200 wl_34 vdd gnd cell_6t
Xbit_r35_c200 bl_200 br_200 wl_35 vdd gnd cell_6t
Xbit_r36_c200 bl_200 br_200 wl_36 vdd gnd cell_6t
Xbit_r37_c200 bl_200 br_200 wl_37 vdd gnd cell_6t
Xbit_r38_c200 bl_200 br_200 wl_38 vdd gnd cell_6t
Xbit_r39_c200 bl_200 br_200 wl_39 vdd gnd cell_6t
Xbit_r40_c200 bl_200 br_200 wl_40 vdd gnd cell_6t
Xbit_r41_c200 bl_200 br_200 wl_41 vdd gnd cell_6t
Xbit_r42_c200 bl_200 br_200 wl_42 vdd gnd cell_6t
Xbit_r43_c200 bl_200 br_200 wl_43 vdd gnd cell_6t
Xbit_r44_c200 bl_200 br_200 wl_44 vdd gnd cell_6t
Xbit_r45_c200 bl_200 br_200 wl_45 vdd gnd cell_6t
Xbit_r46_c200 bl_200 br_200 wl_46 vdd gnd cell_6t
Xbit_r47_c200 bl_200 br_200 wl_47 vdd gnd cell_6t
Xbit_r48_c200 bl_200 br_200 wl_48 vdd gnd cell_6t
Xbit_r49_c200 bl_200 br_200 wl_49 vdd gnd cell_6t
Xbit_r50_c200 bl_200 br_200 wl_50 vdd gnd cell_6t
Xbit_r51_c200 bl_200 br_200 wl_51 vdd gnd cell_6t
Xbit_r52_c200 bl_200 br_200 wl_52 vdd gnd cell_6t
Xbit_r53_c200 bl_200 br_200 wl_53 vdd gnd cell_6t
Xbit_r54_c200 bl_200 br_200 wl_54 vdd gnd cell_6t
Xbit_r55_c200 bl_200 br_200 wl_55 vdd gnd cell_6t
Xbit_r56_c200 bl_200 br_200 wl_56 vdd gnd cell_6t
Xbit_r57_c200 bl_200 br_200 wl_57 vdd gnd cell_6t
Xbit_r58_c200 bl_200 br_200 wl_58 vdd gnd cell_6t
Xbit_r59_c200 bl_200 br_200 wl_59 vdd gnd cell_6t
Xbit_r60_c200 bl_200 br_200 wl_60 vdd gnd cell_6t
Xbit_r61_c200 bl_200 br_200 wl_61 vdd gnd cell_6t
Xbit_r62_c200 bl_200 br_200 wl_62 vdd gnd cell_6t
Xbit_r63_c200 bl_200 br_200 wl_63 vdd gnd cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd cell_6t
Xbit_r1_c201 bl_201 br_201 wl_1 vdd gnd cell_6t
Xbit_r2_c201 bl_201 br_201 wl_2 vdd gnd cell_6t
Xbit_r3_c201 bl_201 br_201 wl_3 vdd gnd cell_6t
Xbit_r4_c201 bl_201 br_201 wl_4 vdd gnd cell_6t
Xbit_r5_c201 bl_201 br_201 wl_5 vdd gnd cell_6t
Xbit_r6_c201 bl_201 br_201 wl_6 vdd gnd cell_6t
Xbit_r7_c201 bl_201 br_201 wl_7 vdd gnd cell_6t
Xbit_r8_c201 bl_201 br_201 wl_8 vdd gnd cell_6t
Xbit_r9_c201 bl_201 br_201 wl_9 vdd gnd cell_6t
Xbit_r10_c201 bl_201 br_201 wl_10 vdd gnd cell_6t
Xbit_r11_c201 bl_201 br_201 wl_11 vdd gnd cell_6t
Xbit_r12_c201 bl_201 br_201 wl_12 vdd gnd cell_6t
Xbit_r13_c201 bl_201 br_201 wl_13 vdd gnd cell_6t
Xbit_r14_c201 bl_201 br_201 wl_14 vdd gnd cell_6t
Xbit_r15_c201 bl_201 br_201 wl_15 vdd gnd cell_6t
Xbit_r16_c201 bl_201 br_201 wl_16 vdd gnd cell_6t
Xbit_r17_c201 bl_201 br_201 wl_17 vdd gnd cell_6t
Xbit_r18_c201 bl_201 br_201 wl_18 vdd gnd cell_6t
Xbit_r19_c201 bl_201 br_201 wl_19 vdd gnd cell_6t
Xbit_r20_c201 bl_201 br_201 wl_20 vdd gnd cell_6t
Xbit_r21_c201 bl_201 br_201 wl_21 vdd gnd cell_6t
Xbit_r22_c201 bl_201 br_201 wl_22 vdd gnd cell_6t
Xbit_r23_c201 bl_201 br_201 wl_23 vdd gnd cell_6t
Xbit_r24_c201 bl_201 br_201 wl_24 vdd gnd cell_6t
Xbit_r25_c201 bl_201 br_201 wl_25 vdd gnd cell_6t
Xbit_r26_c201 bl_201 br_201 wl_26 vdd gnd cell_6t
Xbit_r27_c201 bl_201 br_201 wl_27 vdd gnd cell_6t
Xbit_r28_c201 bl_201 br_201 wl_28 vdd gnd cell_6t
Xbit_r29_c201 bl_201 br_201 wl_29 vdd gnd cell_6t
Xbit_r30_c201 bl_201 br_201 wl_30 vdd gnd cell_6t
Xbit_r31_c201 bl_201 br_201 wl_31 vdd gnd cell_6t
Xbit_r32_c201 bl_201 br_201 wl_32 vdd gnd cell_6t
Xbit_r33_c201 bl_201 br_201 wl_33 vdd gnd cell_6t
Xbit_r34_c201 bl_201 br_201 wl_34 vdd gnd cell_6t
Xbit_r35_c201 bl_201 br_201 wl_35 vdd gnd cell_6t
Xbit_r36_c201 bl_201 br_201 wl_36 vdd gnd cell_6t
Xbit_r37_c201 bl_201 br_201 wl_37 vdd gnd cell_6t
Xbit_r38_c201 bl_201 br_201 wl_38 vdd gnd cell_6t
Xbit_r39_c201 bl_201 br_201 wl_39 vdd gnd cell_6t
Xbit_r40_c201 bl_201 br_201 wl_40 vdd gnd cell_6t
Xbit_r41_c201 bl_201 br_201 wl_41 vdd gnd cell_6t
Xbit_r42_c201 bl_201 br_201 wl_42 vdd gnd cell_6t
Xbit_r43_c201 bl_201 br_201 wl_43 vdd gnd cell_6t
Xbit_r44_c201 bl_201 br_201 wl_44 vdd gnd cell_6t
Xbit_r45_c201 bl_201 br_201 wl_45 vdd gnd cell_6t
Xbit_r46_c201 bl_201 br_201 wl_46 vdd gnd cell_6t
Xbit_r47_c201 bl_201 br_201 wl_47 vdd gnd cell_6t
Xbit_r48_c201 bl_201 br_201 wl_48 vdd gnd cell_6t
Xbit_r49_c201 bl_201 br_201 wl_49 vdd gnd cell_6t
Xbit_r50_c201 bl_201 br_201 wl_50 vdd gnd cell_6t
Xbit_r51_c201 bl_201 br_201 wl_51 vdd gnd cell_6t
Xbit_r52_c201 bl_201 br_201 wl_52 vdd gnd cell_6t
Xbit_r53_c201 bl_201 br_201 wl_53 vdd gnd cell_6t
Xbit_r54_c201 bl_201 br_201 wl_54 vdd gnd cell_6t
Xbit_r55_c201 bl_201 br_201 wl_55 vdd gnd cell_6t
Xbit_r56_c201 bl_201 br_201 wl_56 vdd gnd cell_6t
Xbit_r57_c201 bl_201 br_201 wl_57 vdd gnd cell_6t
Xbit_r58_c201 bl_201 br_201 wl_58 vdd gnd cell_6t
Xbit_r59_c201 bl_201 br_201 wl_59 vdd gnd cell_6t
Xbit_r60_c201 bl_201 br_201 wl_60 vdd gnd cell_6t
Xbit_r61_c201 bl_201 br_201 wl_61 vdd gnd cell_6t
Xbit_r62_c201 bl_201 br_201 wl_62 vdd gnd cell_6t
Xbit_r63_c201 bl_201 br_201 wl_63 vdd gnd cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd cell_6t
Xbit_r1_c202 bl_202 br_202 wl_1 vdd gnd cell_6t
Xbit_r2_c202 bl_202 br_202 wl_2 vdd gnd cell_6t
Xbit_r3_c202 bl_202 br_202 wl_3 vdd gnd cell_6t
Xbit_r4_c202 bl_202 br_202 wl_4 vdd gnd cell_6t
Xbit_r5_c202 bl_202 br_202 wl_5 vdd gnd cell_6t
Xbit_r6_c202 bl_202 br_202 wl_6 vdd gnd cell_6t
Xbit_r7_c202 bl_202 br_202 wl_7 vdd gnd cell_6t
Xbit_r8_c202 bl_202 br_202 wl_8 vdd gnd cell_6t
Xbit_r9_c202 bl_202 br_202 wl_9 vdd gnd cell_6t
Xbit_r10_c202 bl_202 br_202 wl_10 vdd gnd cell_6t
Xbit_r11_c202 bl_202 br_202 wl_11 vdd gnd cell_6t
Xbit_r12_c202 bl_202 br_202 wl_12 vdd gnd cell_6t
Xbit_r13_c202 bl_202 br_202 wl_13 vdd gnd cell_6t
Xbit_r14_c202 bl_202 br_202 wl_14 vdd gnd cell_6t
Xbit_r15_c202 bl_202 br_202 wl_15 vdd gnd cell_6t
Xbit_r16_c202 bl_202 br_202 wl_16 vdd gnd cell_6t
Xbit_r17_c202 bl_202 br_202 wl_17 vdd gnd cell_6t
Xbit_r18_c202 bl_202 br_202 wl_18 vdd gnd cell_6t
Xbit_r19_c202 bl_202 br_202 wl_19 vdd gnd cell_6t
Xbit_r20_c202 bl_202 br_202 wl_20 vdd gnd cell_6t
Xbit_r21_c202 bl_202 br_202 wl_21 vdd gnd cell_6t
Xbit_r22_c202 bl_202 br_202 wl_22 vdd gnd cell_6t
Xbit_r23_c202 bl_202 br_202 wl_23 vdd gnd cell_6t
Xbit_r24_c202 bl_202 br_202 wl_24 vdd gnd cell_6t
Xbit_r25_c202 bl_202 br_202 wl_25 vdd gnd cell_6t
Xbit_r26_c202 bl_202 br_202 wl_26 vdd gnd cell_6t
Xbit_r27_c202 bl_202 br_202 wl_27 vdd gnd cell_6t
Xbit_r28_c202 bl_202 br_202 wl_28 vdd gnd cell_6t
Xbit_r29_c202 bl_202 br_202 wl_29 vdd gnd cell_6t
Xbit_r30_c202 bl_202 br_202 wl_30 vdd gnd cell_6t
Xbit_r31_c202 bl_202 br_202 wl_31 vdd gnd cell_6t
Xbit_r32_c202 bl_202 br_202 wl_32 vdd gnd cell_6t
Xbit_r33_c202 bl_202 br_202 wl_33 vdd gnd cell_6t
Xbit_r34_c202 bl_202 br_202 wl_34 vdd gnd cell_6t
Xbit_r35_c202 bl_202 br_202 wl_35 vdd gnd cell_6t
Xbit_r36_c202 bl_202 br_202 wl_36 vdd gnd cell_6t
Xbit_r37_c202 bl_202 br_202 wl_37 vdd gnd cell_6t
Xbit_r38_c202 bl_202 br_202 wl_38 vdd gnd cell_6t
Xbit_r39_c202 bl_202 br_202 wl_39 vdd gnd cell_6t
Xbit_r40_c202 bl_202 br_202 wl_40 vdd gnd cell_6t
Xbit_r41_c202 bl_202 br_202 wl_41 vdd gnd cell_6t
Xbit_r42_c202 bl_202 br_202 wl_42 vdd gnd cell_6t
Xbit_r43_c202 bl_202 br_202 wl_43 vdd gnd cell_6t
Xbit_r44_c202 bl_202 br_202 wl_44 vdd gnd cell_6t
Xbit_r45_c202 bl_202 br_202 wl_45 vdd gnd cell_6t
Xbit_r46_c202 bl_202 br_202 wl_46 vdd gnd cell_6t
Xbit_r47_c202 bl_202 br_202 wl_47 vdd gnd cell_6t
Xbit_r48_c202 bl_202 br_202 wl_48 vdd gnd cell_6t
Xbit_r49_c202 bl_202 br_202 wl_49 vdd gnd cell_6t
Xbit_r50_c202 bl_202 br_202 wl_50 vdd gnd cell_6t
Xbit_r51_c202 bl_202 br_202 wl_51 vdd gnd cell_6t
Xbit_r52_c202 bl_202 br_202 wl_52 vdd gnd cell_6t
Xbit_r53_c202 bl_202 br_202 wl_53 vdd gnd cell_6t
Xbit_r54_c202 bl_202 br_202 wl_54 vdd gnd cell_6t
Xbit_r55_c202 bl_202 br_202 wl_55 vdd gnd cell_6t
Xbit_r56_c202 bl_202 br_202 wl_56 vdd gnd cell_6t
Xbit_r57_c202 bl_202 br_202 wl_57 vdd gnd cell_6t
Xbit_r58_c202 bl_202 br_202 wl_58 vdd gnd cell_6t
Xbit_r59_c202 bl_202 br_202 wl_59 vdd gnd cell_6t
Xbit_r60_c202 bl_202 br_202 wl_60 vdd gnd cell_6t
Xbit_r61_c202 bl_202 br_202 wl_61 vdd gnd cell_6t
Xbit_r62_c202 bl_202 br_202 wl_62 vdd gnd cell_6t
Xbit_r63_c202 bl_202 br_202 wl_63 vdd gnd cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd cell_6t
Xbit_r1_c203 bl_203 br_203 wl_1 vdd gnd cell_6t
Xbit_r2_c203 bl_203 br_203 wl_2 vdd gnd cell_6t
Xbit_r3_c203 bl_203 br_203 wl_3 vdd gnd cell_6t
Xbit_r4_c203 bl_203 br_203 wl_4 vdd gnd cell_6t
Xbit_r5_c203 bl_203 br_203 wl_5 vdd gnd cell_6t
Xbit_r6_c203 bl_203 br_203 wl_6 vdd gnd cell_6t
Xbit_r7_c203 bl_203 br_203 wl_7 vdd gnd cell_6t
Xbit_r8_c203 bl_203 br_203 wl_8 vdd gnd cell_6t
Xbit_r9_c203 bl_203 br_203 wl_9 vdd gnd cell_6t
Xbit_r10_c203 bl_203 br_203 wl_10 vdd gnd cell_6t
Xbit_r11_c203 bl_203 br_203 wl_11 vdd gnd cell_6t
Xbit_r12_c203 bl_203 br_203 wl_12 vdd gnd cell_6t
Xbit_r13_c203 bl_203 br_203 wl_13 vdd gnd cell_6t
Xbit_r14_c203 bl_203 br_203 wl_14 vdd gnd cell_6t
Xbit_r15_c203 bl_203 br_203 wl_15 vdd gnd cell_6t
Xbit_r16_c203 bl_203 br_203 wl_16 vdd gnd cell_6t
Xbit_r17_c203 bl_203 br_203 wl_17 vdd gnd cell_6t
Xbit_r18_c203 bl_203 br_203 wl_18 vdd gnd cell_6t
Xbit_r19_c203 bl_203 br_203 wl_19 vdd gnd cell_6t
Xbit_r20_c203 bl_203 br_203 wl_20 vdd gnd cell_6t
Xbit_r21_c203 bl_203 br_203 wl_21 vdd gnd cell_6t
Xbit_r22_c203 bl_203 br_203 wl_22 vdd gnd cell_6t
Xbit_r23_c203 bl_203 br_203 wl_23 vdd gnd cell_6t
Xbit_r24_c203 bl_203 br_203 wl_24 vdd gnd cell_6t
Xbit_r25_c203 bl_203 br_203 wl_25 vdd gnd cell_6t
Xbit_r26_c203 bl_203 br_203 wl_26 vdd gnd cell_6t
Xbit_r27_c203 bl_203 br_203 wl_27 vdd gnd cell_6t
Xbit_r28_c203 bl_203 br_203 wl_28 vdd gnd cell_6t
Xbit_r29_c203 bl_203 br_203 wl_29 vdd gnd cell_6t
Xbit_r30_c203 bl_203 br_203 wl_30 vdd gnd cell_6t
Xbit_r31_c203 bl_203 br_203 wl_31 vdd gnd cell_6t
Xbit_r32_c203 bl_203 br_203 wl_32 vdd gnd cell_6t
Xbit_r33_c203 bl_203 br_203 wl_33 vdd gnd cell_6t
Xbit_r34_c203 bl_203 br_203 wl_34 vdd gnd cell_6t
Xbit_r35_c203 bl_203 br_203 wl_35 vdd gnd cell_6t
Xbit_r36_c203 bl_203 br_203 wl_36 vdd gnd cell_6t
Xbit_r37_c203 bl_203 br_203 wl_37 vdd gnd cell_6t
Xbit_r38_c203 bl_203 br_203 wl_38 vdd gnd cell_6t
Xbit_r39_c203 bl_203 br_203 wl_39 vdd gnd cell_6t
Xbit_r40_c203 bl_203 br_203 wl_40 vdd gnd cell_6t
Xbit_r41_c203 bl_203 br_203 wl_41 vdd gnd cell_6t
Xbit_r42_c203 bl_203 br_203 wl_42 vdd gnd cell_6t
Xbit_r43_c203 bl_203 br_203 wl_43 vdd gnd cell_6t
Xbit_r44_c203 bl_203 br_203 wl_44 vdd gnd cell_6t
Xbit_r45_c203 bl_203 br_203 wl_45 vdd gnd cell_6t
Xbit_r46_c203 bl_203 br_203 wl_46 vdd gnd cell_6t
Xbit_r47_c203 bl_203 br_203 wl_47 vdd gnd cell_6t
Xbit_r48_c203 bl_203 br_203 wl_48 vdd gnd cell_6t
Xbit_r49_c203 bl_203 br_203 wl_49 vdd gnd cell_6t
Xbit_r50_c203 bl_203 br_203 wl_50 vdd gnd cell_6t
Xbit_r51_c203 bl_203 br_203 wl_51 vdd gnd cell_6t
Xbit_r52_c203 bl_203 br_203 wl_52 vdd gnd cell_6t
Xbit_r53_c203 bl_203 br_203 wl_53 vdd gnd cell_6t
Xbit_r54_c203 bl_203 br_203 wl_54 vdd gnd cell_6t
Xbit_r55_c203 bl_203 br_203 wl_55 vdd gnd cell_6t
Xbit_r56_c203 bl_203 br_203 wl_56 vdd gnd cell_6t
Xbit_r57_c203 bl_203 br_203 wl_57 vdd gnd cell_6t
Xbit_r58_c203 bl_203 br_203 wl_58 vdd gnd cell_6t
Xbit_r59_c203 bl_203 br_203 wl_59 vdd gnd cell_6t
Xbit_r60_c203 bl_203 br_203 wl_60 vdd gnd cell_6t
Xbit_r61_c203 bl_203 br_203 wl_61 vdd gnd cell_6t
Xbit_r62_c203 bl_203 br_203 wl_62 vdd gnd cell_6t
Xbit_r63_c203 bl_203 br_203 wl_63 vdd gnd cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd cell_6t
Xbit_r1_c204 bl_204 br_204 wl_1 vdd gnd cell_6t
Xbit_r2_c204 bl_204 br_204 wl_2 vdd gnd cell_6t
Xbit_r3_c204 bl_204 br_204 wl_3 vdd gnd cell_6t
Xbit_r4_c204 bl_204 br_204 wl_4 vdd gnd cell_6t
Xbit_r5_c204 bl_204 br_204 wl_5 vdd gnd cell_6t
Xbit_r6_c204 bl_204 br_204 wl_6 vdd gnd cell_6t
Xbit_r7_c204 bl_204 br_204 wl_7 vdd gnd cell_6t
Xbit_r8_c204 bl_204 br_204 wl_8 vdd gnd cell_6t
Xbit_r9_c204 bl_204 br_204 wl_9 vdd gnd cell_6t
Xbit_r10_c204 bl_204 br_204 wl_10 vdd gnd cell_6t
Xbit_r11_c204 bl_204 br_204 wl_11 vdd gnd cell_6t
Xbit_r12_c204 bl_204 br_204 wl_12 vdd gnd cell_6t
Xbit_r13_c204 bl_204 br_204 wl_13 vdd gnd cell_6t
Xbit_r14_c204 bl_204 br_204 wl_14 vdd gnd cell_6t
Xbit_r15_c204 bl_204 br_204 wl_15 vdd gnd cell_6t
Xbit_r16_c204 bl_204 br_204 wl_16 vdd gnd cell_6t
Xbit_r17_c204 bl_204 br_204 wl_17 vdd gnd cell_6t
Xbit_r18_c204 bl_204 br_204 wl_18 vdd gnd cell_6t
Xbit_r19_c204 bl_204 br_204 wl_19 vdd gnd cell_6t
Xbit_r20_c204 bl_204 br_204 wl_20 vdd gnd cell_6t
Xbit_r21_c204 bl_204 br_204 wl_21 vdd gnd cell_6t
Xbit_r22_c204 bl_204 br_204 wl_22 vdd gnd cell_6t
Xbit_r23_c204 bl_204 br_204 wl_23 vdd gnd cell_6t
Xbit_r24_c204 bl_204 br_204 wl_24 vdd gnd cell_6t
Xbit_r25_c204 bl_204 br_204 wl_25 vdd gnd cell_6t
Xbit_r26_c204 bl_204 br_204 wl_26 vdd gnd cell_6t
Xbit_r27_c204 bl_204 br_204 wl_27 vdd gnd cell_6t
Xbit_r28_c204 bl_204 br_204 wl_28 vdd gnd cell_6t
Xbit_r29_c204 bl_204 br_204 wl_29 vdd gnd cell_6t
Xbit_r30_c204 bl_204 br_204 wl_30 vdd gnd cell_6t
Xbit_r31_c204 bl_204 br_204 wl_31 vdd gnd cell_6t
Xbit_r32_c204 bl_204 br_204 wl_32 vdd gnd cell_6t
Xbit_r33_c204 bl_204 br_204 wl_33 vdd gnd cell_6t
Xbit_r34_c204 bl_204 br_204 wl_34 vdd gnd cell_6t
Xbit_r35_c204 bl_204 br_204 wl_35 vdd gnd cell_6t
Xbit_r36_c204 bl_204 br_204 wl_36 vdd gnd cell_6t
Xbit_r37_c204 bl_204 br_204 wl_37 vdd gnd cell_6t
Xbit_r38_c204 bl_204 br_204 wl_38 vdd gnd cell_6t
Xbit_r39_c204 bl_204 br_204 wl_39 vdd gnd cell_6t
Xbit_r40_c204 bl_204 br_204 wl_40 vdd gnd cell_6t
Xbit_r41_c204 bl_204 br_204 wl_41 vdd gnd cell_6t
Xbit_r42_c204 bl_204 br_204 wl_42 vdd gnd cell_6t
Xbit_r43_c204 bl_204 br_204 wl_43 vdd gnd cell_6t
Xbit_r44_c204 bl_204 br_204 wl_44 vdd gnd cell_6t
Xbit_r45_c204 bl_204 br_204 wl_45 vdd gnd cell_6t
Xbit_r46_c204 bl_204 br_204 wl_46 vdd gnd cell_6t
Xbit_r47_c204 bl_204 br_204 wl_47 vdd gnd cell_6t
Xbit_r48_c204 bl_204 br_204 wl_48 vdd gnd cell_6t
Xbit_r49_c204 bl_204 br_204 wl_49 vdd gnd cell_6t
Xbit_r50_c204 bl_204 br_204 wl_50 vdd gnd cell_6t
Xbit_r51_c204 bl_204 br_204 wl_51 vdd gnd cell_6t
Xbit_r52_c204 bl_204 br_204 wl_52 vdd gnd cell_6t
Xbit_r53_c204 bl_204 br_204 wl_53 vdd gnd cell_6t
Xbit_r54_c204 bl_204 br_204 wl_54 vdd gnd cell_6t
Xbit_r55_c204 bl_204 br_204 wl_55 vdd gnd cell_6t
Xbit_r56_c204 bl_204 br_204 wl_56 vdd gnd cell_6t
Xbit_r57_c204 bl_204 br_204 wl_57 vdd gnd cell_6t
Xbit_r58_c204 bl_204 br_204 wl_58 vdd gnd cell_6t
Xbit_r59_c204 bl_204 br_204 wl_59 vdd gnd cell_6t
Xbit_r60_c204 bl_204 br_204 wl_60 vdd gnd cell_6t
Xbit_r61_c204 bl_204 br_204 wl_61 vdd gnd cell_6t
Xbit_r62_c204 bl_204 br_204 wl_62 vdd gnd cell_6t
Xbit_r63_c204 bl_204 br_204 wl_63 vdd gnd cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd cell_6t
Xbit_r1_c205 bl_205 br_205 wl_1 vdd gnd cell_6t
Xbit_r2_c205 bl_205 br_205 wl_2 vdd gnd cell_6t
Xbit_r3_c205 bl_205 br_205 wl_3 vdd gnd cell_6t
Xbit_r4_c205 bl_205 br_205 wl_4 vdd gnd cell_6t
Xbit_r5_c205 bl_205 br_205 wl_5 vdd gnd cell_6t
Xbit_r6_c205 bl_205 br_205 wl_6 vdd gnd cell_6t
Xbit_r7_c205 bl_205 br_205 wl_7 vdd gnd cell_6t
Xbit_r8_c205 bl_205 br_205 wl_8 vdd gnd cell_6t
Xbit_r9_c205 bl_205 br_205 wl_9 vdd gnd cell_6t
Xbit_r10_c205 bl_205 br_205 wl_10 vdd gnd cell_6t
Xbit_r11_c205 bl_205 br_205 wl_11 vdd gnd cell_6t
Xbit_r12_c205 bl_205 br_205 wl_12 vdd gnd cell_6t
Xbit_r13_c205 bl_205 br_205 wl_13 vdd gnd cell_6t
Xbit_r14_c205 bl_205 br_205 wl_14 vdd gnd cell_6t
Xbit_r15_c205 bl_205 br_205 wl_15 vdd gnd cell_6t
Xbit_r16_c205 bl_205 br_205 wl_16 vdd gnd cell_6t
Xbit_r17_c205 bl_205 br_205 wl_17 vdd gnd cell_6t
Xbit_r18_c205 bl_205 br_205 wl_18 vdd gnd cell_6t
Xbit_r19_c205 bl_205 br_205 wl_19 vdd gnd cell_6t
Xbit_r20_c205 bl_205 br_205 wl_20 vdd gnd cell_6t
Xbit_r21_c205 bl_205 br_205 wl_21 vdd gnd cell_6t
Xbit_r22_c205 bl_205 br_205 wl_22 vdd gnd cell_6t
Xbit_r23_c205 bl_205 br_205 wl_23 vdd gnd cell_6t
Xbit_r24_c205 bl_205 br_205 wl_24 vdd gnd cell_6t
Xbit_r25_c205 bl_205 br_205 wl_25 vdd gnd cell_6t
Xbit_r26_c205 bl_205 br_205 wl_26 vdd gnd cell_6t
Xbit_r27_c205 bl_205 br_205 wl_27 vdd gnd cell_6t
Xbit_r28_c205 bl_205 br_205 wl_28 vdd gnd cell_6t
Xbit_r29_c205 bl_205 br_205 wl_29 vdd gnd cell_6t
Xbit_r30_c205 bl_205 br_205 wl_30 vdd gnd cell_6t
Xbit_r31_c205 bl_205 br_205 wl_31 vdd gnd cell_6t
Xbit_r32_c205 bl_205 br_205 wl_32 vdd gnd cell_6t
Xbit_r33_c205 bl_205 br_205 wl_33 vdd gnd cell_6t
Xbit_r34_c205 bl_205 br_205 wl_34 vdd gnd cell_6t
Xbit_r35_c205 bl_205 br_205 wl_35 vdd gnd cell_6t
Xbit_r36_c205 bl_205 br_205 wl_36 vdd gnd cell_6t
Xbit_r37_c205 bl_205 br_205 wl_37 vdd gnd cell_6t
Xbit_r38_c205 bl_205 br_205 wl_38 vdd gnd cell_6t
Xbit_r39_c205 bl_205 br_205 wl_39 vdd gnd cell_6t
Xbit_r40_c205 bl_205 br_205 wl_40 vdd gnd cell_6t
Xbit_r41_c205 bl_205 br_205 wl_41 vdd gnd cell_6t
Xbit_r42_c205 bl_205 br_205 wl_42 vdd gnd cell_6t
Xbit_r43_c205 bl_205 br_205 wl_43 vdd gnd cell_6t
Xbit_r44_c205 bl_205 br_205 wl_44 vdd gnd cell_6t
Xbit_r45_c205 bl_205 br_205 wl_45 vdd gnd cell_6t
Xbit_r46_c205 bl_205 br_205 wl_46 vdd gnd cell_6t
Xbit_r47_c205 bl_205 br_205 wl_47 vdd gnd cell_6t
Xbit_r48_c205 bl_205 br_205 wl_48 vdd gnd cell_6t
Xbit_r49_c205 bl_205 br_205 wl_49 vdd gnd cell_6t
Xbit_r50_c205 bl_205 br_205 wl_50 vdd gnd cell_6t
Xbit_r51_c205 bl_205 br_205 wl_51 vdd gnd cell_6t
Xbit_r52_c205 bl_205 br_205 wl_52 vdd gnd cell_6t
Xbit_r53_c205 bl_205 br_205 wl_53 vdd gnd cell_6t
Xbit_r54_c205 bl_205 br_205 wl_54 vdd gnd cell_6t
Xbit_r55_c205 bl_205 br_205 wl_55 vdd gnd cell_6t
Xbit_r56_c205 bl_205 br_205 wl_56 vdd gnd cell_6t
Xbit_r57_c205 bl_205 br_205 wl_57 vdd gnd cell_6t
Xbit_r58_c205 bl_205 br_205 wl_58 vdd gnd cell_6t
Xbit_r59_c205 bl_205 br_205 wl_59 vdd gnd cell_6t
Xbit_r60_c205 bl_205 br_205 wl_60 vdd gnd cell_6t
Xbit_r61_c205 bl_205 br_205 wl_61 vdd gnd cell_6t
Xbit_r62_c205 bl_205 br_205 wl_62 vdd gnd cell_6t
Xbit_r63_c205 bl_205 br_205 wl_63 vdd gnd cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd cell_6t
Xbit_r1_c206 bl_206 br_206 wl_1 vdd gnd cell_6t
Xbit_r2_c206 bl_206 br_206 wl_2 vdd gnd cell_6t
Xbit_r3_c206 bl_206 br_206 wl_3 vdd gnd cell_6t
Xbit_r4_c206 bl_206 br_206 wl_4 vdd gnd cell_6t
Xbit_r5_c206 bl_206 br_206 wl_5 vdd gnd cell_6t
Xbit_r6_c206 bl_206 br_206 wl_6 vdd gnd cell_6t
Xbit_r7_c206 bl_206 br_206 wl_7 vdd gnd cell_6t
Xbit_r8_c206 bl_206 br_206 wl_8 vdd gnd cell_6t
Xbit_r9_c206 bl_206 br_206 wl_9 vdd gnd cell_6t
Xbit_r10_c206 bl_206 br_206 wl_10 vdd gnd cell_6t
Xbit_r11_c206 bl_206 br_206 wl_11 vdd gnd cell_6t
Xbit_r12_c206 bl_206 br_206 wl_12 vdd gnd cell_6t
Xbit_r13_c206 bl_206 br_206 wl_13 vdd gnd cell_6t
Xbit_r14_c206 bl_206 br_206 wl_14 vdd gnd cell_6t
Xbit_r15_c206 bl_206 br_206 wl_15 vdd gnd cell_6t
Xbit_r16_c206 bl_206 br_206 wl_16 vdd gnd cell_6t
Xbit_r17_c206 bl_206 br_206 wl_17 vdd gnd cell_6t
Xbit_r18_c206 bl_206 br_206 wl_18 vdd gnd cell_6t
Xbit_r19_c206 bl_206 br_206 wl_19 vdd gnd cell_6t
Xbit_r20_c206 bl_206 br_206 wl_20 vdd gnd cell_6t
Xbit_r21_c206 bl_206 br_206 wl_21 vdd gnd cell_6t
Xbit_r22_c206 bl_206 br_206 wl_22 vdd gnd cell_6t
Xbit_r23_c206 bl_206 br_206 wl_23 vdd gnd cell_6t
Xbit_r24_c206 bl_206 br_206 wl_24 vdd gnd cell_6t
Xbit_r25_c206 bl_206 br_206 wl_25 vdd gnd cell_6t
Xbit_r26_c206 bl_206 br_206 wl_26 vdd gnd cell_6t
Xbit_r27_c206 bl_206 br_206 wl_27 vdd gnd cell_6t
Xbit_r28_c206 bl_206 br_206 wl_28 vdd gnd cell_6t
Xbit_r29_c206 bl_206 br_206 wl_29 vdd gnd cell_6t
Xbit_r30_c206 bl_206 br_206 wl_30 vdd gnd cell_6t
Xbit_r31_c206 bl_206 br_206 wl_31 vdd gnd cell_6t
Xbit_r32_c206 bl_206 br_206 wl_32 vdd gnd cell_6t
Xbit_r33_c206 bl_206 br_206 wl_33 vdd gnd cell_6t
Xbit_r34_c206 bl_206 br_206 wl_34 vdd gnd cell_6t
Xbit_r35_c206 bl_206 br_206 wl_35 vdd gnd cell_6t
Xbit_r36_c206 bl_206 br_206 wl_36 vdd gnd cell_6t
Xbit_r37_c206 bl_206 br_206 wl_37 vdd gnd cell_6t
Xbit_r38_c206 bl_206 br_206 wl_38 vdd gnd cell_6t
Xbit_r39_c206 bl_206 br_206 wl_39 vdd gnd cell_6t
Xbit_r40_c206 bl_206 br_206 wl_40 vdd gnd cell_6t
Xbit_r41_c206 bl_206 br_206 wl_41 vdd gnd cell_6t
Xbit_r42_c206 bl_206 br_206 wl_42 vdd gnd cell_6t
Xbit_r43_c206 bl_206 br_206 wl_43 vdd gnd cell_6t
Xbit_r44_c206 bl_206 br_206 wl_44 vdd gnd cell_6t
Xbit_r45_c206 bl_206 br_206 wl_45 vdd gnd cell_6t
Xbit_r46_c206 bl_206 br_206 wl_46 vdd gnd cell_6t
Xbit_r47_c206 bl_206 br_206 wl_47 vdd gnd cell_6t
Xbit_r48_c206 bl_206 br_206 wl_48 vdd gnd cell_6t
Xbit_r49_c206 bl_206 br_206 wl_49 vdd gnd cell_6t
Xbit_r50_c206 bl_206 br_206 wl_50 vdd gnd cell_6t
Xbit_r51_c206 bl_206 br_206 wl_51 vdd gnd cell_6t
Xbit_r52_c206 bl_206 br_206 wl_52 vdd gnd cell_6t
Xbit_r53_c206 bl_206 br_206 wl_53 vdd gnd cell_6t
Xbit_r54_c206 bl_206 br_206 wl_54 vdd gnd cell_6t
Xbit_r55_c206 bl_206 br_206 wl_55 vdd gnd cell_6t
Xbit_r56_c206 bl_206 br_206 wl_56 vdd gnd cell_6t
Xbit_r57_c206 bl_206 br_206 wl_57 vdd gnd cell_6t
Xbit_r58_c206 bl_206 br_206 wl_58 vdd gnd cell_6t
Xbit_r59_c206 bl_206 br_206 wl_59 vdd gnd cell_6t
Xbit_r60_c206 bl_206 br_206 wl_60 vdd gnd cell_6t
Xbit_r61_c206 bl_206 br_206 wl_61 vdd gnd cell_6t
Xbit_r62_c206 bl_206 br_206 wl_62 vdd gnd cell_6t
Xbit_r63_c206 bl_206 br_206 wl_63 vdd gnd cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd cell_6t
Xbit_r1_c207 bl_207 br_207 wl_1 vdd gnd cell_6t
Xbit_r2_c207 bl_207 br_207 wl_2 vdd gnd cell_6t
Xbit_r3_c207 bl_207 br_207 wl_3 vdd gnd cell_6t
Xbit_r4_c207 bl_207 br_207 wl_4 vdd gnd cell_6t
Xbit_r5_c207 bl_207 br_207 wl_5 vdd gnd cell_6t
Xbit_r6_c207 bl_207 br_207 wl_6 vdd gnd cell_6t
Xbit_r7_c207 bl_207 br_207 wl_7 vdd gnd cell_6t
Xbit_r8_c207 bl_207 br_207 wl_8 vdd gnd cell_6t
Xbit_r9_c207 bl_207 br_207 wl_9 vdd gnd cell_6t
Xbit_r10_c207 bl_207 br_207 wl_10 vdd gnd cell_6t
Xbit_r11_c207 bl_207 br_207 wl_11 vdd gnd cell_6t
Xbit_r12_c207 bl_207 br_207 wl_12 vdd gnd cell_6t
Xbit_r13_c207 bl_207 br_207 wl_13 vdd gnd cell_6t
Xbit_r14_c207 bl_207 br_207 wl_14 vdd gnd cell_6t
Xbit_r15_c207 bl_207 br_207 wl_15 vdd gnd cell_6t
Xbit_r16_c207 bl_207 br_207 wl_16 vdd gnd cell_6t
Xbit_r17_c207 bl_207 br_207 wl_17 vdd gnd cell_6t
Xbit_r18_c207 bl_207 br_207 wl_18 vdd gnd cell_6t
Xbit_r19_c207 bl_207 br_207 wl_19 vdd gnd cell_6t
Xbit_r20_c207 bl_207 br_207 wl_20 vdd gnd cell_6t
Xbit_r21_c207 bl_207 br_207 wl_21 vdd gnd cell_6t
Xbit_r22_c207 bl_207 br_207 wl_22 vdd gnd cell_6t
Xbit_r23_c207 bl_207 br_207 wl_23 vdd gnd cell_6t
Xbit_r24_c207 bl_207 br_207 wl_24 vdd gnd cell_6t
Xbit_r25_c207 bl_207 br_207 wl_25 vdd gnd cell_6t
Xbit_r26_c207 bl_207 br_207 wl_26 vdd gnd cell_6t
Xbit_r27_c207 bl_207 br_207 wl_27 vdd gnd cell_6t
Xbit_r28_c207 bl_207 br_207 wl_28 vdd gnd cell_6t
Xbit_r29_c207 bl_207 br_207 wl_29 vdd gnd cell_6t
Xbit_r30_c207 bl_207 br_207 wl_30 vdd gnd cell_6t
Xbit_r31_c207 bl_207 br_207 wl_31 vdd gnd cell_6t
Xbit_r32_c207 bl_207 br_207 wl_32 vdd gnd cell_6t
Xbit_r33_c207 bl_207 br_207 wl_33 vdd gnd cell_6t
Xbit_r34_c207 bl_207 br_207 wl_34 vdd gnd cell_6t
Xbit_r35_c207 bl_207 br_207 wl_35 vdd gnd cell_6t
Xbit_r36_c207 bl_207 br_207 wl_36 vdd gnd cell_6t
Xbit_r37_c207 bl_207 br_207 wl_37 vdd gnd cell_6t
Xbit_r38_c207 bl_207 br_207 wl_38 vdd gnd cell_6t
Xbit_r39_c207 bl_207 br_207 wl_39 vdd gnd cell_6t
Xbit_r40_c207 bl_207 br_207 wl_40 vdd gnd cell_6t
Xbit_r41_c207 bl_207 br_207 wl_41 vdd gnd cell_6t
Xbit_r42_c207 bl_207 br_207 wl_42 vdd gnd cell_6t
Xbit_r43_c207 bl_207 br_207 wl_43 vdd gnd cell_6t
Xbit_r44_c207 bl_207 br_207 wl_44 vdd gnd cell_6t
Xbit_r45_c207 bl_207 br_207 wl_45 vdd gnd cell_6t
Xbit_r46_c207 bl_207 br_207 wl_46 vdd gnd cell_6t
Xbit_r47_c207 bl_207 br_207 wl_47 vdd gnd cell_6t
Xbit_r48_c207 bl_207 br_207 wl_48 vdd gnd cell_6t
Xbit_r49_c207 bl_207 br_207 wl_49 vdd gnd cell_6t
Xbit_r50_c207 bl_207 br_207 wl_50 vdd gnd cell_6t
Xbit_r51_c207 bl_207 br_207 wl_51 vdd gnd cell_6t
Xbit_r52_c207 bl_207 br_207 wl_52 vdd gnd cell_6t
Xbit_r53_c207 bl_207 br_207 wl_53 vdd gnd cell_6t
Xbit_r54_c207 bl_207 br_207 wl_54 vdd gnd cell_6t
Xbit_r55_c207 bl_207 br_207 wl_55 vdd gnd cell_6t
Xbit_r56_c207 bl_207 br_207 wl_56 vdd gnd cell_6t
Xbit_r57_c207 bl_207 br_207 wl_57 vdd gnd cell_6t
Xbit_r58_c207 bl_207 br_207 wl_58 vdd gnd cell_6t
Xbit_r59_c207 bl_207 br_207 wl_59 vdd gnd cell_6t
Xbit_r60_c207 bl_207 br_207 wl_60 vdd gnd cell_6t
Xbit_r61_c207 bl_207 br_207 wl_61 vdd gnd cell_6t
Xbit_r62_c207 bl_207 br_207 wl_62 vdd gnd cell_6t
Xbit_r63_c207 bl_207 br_207 wl_63 vdd gnd cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd cell_6t
Xbit_r1_c208 bl_208 br_208 wl_1 vdd gnd cell_6t
Xbit_r2_c208 bl_208 br_208 wl_2 vdd gnd cell_6t
Xbit_r3_c208 bl_208 br_208 wl_3 vdd gnd cell_6t
Xbit_r4_c208 bl_208 br_208 wl_4 vdd gnd cell_6t
Xbit_r5_c208 bl_208 br_208 wl_5 vdd gnd cell_6t
Xbit_r6_c208 bl_208 br_208 wl_6 vdd gnd cell_6t
Xbit_r7_c208 bl_208 br_208 wl_7 vdd gnd cell_6t
Xbit_r8_c208 bl_208 br_208 wl_8 vdd gnd cell_6t
Xbit_r9_c208 bl_208 br_208 wl_9 vdd gnd cell_6t
Xbit_r10_c208 bl_208 br_208 wl_10 vdd gnd cell_6t
Xbit_r11_c208 bl_208 br_208 wl_11 vdd gnd cell_6t
Xbit_r12_c208 bl_208 br_208 wl_12 vdd gnd cell_6t
Xbit_r13_c208 bl_208 br_208 wl_13 vdd gnd cell_6t
Xbit_r14_c208 bl_208 br_208 wl_14 vdd gnd cell_6t
Xbit_r15_c208 bl_208 br_208 wl_15 vdd gnd cell_6t
Xbit_r16_c208 bl_208 br_208 wl_16 vdd gnd cell_6t
Xbit_r17_c208 bl_208 br_208 wl_17 vdd gnd cell_6t
Xbit_r18_c208 bl_208 br_208 wl_18 vdd gnd cell_6t
Xbit_r19_c208 bl_208 br_208 wl_19 vdd gnd cell_6t
Xbit_r20_c208 bl_208 br_208 wl_20 vdd gnd cell_6t
Xbit_r21_c208 bl_208 br_208 wl_21 vdd gnd cell_6t
Xbit_r22_c208 bl_208 br_208 wl_22 vdd gnd cell_6t
Xbit_r23_c208 bl_208 br_208 wl_23 vdd gnd cell_6t
Xbit_r24_c208 bl_208 br_208 wl_24 vdd gnd cell_6t
Xbit_r25_c208 bl_208 br_208 wl_25 vdd gnd cell_6t
Xbit_r26_c208 bl_208 br_208 wl_26 vdd gnd cell_6t
Xbit_r27_c208 bl_208 br_208 wl_27 vdd gnd cell_6t
Xbit_r28_c208 bl_208 br_208 wl_28 vdd gnd cell_6t
Xbit_r29_c208 bl_208 br_208 wl_29 vdd gnd cell_6t
Xbit_r30_c208 bl_208 br_208 wl_30 vdd gnd cell_6t
Xbit_r31_c208 bl_208 br_208 wl_31 vdd gnd cell_6t
Xbit_r32_c208 bl_208 br_208 wl_32 vdd gnd cell_6t
Xbit_r33_c208 bl_208 br_208 wl_33 vdd gnd cell_6t
Xbit_r34_c208 bl_208 br_208 wl_34 vdd gnd cell_6t
Xbit_r35_c208 bl_208 br_208 wl_35 vdd gnd cell_6t
Xbit_r36_c208 bl_208 br_208 wl_36 vdd gnd cell_6t
Xbit_r37_c208 bl_208 br_208 wl_37 vdd gnd cell_6t
Xbit_r38_c208 bl_208 br_208 wl_38 vdd gnd cell_6t
Xbit_r39_c208 bl_208 br_208 wl_39 vdd gnd cell_6t
Xbit_r40_c208 bl_208 br_208 wl_40 vdd gnd cell_6t
Xbit_r41_c208 bl_208 br_208 wl_41 vdd gnd cell_6t
Xbit_r42_c208 bl_208 br_208 wl_42 vdd gnd cell_6t
Xbit_r43_c208 bl_208 br_208 wl_43 vdd gnd cell_6t
Xbit_r44_c208 bl_208 br_208 wl_44 vdd gnd cell_6t
Xbit_r45_c208 bl_208 br_208 wl_45 vdd gnd cell_6t
Xbit_r46_c208 bl_208 br_208 wl_46 vdd gnd cell_6t
Xbit_r47_c208 bl_208 br_208 wl_47 vdd gnd cell_6t
Xbit_r48_c208 bl_208 br_208 wl_48 vdd gnd cell_6t
Xbit_r49_c208 bl_208 br_208 wl_49 vdd gnd cell_6t
Xbit_r50_c208 bl_208 br_208 wl_50 vdd gnd cell_6t
Xbit_r51_c208 bl_208 br_208 wl_51 vdd gnd cell_6t
Xbit_r52_c208 bl_208 br_208 wl_52 vdd gnd cell_6t
Xbit_r53_c208 bl_208 br_208 wl_53 vdd gnd cell_6t
Xbit_r54_c208 bl_208 br_208 wl_54 vdd gnd cell_6t
Xbit_r55_c208 bl_208 br_208 wl_55 vdd gnd cell_6t
Xbit_r56_c208 bl_208 br_208 wl_56 vdd gnd cell_6t
Xbit_r57_c208 bl_208 br_208 wl_57 vdd gnd cell_6t
Xbit_r58_c208 bl_208 br_208 wl_58 vdd gnd cell_6t
Xbit_r59_c208 bl_208 br_208 wl_59 vdd gnd cell_6t
Xbit_r60_c208 bl_208 br_208 wl_60 vdd gnd cell_6t
Xbit_r61_c208 bl_208 br_208 wl_61 vdd gnd cell_6t
Xbit_r62_c208 bl_208 br_208 wl_62 vdd gnd cell_6t
Xbit_r63_c208 bl_208 br_208 wl_63 vdd gnd cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd cell_6t
Xbit_r1_c209 bl_209 br_209 wl_1 vdd gnd cell_6t
Xbit_r2_c209 bl_209 br_209 wl_2 vdd gnd cell_6t
Xbit_r3_c209 bl_209 br_209 wl_3 vdd gnd cell_6t
Xbit_r4_c209 bl_209 br_209 wl_4 vdd gnd cell_6t
Xbit_r5_c209 bl_209 br_209 wl_5 vdd gnd cell_6t
Xbit_r6_c209 bl_209 br_209 wl_6 vdd gnd cell_6t
Xbit_r7_c209 bl_209 br_209 wl_7 vdd gnd cell_6t
Xbit_r8_c209 bl_209 br_209 wl_8 vdd gnd cell_6t
Xbit_r9_c209 bl_209 br_209 wl_9 vdd gnd cell_6t
Xbit_r10_c209 bl_209 br_209 wl_10 vdd gnd cell_6t
Xbit_r11_c209 bl_209 br_209 wl_11 vdd gnd cell_6t
Xbit_r12_c209 bl_209 br_209 wl_12 vdd gnd cell_6t
Xbit_r13_c209 bl_209 br_209 wl_13 vdd gnd cell_6t
Xbit_r14_c209 bl_209 br_209 wl_14 vdd gnd cell_6t
Xbit_r15_c209 bl_209 br_209 wl_15 vdd gnd cell_6t
Xbit_r16_c209 bl_209 br_209 wl_16 vdd gnd cell_6t
Xbit_r17_c209 bl_209 br_209 wl_17 vdd gnd cell_6t
Xbit_r18_c209 bl_209 br_209 wl_18 vdd gnd cell_6t
Xbit_r19_c209 bl_209 br_209 wl_19 vdd gnd cell_6t
Xbit_r20_c209 bl_209 br_209 wl_20 vdd gnd cell_6t
Xbit_r21_c209 bl_209 br_209 wl_21 vdd gnd cell_6t
Xbit_r22_c209 bl_209 br_209 wl_22 vdd gnd cell_6t
Xbit_r23_c209 bl_209 br_209 wl_23 vdd gnd cell_6t
Xbit_r24_c209 bl_209 br_209 wl_24 vdd gnd cell_6t
Xbit_r25_c209 bl_209 br_209 wl_25 vdd gnd cell_6t
Xbit_r26_c209 bl_209 br_209 wl_26 vdd gnd cell_6t
Xbit_r27_c209 bl_209 br_209 wl_27 vdd gnd cell_6t
Xbit_r28_c209 bl_209 br_209 wl_28 vdd gnd cell_6t
Xbit_r29_c209 bl_209 br_209 wl_29 vdd gnd cell_6t
Xbit_r30_c209 bl_209 br_209 wl_30 vdd gnd cell_6t
Xbit_r31_c209 bl_209 br_209 wl_31 vdd gnd cell_6t
Xbit_r32_c209 bl_209 br_209 wl_32 vdd gnd cell_6t
Xbit_r33_c209 bl_209 br_209 wl_33 vdd gnd cell_6t
Xbit_r34_c209 bl_209 br_209 wl_34 vdd gnd cell_6t
Xbit_r35_c209 bl_209 br_209 wl_35 vdd gnd cell_6t
Xbit_r36_c209 bl_209 br_209 wl_36 vdd gnd cell_6t
Xbit_r37_c209 bl_209 br_209 wl_37 vdd gnd cell_6t
Xbit_r38_c209 bl_209 br_209 wl_38 vdd gnd cell_6t
Xbit_r39_c209 bl_209 br_209 wl_39 vdd gnd cell_6t
Xbit_r40_c209 bl_209 br_209 wl_40 vdd gnd cell_6t
Xbit_r41_c209 bl_209 br_209 wl_41 vdd gnd cell_6t
Xbit_r42_c209 bl_209 br_209 wl_42 vdd gnd cell_6t
Xbit_r43_c209 bl_209 br_209 wl_43 vdd gnd cell_6t
Xbit_r44_c209 bl_209 br_209 wl_44 vdd gnd cell_6t
Xbit_r45_c209 bl_209 br_209 wl_45 vdd gnd cell_6t
Xbit_r46_c209 bl_209 br_209 wl_46 vdd gnd cell_6t
Xbit_r47_c209 bl_209 br_209 wl_47 vdd gnd cell_6t
Xbit_r48_c209 bl_209 br_209 wl_48 vdd gnd cell_6t
Xbit_r49_c209 bl_209 br_209 wl_49 vdd gnd cell_6t
Xbit_r50_c209 bl_209 br_209 wl_50 vdd gnd cell_6t
Xbit_r51_c209 bl_209 br_209 wl_51 vdd gnd cell_6t
Xbit_r52_c209 bl_209 br_209 wl_52 vdd gnd cell_6t
Xbit_r53_c209 bl_209 br_209 wl_53 vdd gnd cell_6t
Xbit_r54_c209 bl_209 br_209 wl_54 vdd gnd cell_6t
Xbit_r55_c209 bl_209 br_209 wl_55 vdd gnd cell_6t
Xbit_r56_c209 bl_209 br_209 wl_56 vdd gnd cell_6t
Xbit_r57_c209 bl_209 br_209 wl_57 vdd gnd cell_6t
Xbit_r58_c209 bl_209 br_209 wl_58 vdd gnd cell_6t
Xbit_r59_c209 bl_209 br_209 wl_59 vdd gnd cell_6t
Xbit_r60_c209 bl_209 br_209 wl_60 vdd gnd cell_6t
Xbit_r61_c209 bl_209 br_209 wl_61 vdd gnd cell_6t
Xbit_r62_c209 bl_209 br_209 wl_62 vdd gnd cell_6t
Xbit_r63_c209 bl_209 br_209 wl_63 vdd gnd cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd cell_6t
Xbit_r1_c210 bl_210 br_210 wl_1 vdd gnd cell_6t
Xbit_r2_c210 bl_210 br_210 wl_2 vdd gnd cell_6t
Xbit_r3_c210 bl_210 br_210 wl_3 vdd gnd cell_6t
Xbit_r4_c210 bl_210 br_210 wl_4 vdd gnd cell_6t
Xbit_r5_c210 bl_210 br_210 wl_5 vdd gnd cell_6t
Xbit_r6_c210 bl_210 br_210 wl_6 vdd gnd cell_6t
Xbit_r7_c210 bl_210 br_210 wl_7 vdd gnd cell_6t
Xbit_r8_c210 bl_210 br_210 wl_8 vdd gnd cell_6t
Xbit_r9_c210 bl_210 br_210 wl_9 vdd gnd cell_6t
Xbit_r10_c210 bl_210 br_210 wl_10 vdd gnd cell_6t
Xbit_r11_c210 bl_210 br_210 wl_11 vdd gnd cell_6t
Xbit_r12_c210 bl_210 br_210 wl_12 vdd gnd cell_6t
Xbit_r13_c210 bl_210 br_210 wl_13 vdd gnd cell_6t
Xbit_r14_c210 bl_210 br_210 wl_14 vdd gnd cell_6t
Xbit_r15_c210 bl_210 br_210 wl_15 vdd gnd cell_6t
Xbit_r16_c210 bl_210 br_210 wl_16 vdd gnd cell_6t
Xbit_r17_c210 bl_210 br_210 wl_17 vdd gnd cell_6t
Xbit_r18_c210 bl_210 br_210 wl_18 vdd gnd cell_6t
Xbit_r19_c210 bl_210 br_210 wl_19 vdd gnd cell_6t
Xbit_r20_c210 bl_210 br_210 wl_20 vdd gnd cell_6t
Xbit_r21_c210 bl_210 br_210 wl_21 vdd gnd cell_6t
Xbit_r22_c210 bl_210 br_210 wl_22 vdd gnd cell_6t
Xbit_r23_c210 bl_210 br_210 wl_23 vdd gnd cell_6t
Xbit_r24_c210 bl_210 br_210 wl_24 vdd gnd cell_6t
Xbit_r25_c210 bl_210 br_210 wl_25 vdd gnd cell_6t
Xbit_r26_c210 bl_210 br_210 wl_26 vdd gnd cell_6t
Xbit_r27_c210 bl_210 br_210 wl_27 vdd gnd cell_6t
Xbit_r28_c210 bl_210 br_210 wl_28 vdd gnd cell_6t
Xbit_r29_c210 bl_210 br_210 wl_29 vdd gnd cell_6t
Xbit_r30_c210 bl_210 br_210 wl_30 vdd gnd cell_6t
Xbit_r31_c210 bl_210 br_210 wl_31 vdd gnd cell_6t
Xbit_r32_c210 bl_210 br_210 wl_32 vdd gnd cell_6t
Xbit_r33_c210 bl_210 br_210 wl_33 vdd gnd cell_6t
Xbit_r34_c210 bl_210 br_210 wl_34 vdd gnd cell_6t
Xbit_r35_c210 bl_210 br_210 wl_35 vdd gnd cell_6t
Xbit_r36_c210 bl_210 br_210 wl_36 vdd gnd cell_6t
Xbit_r37_c210 bl_210 br_210 wl_37 vdd gnd cell_6t
Xbit_r38_c210 bl_210 br_210 wl_38 vdd gnd cell_6t
Xbit_r39_c210 bl_210 br_210 wl_39 vdd gnd cell_6t
Xbit_r40_c210 bl_210 br_210 wl_40 vdd gnd cell_6t
Xbit_r41_c210 bl_210 br_210 wl_41 vdd gnd cell_6t
Xbit_r42_c210 bl_210 br_210 wl_42 vdd gnd cell_6t
Xbit_r43_c210 bl_210 br_210 wl_43 vdd gnd cell_6t
Xbit_r44_c210 bl_210 br_210 wl_44 vdd gnd cell_6t
Xbit_r45_c210 bl_210 br_210 wl_45 vdd gnd cell_6t
Xbit_r46_c210 bl_210 br_210 wl_46 vdd gnd cell_6t
Xbit_r47_c210 bl_210 br_210 wl_47 vdd gnd cell_6t
Xbit_r48_c210 bl_210 br_210 wl_48 vdd gnd cell_6t
Xbit_r49_c210 bl_210 br_210 wl_49 vdd gnd cell_6t
Xbit_r50_c210 bl_210 br_210 wl_50 vdd gnd cell_6t
Xbit_r51_c210 bl_210 br_210 wl_51 vdd gnd cell_6t
Xbit_r52_c210 bl_210 br_210 wl_52 vdd gnd cell_6t
Xbit_r53_c210 bl_210 br_210 wl_53 vdd gnd cell_6t
Xbit_r54_c210 bl_210 br_210 wl_54 vdd gnd cell_6t
Xbit_r55_c210 bl_210 br_210 wl_55 vdd gnd cell_6t
Xbit_r56_c210 bl_210 br_210 wl_56 vdd gnd cell_6t
Xbit_r57_c210 bl_210 br_210 wl_57 vdd gnd cell_6t
Xbit_r58_c210 bl_210 br_210 wl_58 vdd gnd cell_6t
Xbit_r59_c210 bl_210 br_210 wl_59 vdd gnd cell_6t
Xbit_r60_c210 bl_210 br_210 wl_60 vdd gnd cell_6t
Xbit_r61_c210 bl_210 br_210 wl_61 vdd gnd cell_6t
Xbit_r62_c210 bl_210 br_210 wl_62 vdd gnd cell_6t
Xbit_r63_c210 bl_210 br_210 wl_63 vdd gnd cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd cell_6t
Xbit_r1_c211 bl_211 br_211 wl_1 vdd gnd cell_6t
Xbit_r2_c211 bl_211 br_211 wl_2 vdd gnd cell_6t
Xbit_r3_c211 bl_211 br_211 wl_3 vdd gnd cell_6t
Xbit_r4_c211 bl_211 br_211 wl_4 vdd gnd cell_6t
Xbit_r5_c211 bl_211 br_211 wl_5 vdd gnd cell_6t
Xbit_r6_c211 bl_211 br_211 wl_6 vdd gnd cell_6t
Xbit_r7_c211 bl_211 br_211 wl_7 vdd gnd cell_6t
Xbit_r8_c211 bl_211 br_211 wl_8 vdd gnd cell_6t
Xbit_r9_c211 bl_211 br_211 wl_9 vdd gnd cell_6t
Xbit_r10_c211 bl_211 br_211 wl_10 vdd gnd cell_6t
Xbit_r11_c211 bl_211 br_211 wl_11 vdd gnd cell_6t
Xbit_r12_c211 bl_211 br_211 wl_12 vdd gnd cell_6t
Xbit_r13_c211 bl_211 br_211 wl_13 vdd gnd cell_6t
Xbit_r14_c211 bl_211 br_211 wl_14 vdd gnd cell_6t
Xbit_r15_c211 bl_211 br_211 wl_15 vdd gnd cell_6t
Xbit_r16_c211 bl_211 br_211 wl_16 vdd gnd cell_6t
Xbit_r17_c211 bl_211 br_211 wl_17 vdd gnd cell_6t
Xbit_r18_c211 bl_211 br_211 wl_18 vdd gnd cell_6t
Xbit_r19_c211 bl_211 br_211 wl_19 vdd gnd cell_6t
Xbit_r20_c211 bl_211 br_211 wl_20 vdd gnd cell_6t
Xbit_r21_c211 bl_211 br_211 wl_21 vdd gnd cell_6t
Xbit_r22_c211 bl_211 br_211 wl_22 vdd gnd cell_6t
Xbit_r23_c211 bl_211 br_211 wl_23 vdd gnd cell_6t
Xbit_r24_c211 bl_211 br_211 wl_24 vdd gnd cell_6t
Xbit_r25_c211 bl_211 br_211 wl_25 vdd gnd cell_6t
Xbit_r26_c211 bl_211 br_211 wl_26 vdd gnd cell_6t
Xbit_r27_c211 bl_211 br_211 wl_27 vdd gnd cell_6t
Xbit_r28_c211 bl_211 br_211 wl_28 vdd gnd cell_6t
Xbit_r29_c211 bl_211 br_211 wl_29 vdd gnd cell_6t
Xbit_r30_c211 bl_211 br_211 wl_30 vdd gnd cell_6t
Xbit_r31_c211 bl_211 br_211 wl_31 vdd gnd cell_6t
Xbit_r32_c211 bl_211 br_211 wl_32 vdd gnd cell_6t
Xbit_r33_c211 bl_211 br_211 wl_33 vdd gnd cell_6t
Xbit_r34_c211 bl_211 br_211 wl_34 vdd gnd cell_6t
Xbit_r35_c211 bl_211 br_211 wl_35 vdd gnd cell_6t
Xbit_r36_c211 bl_211 br_211 wl_36 vdd gnd cell_6t
Xbit_r37_c211 bl_211 br_211 wl_37 vdd gnd cell_6t
Xbit_r38_c211 bl_211 br_211 wl_38 vdd gnd cell_6t
Xbit_r39_c211 bl_211 br_211 wl_39 vdd gnd cell_6t
Xbit_r40_c211 bl_211 br_211 wl_40 vdd gnd cell_6t
Xbit_r41_c211 bl_211 br_211 wl_41 vdd gnd cell_6t
Xbit_r42_c211 bl_211 br_211 wl_42 vdd gnd cell_6t
Xbit_r43_c211 bl_211 br_211 wl_43 vdd gnd cell_6t
Xbit_r44_c211 bl_211 br_211 wl_44 vdd gnd cell_6t
Xbit_r45_c211 bl_211 br_211 wl_45 vdd gnd cell_6t
Xbit_r46_c211 bl_211 br_211 wl_46 vdd gnd cell_6t
Xbit_r47_c211 bl_211 br_211 wl_47 vdd gnd cell_6t
Xbit_r48_c211 bl_211 br_211 wl_48 vdd gnd cell_6t
Xbit_r49_c211 bl_211 br_211 wl_49 vdd gnd cell_6t
Xbit_r50_c211 bl_211 br_211 wl_50 vdd gnd cell_6t
Xbit_r51_c211 bl_211 br_211 wl_51 vdd gnd cell_6t
Xbit_r52_c211 bl_211 br_211 wl_52 vdd gnd cell_6t
Xbit_r53_c211 bl_211 br_211 wl_53 vdd gnd cell_6t
Xbit_r54_c211 bl_211 br_211 wl_54 vdd gnd cell_6t
Xbit_r55_c211 bl_211 br_211 wl_55 vdd gnd cell_6t
Xbit_r56_c211 bl_211 br_211 wl_56 vdd gnd cell_6t
Xbit_r57_c211 bl_211 br_211 wl_57 vdd gnd cell_6t
Xbit_r58_c211 bl_211 br_211 wl_58 vdd gnd cell_6t
Xbit_r59_c211 bl_211 br_211 wl_59 vdd gnd cell_6t
Xbit_r60_c211 bl_211 br_211 wl_60 vdd gnd cell_6t
Xbit_r61_c211 bl_211 br_211 wl_61 vdd gnd cell_6t
Xbit_r62_c211 bl_211 br_211 wl_62 vdd gnd cell_6t
Xbit_r63_c211 bl_211 br_211 wl_63 vdd gnd cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd cell_6t
Xbit_r1_c212 bl_212 br_212 wl_1 vdd gnd cell_6t
Xbit_r2_c212 bl_212 br_212 wl_2 vdd gnd cell_6t
Xbit_r3_c212 bl_212 br_212 wl_3 vdd gnd cell_6t
Xbit_r4_c212 bl_212 br_212 wl_4 vdd gnd cell_6t
Xbit_r5_c212 bl_212 br_212 wl_5 vdd gnd cell_6t
Xbit_r6_c212 bl_212 br_212 wl_6 vdd gnd cell_6t
Xbit_r7_c212 bl_212 br_212 wl_7 vdd gnd cell_6t
Xbit_r8_c212 bl_212 br_212 wl_8 vdd gnd cell_6t
Xbit_r9_c212 bl_212 br_212 wl_9 vdd gnd cell_6t
Xbit_r10_c212 bl_212 br_212 wl_10 vdd gnd cell_6t
Xbit_r11_c212 bl_212 br_212 wl_11 vdd gnd cell_6t
Xbit_r12_c212 bl_212 br_212 wl_12 vdd gnd cell_6t
Xbit_r13_c212 bl_212 br_212 wl_13 vdd gnd cell_6t
Xbit_r14_c212 bl_212 br_212 wl_14 vdd gnd cell_6t
Xbit_r15_c212 bl_212 br_212 wl_15 vdd gnd cell_6t
Xbit_r16_c212 bl_212 br_212 wl_16 vdd gnd cell_6t
Xbit_r17_c212 bl_212 br_212 wl_17 vdd gnd cell_6t
Xbit_r18_c212 bl_212 br_212 wl_18 vdd gnd cell_6t
Xbit_r19_c212 bl_212 br_212 wl_19 vdd gnd cell_6t
Xbit_r20_c212 bl_212 br_212 wl_20 vdd gnd cell_6t
Xbit_r21_c212 bl_212 br_212 wl_21 vdd gnd cell_6t
Xbit_r22_c212 bl_212 br_212 wl_22 vdd gnd cell_6t
Xbit_r23_c212 bl_212 br_212 wl_23 vdd gnd cell_6t
Xbit_r24_c212 bl_212 br_212 wl_24 vdd gnd cell_6t
Xbit_r25_c212 bl_212 br_212 wl_25 vdd gnd cell_6t
Xbit_r26_c212 bl_212 br_212 wl_26 vdd gnd cell_6t
Xbit_r27_c212 bl_212 br_212 wl_27 vdd gnd cell_6t
Xbit_r28_c212 bl_212 br_212 wl_28 vdd gnd cell_6t
Xbit_r29_c212 bl_212 br_212 wl_29 vdd gnd cell_6t
Xbit_r30_c212 bl_212 br_212 wl_30 vdd gnd cell_6t
Xbit_r31_c212 bl_212 br_212 wl_31 vdd gnd cell_6t
Xbit_r32_c212 bl_212 br_212 wl_32 vdd gnd cell_6t
Xbit_r33_c212 bl_212 br_212 wl_33 vdd gnd cell_6t
Xbit_r34_c212 bl_212 br_212 wl_34 vdd gnd cell_6t
Xbit_r35_c212 bl_212 br_212 wl_35 vdd gnd cell_6t
Xbit_r36_c212 bl_212 br_212 wl_36 vdd gnd cell_6t
Xbit_r37_c212 bl_212 br_212 wl_37 vdd gnd cell_6t
Xbit_r38_c212 bl_212 br_212 wl_38 vdd gnd cell_6t
Xbit_r39_c212 bl_212 br_212 wl_39 vdd gnd cell_6t
Xbit_r40_c212 bl_212 br_212 wl_40 vdd gnd cell_6t
Xbit_r41_c212 bl_212 br_212 wl_41 vdd gnd cell_6t
Xbit_r42_c212 bl_212 br_212 wl_42 vdd gnd cell_6t
Xbit_r43_c212 bl_212 br_212 wl_43 vdd gnd cell_6t
Xbit_r44_c212 bl_212 br_212 wl_44 vdd gnd cell_6t
Xbit_r45_c212 bl_212 br_212 wl_45 vdd gnd cell_6t
Xbit_r46_c212 bl_212 br_212 wl_46 vdd gnd cell_6t
Xbit_r47_c212 bl_212 br_212 wl_47 vdd gnd cell_6t
Xbit_r48_c212 bl_212 br_212 wl_48 vdd gnd cell_6t
Xbit_r49_c212 bl_212 br_212 wl_49 vdd gnd cell_6t
Xbit_r50_c212 bl_212 br_212 wl_50 vdd gnd cell_6t
Xbit_r51_c212 bl_212 br_212 wl_51 vdd gnd cell_6t
Xbit_r52_c212 bl_212 br_212 wl_52 vdd gnd cell_6t
Xbit_r53_c212 bl_212 br_212 wl_53 vdd gnd cell_6t
Xbit_r54_c212 bl_212 br_212 wl_54 vdd gnd cell_6t
Xbit_r55_c212 bl_212 br_212 wl_55 vdd gnd cell_6t
Xbit_r56_c212 bl_212 br_212 wl_56 vdd gnd cell_6t
Xbit_r57_c212 bl_212 br_212 wl_57 vdd gnd cell_6t
Xbit_r58_c212 bl_212 br_212 wl_58 vdd gnd cell_6t
Xbit_r59_c212 bl_212 br_212 wl_59 vdd gnd cell_6t
Xbit_r60_c212 bl_212 br_212 wl_60 vdd gnd cell_6t
Xbit_r61_c212 bl_212 br_212 wl_61 vdd gnd cell_6t
Xbit_r62_c212 bl_212 br_212 wl_62 vdd gnd cell_6t
Xbit_r63_c212 bl_212 br_212 wl_63 vdd gnd cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd cell_6t
Xbit_r1_c213 bl_213 br_213 wl_1 vdd gnd cell_6t
Xbit_r2_c213 bl_213 br_213 wl_2 vdd gnd cell_6t
Xbit_r3_c213 bl_213 br_213 wl_3 vdd gnd cell_6t
Xbit_r4_c213 bl_213 br_213 wl_4 vdd gnd cell_6t
Xbit_r5_c213 bl_213 br_213 wl_5 vdd gnd cell_6t
Xbit_r6_c213 bl_213 br_213 wl_6 vdd gnd cell_6t
Xbit_r7_c213 bl_213 br_213 wl_7 vdd gnd cell_6t
Xbit_r8_c213 bl_213 br_213 wl_8 vdd gnd cell_6t
Xbit_r9_c213 bl_213 br_213 wl_9 vdd gnd cell_6t
Xbit_r10_c213 bl_213 br_213 wl_10 vdd gnd cell_6t
Xbit_r11_c213 bl_213 br_213 wl_11 vdd gnd cell_6t
Xbit_r12_c213 bl_213 br_213 wl_12 vdd gnd cell_6t
Xbit_r13_c213 bl_213 br_213 wl_13 vdd gnd cell_6t
Xbit_r14_c213 bl_213 br_213 wl_14 vdd gnd cell_6t
Xbit_r15_c213 bl_213 br_213 wl_15 vdd gnd cell_6t
Xbit_r16_c213 bl_213 br_213 wl_16 vdd gnd cell_6t
Xbit_r17_c213 bl_213 br_213 wl_17 vdd gnd cell_6t
Xbit_r18_c213 bl_213 br_213 wl_18 vdd gnd cell_6t
Xbit_r19_c213 bl_213 br_213 wl_19 vdd gnd cell_6t
Xbit_r20_c213 bl_213 br_213 wl_20 vdd gnd cell_6t
Xbit_r21_c213 bl_213 br_213 wl_21 vdd gnd cell_6t
Xbit_r22_c213 bl_213 br_213 wl_22 vdd gnd cell_6t
Xbit_r23_c213 bl_213 br_213 wl_23 vdd gnd cell_6t
Xbit_r24_c213 bl_213 br_213 wl_24 vdd gnd cell_6t
Xbit_r25_c213 bl_213 br_213 wl_25 vdd gnd cell_6t
Xbit_r26_c213 bl_213 br_213 wl_26 vdd gnd cell_6t
Xbit_r27_c213 bl_213 br_213 wl_27 vdd gnd cell_6t
Xbit_r28_c213 bl_213 br_213 wl_28 vdd gnd cell_6t
Xbit_r29_c213 bl_213 br_213 wl_29 vdd gnd cell_6t
Xbit_r30_c213 bl_213 br_213 wl_30 vdd gnd cell_6t
Xbit_r31_c213 bl_213 br_213 wl_31 vdd gnd cell_6t
Xbit_r32_c213 bl_213 br_213 wl_32 vdd gnd cell_6t
Xbit_r33_c213 bl_213 br_213 wl_33 vdd gnd cell_6t
Xbit_r34_c213 bl_213 br_213 wl_34 vdd gnd cell_6t
Xbit_r35_c213 bl_213 br_213 wl_35 vdd gnd cell_6t
Xbit_r36_c213 bl_213 br_213 wl_36 vdd gnd cell_6t
Xbit_r37_c213 bl_213 br_213 wl_37 vdd gnd cell_6t
Xbit_r38_c213 bl_213 br_213 wl_38 vdd gnd cell_6t
Xbit_r39_c213 bl_213 br_213 wl_39 vdd gnd cell_6t
Xbit_r40_c213 bl_213 br_213 wl_40 vdd gnd cell_6t
Xbit_r41_c213 bl_213 br_213 wl_41 vdd gnd cell_6t
Xbit_r42_c213 bl_213 br_213 wl_42 vdd gnd cell_6t
Xbit_r43_c213 bl_213 br_213 wl_43 vdd gnd cell_6t
Xbit_r44_c213 bl_213 br_213 wl_44 vdd gnd cell_6t
Xbit_r45_c213 bl_213 br_213 wl_45 vdd gnd cell_6t
Xbit_r46_c213 bl_213 br_213 wl_46 vdd gnd cell_6t
Xbit_r47_c213 bl_213 br_213 wl_47 vdd gnd cell_6t
Xbit_r48_c213 bl_213 br_213 wl_48 vdd gnd cell_6t
Xbit_r49_c213 bl_213 br_213 wl_49 vdd gnd cell_6t
Xbit_r50_c213 bl_213 br_213 wl_50 vdd gnd cell_6t
Xbit_r51_c213 bl_213 br_213 wl_51 vdd gnd cell_6t
Xbit_r52_c213 bl_213 br_213 wl_52 vdd gnd cell_6t
Xbit_r53_c213 bl_213 br_213 wl_53 vdd gnd cell_6t
Xbit_r54_c213 bl_213 br_213 wl_54 vdd gnd cell_6t
Xbit_r55_c213 bl_213 br_213 wl_55 vdd gnd cell_6t
Xbit_r56_c213 bl_213 br_213 wl_56 vdd gnd cell_6t
Xbit_r57_c213 bl_213 br_213 wl_57 vdd gnd cell_6t
Xbit_r58_c213 bl_213 br_213 wl_58 vdd gnd cell_6t
Xbit_r59_c213 bl_213 br_213 wl_59 vdd gnd cell_6t
Xbit_r60_c213 bl_213 br_213 wl_60 vdd gnd cell_6t
Xbit_r61_c213 bl_213 br_213 wl_61 vdd gnd cell_6t
Xbit_r62_c213 bl_213 br_213 wl_62 vdd gnd cell_6t
Xbit_r63_c213 bl_213 br_213 wl_63 vdd gnd cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd cell_6t
Xbit_r1_c214 bl_214 br_214 wl_1 vdd gnd cell_6t
Xbit_r2_c214 bl_214 br_214 wl_2 vdd gnd cell_6t
Xbit_r3_c214 bl_214 br_214 wl_3 vdd gnd cell_6t
Xbit_r4_c214 bl_214 br_214 wl_4 vdd gnd cell_6t
Xbit_r5_c214 bl_214 br_214 wl_5 vdd gnd cell_6t
Xbit_r6_c214 bl_214 br_214 wl_6 vdd gnd cell_6t
Xbit_r7_c214 bl_214 br_214 wl_7 vdd gnd cell_6t
Xbit_r8_c214 bl_214 br_214 wl_8 vdd gnd cell_6t
Xbit_r9_c214 bl_214 br_214 wl_9 vdd gnd cell_6t
Xbit_r10_c214 bl_214 br_214 wl_10 vdd gnd cell_6t
Xbit_r11_c214 bl_214 br_214 wl_11 vdd gnd cell_6t
Xbit_r12_c214 bl_214 br_214 wl_12 vdd gnd cell_6t
Xbit_r13_c214 bl_214 br_214 wl_13 vdd gnd cell_6t
Xbit_r14_c214 bl_214 br_214 wl_14 vdd gnd cell_6t
Xbit_r15_c214 bl_214 br_214 wl_15 vdd gnd cell_6t
Xbit_r16_c214 bl_214 br_214 wl_16 vdd gnd cell_6t
Xbit_r17_c214 bl_214 br_214 wl_17 vdd gnd cell_6t
Xbit_r18_c214 bl_214 br_214 wl_18 vdd gnd cell_6t
Xbit_r19_c214 bl_214 br_214 wl_19 vdd gnd cell_6t
Xbit_r20_c214 bl_214 br_214 wl_20 vdd gnd cell_6t
Xbit_r21_c214 bl_214 br_214 wl_21 vdd gnd cell_6t
Xbit_r22_c214 bl_214 br_214 wl_22 vdd gnd cell_6t
Xbit_r23_c214 bl_214 br_214 wl_23 vdd gnd cell_6t
Xbit_r24_c214 bl_214 br_214 wl_24 vdd gnd cell_6t
Xbit_r25_c214 bl_214 br_214 wl_25 vdd gnd cell_6t
Xbit_r26_c214 bl_214 br_214 wl_26 vdd gnd cell_6t
Xbit_r27_c214 bl_214 br_214 wl_27 vdd gnd cell_6t
Xbit_r28_c214 bl_214 br_214 wl_28 vdd gnd cell_6t
Xbit_r29_c214 bl_214 br_214 wl_29 vdd gnd cell_6t
Xbit_r30_c214 bl_214 br_214 wl_30 vdd gnd cell_6t
Xbit_r31_c214 bl_214 br_214 wl_31 vdd gnd cell_6t
Xbit_r32_c214 bl_214 br_214 wl_32 vdd gnd cell_6t
Xbit_r33_c214 bl_214 br_214 wl_33 vdd gnd cell_6t
Xbit_r34_c214 bl_214 br_214 wl_34 vdd gnd cell_6t
Xbit_r35_c214 bl_214 br_214 wl_35 vdd gnd cell_6t
Xbit_r36_c214 bl_214 br_214 wl_36 vdd gnd cell_6t
Xbit_r37_c214 bl_214 br_214 wl_37 vdd gnd cell_6t
Xbit_r38_c214 bl_214 br_214 wl_38 vdd gnd cell_6t
Xbit_r39_c214 bl_214 br_214 wl_39 vdd gnd cell_6t
Xbit_r40_c214 bl_214 br_214 wl_40 vdd gnd cell_6t
Xbit_r41_c214 bl_214 br_214 wl_41 vdd gnd cell_6t
Xbit_r42_c214 bl_214 br_214 wl_42 vdd gnd cell_6t
Xbit_r43_c214 bl_214 br_214 wl_43 vdd gnd cell_6t
Xbit_r44_c214 bl_214 br_214 wl_44 vdd gnd cell_6t
Xbit_r45_c214 bl_214 br_214 wl_45 vdd gnd cell_6t
Xbit_r46_c214 bl_214 br_214 wl_46 vdd gnd cell_6t
Xbit_r47_c214 bl_214 br_214 wl_47 vdd gnd cell_6t
Xbit_r48_c214 bl_214 br_214 wl_48 vdd gnd cell_6t
Xbit_r49_c214 bl_214 br_214 wl_49 vdd gnd cell_6t
Xbit_r50_c214 bl_214 br_214 wl_50 vdd gnd cell_6t
Xbit_r51_c214 bl_214 br_214 wl_51 vdd gnd cell_6t
Xbit_r52_c214 bl_214 br_214 wl_52 vdd gnd cell_6t
Xbit_r53_c214 bl_214 br_214 wl_53 vdd gnd cell_6t
Xbit_r54_c214 bl_214 br_214 wl_54 vdd gnd cell_6t
Xbit_r55_c214 bl_214 br_214 wl_55 vdd gnd cell_6t
Xbit_r56_c214 bl_214 br_214 wl_56 vdd gnd cell_6t
Xbit_r57_c214 bl_214 br_214 wl_57 vdd gnd cell_6t
Xbit_r58_c214 bl_214 br_214 wl_58 vdd gnd cell_6t
Xbit_r59_c214 bl_214 br_214 wl_59 vdd gnd cell_6t
Xbit_r60_c214 bl_214 br_214 wl_60 vdd gnd cell_6t
Xbit_r61_c214 bl_214 br_214 wl_61 vdd gnd cell_6t
Xbit_r62_c214 bl_214 br_214 wl_62 vdd gnd cell_6t
Xbit_r63_c214 bl_214 br_214 wl_63 vdd gnd cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd cell_6t
Xbit_r1_c215 bl_215 br_215 wl_1 vdd gnd cell_6t
Xbit_r2_c215 bl_215 br_215 wl_2 vdd gnd cell_6t
Xbit_r3_c215 bl_215 br_215 wl_3 vdd gnd cell_6t
Xbit_r4_c215 bl_215 br_215 wl_4 vdd gnd cell_6t
Xbit_r5_c215 bl_215 br_215 wl_5 vdd gnd cell_6t
Xbit_r6_c215 bl_215 br_215 wl_6 vdd gnd cell_6t
Xbit_r7_c215 bl_215 br_215 wl_7 vdd gnd cell_6t
Xbit_r8_c215 bl_215 br_215 wl_8 vdd gnd cell_6t
Xbit_r9_c215 bl_215 br_215 wl_9 vdd gnd cell_6t
Xbit_r10_c215 bl_215 br_215 wl_10 vdd gnd cell_6t
Xbit_r11_c215 bl_215 br_215 wl_11 vdd gnd cell_6t
Xbit_r12_c215 bl_215 br_215 wl_12 vdd gnd cell_6t
Xbit_r13_c215 bl_215 br_215 wl_13 vdd gnd cell_6t
Xbit_r14_c215 bl_215 br_215 wl_14 vdd gnd cell_6t
Xbit_r15_c215 bl_215 br_215 wl_15 vdd gnd cell_6t
Xbit_r16_c215 bl_215 br_215 wl_16 vdd gnd cell_6t
Xbit_r17_c215 bl_215 br_215 wl_17 vdd gnd cell_6t
Xbit_r18_c215 bl_215 br_215 wl_18 vdd gnd cell_6t
Xbit_r19_c215 bl_215 br_215 wl_19 vdd gnd cell_6t
Xbit_r20_c215 bl_215 br_215 wl_20 vdd gnd cell_6t
Xbit_r21_c215 bl_215 br_215 wl_21 vdd gnd cell_6t
Xbit_r22_c215 bl_215 br_215 wl_22 vdd gnd cell_6t
Xbit_r23_c215 bl_215 br_215 wl_23 vdd gnd cell_6t
Xbit_r24_c215 bl_215 br_215 wl_24 vdd gnd cell_6t
Xbit_r25_c215 bl_215 br_215 wl_25 vdd gnd cell_6t
Xbit_r26_c215 bl_215 br_215 wl_26 vdd gnd cell_6t
Xbit_r27_c215 bl_215 br_215 wl_27 vdd gnd cell_6t
Xbit_r28_c215 bl_215 br_215 wl_28 vdd gnd cell_6t
Xbit_r29_c215 bl_215 br_215 wl_29 vdd gnd cell_6t
Xbit_r30_c215 bl_215 br_215 wl_30 vdd gnd cell_6t
Xbit_r31_c215 bl_215 br_215 wl_31 vdd gnd cell_6t
Xbit_r32_c215 bl_215 br_215 wl_32 vdd gnd cell_6t
Xbit_r33_c215 bl_215 br_215 wl_33 vdd gnd cell_6t
Xbit_r34_c215 bl_215 br_215 wl_34 vdd gnd cell_6t
Xbit_r35_c215 bl_215 br_215 wl_35 vdd gnd cell_6t
Xbit_r36_c215 bl_215 br_215 wl_36 vdd gnd cell_6t
Xbit_r37_c215 bl_215 br_215 wl_37 vdd gnd cell_6t
Xbit_r38_c215 bl_215 br_215 wl_38 vdd gnd cell_6t
Xbit_r39_c215 bl_215 br_215 wl_39 vdd gnd cell_6t
Xbit_r40_c215 bl_215 br_215 wl_40 vdd gnd cell_6t
Xbit_r41_c215 bl_215 br_215 wl_41 vdd gnd cell_6t
Xbit_r42_c215 bl_215 br_215 wl_42 vdd gnd cell_6t
Xbit_r43_c215 bl_215 br_215 wl_43 vdd gnd cell_6t
Xbit_r44_c215 bl_215 br_215 wl_44 vdd gnd cell_6t
Xbit_r45_c215 bl_215 br_215 wl_45 vdd gnd cell_6t
Xbit_r46_c215 bl_215 br_215 wl_46 vdd gnd cell_6t
Xbit_r47_c215 bl_215 br_215 wl_47 vdd gnd cell_6t
Xbit_r48_c215 bl_215 br_215 wl_48 vdd gnd cell_6t
Xbit_r49_c215 bl_215 br_215 wl_49 vdd gnd cell_6t
Xbit_r50_c215 bl_215 br_215 wl_50 vdd gnd cell_6t
Xbit_r51_c215 bl_215 br_215 wl_51 vdd gnd cell_6t
Xbit_r52_c215 bl_215 br_215 wl_52 vdd gnd cell_6t
Xbit_r53_c215 bl_215 br_215 wl_53 vdd gnd cell_6t
Xbit_r54_c215 bl_215 br_215 wl_54 vdd gnd cell_6t
Xbit_r55_c215 bl_215 br_215 wl_55 vdd gnd cell_6t
Xbit_r56_c215 bl_215 br_215 wl_56 vdd gnd cell_6t
Xbit_r57_c215 bl_215 br_215 wl_57 vdd gnd cell_6t
Xbit_r58_c215 bl_215 br_215 wl_58 vdd gnd cell_6t
Xbit_r59_c215 bl_215 br_215 wl_59 vdd gnd cell_6t
Xbit_r60_c215 bl_215 br_215 wl_60 vdd gnd cell_6t
Xbit_r61_c215 bl_215 br_215 wl_61 vdd gnd cell_6t
Xbit_r62_c215 bl_215 br_215 wl_62 vdd gnd cell_6t
Xbit_r63_c215 bl_215 br_215 wl_63 vdd gnd cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd cell_6t
Xbit_r1_c216 bl_216 br_216 wl_1 vdd gnd cell_6t
Xbit_r2_c216 bl_216 br_216 wl_2 vdd gnd cell_6t
Xbit_r3_c216 bl_216 br_216 wl_3 vdd gnd cell_6t
Xbit_r4_c216 bl_216 br_216 wl_4 vdd gnd cell_6t
Xbit_r5_c216 bl_216 br_216 wl_5 vdd gnd cell_6t
Xbit_r6_c216 bl_216 br_216 wl_6 vdd gnd cell_6t
Xbit_r7_c216 bl_216 br_216 wl_7 vdd gnd cell_6t
Xbit_r8_c216 bl_216 br_216 wl_8 vdd gnd cell_6t
Xbit_r9_c216 bl_216 br_216 wl_9 vdd gnd cell_6t
Xbit_r10_c216 bl_216 br_216 wl_10 vdd gnd cell_6t
Xbit_r11_c216 bl_216 br_216 wl_11 vdd gnd cell_6t
Xbit_r12_c216 bl_216 br_216 wl_12 vdd gnd cell_6t
Xbit_r13_c216 bl_216 br_216 wl_13 vdd gnd cell_6t
Xbit_r14_c216 bl_216 br_216 wl_14 vdd gnd cell_6t
Xbit_r15_c216 bl_216 br_216 wl_15 vdd gnd cell_6t
Xbit_r16_c216 bl_216 br_216 wl_16 vdd gnd cell_6t
Xbit_r17_c216 bl_216 br_216 wl_17 vdd gnd cell_6t
Xbit_r18_c216 bl_216 br_216 wl_18 vdd gnd cell_6t
Xbit_r19_c216 bl_216 br_216 wl_19 vdd gnd cell_6t
Xbit_r20_c216 bl_216 br_216 wl_20 vdd gnd cell_6t
Xbit_r21_c216 bl_216 br_216 wl_21 vdd gnd cell_6t
Xbit_r22_c216 bl_216 br_216 wl_22 vdd gnd cell_6t
Xbit_r23_c216 bl_216 br_216 wl_23 vdd gnd cell_6t
Xbit_r24_c216 bl_216 br_216 wl_24 vdd gnd cell_6t
Xbit_r25_c216 bl_216 br_216 wl_25 vdd gnd cell_6t
Xbit_r26_c216 bl_216 br_216 wl_26 vdd gnd cell_6t
Xbit_r27_c216 bl_216 br_216 wl_27 vdd gnd cell_6t
Xbit_r28_c216 bl_216 br_216 wl_28 vdd gnd cell_6t
Xbit_r29_c216 bl_216 br_216 wl_29 vdd gnd cell_6t
Xbit_r30_c216 bl_216 br_216 wl_30 vdd gnd cell_6t
Xbit_r31_c216 bl_216 br_216 wl_31 vdd gnd cell_6t
Xbit_r32_c216 bl_216 br_216 wl_32 vdd gnd cell_6t
Xbit_r33_c216 bl_216 br_216 wl_33 vdd gnd cell_6t
Xbit_r34_c216 bl_216 br_216 wl_34 vdd gnd cell_6t
Xbit_r35_c216 bl_216 br_216 wl_35 vdd gnd cell_6t
Xbit_r36_c216 bl_216 br_216 wl_36 vdd gnd cell_6t
Xbit_r37_c216 bl_216 br_216 wl_37 vdd gnd cell_6t
Xbit_r38_c216 bl_216 br_216 wl_38 vdd gnd cell_6t
Xbit_r39_c216 bl_216 br_216 wl_39 vdd gnd cell_6t
Xbit_r40_c216 bl_216 br_216 wl_40 vdd gnd cell_6t
Xbit_r41_c216 bl_216 br_216 wl_41 vdd gnd cell_6t
Xbit_r42_c216 bl_216 br_216 wl_42 vdd gnd cell_6t
Xbit_r43_c216 bl_216 br_216 wl_43 vdd gnd cell_6t
Xbit_r44_c216 bl_216 br_216 wl_44 vdd gnd cell_6t
Xbit_r45_c216 bl_216 br_216 wl_45 vdd gnd cell_6t
Xbit_r46_c216 bl_216 br_216 wl_46 vdd gnd cell_6t
Xbit_r47_c216 bl_216 br_216 wl_47 vdd gnd cell_6t
Xbit_r48_c216 bl_216 br_216 wl_48 vdd gnd cell_6t
Xbit_r49_c216 bl_216 br_216 wl_49 vdd gnd cell_6t
Xbit_r50_c216 bl_216 br_216 wl_50 vdd gnd cell_6t
Xbit_r51_c216 bl_216 br_216 wl_51 vdd gnd cell_6t
Xbit_r52_c216 bl_216 br_216 wl_52 vdd gnd cell_6t
Xbit_r53_c216 bl_216 br_216 wl_53 vdd gnd cell_6t
Xbit_r54_c216 bl_216 br_216 wl_54 vdd gnd cell_6t
Xbit_r55_c216 bl_216 br_216 wl_55 vdd gnd cell_6t
Xbit_r56_c216 bl_216 br_216 wl_56 vdd gnd cell_6t
Xbit_r57_c216 bl_216 br_216 wl_57 vdd gnd cell_6t
Xbit_r58_c216 bl_216 br_216 wl_58 vdd gnd cell_6t
Xbit_r59_c216 bl_216 br_216 wl_59 vdd gnd cell_6t
Xbit_r60_c216 bl_216 br_216 wl_60 vdd gnd cell_6t
Xbit_r61_c216 bl_216 br_216 wl_61 vdd gnd cell_6t
Xbit_r62_c216 bl_216 br_216 wl_62 vdd gnd cell_6t
Xbit_r63_c216 bl_216 br_216 wl_63 vdd gnd cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd cell_6t
Xbit_r1_c217 bl_217 br_217 wl_1 vdd gnd cell_6t
Xbit_r2_c217 bl_217 br_217 wl_2 vdd gnd cell_6t
Xbit_r3_c217 bl_217 br_217 wl_3 vdd gnd cell_6t
Xbit_r4_c217 bl_217 br_217 wl_4 vdd gnd cell_6t
Xbit_r5_c217 bl_217 br_217 wl_5 vdd gnd cell_6t
Xbit_r6_c217 bl_217 br_217 wl_6 vdd gnd cell_6t
Xbit_r7_c217 bl_217 br_217 wl_7 vdd gnd cell_6t
Xbit_r8_c217 bl_217 br_217 wl_8 vdd gnd cell_6t
Xbit_r9_c217 bl_217 br_217 wl_9 vdd gnd cell_6t
Xbit_r10_c217 bl_217 br_217 wl_10 vdd gnd cell_6t
Xbit_r11_c217 bl_217 br_217 wl_11 vdd gnd cell_6t
Xbit_r12_c217 bl_217 br_217 wl_12 vdd gnd cell_6t
Xbit_r13_c217 bl_217 br_217 wl_13 vdd gnd cell_6t
Xbit_r14_c217 bl_217 br_217 wl_14 vdd gnd cell_6t
Xbit_r15_c217 bl_217 br_217 wl_15 vdd gnd cell_6t
Xbit_r16_c217 bl_217 br_217 wl_16 vdd gnd cell_6t
Xbit_r17_c217 bl_217 br_217 wl_17 vdd gnd cell_6t
Xbit_r18_c217 bl_217 br_217 wl_18 vdd gnd cell_6t
Xbit_r19_c217 bl_217 br_217 wl_19 vdd gnd cell_6t
Xbit_r20_c217 bl_217 br_217 wl_20 vdd gnd cell_6t
Xbit_r21_c217 bl_217 br_217 wl_21 vdd gnd cell_6t
Xbit_r22_c217 bl_217 br_217 wl_22 vdd gnd cell_6t
Xbit_r23_c217 bl_217 br_217 wl_23 vdd gnd cell_6t
Xbit_r24_c217 bl_217 br_217 wl_24 vdd gnd cell_6t
Xbit_r25_c217 bl_217 br_217 wl_25 vdd gnd cell_6t
Xbit_r26_c217 bl_217 br_217 wl_26 vdd gnd cell_6t
Xbit_r27_c217 bl_217 br_217 wl_27 vdd gnd cell_6t
Xbit_r28_c217 bl_217 br_217 wl_28 vdd gnd cell_6t
Xbit_r29_c217 bl_217 br_217 wl_29 vdd gnd cell_6t
Xbit_r30_c217 bl_217 br_217 wl_30 vdd gnd cell_6t
Xbit_r31_c217 bl_217 br_217 wl_31 vdd gnd cell_6t
Xbit_r32_c217 bl_217 br_217 wl_32 vdd gnd cell_6t
Xbit_r33_c217 bl_217 br_217 wl_33 vdd gnd cell_6t
Xbit_r34_c217 bl_217 br_217 wl_34 vdd gnd cell_6t
Xbit_r35_c217 bl_217 br_217 wl_35 vdd gnd cell_6t
Xbit_r36_c217 bl_217 br_217 wl_36 vdd gnd cell_6t
Xbit_r37_c217 bl_217 br_217 wl_37 vdd gnd cell_6t
Xbit_r38_c217 bl_217 br_217 wl_38 vdd gnd cell_6t
Xbit_r39_c217 bl_217 br_217 wl_39 vdd gnd cell_6t
Xbit_r40_c217 bl_217 br_217 wl_40 vdd gnd cell_6t
Xbit_r41_c217 bl_217 br_217 wl_41 vdd gnd cell_6t
Xbit_r42_c217 bl_217 br_217 wl_42 vdd gnd cell_6t
Xbit_r43_c217 bl_217 br_217 wl_43 vdd gnd cell_6t
Xbit_r44_c217 bl_217 br_217 wl_44 vdd gnd cell_6t
Xbit_r45_c217 bl_217 br_217 wl_45 vdd gnd cell_6t
Xbit_r46_c217 bl_217 br_217 wl_46 vdd gnd cell_6t
Xbit_r47_c217 bl_217 br_217 wl_47 vdd gnd cell_6t
Xbit_r48_c217 bl_217 br_217 wl_48 vdd gnd cell_6t
Xbit_r49_c217 bl_217 br_217 wl_49 vdd gnd cell_6t
Xbit_r50_c217 bl_217 br_217 wl_50 vdd gnd cell_6t
Xbit_r51_c217 bl_217 br_217 wl_51 vdd gnd cell_6t
Xbit_r52_c217 bl_217 br_217 wl_52 vdd gnd cell_6t
Xbit_r53_c217 bl_217 br_217 wl_53 vdd gnd cell_6t
Xbit_r54_c217 bl_217 br_217 wl_54 vdd gnd cell_6t
Xbit_r55_c217 bl_217 br_217 wl_55 vdd gnd cell_6t
Xbit_r56_c217 bl_217 br_217 wl_56 vdd gnd cell_6t
Xbit_r57_c217 bl_217 br_217 wl_57 vdd gnd cell_6t
Xbit_r58_c217 bl_217 br_217 wl_58 vdd gnd cell_6t
Xbit_r59_c217 bl_217 br_217 wl_59 vdd gnd cell_6t
Xbit_r60_c217 bl_217 br_217 wl_60 vdd gnd cell_6t
Xbit_r61_c217 bl_217 br_217 wl_61 vdd gnd cell_6t
Xbit_r62_c217 bl_217 br_217 wl_62 vdd gnd cell_6t
Xbit_r63_c217 bl_217 br_217 wl_63 vdd gnd cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd cell_6t
Xbit_r1_c218 bl_218 br_218 wl_1 vdd gnd cell_6t
Xbit_r2_c218 bl_218 br_218 wl_2 vdd gnd cell_6t
Xbit_r3_c218 bl_218 br_218 wl_3 vdd gnd cell_6t
Xbit_r4_c218 bl_218 br_218 wl_4 vdd gnd cell_6t
Xbit_r5_c218 bl_218 br_218 wl_5 vdd gnd cell_6t
Xbit_r6_c218 bl_218 br_218 wl_6 vdd gnd cell_6t
Xbit_r7_c218 bl_218 br_218 wl_7 vdd gnd cell_6t
Xbit_r8_c218 bl_218 br_218 wl_8 vdd gnd cell_6t
Xbit_r9_c218 bl_218 br_218 wl_9 vdd gnd cell_6t
Xbit_r10_c218 bl_218 br_218 wl_10 vdd gnd cell_6t
Xbit_r11_c218 bl_218 br_218 wl_11 vdd gnd cell_6t
Xbit_r12_c218 bl_218 br_218 wl_12 vdd gnd cell_6t
Xbit_r13_c218 bl_218 br_218 wl_13 vdd gnd cell_6t
Xbit_r14_c218 bl_218 br_218 wl_14 vdd gnd cell_6t
Xbit_r15_c218 bl_218 br_218 wl_15 vdd gnd cell_6t
Xbit_r16_c218 bl_218 br_218 wl_16 vdd gnd cell_6t
Xbit_r17_c218 bl_218 br_218 wl_17 vdd gnd cell_6t
Xbit_r18_c218 bl_218 br_218 wl_18 vdd gnd cell_6t
Xbit_r19_c218 bl_218 br_218 wl_19 vdd gnd cell_6t
Xbit_r20_c218 bl_218 br_218 wl_20 vdd gnd cell_6t
Xbit_r21_c218 bl_218 br_218 wl_21 vdd gnd cell_6t
Xbit_r22_c218 bl_218 br_218 wl_22 vdd gnd cell_6t
Xbit_r23_c218 bl_218 br_218 wl_23 vdd gnd cell_6t
Xbit_r24_c218 bl_218 br_218 wl_24 vdd gnd cell_6t
Xbit_r25_c218 bl_218 br_218 wl_25 vdd gnd cell_6t
Xbit_r26_c218 bl_218 br_218 wl_26 vdd gnd cell_6t
Xbit_r27_c218 bl_218 br_218 wl_27 vdd gnd cell_6t
Xbit_r28_c218 bl_218 br_218 wl_28 vdd gnd cell_6t
Xbit_r29_c218 bl_218 br_218 wl_29 vdd gnd cell_6t
Xbit_r30_c218 bl_218 br_218 wl_30 vdd gnd cell_6t
Xbit_r31_c218 bl_218 br_218 wl_31 vdd gnd cell_6t
Xbit_r32_c218 bl_218 br_218 wl_32 vdd gnd cell_6t
Xbit_r33_c218 bl_218 br_218 wl_33 vdd gnd cell_6t
Xbit_r34_c218 bl_218 br_218 wl_34 vdd gnd cell_6t
Xbit_r35_c218 bl_218 br_218 wl_35 vdd gnd cell_6t
Xbit_r36_c218 bl_218 br_218 wl_36 vdd gnd cell_6t
Xbit_r37_c218 bl_218 br_218 wl_37 vdd gnd cell_6t
Xbit_r38_c218 bl_218 br_218 wl_38 vdd gnd cell_6t
Xbit_r39_c218 bl_218 br_218 wl_39 vdd gnd cell_6t
Xbit_r40_c218 bl_218 br_218 wl_40 vdd gnd cell_6t
Xbit_r41_c218 bl_218 br_218 wl_41 vdd gnd cell_6t
Xbit_r42_c218 bl_218 br_218 wl_42 vdd gnd cell_6t
Xbit_r43_c218 bl_218 br_218 wl_43 vdd gnd cell_6t
Xbit_r44_c218 bl_218 br_218 wl_44 vdd gnd cell_6t
Xbit_r45_c218 bl_218 br_218 wl_45 vdd gnd cell_6t
Xbit_r46_c218 bl_218 br_218 wl_46 vdd gnd cell_6t
Xbit_r47_c218 bl_218 br_218 wl_47 vdd gnd cell_6t
Xbit_r48_c218 bl_218 br_218 wl_48 vdd gnd cell_6t
Xbit_r49_c218 bl_218 br_218 wl_49 vdd gnd cell_6t
Xbit_r50_c218 bl_218 br_218 wl_50 vdd gnd cell_6t
Xbit_r51_c218 bl_218 br_218 wl_51 vdd gnd cell_6t
Xbit_r52_c218 bl_218 br_218 wl_52 vdd gnd cell_6t
Xbit_r53_c218 bl_218 br_218 wl_53 vdd gnd cell_6t
Xbit_r54_c218 bl_218 br_218 wl_54 vdd gnd cell_6t
Xbit_r55_c218 bl_218 br_218 wl_55 vdd gnd cell_6t
Xbit_r56_c218 bl_218 br_218 wl_56 vdd gnd cell_6t
Xbit_r57_c218 bl_218 br_218 wl_57 vdd gnd cell_6t
Xbit_r58_c218 bl_218 br_218 wl_58 vdd gnd cell_6t
Xbit_r59_c218 bl_218 br_218 wl_59 vdd gnd cell_6t
Xbit_r60_c218 bl_218 br_218 wl_60 vdd gnd cell_6t
Xbit_r61_c218 bl_218 br_218 wl_61 vdd gnd cell_6t
Xbit_r62_c218 bl_218 br_218 wl_62 vdd gnd cell_6t
Xbit_r63_c218 bl_218 br_218 wl_63 vdd gnd cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd cell_6t
Xbit_r1_c219 bl_219 br_219 wl_1 vdd gnd cell_6t
Xbit_r2_c219 bl_219 br_219 wl_2 vdd gnd cell_6t
Xbit_r3_c219 bl_219 br_219 wl_3 vdd gnd cell_6t
Xbit_r4_c219 bl_219 br_219 wl_4 vdd gnd cell_6t
Xbit_r5_c219 bl_219 br_219 wl_5 vdd gnd cell_6t
Xbit_r6_c219 bl_219 br_219 wl_6 vdd gnd cell_6t
Xbit_r7_c219 bl_219 br_219 wl_7 vdd gnd cell_6t
Xbit_r8_c219 bl_219 br_219 wl_8 vdd gnd cell_6t
Xbit_r9_c219 bl_219 br_219 wl_9 vdd gnd cell_6t
Xbit_r10_c219 bl_219 br_219 wl_10 vdd gnd cell_6t
Xbit_r11_c219 bl_219 br_219 wl_11 vdd gnd cell_6t
Xbit_r12_c219 bl_219 br_219 wl_12 vdd gnd cell_6t
Xbit_r13_c219 bl_219 br_219 wl_13 vdd gnd cell_6t
Xbit_r14_c219 bl_219 br_219 wl_14 vdd gnd cell_6t
Xbit_r15_c219 bl_219 br_219 wl_15 vdd gnd cell_6t
Xbit_r16_c219 bl_219 br_219 wl_16 vdd gnd cell_6t
Xbit_r17_c219 bl_219 br_219 wl_17 vdd gnd cell_6t
Xbit_r18_c219 bl_219 br_219 wl_18 vdd gnd cell_6t
Xbit_r19_c219 bl_219 br_219 wl_19 vdd gnd cell_6t
Xbit_r20_c219 bl_219 br_219 wl_20 vdd gnd cell_6t
Xbit_r21_c219 bl_219 br_219 wl_21 vdd gnd cell_6t
Xbit_r22_c219 bl_219 br_219 wl_22 vdd gnd cell_6t
Xbit_r23_c219 bl_219 br_219 wl_23 vdd gnd cell_6t
Xbit_r24_c219 bl_219 br_219 wl_24 vdd gnd cell_6t
Xbit_r25_c219 bl_219 br_219 wl_25 vdd gnd cell_6t
Xbit_r26_c219 bl_219 br_219 wl_26 vdd gnd cell_6t
Xbit_r27_c219 bl_219 br_219 wl_27 vdd gnd cell_6t
Xbit_r28_c219 bl_219 br_219 wl_28 vdd gnd cell_6t
Xbit_r29_c219 bl_219 br_219 wl_29 vdd gnd cell_6t
Xbit_r30_c219 bl_219 br_219 wl_30 vdd gnd cell_6t
Xbit_r31_c219 bl_219 br_219 wl_31 vdd gnd cell_6t
Xbit_r32_c219 bl_219 br_219 wl_32 vdd gnd cell_6t
Xbit_r33_c219 bl_219 br_219 wl_33 vdd gnd cell_6t
Xbit_r34_c219 bl_219 br_219 wl_34 vdd gnd cell_6t
Xbit_r35_c219 bl_219 br_219 wl_35 vdd gnd cell_6t
Xbit_r36_c219 bl_219 br_219 wl_36 vdd gnd cell_6t
Xbit_r37_c219 bl_219 br_219 wl_37 vdd gnd cell_6t
Xbit_r38_c219 bl_219 br_219 wl_38 vdd gnd cell_6t
Xbit_r39_c219 bl_219 br_219 wl_39 vdd gnd cell_6t
Xbit_r40_c219 bl_219 br_219 wl_40 vdd gnd cell_6t
Xbit_r41_c219 bl_219 br_219 wl_41 vdd gnd cell_6t
Xbit_r42_c219 bl_219 br_219 wl_42 vdd gnd cell_6t
Xbit_r43_c219 bl_219 br_219 wl_43 vdd gnd cell_6t
Xbit_r44_c219 bl_219 br_219 wl_44 vdd gnd cell_6t
Xbit_r45_c219 bl_219 br_219 wl_45 vdd gnd cell_6t
Xbit_r46_c219 bl_219 br_219 wl_46 vdd gnd cell_6t
Xbit_r47_c219 bl_219 br_219 wl_47 vdd gnd cell_6t
Xbit_r48_c219 bl_219 br_219 wl_48 vdd gnd cell_6t
Xbit_r49_c219 bl_219 br_219 wl_49 vdd gnd cell_6t
Xbit_r50_c219 bl_219 br_219 wl_50 vdd gnd cell_6t
Xbit_r51_c219 bl_219 br_219 wl_51 vdd gnd cell_6t
Xbit_r52_c219 bl_219 br_219 wl_52 vdd gnd cell_6t
Xbit_r53_c219 bl_219 br_219 wl_53 vdd gnd cell_6t
Xbit_r54_c219 bl_219 br_219 wl_54 vdd gnd cell_6t
Xbit_r55_c219 bl_219 br_219 wl_55 vdd gnd cell_6t
Xbit_r56_c219 bl_219 br_219 wl_56 vdd gnd cell_6t
Xbit_r57_c219 bl_219 br_219 wl_57 vdd gnd cell_6t
Xbit_r58_c219 bl_219 br_219 wl_58 vdd gnd cell_6t
Xbit_r59_c219 bl_219 br_219 wl_59 vdd gnd cell_6t
Xbit_r60_c219 bl_219 br_219 wl_60 vdd gnd cell_6t
Xbit_r61_c219 bl_219 br_219 wl_61 vdd gnd cell_6t
Xbit_r62_c219 bl_219 br_219 wl_62 vdd gnd cell_6t
Xbit_r63_c219 bl_219 br_219 wl_63 vdd gnd cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd cell_6t
Xbit_r1_c220 bl_220 br_220 wl_1 vdd gnd cell_6t
Xbit_r2_c220 bl_220 br_220 wl_2 vdd gnd cell_6t
Xbit_r3_c220 bl_220 br_220 wl_3 vdd gnd cell_6t
Xbit_r4_c220 bl_220 br_220 wl_4 vdd gnd cell_6t
Xbit_r5_c220 bl_220 br_220 wl_5 vdd gnd cell_6t
Xbit_r6_c220 bl_220 br_220 wl_6 vdd gnd cell_6t
Xbit_r7_c220 bl_220 br_220 wl_7 vdd gnd cell_6t
Xbit_r8_c220 bl_220 br_220 wl_8 vdd gnd cell_6t
Xbit_r9_c220 bl_220 br_220 wl_9 vdd gnd cell_6t
Xbit_r10_c220 bl_220 br_220 wl_10 vdd gnd cell_6t
Xbit_r11_c220 bl_220 br_220 wl_11 vdd gnd cell_6t
Xbit_r12_c220 bl_220 br_220 wl_12 vdd gnd cell_6t
Xbit_r13_c220 bl_220 br_220 wl_13 vdd gnd cell_6t
Xbit_r14_c220 bl_220 br_220 wl_14 vdd gnd cell_6t
Xbit_r15_c220 bl_220 br_220 wl_15 vdd gnd cell_6t
Xbit_r16_c220 bl_220 br_220 wl_16 vdd gnd cell_6t
Xbit_r17_c220 bl_220 br_220 wl_17 vdd gnd cell_6t
Xbit_r18_c220 bl_220 br_220 wl_18 vdd gnd cell_6t
Xbit_r19_c220 bl_220 br_220 wl_19 vdd gnd cell_6t
Xbit_r20_c220 bl_220 br_220 wl_20 vdd gnd cell_6t
Xbit_r21_c220 bl_220 br_220 wl_21 vdd gnd cell_6t
Xbit_r22_c220 bl_220 br_220 wl_22 vdd gnd cell_6t
Xbit_r23_c220 bl_220 br_220 wl_23 vdd gnd cell_6t
Xbit_r24_c220 bl_220 br_220 wl_24 vdd gnd cell_6t
Xbit_r25_c220 bl_220 br_220 wl_25 vdd gnd cell_6t
Xbit_r26_c220 bl_220 br_220 wl_26 vdd gnd cell_6t
Xbit_r27_c220 bl_220 br_220 wl_27 vdd gnd cell_6t
Xbit_r28_c220 bl_220 br_220 wl_28 vdd gnd cell_6t
Xbit_r29_c220 bl_220 br_220 wl_29 vdd gnd cell_6t
Xbit_r30_c220 bl_220 br_220 wl_30 vdd gnd cell_6t
Xbit_r31_c220 bl_220 br_220 wl_31 vdd gnd cell_6t
Xbit_r32_c220 bl_220 br_220 wl_32 vdd gnd cell_6t
Xbit_r33_c220 bl_220 br_220 wl_33 vdd gnd cell_6t
Xbit_r34_c220 bl_220 br_220 wl_34 vdd gnd cell_6t
Xbit_r35_c220 bl_220 br_220 wl_35 vdd gnd cell_6t
Xbit_r36_c220 bl_220 br_220 wl_36 vdd gnd cell_6t
Xbit_r37_c220 bl_220 br_220 wl_37 vdd gnd cell_6t
Xbit_r38_c220 bl_220 br_220 wl_38 vdd gnd cell_6t
Xbit_r39_c220 bl_220 br_220 wl_39 vdd gnd cell_6t
Xbit_r40_c220 bl_220 br_220 wl_40 vdd gnd cell_6t
Xbit_r41_c220 bl_220 br_220 wl_41 vdd gnd cell_6t
Xbit_r42_c220 bl_220 br_220 wl_42 vdd gnd cell_6t
Xbit_r43_c220 bl_220 br_220 wl_43 vdd gnd cell_6t
Xbit_r44_c220 bl_220 br_220 wl_44 vdd gnd cell_6t
Xbit_r45_c220 bl_220 br_220 wl_45 vdd gnd cell_6t
Xbit_r46_c220 bl_220 br_220 wl_46 vdd gnd cell_6t
Xbit_r47_c220 bl_220 br_220 wl_47 vdd gnd cell_6t
Xbit_r48_c220 bl_220 br_220 wl_48 vdd gnd cell_6t
Xbit_r49_c220 bl_220 br_220 wl_49 vdd gnd cell_6t
Xbit_r50_c220 bl_220 br_220 wl_50 vdd gnd cell_6t
Xbit_r51_c220 bl_220 br_220 wl_51 vdd gnd cell_6t
Xbit_r52_c220 bl_220 br_220 wl_52 vdd gnd cell_6t
Xbit_r53_c220 bl_220 br_220 wl_53 vdd gnd cell_6t
Xbit_r54_c220 bl_220 br_220 wl_54 vdd gnd cell_6t
Xbit_r55_c220 bl_220 br_220 wl_55 vdd gnd cell_6t
Xbit_r56_c220 bl_220 br_220 wl_56 vdd gnd cell_6t
Xbit_r57_c220 bl_220 br_220 wl_57 vdd gnd cell_6t
Xbit_r58_c220 bl_220 br_220 wl_58 vdd gnd cell_6t
Xbit_r59_c220 bl_220 br_220 wl_59 vdd gnd cell_6t
Xbit_r60_c220 bl_220 br_220 wl_60 vdd gnd cell_6t
Xbit_r61_c220 bl_220 br_220 wl_61 vdd gnd cell_6t
Xbit_r62_c220 bl_220 br_220 wl_62 vdd gnd cell_6t
Xbit_r63_c220 bl_220 br_220 wl_63 vdd gnd cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd cell_6t
Xbit_r1_c221 bl_221 br_221 wl_1 vdd gnd cell_6t
Xbit_r2_c221 bl_221 br_221 wl_2 vdd gnd cell_6t
Xbit_r3_c221 bl_221 br_221 wl_3 vdd gnd cell_6t
Xbit_r4_c221 bl_221 br_221 wl_4 vdd gnd cell_6t
Xbit_r5_c221 bl_221 br_221 wl_5 vdd gnd cell_6t
Xbit_r6_c221 bl_221 br_221 wl_6 vdd gnd cell_6t
Xbit_r7_c221 bl_221 br_221 wl_7 vdd gnd cell_6t
Xbit_r8_c221 bl_221 br_221 wl_8 vdd gnd cell_6t
Xbit_r9_c221 bl_221 br_221 wl_9 vdd gnd cell_6t
Xbit_r10_c221 bl_221 br_221 wl_10 vdd gnd cell_6t
Xbit_r11_c221 bl_221 br_221 wl_11 vdd gnd cell_6t
Xbit_r12_c221 bl_221 br_221 wl_12 vdd gnd cell_6t
Xbit_r13_c221 bl_221 br_221 wl_13 vdd gnd cell_6t
Xbit_r14_c221 bl_221 br_221 wl_14 vdd gnd cell_6t
Xbit_r15_c221 bl_221 br_221 wl_15 vdd gnd cell_6t
Xbit_r16_c221 bl_221 br_221 wl_16 vdd gnd cell_6t
Xbit_r17_c221 bl_221 br_221 wl_17 vdd gnd cell_6t
Xbit_r18_c221 bl_221 br_221 wl_18 vdd gnd cell_6t
Xbit_r19_c221 bl_221 br_221 wl_19 vdd gnd cell_6t
Xbit_r20_c221 bl_221 br_221 wl_20 vdd gnd cell_6t
Xbit_r21_c221 bl_221 br_221 wl_21 vdd gnd cell_6t
Xbit_r22_c221 bl_221 br_221 wl_22 vdd gnd cell_6t
Xbit_r23_c221 bl_221 br_221 wl_23 vdd gnd cell_6t
Xbit_r24_c221 bl_221 br_221 wl_24 vdd gnd cell_6t
Xbit_r25_c221 bl_221 br_221 wl_25 vdd gnd cell_6t
Xbit_r26_c221 bl_221 br_221 wl_26 vdd gnd cell_6t
Xbit_r27_c221 bl_221 br_221 wl_27 vdd gnd cell_6t
Xbit_r28_c221 bl_221 br_221 wl_28 vdd gnd cell_6t
Xbit_r29_c221 bl_221 br_221 wl_29 vdd gnd cell_6t
Xbit_r30_c221 bl_221 br_221 wl_30 vdd gnd cell_6t
Xbit_r31_c221 bl_221 br_221 wl_31 vdd gnd cell_6t
Xbit_r32_c221 bl_221 br_221 wl_32 vdd gnd cell_6t
Xbit_r33_c221 bl_221 br_221 wl_33 vdd gnd cell_6t
Xbit_r34_c221 bl_221 br_221 wl_34 vdd gnd cell_6t
Xbit_r35_c221 bl_221 br_221 wl_35 vdd gnd cell_6t
Xbit_r36_c221 bl_221 br_221 wl_36 vdd gnd cell_6t
Xbit_r37_c221 bl_221 br_221 wl_37 vdd gnd cell_6t
Xbit_r38_c221 bl_221 br_221 wl_38 vdd gnd cell_6t
Xbit_r39_c221 bl_221 br_221 wl_39 vdd gnd cell_6t
Xbit_r40_c221 bl_221 br_221 wl_40 vdd gnd cell_6t
Xbit_r41_c221 bl_221 br_221 wl_41 vdd gnd cell_6t
Xbit_r42_c221 bl_221 br_221 wl_42 vdd gnd cell_6t
Xbit_r43_c221 bl_221 br_221 wl_43 vdd gnd cell_6t
Xbit_r44_c221 bl_221 br_221 wl_44 vdd gnd cell_6t
Xbit_r45_c221 bl_221 br_221 wl_45 vdd gnd cell_6t
Xbit_r46_c221 bl_221 br_221 wl_46 vdd gnd cell_6t
Xbit_r47_c221 bl_221 br_221 wl_47 vdd gnd cell_6t
Xbit_r48_c221 bl_221 br_221 wl_48 vdd gnd cell_6t
Xbit_r49_c221 bl_221 br_221 wl_49 vdd gnd cell_6t
Xbit_r50_c221 bl_221 br_221 wl_50 vdd gnd cell_6t
Xbit_r51_c221 bl_221 br_221 wl_51 vdd gnd cell_6t
Xbit_r52_c221 bl_221 br_221 wl_52 vdd gnd cell_6t
Xbit_r53_c221 bl_221 br_221 wl_53 vdd gnd cell_6t
Xbit_r54_c221 bl_221 br_221 wl_54 vdd gnd cell_6t
Xbit_r55_c221 bl_221 br_221 wl_55 vdd gnd cell_6t
Xbit_r56_c221 bl_221 br_221 wl_56 vdd gnd cell_6t
Xbit_r57_c221 bl_221 br_221 wl_57 vdd gnd cell_6t
Xbit_r58_c221 bl_221 br_221 wl_58 vdd gnd cell_6t
Xbit_r59_c221 bl_221 br_221 wl_59 vdd gnd cell_6t
Xbit_r60_c221 bl_221 br_221 wl_60 vdd gnd cell_6t
Xbit_r61_c221 bl_221 br_221 wl_61 vdd gnd cell_6t
Xbit_r62_c221 bl_221 br_221 wl_62 vdd gnd cell_6t
Xbit_r63_c221 bl_221 br_221 wl_63 vdd gnd cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd cell_6t
Xbit_r1_c222 bl_222 br_222 wl_1 vdd gnd cell_6t
Xbit_r2_c222 bl_222 br_222 wl_2 vdd gnd cell_6t
Xbit_r3_c222 bl_222 br_222 wl_3 vdd gnd cell_6t
Xbit_r4_c222 bl_222 br_222 wl_4 vdd gnd cell_6t
Xbit_r5_c222 bl_222 br_222 wl_5 vdd gnd cell_6t
Xbit_r6_c222 bl_222 br_222 wl_6 vdd gnd cell_6t
Xbit_r7_c222 bl_222 br_222 wl_7 vdd gnd cell_6t
Xbit_r8_c222 bl_222 br_222 wl_8 vdd gnd cell_6t
Xbit_r9_c222 bl_222 br_222 wl_9 vdd gnd cell_6t
Xbit_r10_c222 bl_222 br_222 wl_10 vdd gnd cell_6t
Xbit_r11_c222 bl_222 br_222 wl_11 vdd gnd cell_6t
Xbit_r12_c222 bl_222 br_222 wl_12 vdd gnd cell_6t
Xbit_r13_c222 bl_222 br_222 wl_13 vdd gnd cell_6t
Xbit_r14_c222 bl_222 br_222 wl_14 vdd gnd cell_6t
Xbit_r15_c222 bl_222 br_222 wl_15 vdd gnd cell_6t
Xbit_r16_c222 bl_222 br_222 wl_16 vdd gnd cell_6t
Xbit_r17_c222 bl_222 br_222 wl_17 vdd gnd cell_6t
Xbit_r18_c222 bl_222 br_222 wl_18 vdd gnd cell_6t
Xbit_r19_c222 bl_222 br_222 wl_19 vdd gnd cell_6t
Xbit_r20_c222 bl_222 br_222 wl_20 vdd gnd cell_6t
Xbit_r21_c222 bl_222 br_222 wl_21 vdd gnd cell_6t
Xbit_r22_c222 bl_222 br_222 wl_22 vdd gnd cell_6t
Xbit_r23_c222 bl_222 br_222 wl_23 vdd gnd cell_6t
Xbit_r24_c222 bl_222 br_222 wl_24 vdd gnd cell_6t
Xbit_r25_c222 bl_222 br_222 wl_25 vdd gnd cell_6t
Xbit_r26_c222 bl_222 br_222 wl_26 vdd gnd cell_6t
Xbit_r27_c222 bl_222 br_222 wl_27 vdd gnd cell_6t
Xbit_r28_c222 bl_222 br_222 wl_28 vdd gnd cell_6t
Xbit_r29_c222 bl_222 br_222 wl_29 vdd gnd cell_6t
Xbit_r30_c222 bl_222 br_222 wl_30 vdd gnd cell_6t
Xbit_r31_c222 bl_222 br_222 wl_31 vdd gnd cell_6t
Xbit_r32_c222 bl_222 br_222 wl_32 vdd gnd cell_6t
Xbit_r33_c222 bl_222 br_222 wl_33 vdd gnd cell_6t
Xbit_r34_c222 bl_222 br_222 wl_34 vdd gnd cell_6t
Xbit_r35_c222 bl_222 br_222 wl_35 vdd gnd cell_6t
Xbit_r36_c222 bl_222 br_222 wl_36 vdd gnd cell_6t
Xbit_r37_c222 bl_222 br_222 wl_37 vdd gnd cell_6t
Xbit_r38_c222 bl_222 br_222 wl_38 vdd gnd cell_6t
Xbit_r39_c222 bl_222 br_222 wl_39 vdd gnd cell_6t
Xbit_r40_c222 bl_222 br_222 wl_40 vdd gnd cell_6t
Xbit_r41_c222 bl_222 br_222 wl_41 vdd gnd cell_6t
Xbit_r42_c222 bl_222 br_222 wl_42 vdd gnd cell_6t
Xbit_r43_c222 bl_222 br_222 wl_43 vdd gnd cell_6t
Xbit_r44_c222 bl_222 br_222 wl_44 vdd gnd cell_6t
Xbit_r45_c222 bl_222 br_222 wl_45 vdd gnd cell_6t
Xbit_r46_c222 bl_222 br_222 wl_46 vdd gnd cell_6t
Xbit_r47_c222 bl_222 br_222 wl_47 vdd gnd cell_6t
Xbit_r48_c222 bl_222 br_222 wl_48 vdd gnd cell_6t
Xbit_r49_c222 bl_222 br_222 wl_49 vdd gnd cell_6t
Xbit_r50_c222 bl_222 br_222 wl_50 vdd gnd cell_6t
Xbit_r51_c222 bl_222 br_222 wl_51 vdd gnd cell_6t
Xbit_r52_c222 bl_222 br_222 wl_52 vdd gnd cell_6t
Xbit_r53_c222 bl_222 br_222 wl_53 vdd gnd cell_6t
Xbit_r54_c222 bl_222 br_222 wl_54 vdd gnd cell_6t
Xbit_r55_c222 bl_222 br_222 wl_55 vdd gnd cell_6t
Xbit_r56_c222 bl_222 br_222 wl_56 vdd gnd cell_6t
Xbit_r57_c222 bl_222 br_222 wl_57 vdd gnd cell_6t
Xbit_r58_c222 bl_222 br_222 wl_58 vdd gnd cell_6t
Xbit_r59_c222 bl_222 br_222 wl_59 vdd gnd cell_6t
Xbit_r60_c222 bl_222 br_222 wl_60 vdd gnd cell_6t
Xbit_r61_c222 bl_222 br_222 wl_61 vdd gnd cell_6t
Xbit_r62_c222 bl_222 br_222 wl_62 vdd gnd cell_6t
Xbit_r63_c222 bl_222 br_222 wl_63 vdd gnd cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd cell_6t
Xbit_r1_c223 bl_223 br_223 wl_1 vdd gnd cell_6t
Xbit_r2_c223 bl_223 br_223 wl_2 vdd gnd cell_6t
Xbit_r3_c223 bl_223 br_223 wl_3 vdd gnd cell_6t
Xbit_r4_c223 bl_223 br_223 wl_4 vdd gnd cell_6t
Xbit_r5_c223 bl_223 br_223 wl_5 vdd gnd cell_6t
Xbit_r6_c223 bl_223 br_223 wl_6 vdd gnd cell_6t
Xbit_r7_c223 bl_223 br_223 wl_7 vdd gnd cell_6t
Xbit_r8_c223 bl_223 br_223 wl_8 vdd gnd cell_6t
Xbit_r9_c223 bl_223 br_223 wl_9 vdd gnd cell_6t
Xbit_r10_c223 bl_223 br_223 wl_10 vdd gnd cell_6t
Xbit_r11_c223 bl_223 br_223 wl_11 vdd gnd cell_6t
Xbit_r12_c223 bl_223 br_223 wl_12 vdd gnd cell_6t
Xbit_r13_c223 bl_223 br_223 wl_13 vdd gnd cell_6t
Xbit_r14_c223 bl_223 br_223 wl_14 vdd gnd cell_6t
Xbit_r15_c223 bl_223 br_223 wl_15 vdd gnd cell_6t
Xbit_r16_c223 bl_223 br_223 wl_16 vdd gnd cell_6t
Xbit_r17_c223 bl_223 br_223 wl_17 vdd gnd cell_6t
Xbit_r18_c223 bl_223 br_223 wl_18 vdd gnd cell_6t
Xbit_r19_c223 bl_223 br_223 wl_19 vdd gnd cell_6t
Xbit_r20_c223 bl_223 br_223 wl_20 vdd gnd cell_6t
Xbit_r21_c223 bl_223 br_223 wl_21 vdd gnd cell_6t
Xbit_r22_c223 bl_223 br_223 wl_22 vdd gnd cell_6t
Xbit_r23_c223 bl_223 br_223 wl_23 vdd gnd cell_6t
Xbit_r24_c223 bl_223 br_223 wl_24 vdd gnd cell_6t
Xbit_r25_c223 bl_223 br_223 wl_25 vdd gnd cell_6t
Xbit_r26_c223 bl_223 br_223 wl_26 vdd gnd cell_6t
Xbit_r27_c223 bl_223 br_223 wl_27 vdd gnd cell_6t
Xbit_r28_c223 bl_223 br_223 wl_28 vdd gnd cell_6t
Xbit_r29_c223 bl_223 br_223 wl_29 vdd gnd cell_6t
Xbit_r30_c223 bl_223 br_223 wl_30 vdd gnd cell_6t
Xbit_r31_c223 bl_223 br_223 wl_31 vdd gnd cell_6t
Xbit_r32_c223 bl_223 br_223 wl_32 vdd gnd cell_6t
Xbit_r33_c223 bl_223 br_223 wl_33 vdd gnd cell_6t
Xbit_r34_c223 bl_223 br_223 wl_34 vdd gnd cell_6t
Xbit_r35_c223 bl_223 br_223 wl_35 vdd gnd cell_6t
Xbit_r36_c223 bl_223 br_223 wl_36 vdd gnd cell_6t
Xbit_r37_c223 bl_223 br_223 wl_37 vdd gnd cell_6t
Xbit_r38_c223 bl_223 br_223 wl_38 vdd gnd cell_6t
Xbit_r39_c223 bl_223 br_223 wl_39 vdd gnd cell_6t
Xbit_r40_c223 bl_223 br_223 wl_40 vdd gnd cell_6t
Xbit_r41_c223 bl_223 br_223 wl_41 vdd gnd cell_6t
Xbit_r42_c223 bl_223 br_223 wl_42 vdd gnd cell_6t
Xbit_r43_c223 bl_223 br_223 wl_43 vdd gnd cell_6t
Xbit_r44_c223 bl_223 br_223 wl_44 vdd gnd cell_6t
Xbit_r45_c223 bl_223 br_223 wl_45 vdd gnd cell_6t
Xbit_r46_c223 bl_223 br_223 wl_46 vdd gnd cell_6t
Xbit_r47_c223 bl_223 br_223 wl_47 vdd gnd cell_6t
Xbit_r48_c223 bl_223 br_223 wl_48 vdd gnd cell_6t
Xbit_r49_c223 bl_223 br_223 wl_49 vdd gnd cell_6t
Xbit_r50_c223 bl_223 br_223 wl_50 vdd gnd cell_6t
Xbit_r51_c223 bl_223 br_223 wl_51 vdd gnd cell_6t
Xbit_r52_c223 bl_223 br_223 wl_52 vdd gnd cell_6t
Xbit_r53_c223 bl_223 br_223 wl_53 vdd gnd cell_6t
Xbit_r54_c223 bl_223 br_223 wl_54 vdd gnd cell_6t
Xbit_r55_c223 bl_223 br_223 wl_55 vdd gnd cell_6t
Xbit_r56_c223 bl_223 br_223 wl_56 vdd gnd cell_6t
Xbit_r57_c223 bl_223 br_223 wl_57 vdd gnd cell_6t
Xbit_r58_c223 bl_223 br_223 wl_58 vdd gnd cell_6t
Xbit_r59_c223 bl_223 br_223 wl_59 vdd gnd cell_6t
Xbit_r60_c223 bl_223 br_223 wl_60 vdd gnd cell_6t
Xbit_r61_c223 bl_223 br_223 wl_61 vdd gnd cell_6t
Xbit_r62_c223 bl_223 br_223 wl_62 vdd gnd cell_6t
Xbit_r63_c223 bl_223 br_223 wl_63 vdd gnd cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd cell_6t
Xbit_r1_c224 bl_224 br_224 wl_1 vdd gnd cell_6t
Xbit_r2_c224 bl_224 br_224 wl_2 vdd gnd cell_6t
Xbit_r3_c224 bl_224 br_224 wl_3 vdd gnd cell_6t
Xbit_r4_c224 bl_224 br_224 wl_4 vdd gnd cell_6t
Xbit_r5_c224 bl_224 br_224 wl_5 vdd gnd cell_6t
Xbit_r6_c224 bl_224 br_224 wl_6 vdd gnd cell_6t
Xbit_r7_c224 bl_224 br_224 wl_7 vdd gnd cell_6t
Xbit_r8_c224 bl_224 br_224 wl_8 vdd gnd cell_6t
Xbit_r9_c224 bl_224 br_224 wl_9 vdd gnd cell_6t
Xbit_r10_c224 bl_224 br_224 wl_10 vdd gnd cell_6t
Xbit_r11_c224 bl_224 br_224 wl_11 vdd gnd cell_6t
Xbit_r12_c224 bl_224 br_224 wl_12 vdd gnd cell_6t
Xbit_r13_c224 bl_224 br_224 wl_13 vdd gnd cell_6t
Xbit_r14_c224 bl_224 br_224 wl_14 vdd gnd cell_6t
Xbit_r15_c224 bl_224 br_224 wl_15 vdd gnd cell_6t
Xbit_r16_c224 bl_224 br_224 wl_16 vdd gnd cell_6t
Xbit_r17_c224 bl_224 br_224 wl_17 vdd gnd cell_6t
Xbit_r18_c224 bl_224 br_224 wl_18 vdd gnd cell_6t
Xbit_r19_c224 bl_224 br_224 wl_19 vdd gnd cell_6t
Xbit_r20_c224 bl_224 br_224 wl_20 vdd gnd cell_6t
Xbit_r21_c224 bl_224 br_224 wl_21 vdd gnd cell_6t
Xbit_r22_c224 bl_224 br_224 wl_22 vdd gnd cell_6t
Xbit_r23_c224 bl_224 br_224 wl_23 vdd gnd cell_6t
Xbit_r24_c224 bl_224 br_224 wl_24 vdd gnd cell_6t
Xbit_r25_c224 bl_224 br_224 wl_25 vdd gnd cell_6t
Xbit_r26_c224 bl_224 br_224 wl_26 vdd gnd cell_6t
Xbit_r27_c224 bl_224 br_224 wl_27 vdd gnd cell_6t
Xbit_r28_c224 bl_224 br_224 wl_28 vdd gnd cell_6t
Xbit_r29_c224 bl_224 br_224 wl_29 vdd gnd cell_6t
Xbit_r30_c224 bl_224 br_224 wl_30 vdd gnd cell_6t
Xbit_r31_c224 bl_224 br_224 wl_31 vdd gnd cell_6t
Xbit_r32_c224 bl_224 br_224 wl_32 vdd gnd cell_6t
Xbit_r33_c224 bl_224 br_224 wl_33 vdd gnd cell_6t
Xbit_r34_c224 bl_224 br_224 wl_34 vdd gnd cell_6t
Xbit_r35_c224 bl_224 br_224 wl_35 vdd gnd cell_6t
Xbit_r36_c224 bl_224 br_224 wl_36 vdd gnd cell_6t
Xbit_r37_c224 bl_224 br_224 wl_37 vdd gnd cell_6t
Xbit_r38_c224 bl_224 br_224 wl_38 vdd gnd cell_6t
Xbit_r39_c224 bl_224 br_224 wl_39 vdd gnd cell_6t
Xbit_r40_c224 bl_224 br_224 wl_40 vdd gnd cell_6t
Xbit_r41_c224 bl_224 br_224 wl_41 vdd gnd cell_6t
Xbit_r42_c224 bl_224 br_224 wl_42 vdd gnd cell_6t
Xbit_r43_c224 bl_224 br_224 wl_43 vdd gnd cell_6t
Xbit_r44_c224 bl_224 br_224 wl_44 vdd gnd cell_6t
Xbit_r45_c224 bl_224 br_224 wl_45 vdd gnd cell_6t
Xbit_r46_c224 bl_224 br_224 wl_46 vdd gnd cell_6t
Xbit_r47_c224 bl_224 br_224 wl_47 vdd gnd cell_6t
Xbit_r48_c224 bl_224 br_224 wl_48 vdd gnd cell_6t
Xbit_r49_c224 bl_224 br_224 wl_49 vdd gnd cell_6t
Xbit_r50_c224 bl_224 br_224 wl_50 vdd gnd cell_6t
Xbit_r51_c224 bl_224 br_224 wl_51 vdd gnd cell_6t
Xbit_r52_c224 bl_224 br_224 wl_52 vdd gnd cell_6t
Xbit_r53_c224 bl_224 br_224 wl_53 vdd gnd cell_6t
Xbit_r54_c224 bl_224 br_224 wl_54 vdd gnd cell_6t
Xbit_r55_c224 bl_224 br_224 wl_55 vdd gnd cell_6t
Xbit_r56_c224 bl_224 br_224 wl_56 vdd gnd cell_6t
Xbit_r57_c224 bl_224 br_224 wl_57 vdd gnd cell_6t
Xbit_r58_c224 bl_224 br_224 wl_58 vdd gnd cell_6t
Xbit_r59_c224 bl_224 br_224 wl_59 vdd gnd cell_6t
Xbit_r60_c224 bl_224 br_224 wl_60 vdd gnd cell_6t
Xbit_r61_c224 bl_224 br_224 wl_61 vdd gnd cell_6t
Xbit_r62_c224 bl_224 br_224 wl_62 vdd gnd cell_6t
Xbit_r63_c224 bl_224 br_224 wl_63 vdd gnd cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd cell_6t
Xbit_r1_c225 bl_225 br_225 wl_1 vdd gnd cell_6t
Xbit_r2_c225 bl_225 br_225 wl_2 vdd gnd cell_6t
Xbit_r3_c225 bl_225 br_225 wl_3 vdd gnd cell_6t
Xbit_r4_c225 bl_225 br_225 wl_4 vdd gnd cell_6t
Xbit_r5_c225 bl_225 br_225 wl_5 vdd gnd cell_6t
Xbit_r6_c225 bl_225 br_225 wl_6 vdd gnd cell_6t
Xbit_r7_c225 bl_225 br_225 wl_7 vdd gnd cell_6t
Xbit_r8_c225 bl_225 br_225 wl_8 vdd gnd cell_6t
Xbit_r9_c225 bl_225 br_225 wl_9 vdd gnd cell_6t
Xbit_r10_c225 bl_225 br_225 wl_10 vdd gnd cell_6t
Xbit_r11_c225 bl_225 br_225 wl_11 vdd gnd cell_6t
Xbit_r12_c225 bl_225 br_225 wl_12 vdd gnd cell_6t
Xbit_r13_c225 bl_225 br_225 wl_13 vdd gnd cell_6t
Xbit_r14_c225 bl_225 br_225 wl_14 vdd gnd cell_6t
Xbit_r15_c225 bl_225 br_225 wl_15 vdd gnd cell_6t
Xbit_r16_c225 bl_225 br_225 wl_16 vdd gnd cell_6t
Xbit_r17_c225 bl_225 br_225 wl_17 vdd gnd cell_6t
Xbit_r18_c225 bl_225 br_225 wl_18 vdd gnd cell_6t
Xbit_r19_c225 bl_225 br_225 wl_19 vdd gnd cell_6t
Xbit_r20_c225 bl_225 br_225 wl_20 vdd gnd cell_6t
Xbit_r21_c225 bl_225 br_225 wl_21 vdd gnd cell_6t
Xbit_r22_c225 bl_225 br_225 wl_22 vdd gnd cell_6t
Xbit_r23_c225 bl_225 br_225 wl_23 vdd gnd cell_6t
Xbit_r24_c225 bl_225 br_225 wl_24 vdd gnd cell_6t
Xbit_r25_c225 bl_225 br_225 wl_25 vdd gnd cell_6t
Xbit_r26_c225 bl_225 br_225 wl_26 vdd gnd cell_6t
Xbit_r27_c225 bl_225 br_225 wl_27 vdd gnd cell_6t
Xbit_r28_c225 bl_225 br_225 wl_28 vdd gnd cell_6t
Xbit_r29_c225 bl_225 br_225 wl_29 vdd gnd cell_6t
Xbit_r30_c225 bl_225 br_225 wl_30 vdd gnd cell_6t
Xbit_r31_c225 bl_225 br_225 wl_31 vdd gnd cell_6t
Xbit_r32_c225 bl_225 br_225 wl_32 vdd gnd cell_6t
Xbit_r33_c225 bl_225 br_225 wl_33 vdd gnd cell_6t
Xbit_r34_c225 bl_225 br_225 wl_34 vdd gnd cell_6t
Xbit_r35_c225 bl_225 br_225 wl_35 vdd gnd cell_6t
Xbit_r36_c225 bl_225 br_225 wl_36 vdd gnd cell_6t
Xbit_r37_c225 bl_225 br_225 wl_37 vdd gnd cell_6t
Xbit_r38_c225 bl_225 br_225 wl_38 vdd gnd cell_6t
Xbit_r39_c225 bl_225 br_225 wl_39 vdd gnd cell_6t
Xbit_r40_c225 bl_225 br_225 wl_40 vdd gnd cell_6t
Xbit_r41_c225 bl_225 br_225 wl_41 vdd gnd cell_6t
Xbit_r42_c225 bl_225 br_225 wl_42 vdd gnd cell_6t
Xbit_r43_c225 bl_225 br_225 wl_43 vdd gnd cell_6t
Xbit_r44_c225 bl_225 br_225 wl_44 vdd gnd cell_6t
Xbit_r45_c225 bl_225 br_225 wl_45 vdd gnd cell_6t
Xbit_r46_c225 bl_225 br_225 wl_46 vdd gnd cell_6t
Xbit_r47_c225 bl_225 br_225 wl_47 vdd gnd cell_6t
Xbit_r48_c225 bl_225 br_225 wl_48 vdd gnd cell_6t
Xbit_r49_c225 bl_225 br_225 wl_49 vdd gnd cell_6t
Xbit_r50_c225 bl_225 br_225 wl_50 vdd gnd cell_6t
Xbit_r51_c225 bl_225 br_225 wl_51 vdd gnd cell_6t
Xbit_r52_c225 bl_225 br_225 wl_52 vdd gnd cell_6t
Xbit_r53_c225 bl_225 br_225 wl_53 vdd gnd cell_6t
Xbit_r54_c225 bl_225 br_225 wl_54 vdd gnd cell_6t
Xbit_r55_c225 bl_225 br_225 wl_55 vdd gnd cell_6t
Xbit_r56_c225 bl_225 br_225 wl_56 vdd gnd cell_6t
Xbit_r57_c225 bl_225 br_225 wl_57 vdd gnd cell_6t
Xbit_r58_c225 bl_225 br_225 wl_58 vdd gnd cell_6t
Xbit_r59_c225 bl_225 br_225 wl_59 vdd gnd cell_6t
Xbit_r60_c225 bl_225 br_225 wl_60 vdd gnd cell_6t
Xbit_r61_c225 bl_225 br_225 wl_61 vdd gnd cell_6t
Xbit_r62_c225 bl_225 br_225 wl_62 vdd gnd cell_6t
Xbit_r63_c225 bl_225 br_225 wl_63 vdd gnd cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd cell_6t
Xbit_r1_c226 bl_226 br_226 wl_1 vdd gnd cell_6t
Xbit_r2_c226 bl_226 br_226 wl_2 vdd gnd cell_6t
Xbit_r3_c226 bl_226 br_226 wl_3 vdd gnd cell_6t
Xbit_r4_c226 bl_226 br_226 wl_4 vdd gnd cell_6t
Xbit_r5_c226 bl_226 br_226 wl_5 vdd gnd cell_6t
Xbit_r6_c226 bl_226 br_226 wl_6 vdd gnd cell_6t
Xbit_r7_c226 bl_226 br_226 wl_7 vdd gnd cell_6t
Xbit_r8_c226 bl_226 br_226 wl_8 vdd gnd cell_6t
Xbit_r9_c226 bl_226 br_226 wl_9 vdd gnd cell_6t
Xbit_r10_c226 bl_226 br_226 wl_10 vdd gnd cell_6t
Xbit_r11_c226 bl_226 br_226 wl_11 vdd gnd cell_6t
Xbit_r12_c226 bl_226 br_226 wl_12 vdd gnd cell_6t
Xbit_r13_c226 bl_226 br_226 wl_13 vdd gnd cell_6t
Xbit_r14_c226 bl_226 br_226 wl_14 vdd gnd cell_6t
Xbit_r15_c226 bl_226 br_226 wl_15 vdd gnd cell_6t
Xbit_r16_c226 bl_226 br_226 wl_16 vdd gnd cell_6t
Xbit_r17_c226 bl_226 br_226 wl_17 vdd gnd cell_6t
Xbit_r18_c226 bl_226 br_226 wl_18 vdd gnd cell_6t
Xbit_r19_c226 bl_226 br_226 wl_19 vdd gnd cell_6t
Xbit_r20_c226 bl_226 br_226 wl_20 vdd gnd cell_6t
Xbit_r21_c226 bl_226 br_226 wl_21 vdd gnd cell_6t
Xbit_r22_c226 bl_226 br_226 wl_22 vdd gnd cell_6t
Xbit_r23_c226 bl_226 br_226 wl_23 vdd gnd cell_6t
Xbit_r24_c226 bl_226 br_226 wl_24 vdd gnd cell_6t
Xbit_r25_c226 bl_226 br_226 wl_25 vdd gnd cell_6t
Xbit_r26_c226 bl_226 br_226 wl_26 vdd gnd cell_6t
Xbit_r27_c226 bl_226 br_226 wl_27 vdd gnd cell_6t
Xbit_r28_c226 bl_226 br_226 wl_28 vdd gnd cell_6t
Xbit_r29_c226 bl_226 br_226 wl_29 vdd gnd cell_6t
Xbit_r30_c226 bl_226 br_226 wl_30 vdd gnd cell_6t
Xbit_r31_c226 bl_226 br_226 wl_31 vdd gnd cell_6t
Xbit_r32_c226 bl_226 br_226 wl_32 vdd gnd cell_6t
Xbit_r33_c226 bl_226 br_226 wl_33 vdd gnd cell_6t
Xbit_r34_c226 bl_226 br_226 wl_34 vdd gnd cell_6t
Xbit_r35_c226 bl_226 br_226 wl_35 vdd gnd cell_6t
Xbit_r36_c226 bl_226 br_226 wl_36 vdd gnd cell_6t
Xbit_r37_c226 bl_226 br_226 wl_37 vdd gnd cell_6t
Xbit_r38_c226 bl_226 br_226 wl_38 vdd gnd cell_6t
Xbit_r39_c226 bl_226 br_226 wl_39 vdd gnd cell_6t
Xbit_r40_c226 bl_226 br_226 wl_40 vdd gnd cell_6t
Xbit_r41_c226 bl_226 br_226 wl_41 vdd gnd cell_6t
Xbit_r42_c226 bl_226 br_226 wl_42 vdd gnd cell_6t
Xbit_r43_c226 bl_226 br_226 wl_43 vdd gnd cell_6t
Xbit_r44_c226 bl_226 br_226 wl_44 vdd gnd cell_6t
Xbit_r45_c226 bl_226 br_226 wl_45 vdd gnd cell_6t
Xbit_r46_c226 bl_226 br_226 wl_46 vdd gnd cell_6t
Xbit_r47_c226 bl_226 br_226 wl_47 vdd gnd cell_6t
Xbit_r48_c226 bl_226 br_226 wl_48 vdd gnd cell_6t
Xbit_r49_c226 bl_226 br_226 wl_49 vdd gnd cell_6t
Xbit_r50_c226 bl_226 br_226 wl_50 vdd gnd cell_6t
Xbit_r51_c226 bl_226 br_226 wl_51 vdd gnd cell_6t
Xbit_r52_c226 bl_226 br_226 wl_52 vdd gnd cell_6t
Xbit_r53_c226 bl_226 br_226 wl_53 vdd gnd cell_6t
Xbit_r54_c226 bl_226 br_226 wl_54 vdd gnd cell_6t
Xbit_r55_c226 bl_226 br_226 wl_55 vdd gnd cell_6t
Xbit_r56_c226 bl_226 br_226 wl_56 vdd gnd cell_6t
Xbit_r57_c226 bl_226 br_226 wl_57 vdd gnd cell_6t
Xbit_r58_c226 bl_226 br_226 wl_58 vdd gnd cell_6t
Xbit_r59_c226 bl_226 br_226 wl_59 vdd gnd cell_6t
Xbit_r60_c226 bl_226 br_226 wl_60 vdd gnd cell_6t
Xbit_r61_c226 bl_226 br_226 wl_61 vdd gnd cell_6t
Xbit_r62_c226 bl_226 br_226 wl_62 vdd gnd cell_6t
Xbit_r63_c226 bl_226 br_226 wl_63 vdd gnd cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd cell_6t
Xbit_r1_c227 bl_227 br_227 wl_1 vdd gnd cell_6t
Xbit_r2_c227 bl_227 br_227 wl_2 vdd gnd cell_6t
Xbit_r3_c227 bl_227 br_227 wl_3 vdd gnd cell_6t
Xbit_r4_c227 bl_227 br_227 wl_4 vdd gnd cell_6t
Xbit_r5_c227 bl_227 br_227 wl_5 vdd gnd cell_6t
Xbit_r6_c227 bl_227 br_227 wl_6 vdd gnd cell_6t
Xbit_r7_c227 bl_227 br_227 wl_7 vdd gnd cell_6t
Xbit_r8_c227 bl_227 br_227 wl_8 vdd gnd cell_6t
Xbit_r9_c227 bl_227 br_227 wl_9 vdd gnd cell_6t
Xbit_r10_c227 bl_227 br_227 wl_10 vdd gnd cell_6t
Xbit_r11_c227 bl_227 br_227 wl_11 vdd gnd cell_6t
Xbit_r12_c227 bl_227 br_227 wl_12 vdd gnd cell_6t
Xbit_r13_c227 bl_227 br_227 wl_13 vdd gnd cell_6t
Xbit_r14_c227 bl_227 br_227 wl_14 vdd gnd cell_6t
Xbit_r15_c227 bl_227 br_227 wl_15 vdd gnd cell_6t
Xbit_r16_c227 bl_227 br_227 wl_16 vdd gnd cell_6t
Xbit_r17_c227 bl_227 br_227 wl_17 vdd gnd cell_6t
Xbit_r18_c227 bl_227 br_227 wl_18 vdd gnd cell_6t
Xbit_r19_c227 bl_227 br_227 wl_19 vdd gnd cell_6t
Xbit_r20_c227 bl_227 br_227 wl_20 vdd gnd cell_6t
Xbit_r21_c227 bl_227 br_227 wl_21 vdd gnd cell_6t
Xbit_r22_c227 bl_227 br_227 wl_22 vdd gnd cell_6t
Xbit_r23_c227 bl_227 br_227 wl_23 vdd gnd cell_6t
Xbit_r24_c227 bl_227 br_227 wl_24 vdd gnd cell_6t
Xbit_r25_c227 bl_227 br_227 wl_25 vdd gnd cell_6t
Xbit_r26_c227 bl_227 br_227 wl_26 vdd gnd cell_6t
Xbit_r27_c227 bl_227 br_227 wl_27 vdd gnd cell_6t
Xbit_r28_c227 bl_227 br_227 wl_28 vdd gnd cell_6t
Xbit_r29_c227 bl_227 br_227 wl_29 vdd gnd cell_6t
Xbit_r30_c227 bl_227 br_227 wl_30 vdd gnd cell_6t
Xbit_r31_c227 bl_227 br_227 wl_31 vdd gnd cell_6t
Xbit_r32_c227 bl_227 br_227 wl_32 vdd gnd cell_6t
Xbit_r33_c227 bl_227 br_227 wl_33 vdd gnd cell_6t
Xbit_r34_c227 bl_227 br_227 wl_34 vdd gnd cell_6t
Xbit_r35_c227 bl_227 br_227 wl_35 vdd gnd cell_6t
Xbit_r36_c227 bl_227 br_227 wl_36 vdd gnd cell_6t
Xbit_r37_c227 bl_227 br_227 wl_37 vdd gnd cell_6t
Xbit_r38_c227 bl_227 br_227 wl_38 vdd gnd cell_6t
Xbit_r39_c227 bl_227 br_227 wl_39 vdd gnd cell_6t
Xbit_r40_c227 bl_227 br_227 wl_40 vdd gnd cell_6t
Xbit_r41_c227 bl_227 br_227 wl_41 vdd gnd cell_6t
Xbit_r42_c227 bl_227 br_227 wl_42 vdd gnd cell_6t
Xbit_r43_c227 bl_227 br_227 wl_43 vdd gnd cell_6t
Xbit_r44_c227 bl_227 br_227 wl_44 vdd gnd cell_6t
Xbit_r45_c227 bl_227 br_227 wl_45 vdd gnd cell_6t
Xbit_r46_c227 bl_227 br_227 wl_46 vdd gnd cell_6t
Xbit_r47_c227 bl_227 br_227 wl_47 vdd gnd cell_6t
Xbit_r48_c227 bl_227 br_227 wl_48 vdd gnd cell_6t
Xbit_r49_c227 bl_227 br_227 wl_49 vdd gnd cell_6t
Xbit_r50_c227 bl_227 br_227 wl_50 vdd gnd cell_6t
Xbit_r51_c227 bl_227 br_227 wl_51 vdd gnd cell_6t
Xbit_r52_c227 bl_227 br_227 wl_52 vdd gnd cell_6t
Xbit_r53_c227 bl_227 br_227 wl_53 vdd gnd cell_6t
Xbit_r54_c227 bl_227 br_227 wl_54 vdd gnd cell_6t
Xbit_r55_c227 bl_227 br_227 wl_55 vdd gnd cell_6t
Xbit_r56_c227 bl_227 br_227 wl_56 vdd gnd cell_6t
Xbit_r57_c227 bl_227 br_227 wl_57 vdd gnd cell_6t
Xbit_r58_c227 bl_227 br_227 wl_58 vdd gnd cell_6t
Xbit_r59_c227 bl_227 br_227 wl_59 vdd gnd cell_6t
Xbit_r60_c227 bl_227 br_227 wl_60 vdd gnd cell_6t
Xbit_r61_c227 bl_227 br_227 wl_61 vdd gnd cell_6t
Xbit_r62_c227 bl_227 br_227 wl_62 vdd gnd cell_6t
Xbit_r63_c227 bl_227 br_227 wl_63 vdd gnd cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd cell_6t
Xbit_r1_c228 bl_228 br_228 wl_1 vdd gnd cell_6t
Xbit_r2_c228 bl_228 br_228 wl_2 vdd gnd cell_6t
Xbit_r3_c228 bl_228 br_228 wl_3 vdd gnd cell_6t
Xbit_r4_c228 bl_228 br_228 wl_4 vdd gnd cell_6t
Xbit_r5_c228 bl_228 br_228 wl_5 vdd gnd cell_6t
Xbit_r6_c228 bl_228 br_228 wl_6 vdd gnd cell_6t
Xbit_r7_c228 bl_228 br_228 wl_7 vdd gnd cell_6t
Xbit_r8_c228 bl_228 br_228 wl_8 vdd gnd cell_6t
Xbit_r9_c228 bl_228 br_228 wl_9 vdd gnd cell_6t
Xbit_r10_c228 bl_228 br_228 wl_10 vdd gnd cell_6t
Xbit_r11_c228 bl_228 br_228 wl_11 vdd gnd cell_6t
Xbit_r12_c228 bl_228 br_228 wl_12 vdd gnd cell_6t
Xbit_r13_c228 bl_228 br_228 wl_13 vdd gnd cell_6t
Xbit_r14_c228 bl_228 br_228 wl_14 vdd gnd cell_6t
Xbit_r15_c228 bl_228 br_228 wl_15 vdd gnd cell_6t
Xbit_r16_c228 bl_228 br_228 wl_16 vdd gnd cell_6t
Xbit_r17_c228 bl_228 br_228 wl_17 vdd gnd cell_6t
Xbit_r18_c228 bl_228 br_228 wl_18 vdd gnd cell_6t
Xbit_r19_c228 bl_228 br_228 wl_19 vdd gnd cell_6t
Xbit_r20_c228 bl_228 br_228 wl_20 vdd gnd cell_6t
Xbit_r21_c228 bl_228 br_228 wl_21 vdd gnd cell_6t
Xbit_r22_c228 bl_228 br_228 wl_22 vdd gnd cell_6t
Xbit_r23_c228 bl_228 br_228 wl_23 vdd gnd cell_6t
Xbit_r24_c228 bl_228 br_228 wl_24 vdd gnd cell_6t
Xbit_r25_c228 bl_228 br_228 wl_25 vdd gnd cell_6t
Xbit_r26_c228 bl_228 br_228 wl_26 vdd gnd cell_6t
Xbit_r27_c228 bl_228 br_228 wl_27 vdd gnd cell_6t
Xbit_r28_c228 bl_228 br_228 wl_28 vdd gnd cell_6t
Xbit_r29_c228 bl_228 br_228 wl_29 vdd gnd cell_6t
Xbit_r30_c228 bl_228 br_228 wl_30 vdd gnd cell_6t
Xbit_r31_c228 bl_228 br_228 wl_31 vdd gnd cell_6t
Xbit_r32_c228 bl_228 br_228 wl_32 vdd gnd cell_6t
Xbit_r33_c228 bl_228 br_228 wl_33 vdd gnd cell_6t
Xbit_r34_c228 bl_228 br_228 wl_34 vdd gnd cell_6t
Xbit_r35_c228 bl_228 br_228 wl_35 vdd gnd cell_6t
Xbit_r36_c228 bl_228 br_228 wl_36 vdd gnd cell_6t
Xbit_r37_c228 bl_228 br_228 wl_37 vdd gnd cell_6t
Xbit_r38_c228 bl_228 br_228 wl_38 vdd gnd cell_6t
Xbit_r39_c228 bl_228 br_228 wl_39 vdd gnd cell_6t
Xbit_r40_c228 bl_228 br_228 wl_40 vdd gnd cell_6t
Xbit_r41_c228 bl_228 br_228 wl_41 vdd gnd cell_6t
Xbit_r42_c228 bl_228 br_228 wl_42 vdd gnd cell_6t
Xbit_r43_c228 bl_228 br_228 wl_43 vdd gnd cell_6t
Xbit_r44_c228 bl_228 br_228 wl_44 vdd gnd cell_6t
Xbit_r45_c228 bl_228 br_228 wl_45 vdd gnd cell_6t
Xbit_r46_c228 bl_228 br_228 wl_46 vdd gnd cell_6t
Xbit_r47_c228 bl_228 br_228 wl_47 vdd gnd cell_6t
Xbit_r48_c228 bl_228 br_228 wl_48 vdd gnd cell_6t
Xbit_r49_c228 bl_228 br_228 wl_49 vdd gnd cell_6t
Xbit_r50_c228 bl_228 br_228 wl_50 vdd gnd cell_6t
Xbit_r51_c228 bl_228 br_228 wl_51 vdd gnd cell_6t
Xbit_r52_c228 bl_228 br_228 wl_52 vdd gnd cell_6t
Xbit_r53_c228 bl_228 br_228 wl_53 vdd gnd cell_6t
Xbit_r54_c228 bl_228 br_228 wl_54 vdd gnd cell_6t
Xbit_r55_c228 bl_228 br_228 wl_55 vdd gnd cell_6t
Xbit_r56_c228 bl_228 br_228 wl_56 vdd gnd cell_6t
Xbit_r57_c228 bl_228 br_228 wl_57 vdd gnd cell_6t
Xbit_r58_c228 bl_228 br_228 wl_58 vdd gnd cell_6t
Xbit_r59_c228 bl_228 br_228 wl_59 vdd gnd cell_6t
Xbit_r60_c228 bl_228 br_228 wl_60 vdd gnd cell_6t
Xbit_r61_c228 bl_228 br_228 wl_61 vdd gnd cell_6t
Xbit_r62_c228 bl_228 br_228 wl_62 vdd gnd cell_6t
Xbit_r63_c228 bl_228 br_228 wl_63 vdd gnd cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd cell_6t
Xbit_r1_c229 bl_229 br_229 wl_1 vdd gnd cell_6t
Xbit_r2_c229 bl_229 br_229 wl_2 vdd gnd cell_6t
Xbit_r3_c229 bl_229 br_229 wl_3 vdd gnd cell_6t
Xbit_r4_c229 bl_229 br_229 wl_4 vdd gnd cell_6t
Xbit_r5_c229 bl_229 br_229 wl_5 vdd gnd cell_6t
Xbit_r6_c229 bl_229 br_229 wl_6 vdd gnd cell_6t
Xbit_r7_c229 bl_229 br_229 wl_7 vdd gnd cell_6t
Xbit_r8_c229 bl_229 br_229 wl_8 vdd gnd cell_6t
Xbit_r9_c229 bl_229 br_229 wl_9 vdd gnd cell_6t
Xbit_r10_c229 bl_229 br_229 wl_10 vdd gnd cell_6t
Xbit_r11_c229 bl_229 br_229 wl_11 vdd gnd cell_6t
Xbit_r12_c229 bl_229 br_229 wl_12 vdd gnd cell_6t
Xbit_r13_c229 bl_229 br_229 wl_13 vdd gnd cell_6t
Xbit_r14_c229 bl_229 br_229 wl_14 vdd gnd cell_6t
Xbit_r15_c229 bl_229 br_229 wl_15 vdd gnd cell_6t
Xbit_r16_c229 bl_229 br_229 wl_16 vdd gnd cell_6t
Xbit_r17_c229 bl_229 br_229 wl_17 vdd gnd cell_6t
Xbit_r18_c229 bl_229 br_229 wl_18 vdd gnd cell_6t
Xbit_r19_c229 bl_229 br_229 wl_19 vdd gnd cell_6t
Xbit_r20_c229 bl_229 br_229 wl_20 vdd gnd cell_6t
Xbit_r21_c229 bl_229 br_229 wl_21 vdd gnd cell_6t
Xbit_r22_c229 bl_229 br_229 wl_22 vdd gnd cell_6t
Xbit_r23_c229 bl_229 br_229 wl_23 vdd gnd cell_6t
Xbit_r24_c229 bl_229 br_229 wl_24 vdd gnd cell_6t
Xbit_r25_c229 bl_229 br_229 wl_25 vdd gnd cell_6t
Xbit_r26_c229 bl_229 br_229 wl_26 vdd gnd cell_6t
Xbit_r27_c229 bl_229 br_229 wl_27 vdd gnd cell_6t
Xbit_r28_c229 bl_229 br_229 wl_28 vdd gnd cell_6t
Xbit_r29_c229 bl_229 br_229 wl_29 vdd gnd cell_6t
Xbit_r30_c229 bl_229 br_229 wl_30 vdd gnd cell_6t
Xbit_r31_c229 bl_229 br_229 wl_31 vdd gnd cell_6t
Xbit_r32_c229 bl_229 br_229 wl_32 vdd gnd cell_6t
Xbit_r33_c229 bl_229 br_229 wl_33 vdd gnd cell_6t
Xbit_r34_c229 bl_229 br_229 wl_34 vdd gnd cell_6t
Xbit_r35_c229 bl_229 br_229 wl_35 vdd gnd cell_6t
Xbit_r36_c229 bl_229 br_229 wl_36 vdd gnd cell_6t
Xbit_r37_c229 bl_229 br_229 wl_37 vdd gnd cell_6t
Xbit_r38_c229 bl_229 br_229 wl_38 vdd gnd cell_6t
Xbit_r39_c229 bl_229 br_229 wl_39 vdd gnd cell_6t
Xbit_r40_c229 bl_229 br_229 wl_40 vdd gnd cell_6t
Xbit_r41_c229 bl_229 br_229 wl_41 vdd gnd cell_6t
Xbit_r42_c229 bl_229 br_229 wl_42 vdd gnd cell_6t
Xbit_r43_c229 bl_229 br_229 wl_43 vdd gnd cell_6t
Xbit_r44_c229 bl_229 br_229 wl_44 vdd gnd cell_6t
Xbit_r45_c229 bl_229 br_229 wl_45 vdd gnd cell_6t
Xbit_r46_c229 bl_229 br_229 wl_46 vdd gnd cell_6t
Xbit_r47_c229 bl_229 br_229 wl_47 vdd gnd cell_6t
Xbit_r48_c229 bl_229 br_229 wl_48 vdd gnd cell_6t
Xbit_r49_c229 bl_229 br_229 wl_49 vdd gnd cell_6t
Xbit_r50_c229 bl_229 br_229 wl_50 vdd gnd cell_6t
Xbit_r51_c229 bl_229 br_229 wl_51 vdd gnd cell_6t
Xbit_r52_c229 bl_229 br_229 wl_52 vdd gnd cell_6t
Xbit_r53_c229 bl_229 br_229 wl_53 vdd gnd cell_6t
Xbit_r54_c229 bl_229 br_229 wl_54 vdd gnd cell_6t
Xbit_r55_c229 bl_229 br_229 wl_55 vdd gnd cell_6t
Xbit_r56_c229 bl_229 br_229 wl_56 vdd gnd cell_6t
Xbit_r57_c229 bl_229 br_229 wl_57 vdd gnd cell_6t
Xbit_r58_c229 bl_229 br_229 wl_58 vdd gnd cell_6t
Xbit_r59_c229 bl_229 br_229 wl_59 vdd gnd cell_6t
Xbit_r60_c229 bl_229 br_229 wl_60 vdd gnd cell_6t
Xbit_r61_c229 bl_229 br_229 wl_61 vdd gnd cell_6t
Xbit_r62_c229 bl_229 br_229 wl_62 vdd gnd cell_6t
Xbit_r63_c229 bl_229 br_229 wl_63 vdd gnd cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd cell_6t
Xbit_r1_c230 bl_230 br_230 wl_1 vdd gnd cell_6t
Xbit_r2_c230 bl_230 br_230 wl_2 vdd gnd cell_6t
Xbit_r3_c230 bl_230 br_230 wl_3 vdd gnd cell_6t
Xbit_r4_c230 bl_230 br_230 wl_4 vdd gnd cell_6t
Xbit_r5_c230 bl_230 br_230 wl_5 vdd gnd cell_6t
Xbit_r6_c230 bl_230 br_230 wl_6 vdd gnd cell_6t
Xbit_r7_c230 bl_230 br_230 wl_7 vdd gnd cell_6t
Xbit_r8_c230 bl_230 br_230 wl_8 vdd gnd cell_6t
Xbit_r9_c230 bl_230 br_230 wl_9 vdd gnd cell_6t
Xbit_r10_c230 bl_230 br_230 wl_10 vdd gnd cell_6t
Xbit_r11_c230 bl_230 br_230 wl_11 vdd gnd cell_6t
Xbit_r12_c230 bl_230 br_230 wl_12 vdd gnd cell_6t
Xbit_r13_c230 bl_230 br_230 wl_13 vdd gnd cell_6t
Xbit_r14_c230 bl_230 br_230 wl_14 vdd gnd cell_6t
Xbit_r15_c230 bl_230 br_230 wl_15 vdd gnd cell_6t
Xbit_r16_c230 bl_230 br_230 wl_16 vdd gnd cell_6t
Xbit_r17_c230 bl_230 br_230 wl_17 vdd gnd cell_6t
Xbit_r18_c230 bl_230 br_230 wl_18 vdd gnd cell_6t
Xbit_r19_c230 bl_230 br_230 wl_19 vdd gnd cell_6t
Xbit_r20_c230 bl_230 br_230 wl_20 vdd gnd cell_6t
Xbit_r21_c230 bl_230 br_230 wl_21 vdd gnd cell_6t
Xbit_r22_c230 bl_230 br_230 wl_22 vdd gnd cell_6t
Xbit_r23_c230 bl_230 br_230 wl_23 vdd gnd cell_6t
Xbit_r24_c230 bl_230 br_230 wl_24 vdd gnd cell_6t
Xbit_r25_c230 bl_230 br_230 wl_25 vdd gnd cell_6t
Xbit_r26_c230 bl_230 br_230 wl_26 vdd gnd cell_6t
Xbit_r27_c230 bl_230 br_230 wl_27 vdd gnd cell_6t
Xbit_r28_c230 bl_230 br_230 wl_28 vdd gnd cell_6t
Xbit_r29_c230 bl_230 br_230 wl_29 vdd gnd cell_6t
Xbit_r30_c230 bl_230 br_230 wl_30 vdd gnd cell_6t
Xbit_r31_c230 bl_230 br_230 wl_31 vdd gnd cell_6t
Xbit_r32_c230 bl_230 br_230 wl_32 vdd gnd cell_6t
Xbit_r33_c230 bl_230 br_230 wl_33 vdd gnd cell_6t
Xbit_r34_c230 bl_230 br_230 wl_34 vdd gnd cell_6t
Xbit_r35_c230 bl_230 br_230 wl_35 vdd gnd cell_6t
Xbit_r36_c230 bl_230 br_230 wl_36 vdd gnd cell_6t
Xbit_r37_c230 bl_230 br_230 wl_37 vdd gnd cell_6t
Xbit_r38_c230 bl_230 br_230 wl_38 vdd gnd cell_6t
Xbit_r39_c230 bl_230 br_230 wl_39 vdd gnd cell_6t
Xbit_r40_c230 bl_230 br_230 wl_40 vdd gnd cell_6t
Xbit_r41_c230 bl_230 br_230 wl_41 vdd gnd cell_6t
Xbit_r42_c230 bl_230 br_230 wl_42 vdd gnd cell_6t
Xbit_r43_c230 bl_230 br_230 wl_43 vdd gnd cell_6t
Xbit_r44_c230 bl_230 br_230 wl_44 vdd gnd cell_6t
Xbit_r45_c230 bl_230 br_230 wl_45 vdd gnd cell_6t
Xbit_r46_c230 bl_230 br_230 wl_46 vdd gnd cell_6t
Xbit_r47_c230 bl_230 br_230 wl_47 vdd gnd cell_6t
Xbit_r48_c230 bl_230 br_230 wl_48 vdd gnd cell_6t
Xbit_r49_c230 bl_230 br_230 wl_49 vdd gnd cell_6t
Xbit_r50_c230 bl_230 br_230 wl_50 vdd gnd cell_6t
Xbit_r51_c230 bl_230 br_230 wl_51 vdd gnd cell_6t
Xbit_r52_c230 bl_230 br_230 wl_52 vdd gnd cell_6t
Xbit_r53_c230 bl_230 br_230 wl_53 vdd gnd cell_6t
Xbit_r54_c230 bl_230 br_230 wl_54 vdd gnd cell_6t
Xbit_r55_c230 bl_230 br_230 wl_55 vdd gnd cell_6t
Xbit_r56_c230 bl_230 br_230 wl_56 vdd gnd cell_6t
Xbit_r57_c230 bl_230 br_230 wl_57 vdd gnd cell_6t
Xbit_r58_c230 bl_230 br_230 wl_58 vdd gnd cell_6t
Xbit_r59_c230 bl_230 br_230 wl_59 vdd gnd cell_6t
Xbit_r60_c230 bl_230 br_230 wl_60 vdd gnd cell_6t
Xbit_r61_c230 bl_230 br_230 wl_61 vdd gnd cell_6t
Xbit_r62_c230 bl_230 br_230 wl_62 vdd gnd cell_6t
Xbit_r63_c230 bl_230 br_230 wl_63 vdd gnd cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd cell_6t
Xbit_r1_c231 bl_231 br_231 wl_1 vdd gnd cell_6t
Xbit_r2_c231 bl_231 br_231 wl_2 vdd gnd cell_6t
Xbit_r3_c231 bl_231 br_231 wl_3 vdd gnd cell_6t
Xbit_r4_c231 bl_231 br_231 wl_4 vdd gnd cell_6t
Xbit_r5_c231 bl_231 br_231 wl_5 vdd gnd cell_6t
Xbit_r6_c231 bl_231 br_231 wl_6 vdd gnd cell_6t
Xbit_r7_c231 bl_231 br_231 wl_7 vdd gnd cell_6t
Xbit_r8_c231 bl_231 br_231 wl_8 vdd gnd cell_6t
Xbit_r9_c231 bl_231 br_231 wl_9 vdd gnd cell_6t
Xbit_r10_c231 bl_231 br_231 wl_10 vdd gnd cell_6t
Xbit_r11_c231 bl_231 br_231 wl_11 vdd gnd cell_6t
Xbit_r12_c231 bl_231 br_231 wl_12 vdd gnd cell_6t
Xbit_r13_c231 bl_231 br_231 wl_13 vdd gnd cell_6t
Xbit_r14_c231 bl_231 br_231 wl_14 vdd gnd cell_6t
Xbit_r15_c231 bl_231 br_231 wl_15 vdd gnd cell_6t
Xbit_r16_c231 bl_231 br_231 wl_16 vdd gnd cell_6t
Xbit_r17_c231 bl_231 br_231 wl_17 vdd gnd cell_6t
Xbit_r18_c231 bl_231 br_231 wl_18 vdd gnd cell_6t
Xbit_r19_c231 bl_231 br_231 wl_19 vdd gnd cell_6t
Xbit_r20_c231 bl_231 br_231 wl_20 vdd gnd cell_6t
Xbit_r21_c231 bl_231 br_231 wl_21 vdd gnd cell_6t
Xbit_r22_c231 bl_231 br_231 wl_22 vdd gnd cell_6t
Xbit_r23_c231 bl_231 br_231 wl_23 vdd gnd cell_6t
Xbit_r24_c231 bl_231 br_231 wl_24 vdd gnd cell_6t
Xbit_r25_c231 bl_231 br_231 wl_25 vdd gnd cell_6t
Xbit_r26_c231 bl_231 br_231 wl_26 vdd gnd cell_6t
Xbit_r27_c231 bl_231 br_231 wl_27 vdd gnd cell_6t
Xbit_r28_c231 bl_231 br_231 wl_28 vdd gnd cell_6t
Xbit_r29_c231 bl_231 br_231 wl_29 vdd gnd cell_6t
Xbit_r30_c231 bl_231 br_231 wl_30 vdd gnd cell_6t
Xbit_r31_c231 bl_231 br_231 wl_31 vdd gnd cell_6t
Xbit_r32_c231 bl_231 br_231 wl_32 vdd gnd cell_6t
Xbit_r33_c231 bl_231 br_231 wl_33 vdd gnd cell_6t
Xbit_r34_c231 bl_231 br_231 wl_34 vdd gnd cell_6t
Xbit_r35_c231 bl_231 br_231 wl_35 vdd gnd cell_6t
Xbit_r36_c231 bl_231 br_231 wl_36 vdd gnd cell_6t
Xbit_r37_c231 bl_231 br_231 wl_37 vdd gnd cell_6t
Xbit_r38_c231 bl_231 br_231 wl_38 vdd gnd cell_6t
Xbit_r39_c231 bl_231 br_231 wl_39 vdd gnd cell_6t
Xbit_r40_c231 bl_231 br_231 wl_40 vdd gnd cell_6t
Xbit_r41_c231 bl_231 br_231 wl_41 vdd gnd cell_6t
Xbit_r42_c231 bl_231 br_231 wl_42 vdd gnd cell_6t
Xbit_r43_c231 bl_231 br_231 wl_43 vdd gnd cell_6t
Xbit_r44_c231 bl_231 br_231 wl_44 vdd gnd cell_6t
Xbit_r45_c231 bl_231 br_231 wl_45 vdd gnd cell_6t
Xbit_r46_c231 bl_231 br_231 wl_46 vdd gnd cell_6t
Xbit_r47_c231 bl_231 br_231 wl_47 vdd gnd cell_6t
Xbit_r48_c231 bl_231 br_231 wl_48 vdd gnd cell_6t
Xbit_r49_c231 bl_231 br_231 wl_49 vdd gnd cell_6t
Xbit_r50_c231 bl_231 br_231 wl_50 vdd gnd cell_6t
Xbit_r51_c231 bl_231 br_231 wl_51 vdd gnd cell_6t
Xbit_r52_c231 bl_231 br_231 wl_52 vdd gnd cell_6t
Xbit_r53_c231 bl_231 br_231 wl_53 vdd gnd cell_6t
Xbit_r54_c231 bl_231 br_231 wl_54 vdd gnd cell_6t
Xbit_r55_c231 bl_231 br_231 wl_55 vdd gnd cell_6t
Xbit_r56_c231 bl_231 br_231 wl_56 vdd gnd cell_6t
Xbit_r57_c231 bl_231 br_231 wl_57 vdd gnd cell_6t
Xbit_r58_c231 bl_231 br_231 wl_58 vdd gnd cell_6t
Xbit_r59_c231 bl_231 br_231 wl_59 vdd gnd cell_6t
Xbit_r60_c231 bl_231 br_231 wl_60 vdd gnd cell_6t
Xbit_r61_c231 bl_231 br_231 wl_61 vdd gnd cell_6t
Xbit_r62_c231 bl_231 br_231 wl_62 vdd gnd cell_6t
Xbit_r63_c231 bl_231 br_231 wl_63 vdd gnd cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd cell_6t
Xbit_r1_c232 bl_232 br_232 wl_1 vdd gnd cell_6t
Xbit_r2_c232 bl_232 br_232 wl_2 vdd gnd cell_6t
Xbit_r3_c232 bl_232 br_232 wl_3 vdd gnd cell_6t
Xbit_r4_c232 bl_232 br_232 wl_4 vdd gnd cell_6t
Xbit_r5_c232 bl_232 br_232 wl_5 vdd gnd cell_6t
Xbit_r6_c232 bl_232 br_232 wl_6 vdd gnd cell_6t
Xbit_r7_c232 bl_232 br_232 wl_7 vdd gnd cell_6t
Xbit_r8_c232 bl_232 br_232 wl_8 vdd gnd cell_6t
Xbit_r9_c232 bl_232 br_232 wl_9 vdd gnd cell_6t
Xbit_r10_c232 bl_232 br_232 wl_10 vdd gnd cell_6t
Xbit_r11_c232 bl_232 br_232 wl_11 vdd gnd cell_6t
Xbit_r12_c232 bl_232 br_232 wl_12 vdd gnd cell_6t
Xbit_r13_c232 bl_232 br_232 wl_13 vdd gnd cell_6t
Xbit_r14_c232 bl_232 br_232 wl_14 vdd gnd cell_6t
Xbit_r15_c232 bl_232 br_232 wl_15 vdd gnd cell_6t
Xbit_r16_c232 bl_232 br_232 wl_16 vdd gnd cell_6t
Xbit_r17_c232 bl_232 br_232 wl_17 vdd gnd cell_6t
Xbit_r18_c232 bl_232 br_232 wl_18 vdd gnd cell_6t
Xbit_r19_c232 bl_232 br_232 wl_19 vdd gnd cell_6t
Xbit_r20_c232 bl_232 br_232 wl_20 vdd gnd cell_6t
Xbit_r21_c232 bl_232 br_232 wl_21 vdd gnd cell_6t
Xbit_r22_c232 bl_232 br_232 wl_22 vdd gnd cell_6t
Xbit_r23_c232 bl_232 br_232 wl_23 vdd gnd cell_6t
Xbit_r24_c232 bl_232 br_232 wl_24 vdd gnd cell_6t
Xbit_r25_c232 bl_232 br_232 wl_25 vdd gnd cell_6t
Xbit_r26_c232 bl_232 br_232 wl_26 vdd gnd cell_6t
Xbit_r27_c232 bl_232 br_232 wl_27 vdd gnd cell_6t
Xbit_r28_c232 bl_232 br_232 wl_28 vdd gnd cell_6t
Xbit_r29_c232 bl_232 br_232 wl_29 vdd gnd cell_6t
Xbit_r30_c232 bl_232 br_232 wl_30 vdd gnd cell_6t
Xbit_r31_c232 bl_232 br_232 wl_31 vdd gnd cell_6t
Xbit_r32_c232 bl_232 br_232 wl_32 vdd gnd cell_6t
Xbit_r33_c232 bl_232 br_232 wl_33 vdd gnd cell_6t
Xbit_r34_c232 bl_232 br_232 wl_34 vdd gnd cell_6t
Xbit_r35_c232 bl_232 br_232 wl_35 vdd gnd cell_6t
Xbit_r36_c232 bl_232 br_232 wl_36 vdd gnd cell_6t
Xbit_r37_c232 bl_232 br_232 wl_37 vdd gnd cell_6t
Xbit_r38_c232 bl_232 br_232 wl_38 vdd gnd cell_6t
Xbit_r39_c232 bl_232 br_232 wl_39 vdd gnd cell_6t
Xbit_r40_c232 bl_232 br_232 wl_40 vdd gnd cell_6t
Xbit_r41_c232 bl_232 br_232 wl_41 vdd gnd cell_6t
Xbit_r42_c232 bl_232 br_232 wl_42 vdd gnd cell_6t
Xbit_r43_c232 bl_232 br_232 wl_43 vdd gnd cell_6t
Xbit_r44_c232 bl_232 br_232 wl_44 vdd gnd cell_6t
Xbit_r45_c232 bl_232 br_232 wl_45 vdd gnd cell_6t
Xbit_r46_c232 bl_232 br_232 wl_46 vdd gnd cell_6t
Xbit_r47_c232 bl_232 br_232 wl_47 vdd gnd cell_6t
Xbit_r48_c232 bl_232 br_232 wl_48 vdd gnd cell_6t
Xbit_r49_c232 bl_232 br_232 wl_49 vdd gnd cell_6t
Xbit_r50_c232 bl_232 br_232 wl_50 vdd gnd cell_6t
Xbit_r51_c232 bl_232 br_232 wl_51 vdd gnd cell_6t
Xbit_r52_c232 bl_232 br_232 wl_52 vdd gnd cell_6t
Xbit_r53_c232 bl_232 br_232 wl_53 vdd gnd cell_6t
Xbit_r54_c232 bl_232 br_232 wl_54 vdd gnd cell_6t
Xbit_r55_c232 bl_232 br_232 wl_55 vdd gnd cell_6t
Xbit_r56_c232 bl_232 br_232 wl_56 vdd gnd cell_6t
Xbit_r57_c232 bl_232 br_232 wl_57 vdd gnd cell_6t
Xbit_r58_c232 bl_232 br_232 wl_58 vdd gnd cell_6t
Xbit_r59_c232 bl_232 br_232 wl_59 vdd gnd cell_6t
Xbit_r60_c232 bl_232 br_232 wl_60 vdd gnd cell_6t
Xbit_r61_c232 bl_232 br_232 wl_61 vdd gnd cell_6t
Xbit_r62_c232 bl_232 br_232 wl_62 vdd gnd cell_6t
Xbit_r63_c232 bl_232 br_232 wl_63 vdd gnd cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd cell_6t
Xbit_r1_c233 bl_233 br_233 wl_1 vdd gnd cell_6t
Xbit_r2_c233 bl_233 br_233 wl_2 vdd gnd cell_6t
Xbit_r3_c233 bl_233 br_233 wl_3 vdd gnd cell_6t
Xbit_r4_c233 bl_233 br_233 wl_4 vdd gnd cell_6t
Xbit_r5_c233 bl_233 br_233 wl_5 vdd gnd cell_6t
Xbit_r6_c233 bl_233 br_233 wl_6 vdd gnd cell_6t
Xbit_r7_c233 bl_233 br_233 wl_7 vdd gnd cell_6t
Xbit_r8_c233 bl_233 br_233 wl_8 vdd gnd cell_6t
Xbit_r9_c233 bl_233 br_233 wl_9 vdd gnd cell_6t
Xbit_r10_c233 bl_233 br_233 wl_10 vdd gnd cell_6t
Xbit_r11_c233 bl_233 br_233 wl_11 vdd gnd cell_6t
Xbit_r12_c233 bl_233 br_233 wl_12 vdd gnd cell_6t
Xbit_r13_c233 bl_233 br_233 wl_13 vdd gnd cell_6t
Xbit_r14_c233 bl_233 br_233 wl_14 vdd gnd cell_6t
Xbit_r15_c233 bl_233 br_233 wl_15 vdd gnd cell_6t
Xbit_r16_c233 bl_233 br_233 wl_16 vdd gnd cell_6t
Xbit_r17_c233 bl_233 br_233 wl_17 vdd gnd cell_6t
Xbit_r18_c233 bl_233 br_233 wl_18 vdd gnd cell_6t
Xbit_r19_c233 bl_233 br_233 wl_19 vdd gnd cell_6t
Xbit_r20_c233 bl_233 br_233 wl_20 vdd gnd cell_6t
Xbit_r21_c233 bl_233 br_233 wl_21 vdd gnd cell_6t
Xbit_r22_c233 bl_233 br_233 wl_22 vdd gnd cell_6t
Xbit_r23_c233 bl_233 br_233 wl_23 vdd gnd cell_6t
Xbit_r24_c233 bl_233 br_233 wl_24 vdd gnd cell_6t
Xbit_r25_c233 bl_233 br_233 wl_25 vdd gnd cell_6t
Xbit_r26_c233 bl_233 br_233 wl_26 vdd gnd cell_6t
Xbit_r27_c233 bl_233 br_233 wl_27 vdd gnd cell_6t
Xbit_r28_c233 bl_233 br_233 wl_28 vdd gnd cell_6t
Xbit_r29_c233 bl_233 br_233 wl_29 vdd gnd cell_6t
Xbit_r30_c233 bl_233 br_233 wl_30 vdd gnd cell_6t
Xbit_r31_c233 bl_233 br_233 wl_31 vdd gnd cell_6t
Xbit_r32_c233 bl_233 br_233 wl_32 vdd gnd cell_6t
Xbit_r33_c233 bl_233 br_233 wl_33 vdd gnd cell_6t
Xbit_r34_c233 bl_233 br_233 wl_34 vdd gnd cell_6t
Xbit_r35_c233 bl_233 br_233 wl_35 vdd gnd cell_6t
Xbit_r36_c233 bl_233 br_233 wl_36 vdd gnd cell_6t
Xbit_r37_c233 bl_233 br_233 wl_37 vdd gnd cell_6t
Xbit_r38_c233 bl_233 br_233 wl_38 vdd gnd cell_6t
Xbit_r39_c233 bl_233 br_233 wl_39 vdd gnd cell_6t
Xbit_r40_c233 bl_233 br_233 wl_40 vdd gnd cell_6t
Xbit_r41_c233 bl_233 br_233 wl_41 vdd gnd cell_6t
Xbit_r42_c233 bl_233 br_233 wl_42 vdd gnd cell_6t
Xbit_r43_c233 bl_233 br_233 wl_43 vdd gnd cell_6t
Xbit_r44_c233 bl_233 br_233 wl_44 vdd gnd cell_6t
Xbit_r45_c233 bl_233 br_233 wl_45 vdd gnd cell_6t
Xbit_r46_c233 bl_233 br_233 wl_46 vdd gnd cell_6t
Xbit_r47_c233 bl_233 br_233 wl_47 vdd gnd cell_6t
Xbit_r48_c233 bl_233 br_233 wl_48 vdd gnd cell_6t
Xbit_r49_c233 bl_233 br_233 wl_49 vdd gnd cell_6t
Xbit_r50_c233 bl_233 br_233 wl_50 vdd gnd cell_6t
Xbit_r51_c233 bl_233 br_233 wl_51 vdd gnd cell_6t
Xbit_r52_c233 bl_233 br_233 wl_52 vdd gnd cell_6t
Xbit_r53_c233 bl_233 br_233 wl_53 vdd gnd cell_6t
Xbit_r54_c233 bl_233 br_233 wl_54 vdd gnd cell_6t
Xbit_r55_c233 bl_233 br_233 wl_55 vdd gnd cell_6t
Xbit_r56_c233 bl_233 br_233 wl_56 vdd gnd cell_6t
Xbit_r57_c233 bl_233 br_233 wl_57 vdd gnd cell_6t
Xbit_r58_c233 bl_233 br_233 wl_58 vdd gnd cell_6t
Xbit_r59_c233 bl_233 br_233 wl_59 vdd gnd cell_6t
Xbit_r60_c233 bl_233 br_233 wl_60 vdd gnd cell_6t
Xbit_r61_c233 bl_233 br_233 wl_61 vdd gnd cell_6t
Xbit_r62_c233 bl_233 br_233 wl_62 vdd gnd cell_6t
Xbit_r63_c233 bl_233 br_233 wl_63 vdd gnd cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd cell_6t
Xbit_r1_c234 bl_234 br_234 wl_1 vdd gnd cell_6t
Xbit_r2_c234 bl_234 br_234 wl_2 vdd gnd cell_6t
Xbit_r3_c234 bl_234 br_234 wl_3 vdd gnd cell_6t
Xbit_r4_c234 bl_234 br_234 wl_4 vdd gnd cell_6t
Xbit_r5_c234 bl_234 br_234 wl_5 vdd gnd cell_6t
Xbit_r6_c234 bl_234 br_234 wl_6 vdd gnd cell_6t
Xbit_r7_c234 bl_234 br_234 wl_7 vdd gnd cell_6t
Xbit_r8_c234 bl_234 br_234 wl_8 vdd gnd cell_6t
Xbit_r9_c234 bl_234 br_234 wl_9 vdd gnd cell_6t
Xbit_r10_c234 bl_234 br_234 wl_10 vdd gnd cell_6t
Xbit_r11_c234 bl_234 br_234 wl_11 vdd gnd cell_6t
Xbit_r12_c234 bl_234 br_234 wl_12 vdd gnd cell_6t
Xbit_r13_c234 bl_234 br_234 wl_13 vdd gnd cell_6t
Xbit_r14_c234 bl_234 br_234 wl_14 vdd gnd cell_6t
Xbit_r15_c234 bl_234 br_234 wl_15 vdd gnd cell_6t
Xbit_r16_c234 bl_234 br_234 wl_16 vdd gnd cell_6t
Xbit_r17_c234 bl_234 br_234 wl_17 vdd gnd cell_6t
Xbit_r18_c234 bl_234 br_234 wl_18 vdd gnd cell_6t
Xbit_r19_c234 bl_234 br_234 wl_19 vdd gnd cell_6t
Xbit_r20_c234 bl_234 br_234 wl_20 vdd gnd cell_6t
Xbit_r21_c234 bl_234 br_234 wl_21 vdd gnd cell_6t
Xbit_r22_c234 bl_234 br_234 wl_22 vdd gnd cell_6t
Xbit_r23_c234 bl_234 br_234 wl_23 vdd gnd cell_6t
Xbit_r24_c234 bl_234 br_234 wl_24 vdd gnd cell_6t
Xbit_r25_c234 bl_234 br_234 wl_25 vdd gnd cell_6t
Xbit_r26_c234 bl_234 br_234 wl_26 vdd gnd cell_6t
Xbit_r27_c234 bl_234 br_234 wl_27 vdd gnd cell_6t
Xbit_r28_c234 bl_234 br_234 wl_28 vdd gnd cell_6t
Xbit_r29_c234 bl_234 br_234 wl_29 vdd gnd cell_6t
Xbit_r30_c234 bl_234 br_234 wl_30 vdd gnd cell_6t
Xbit_r31_c234 bl_234 br_234 wl_31 vdd gnd cell_6t
Xbit_r32_c234 bl_234 br_234 wl_32 vdd gnd cell_6t
Xbit_r33_c234 bl_234 br_234 wl_33 vdd gnd cell_6t
Xbit_r34_c234 bl_234 br_234 wl_34 vdd gnd cell_6t
Xbit_r35_c234 bl_234 br_234 wl_35 vdd gnd cell_6t
Xbit_r36_c234 bl_234 br_234 wl_36 vdd gnd cell_6t
Xbit_r37_c234 bl_234 br_234 wl_37 vdd gnd cell_6t
Xbit_r38_c234 bl_234 br_234 wl_38 vdd gnd cell_6t
Xbit_r39_c234 bl_234 br_234 wl_39 vdd gnd cell_6t
Xbit_r40_c234 bl_234 br_234 wl_40 vdd gnd cell_6t
Xbit_r41_c234 bl_234 br_234 wl_41 vdd gnd cell_6t
Xbit_r42_c234 bl_234 br_234 wl_42 vdd gnd cell_6t
Xbit_r43_c234 bl_234 br_234 wl_43 vdd gnd cell_6t
Xbit_r44_c234 bl_234 br_234 wl_44 vdd gnd cell_6t
Xbit_r45_c234 bl_234 br_234 wl_45 vdd gnd cell_6t
Xbit_r46_c234 bl_234 br_234 wl_46 vdd gnd cell_6t
Xbit_r47_c234 bl_234 br_234 wl_47 vdd gnd cell_6t
Xbit_r48_c234 bl_234 br_234 wl_48 vdd gnd cell_6t
Xbit_r49_c234 bl_234 br_234 wl_49 vdd gnd cell_6t
Xbit_r50_c234 bl_234 br_234 wl_50 vdd gnd cell_6t
Xbit_r51_c234 bl_234 br_234 wl_51 vdd gnd cell_6t
Xbit_r52_c234 bl_234 br_234 wl_52 vdd gnd cell_6t
Xbit_r53_c234 bl_234 br_234 wl_53 vdd gnd cell_6t
Xbit_r54_c234 bl_234 br_234 wl_54 vdd gnd cell_6t
Xbit_r55_c234 bl_234 br_234 wl_55 vdd gnd cell_6t
Xbit_r56_c234 bl_234 br_234 wl_56 vdd gnd cell_6t
Xbit_r57_c234 bl_234 br_234 wl_57 vdd gnd cell_6t
Xbit_r58_c234 bl_234 br_234 wl_58 vdd gnd cell_6t
Xbit_r59_c234 bl_234 br_234 wl_59 vdd gnd cell_6t
Xbit_r60_c234 bl_234 br_234 wl_60 vdd gnd cell_6t
Xbit_r61_c234 bl_234 br_234 wl_61 vdd gnd cell_6t
Xbit_r62_c234 bl_234 br_234 wl_62 vdd gnd cell_6t
Xbit_r63_c234 bl_234 br_234 wl_63 vdd gnd cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd cell_6t
Xbit_r1_c235 bl_235 br_235 wl_1 vdd gnd cell_6t
Xbit_r2_c235 bl_235 br_235 wl_2 vdd gnd cell_6t
Xbit_r3_c235 bl_235 br_235 wl_3 vdd gnd cell_6t
Xbit_r4_c235 bl_235 br_235 wl_4 vdd gnd cell_6t
Xbit_r5_c235 bl_235 br_235 wl_5 vdd gnd cell_6t
Xbit_r6_c235 bl_235 br_235 wl_6 vdd gnd cell_6t
Xbit_r7_c235 bl_235 br_235 wl_7 vdd gnd cell_6t
Xbit_r8_c235 bl_235 br_235 wl_8 vdd gnd cell_6t
Xbit_r9_c235 bl_235 br_235 wl_9 vdd gnd cell_6t
Xbit_r10_c235 bl_235 br_235 wl_10 vdd gnd cell_6t
Xbit_r11_c235 bl_235 br_235 wl_11 vdd gnd cell_6t
Xbit_r12_c235 bl_235 br_235 wl_12 vdd gnd cell_6t
Xbit_r13_c235 bl_235 br_235 wl_13 vdd gnd cell_6t
Xbit_r14_c235 bl_235 br_235 wl_14 vdd gnd cell_6t
Xbit_r15_c235 bl_235 br_235 wl_15 vdd gnd cell_6t
Xbit_r16_c235 bl_235 br_235 wl_16 vdd gnd cell_6t
Xbit_r17_c235 bl_235 br_235 wl_17 vdd gnd cell_6t
Xbit_r18_c235 bl_235 br_235 wl_18 vdd gnd cell_6t
Xbit_r19_c235 bl_235 br_235 wl_19 vdd gnd cell_6t
Xbit_r20_c235 bl_235 br_235 wl_20 vdd gnd cell_6t
Xbit_r21_c235 bl_235 br_235 wl_21 vdd gnd cell_6t
Xbit_r22_c235 bl_235 br_235 wl_22 vdd gnd cell_6t
Xbit_r23_c235 bl_235 br_235 wl_23 vdd gnd cell_6t
Xbit_r24_c235 bl_235 br_235 wl_24 vdd gnd cell_6t
Xbit_r25_c235 bl_235 br_235 wl_25 vdd gnd cell_6t
Xbit_r26_c235 bl_235 br_235 wl_26 vdd gnd cell_6t
Xbit_r27_c235 bl_235 br_235 wl_27 vdd gnd cell_6t
Xbit_r28_c235 bl_235 br_235 wl_28 vdd gnd cell_6t
Xbit_r29_c235 bl_235 br_235 wl_29 vdd gnd cell_6t
Xbit_r30_c235 bl_235 br_235 wl_30 vdd gnd cell_6t
Xbit_r31_c235 bl_235 br_235 wl_31 vdd gnd cell_6t
Xbit_r32_c235 bl_235 br_235 wl_32 vdd gnd cell_6t
Xbit_r33_c235 bl_235 br_235 wl_33 vdd gnd cell_6t
Xbit_r34_c235 bl_235 br_235 wl_34 vdd gnd cell_6t
Xbit_r35_c235 bl_235 br_235 wl_35 vdd gnd cell_6t
Xbit_r36_c235 bl_235 br_235 wl_36 vdd gnd cell_6t
Xbit_r37_c235 bl_235 br_235 wl_37 vdd gnd cell_6t
Xbit_r38_c235 bl_235 br_235 wl_38 vdd gnd cell_6t
Xbit_r39_c235 bl_235 br_235 wl_39 vdd gnd cell_6t
Xbit_r40_c235 bl_235 br_235 wl_40 vdd gnd cell_6t
Xbit_r41_c235 bl_235 br_235 wl_41 vdd gnd cell_6t
Xbit_r42_c235 bl_235 br_235 wl_42 vdd gnd cell_6t
Xbit_r43_c235 bl_235 br_235 wl_43 vdd gnd cell_6t
Xbit_r44_c235 bl_235 br_235 wl_44 vdd gnd cell_6t
Xbit_r45_c235 bl_235 br_235 wl_45 vdd gnd cell_6t
Xbit_r46_c235 bl_235 br_235 wl_46 vdd gnd cell_6t
Xbit_r47_c235 bl_235 br_235 wl_47 vdd gnd cell_6t
Xbit_r48_c235 bl_235 br_235 wl_48 vdd gnd cell_6t
Xbit_r49_c235 bl_235 br_235 wl_49 vdd gnd cell_6t
Xbit_r50_c235 bl_235 br_235 wl_50 vdd gnd cell_6t
Xbit_r51_c235 bl_235 br_235 wl_51 vdd gnd cell_6t
Xbit_r52_c235 bl_235 br_235 wl_52 vdd gnd cell_6t
Xbit_r53_c235 bl_235 br_235 wl_53 vdd gnd cell_6t
Xbit_r54_c235 bl_235 br_235 wl_54 vdd gnd cell_6t
Xbit_r55_c235 bl_235 br_235 wl_55 vdd gnd cell_6t
Xbit_r56_c235 bl_235 br_235 wl_56 vdd gnd cell_6t
Xbit_r57_c235 bl_235 br_235 wl_57 vdd gnd cell_6t
Xbit_r58_c235 bl_235 br_235 wl_58 vdd gnd cell_6t
Xbit_r59_c235 bl_235 br_235 wl_59 vdd gnd cell_6t
Xbit_r60_c235 bl_235 br_235 wl_60 vdd gnd cell_6t
Xbit_r61_c235 bl_235 br_235 wl_61 vdd gnd cell_6t
Xbit_r62_c235 bl_235 br_235 wl_62 vdd gnd cell_6t
Xbit_r63_c235 bl_235 br_235 wl_63 vdd gnd cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd cell_6t
Xbit_r1_c236 bl_236 br_236 wl_1 vdd gnd cell_6t
Xbit_r2_c236 bl_236 br_236 wl_2 vdd gnd cell_6t
Xbit_r3_c236 bl_236 br_236 wl_3 vdd gnd cell_6t
Xbit_r4_c236 bl_236 br_236 wl_4 vdd gnd cell_6t
Xbit_r5_c236 bl_236 br_236 wl_5 vdd gnd cell_6t
Xbit_r6_c236 bl_236 br_236 wl_6 vdd gnd cell_6t
Xbit_r7_c236 bl_236 br_236 wl_7 vdd gnd cell_6t
Xbit_r8_c236 bl_236 br_236 wl_8 vdd gnd cell_6t
Xbit_r9_c236 bl_236 br_236 wl_9 vdd gnd cell_6t
Xbit_r10_c236 bl_236 br_236 wl_10 vdd gnd cell_6t
Xbit_r11_c236 bl_236 br_236 wl_11 vdd gnd cell_6t
Xbit_r12_c236 bl_236 br_236 wl_12 vdd gnd cell_6t
Xbit_r13_c236 bl_236 br_236 wl_13 vdd gnd cell_6t
Xbit_r14_c236 bl_236 br_236 wl_14 vdd gnd cell_6t
Xbit_r15_c236 bl_236 br_236 wl_15 vdd gnd cell_6t
Xbit_r16_c236 bl_236 br_236 wl_16 vdd gnd cell_6t
Xbit_r17_c236 bl_236 br_236 wl_17 vdd gnd cell_6t
Xbit_r18_c236 bl_236 br_236 wl_18 vdd gnd cell_6t
Xbit_r19_c236 bl_236 br_236 wl_19 vdd gnd cell_6t
Xbit_r20_c236 bl_236 br_236 wl_20 vdd gnd cell_6t
Xbit_r21_c236 bl_236 br_236 wl_21 vdd gnd cell_6t
Xbit_r22_c236 bl_236 br_236 wl_22 vdd gnd cell_6t
Xbit_r23_c236 bl_236 br_236 wl_23 vdd gnd cell_6t
Xbit_r24_c236 bl_236 br_236 wl_24 vdd gnd cell_6t
Xbit_r25_c236 bl_236 br_236 wl_25 vdd gnd cell_6t
Xbit_r26_c236 bl_236 br_236 wl_26 vdd gnd cell_6t
Xbit_r27_c236 bl_236 br_236 wl_27 vdd gnd cell_6t
Xbit_r28_c236 bl_236 br_236 wl_28 vdd gnd cell_6t
Xbit_r29_c236 bl_236 br_236 wl_29 vdd gnd cell_6t
Xbit_r30_c236 bl_236 br_236 wl_30 vdd gnd cell_6t
Xbit_r31_c236 bl_236 br_236 wl_31 vdd gnd cell_6t
Xbit_r32_c236 bl_236 br_236 wl_32 vdd gnd cell_6t
Xbit_r33_c236 bl_236 br_236 wl_33 vdd gnd cell_6t
Xbit_r34_c236 bl_236 br_236 wl_34 vdd gnd cell_6t
Xbit_r35_c236 bl_236 br_236 wl_35 vdd gnd cell_6t
Xbit_r36_c236 bl_236 br_236 wl_36 vdd gnd cell_6t
Xbit_r37_c236 bl_236 br_236 wl_37 vdd gnd cell_6t
Xbit_r38_c236 bl_236 br_236 wl_38 vdd gnd cell_6t
Xbit_r39_c236 bl_236 br_236 wl_39 vdd gnd cell_6t
Xbit_r40_c236 bl_236 br_236 wl_40 vdd gnd cell_6t
Xbit_r41_c236 bl_236 br_236 wl_41 vdd gnd cell_6t
Xbit_r42_c236 bl_236 br_236 wl_42 vdd gnd cell_6t
Xbit_r43_c236 bl_236 br_236 wl_43 vdd gnd cell_6t
Xbit_r44_c236 bl_236 br_236 wl_44 vdd gnd cell_6t
Xbit_r45_c236 bl_236 br_236 wl_45 vdd gnd cell_6t
Xbit_r46_c236 bl_236 br_236 wl_46 vdd gnd cell_6t
Xbit_r47_c236 bl_236 br_236 wl_47 vdd gnd cell_6t
Xbit_r48_c236 bl_236 br_236 wl_48 vdd gnd cell_6t
Xbit_r49_c236 bl_236 br_236 wl_49 vdd gnd cell_6t
Xbit_r50_c236 bl_236 br_236 wl_50 vdd gnd cell_6t
Xbit_r51_c236 bl_236 br_236 wl_51 vdd gnd cell_6t
Xbit_r52_c236 bl_236 br_236 wl_52 vdd gnd cell_6t
Xbit_r53_c236 bl_236 br_236 wl_53 vdd gnd cell_6t
Xbit_r54_c236 bl_236 br_236 wl_54 vdd gnd cell_6t
Xbit_r55_c236 bl_236 br_236 wl_55 vdd gnd cell_6t
Xbit_r56_c236 bl_236 br_236 wl_56 vdd gnd cell_6t
Xbit_r57_c236 bl_236 br_236 wl_57 vdd gnd cell_6t
Xbit_r58_c236 bl_236 br_236 wl_58 vdd gnd cell_6t
Xbit_r59_c236 bl_236 br_236 wl_59 vdd gnd cell_6t
Xbit_r60_c236 bl_236 br_236 wl_60 vdd gnd cell_6t
Xbit_r61_c236 bl_236 br_236 wl_61 vdd gnd cell_6t
Xbit_r62_c236 bl_236 br_236 wl_62 vdd gnd cell_6t
Xbit_r63_c236 bl_236 br_236 wl_63 vdd gnd cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd cell_6t
Xbit_r1_c237 bl_237 br_237 wl_1 vdd gnd cell_6t
Xbit_r2_c237 bl_237 br_237 wl_2 vdd gnd cell_6t
Xbit_r3_c237 bl_237 br_237 wl_3 vdd gnd cell_6t
Xbit_r4_c237 bl_237 br_237 wl_4 vdd gnd cell_6t
Xbit_r5_c237 bl_237 br_237 wl_5 vdd gnd cell_6t
Xbit_r6_c237 bl_237 br_237 wl_6 vdd gnd cell_6t
Xbit_r7_c237 bl_237 br_237 wl_7 vdd gnd cell_6t
Xbit_r8_c237 bl_237 br_237 wl_8 vdd gnd cell_6t
Xbit_r9_c237 bl_237 br_237 wl_9 vdd gnd cell_6t
Xbit_r10_c237 bl_237 br_237 wl_10 vdd gnd cell_6t
Xbit_r11_c237 bl_237 br_237 wl_11 vdd gnd cell_6t
Xbit_r12_c237 bl_237 br_237 wl_12 vdd gnd cell_6t
Xbit_r13_c237 bl_237 br_237 wl_13 vdd gnd cell_6t
Xbit_r14_c237 bl_237 br_237 wl_14 vdd gnd cell_6t
Xbit_r15_c237 bl_237 br_237 wl_15 vdd gnd cell_6t
Xbit_r16_c237 bl_237 br_237 wl_16 vdd gnd cell_6t
Xbit_r17_c237 bl_237 br_237 wl_17 vdd gnd cell_6t
Xbit_r18_c237 bl_237 br_237 wl_18 vdd gnd cell_6t
Xbit_r19_c237 bl_237 br_237 wl_19 vdd gnd cell_6t
Xbit_r20_c237 bl_237 br_237 wl_20 vdd gnd cell_6t
Xbit_r21_c237 bl_237 br_237 wl_21 vdd gnd cell_6t
Xbit_r22_c237 bl_237 br_237 wl_22 vdd gnd cell_6t
Xbit_r23_c237 bl_237 br_237 wl_23 vdd gnd cell_6t
Xbit_r24_c237 bl_237 br_237 wl_24 vdd gnd cell_6t
Xbit_r25_c237 bl_237 br_237 wl_25 vdd gnd cell_6t
Xbit_r26_c237 bl_237 br_237 wl_26 vdd gnd cell_6t
Xbit_r27_c237 bl_237 br_237 wl_27 vdd gnd cell_6t
Xbit_r28_c237 bl_237 br_237 wl_28 vdd gnd cell_6t
Xbit_r29_c237 bl_237 br_237 wl_29 vdd gnd cell_6t
Xbit_r30_c237 bl_237 br_237 wl_30 vdd gnd cell_6t
Xbit_r31_c237 bl_237 br_237 wl_31 vdd gnd cell_6t
Xbit_r32_c237 bl_237 br_237 wl_32 vdd gnd cell_6t
Xbit_r33_c237 bl_237 br_237 wl_33 vdd gnd cell_6t
Xbit_r34_c237 bl_237 br_237 wl_34 vdd gnd cell_6t
Xbit_r35_c237 bl_237 br_237 wl_35 vdd gnd cell_6t
Xbit_r36_c237 bl_237 br_237 wl_36 vdd gnd cell_6t
Xbit_r37_c237 bl_237 br_237 wl_37 vdd gnd cell_6t
Xbit_r38_c237 bl_237 br_237 wl_38 vdd gnd cell_6t
Xbit_r39_c237 bl_237 br_237 wl_39 vdd gnd cell_6t
Xbit_r40_c237 bl_237 br_237 wl_40 vdd gnd cell_6t
Xbit_r41_c237 bl_237 br_237 wl_41 vdd gnd cell_6t
Xbit_r42_c237 bl_237 br_237 wl_42 vdd gnd cell_6t
Xbit_r43_c237 bl_237 br_237 wl_43 vdd gnd cell_6t
Xbit_r44_c237 bl_237 br_237 wl_44 vdd gnd cell_6t
Xbit_r45_c237 bl_237 br_237 wl_45 vdd gnd cell_6t
Xbit_r46_c237 bl_237 br_237 wl_46 vdd gnd cell_6t
Xbit_r47_c237 bl_237 br_237 wl_47 vdd gnd cell_6t
Xbit_r48_c237 bl_237 br_237 wl_48 vdd gnd cell_6t
Xbit_r49_c237 bl_237 br_237 wl_49 vdd gnd cell_6t
Xbit_r50_c237 bl_237 br_237 wl_50 vdd gnd cell_6t
Xbit_r51_c237 bl_237 br_237 wl_51 vdd gnd cell_6t
Xbit_r52_c237 bl_237 br_237 wl_52 vdd gnd cell_6t
Xbit_r53_c237 bl_237 br_237 wl_53 vdd gnd cell_6t
Xbit_r54_c237 bl_237 br_237 wl_54 vdd gnd cell_6t
Xbit_r55_c237 bl_237 br_237 wl_55 vdd gnd cell_6t
Xbit_r56_c237 bl_237 br_237 wl_56 vdd gnd cell_6t
Xbit_r57_c237 bl_237 br_237 wl_57 vdd gnd cell_6t
Xbit_r58_c237 bl_237 br_237 wl_58 vdd gnd cell_6t
Xbit_r59_c237 bl_237 br_237 wl_59 vdd gnd cell_6t
Xbit_r60_c237 bl_237 br_237 wl_60 vdd gnd cell_6t
Xbit_r61_c237 bl_237 br_237 wl_61 vdd gnd cell_6t
Xbit_r62_c237 bl_237 br_237 wl_62 vdd gnd cell_6t
Xbit_r63_c237 bl_237 br_237 wl_63 vdd gnd cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd cell_6t
Xbit_r1_c238 bl_238 br_238 wl_1 vdd gnd cell_6t
Xbit_r2_c238 bl_238 br_238 wl_2 vdd gnd cell_6t
Xbit_r3_c238 bl_238 br_238 wl_3 vdd gnd cell_6t
Xbit_r4_c238 bl_238 br_238 wl_4 vdd gnd cell_6t
Xbit_r5_c238 bl_238 br_238 wl_5 vdd gnd cell_6t
Xbit_r6_c238 bl_238 br_238 wl_6 vdd gnd cell_6t
Xbit_r7_c238 bl_238 br_238 wl_7 vdd gnd cell_6t
Xbit_r8_c238 bl_238 br_238 wl_8 vdd gnd cell_6t
Xbit_r9_c238 bl_238 br_238 wl_9 vdd gnd cell_6t
Xbit_r10_c238 bl_238 br_238 wl_10 vdd gnd cell_6t
Xbit_r11_c238 bl_238 br_238 wl_11 vdd gnd cell_6t
Xbit_r12_c238 bl_238 br_238 wl_12 vdd gnd cell_6t
Xbit_r13_c238 bl_238 br_238 wl_13 vdd gnd cell_6t
Xbit_r14_c238 bl_238 br_238 wl_14 vdd gnd cell_6t
Xbit_r15_c238 bl_238 br_238 wl_15 vdd gnd cell_6t
Xbit_r16_c238 bl_238 br_238 wl_16 vdd gnd cell_6t
Xbit_r17_c238 bl_238 br_238 wl_17 vdd gnd cell_6t
Xbit_r18_c238 bl_238 br_238 wl_18 vdd gnd cell_6t
Xbit_r19_c238 bl_238 br_238 wl_19 vdd gnd cell_6t
Xbit_r20_c238 bl_238 br_238 wl_20 vdd gnd cell_6t
Xbit_r21_c238 bl_238 br_238 wl_21 vdd gnd cell_6t
Xbit_r22_c238 bl_238 br_238 wl_22 vdd gnd cell_6t
Xbit_r23_c238 bl_238 br_238 wl_23 vdd gnd cell_6t
Xbit_r24_c238 bl_238 br_238 wl_24 vdd gnd cell_6t
Xbit_r25_c238 bl_238 br_238 wl_25 vdd gnd cell_6t
Xbit_r26_c238 bl_238 br_238 wl_26 vdd gnd cell_6t
Xbit_r27_c238 bl_238 br_238 wl_27 vdd gnd cell_6t
Xbit_r28_c238 bl_238 br_238 wl_28 vdd gnd cell_6t
Xbit_r29_c238 bl_238 br_238 wl_29 vdd gnd cell_6t
Xbit_r30_c238 bl_238 br_238 wl_30 vdd gnd cell_6t
Xbit_r31_c238 bl_238 br_238 wl_31 vdd gnd cell_6t
Xbit_r32_c238 bl_238 br_238 wl_32 vdd gnd cell_6t
Xbit_r33_c238 bl_238 br_238 wl_33 vdd gnd cell_6t
Xbit_r34_c238 bl_238 br_238 wl_34 vdd gnd cell_6t
Xbit_r35_c238 bl_238 br_238 wl_35 vdd gnd cell_6t
Xbit_r36_c238 bl_238 br_238 wl_36 vdd gnd cell_6t
Xbit_r37_c238 bl_238 br_238 wl_37 vdd gnd cell_6t
Xbit_r38_c238 bl_238 br_238 wl_38 vdd gnd cell_6t
Xbit_r39_c238 bl_238 br_238 wl_39 vdd gnd cell_6t
Xbit_r40_c238 bl_238 br_238 wl_40 vdd gnd cell_6t
Xbit_r41_c238 bl_238 br_238 wl_41 vdd gnd cell_6t
Xbit_r42_c238 bl_238 br_238 wl_42 vdd gnd cell_6t
Xbit_r43_c238 bl_238 br_238 wl_43 vdd gnd cell_6t
Xbit_r44_c238 bl_238 br_238 wl_44 vdd gnd cell_6t
Xbit_r45_c238 bl_238 br_238 wl_45 vdd gnd cell_6t
Xbit_r46_c238 bl_238 br_238 wl_46 vdd gnd cell_6t
Xbit_r47_c238 bl_238 br_238 wl_47 vdd gnd cell_6t
Xbit_r48_c238 bl_238 br_238 wl_48 vdd gnd cell_6t
Xbit_r49_c238 bl_238 br_238 wl_49 vdd gnd cell_6t
Xbit_r50_c238 bl_238 br_238 wl_50 vdd gnd cell_6t
Xbit_r51_c238 bl_238 br_238 wl_51 vdd gnd cell_6t
Xbit_r52_c238 bl_238 br_238 wl_52 vdd gnd cell_6t
Xbit_r53_c238 bl_238 br_238 wl_53 vdd gnd cell_6t
Xbit_r54_c238 bl_238 br_238 wl_54 vdd gnd cell_6t
Xbit_r55_c238 bl_238 br_238 wl_55 vdd gnd cell_6t
Xbit_r56_c238 bl_238 br_238 wl_56 vdd gnd cell_6t
Xbit_r57_c238 bl_238 br_238 wl_57 vdd gnd cell_6t
Xbit_r58_c238 bl_238 br_238 wl_58 vdd gnd cell_6t
Xbit_r59_c238 bl_238 br_238 wl_59 vdd gnd cell_6t
Xbit_r60_c238 bl_238 br_238 wl_60 vdd gnd cell_6t
Xbit_r61_c238 bl_238 br_238 wl_61 vdd gnd cell_6t
Xbit_r62_c238 bl_238 br_238 wl_62 vdd gnd cell_6t
Xbit_r63_c238 bl_238 br_238 wl_63 vdd gnd cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd cell_6t
Xbit_r1_c239 bl_239 br_239 wl_1 vdd gnd cell_6t
Xbit_r2_c239 bl_239 br_239 wl_2 vdd gnd cell_6t
Xbit_r3_c239 bl_239 br_239 wl_3 vdd gnd cell_6t
Xbit_r4_c239 bl_239 br_239 wl_4 vdd gnd cell_6t
Xbit_r5_c239 bl_239 br_239 wl_5 vdd gnd cell_6t
Xbit_r6_c239 bl_239 br_239 wl_6 vdd gnd cell_6t
Xbit_r7_c239 bl_239 br_239 wl_7 vdd gnd cell_6t
Xbit_r8_c239 bl_239 br_239 wl_8 vdd gnd cell_6t
Xbit_r9_c239 bl_239 br_239 wl_9 vdd gnd cell_6t
Xbit_r10_c239 bl_239 br_239 wl_10 vdd gnd cell_6t
Xbit_r11_c239 bl_239 br_239 wl_11 vdd gnd cell_6t
Xbit_r12_c239 bl_239 br_239 wl_12 vdd gnd cell_6t
Xbit_r13_c239 bl_239 br_239 wl_13 vdd gnd cell_6t
Xbit_r14_c239 bl_239 br_239 wl_14 vdd gnd cell_6t
Xbit_r15_c239 bl_239 br_239 wl_15 vdd gnd cell_6t
Xbit_r16_c239 bl_239 br_239 wl_16 vdd gnd cell_6t
Xbit_r17_c239 bl_239 br_239 wl_17 vdd gnd cell_6t
Xbit_r18_c239 bl_239 br_239 wl_18 vdd gnd cell_6t
Xbit_r19_c239 bl_239 br_239 wl_19 vdd gnd cell_6t
Xbit_r20_c239 bl_239 br_239 wl_20 vdd gnd cell_6t
Xbit_r21_c239 bl_239 br_239 wl_21 vdd gnd cell_6t
Xbit_r22_c239 bl_239 br_239 wl_22 vdd gnd cell_6t
Xbit_r23_c239 bl_239 br_239 wl_23 vdd gnd cell_6t
Xbit_r24_c239 bl_239 br_239 wl_24 vdd gnd cell_6t
Xbit_r25_c239 bl_239 br_239 wl_25 vdd gnd cell_6t
Xbit_r26_c239 bl_239 br_239 wl_26 vdd gnd cell_6t
Xbit_r27_c239 bl_239 br_239 wl_27 vdd gnd cell_6t
Xbit_r28_c239 bl_239 br_239 wl_28 vdd gnd cell_6t
Xbit_r29_c239 bl_239 br_239 wl_29 vdd gnd cell_6t
Xbit_r30_c239 bl_239 br_239 wl_30 vdd gnd cell_6t
Xbit_r31_c239 bl_239 br_239 wl_31 vdd gnd cell_6t
Xbit_r32_c239 bl_239 br_239 wl_32 vdd gnd cell_6t
Xbit_r33_c239 bl_239 br_239 wl_33 vdd gnd cell_6t
Xbit_r34_c239 bl_239 br_239 wl_34 vdd gnd cell_6t
Xbit_r35_c239 bl_239 br_239 wl_35 vdd gnd cell_6t
Xbit_r36_c239 bl_239 br_239 wl_36 vdd gnd cell_6t
Xbit_r37_c239 bl_239 br_239 wl_37 vdd gnd cell_6t
Xbit_r38_c239 bl_239 br_239 wl_38 vdd gnd cell_6t
Xbit_r39_c239 bl_239 br_239 wl_39 vdd gnd cell_6t
Xbit_r40_c239 bl_239 br_239 wl_40 vdd gnd cell_6t
Xbit_r41_c239 bl_239 br_239 wl_41 vdd gnd cell_6t
Xbit_r42_c239 bl_239 br_239 wl_42 vdd gnd cell_6t
Xbit_r43_c239 bl_239 br_239 wl_43 vdd gnd cell_6t
Xbit_r44_c239 bl_239 br_239 wl_44 vdd gnd cell_6t
Xbit_r45_c239 bl_239 br_239 wl_45 vdd gnd cell_6t
Xbit_r46_c239 bl_239 br_239 wl_46 vdd gnd cell_6t
Xbit_r47_c239 bl_239 br_239 wl_47 vdd gnd cell_6t
Xbit_r48_c239 bl_239 br_239 wl_48 vdd gnd cell_6t
Xbit_r49_c239 bl_239 br_239 wl_49 vdd gnd cell_6t
Xbit_r50_c239 bl_239 br_239 wl_50 vdd gnd cell_6t
Xbit_r51_c239 bl_239 br_239 wl_51 vdd gnd cell_6t
Xbit_r52_c239 bl_239 br_239 wl_52 vdd gnd cell_6t
Xbit_r53_c239 bl_239 br_239 wl_53 vdd gnd cell_6t
Xbit_r54_c239 bl_239 br_239 wl_54 vdd gnd cell_6t
Xbit_r55_c239 bl_239 br_239 wl_55 vdd gnd cell_6t
Xbit_r56_c239 bl_239 br_239 wl_56 vdd gnd cell_6t
Xbit_r57_c239 bl_239 br_239 wl_57 vdd gnd cell_6t
Xbit_r58_c239 bl_239 br_239 wl_58 vdd gnd cell_6t
Xbit_r59_c239 bl_239 br_239 wl_59 vdd gnd cell_6t
Xbit_r60_c239 bl_239 br_239 wl_60 vdd gnd cell_6t
Xbit_r61_c239 bl_239 br_239 wl_61 vdd gnd cell_6t
Xbit_r62_c239 bl_239 br_239 wl_62 vdd gnd cell_6t
Xbit_r63_c239 bl_239 br_239 wl_63 vdd gnd cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd cell_6t
Xbit_r1_c240 bl_240 br_240 wl_1 vdd gnd cell_6t
Xbit_r2_c240 bl_240 br_240 wl_2 vdd gnd cell_6t
Xbit_r3_c240 bl_240 br_240 wl_3 vdd gnd cell_6t
Xbit_r4_c240 bl_240 br_240 wl_4 vdd gnd cell_6t
Xbit_r5_c240 bl_240 br_240 wl_5 vdd gnd cell_6t
Xbit_r6_c240 bl_240 br_240 wl_6 vdd gnd cell_6t
Xbit_r7_c240 bl_240 br_240 wl_7 vdd gnd cell_6t
Xbit_r8_c240 bl_240 br_240 wl_8 vdd gnd cell_6t
Xbit_r9_c240 bl_240 br_240 wl_9 vdd gnd cell_6t
Xbit_r10_c240 bl_240 br_240 wl_10 vdd gnd cell_6t
Xbit_r11_c240 bl_240 br_240 wl_11 vdd gnd cell_6t
Xbit_r12_c240 bl_240 br_240 wl_12 vdd gnd cell_6t
Xbit_r13_c240 bl_240 br_240 wl_13 vdd gnd cell_6t
Xbit_r14_c240 bl_240 br_240 wl_14 vdd gnd cell_6t
Xbit_r15_c240 bl_240 br_240 wl_15 vdd gnd cell_6t
Xbit_r16_c240 bl_240 br_240 wl_16 vdd gnd cell_6t
Xbit_r17_c240 bl_240 br_240 wl_17 vdd gnd cell_6t
Xbit_r18_c240 bl_240 br_240 wl_18 vdd gnd cell_6t
Xbit_r19_c240 bl_240 br_240 wl_19 vdd gnd cell_6t
Xbit_r20_c240 bl_240 br_240 wl_20 vdd gnd cell_6t
Xbit_r21_c240 bl_240 br_240 wl_21 vdd gnd cell_6t
Xbit_r22_c240 bl_240 br_240 wl_22 vdd gnd cell_6t
Xbit_r23_c240 bl_240 br_240 wl_23 vdd gnd cell_6t
Xbit_r24_c240 bl_240 br_240 wl_24 vdd gnd cell_6t
Xbit_r25_c240 bl_240 br_240 wl_25 vdd gnd cell_6t
Xbit_r26_c240 bl_240 br_240 wl_26 vdd gnd cell_6t
Xbit_r27_c240 bl_240 br_240 wl_27 vdd gnd cell_6t
Xbit_r28_c240 bl_240 br_240 wl_28 vdd gnd cell_6t
Xbit_r29_c240 bl_240 br_240 wl_29 vdd gnd cell_6t
Xbit_r30_c240 bl_240 br_240 wl_30 vdd gnd cell_6t
Xbit_r31_c240 bl_240 br_240 wl_31 vdd gnd cell_6t
Xbit_r32_c240 bl_240 br_240 wl_32 vdd gnd cell_6t
Xbit_r33_c240 bl_240 br_240 wl_33 vdd gnd cell_6t
Xbit_r34_c240 bl_240 br_240 wl_34 vdd gnd cell_6t
Xbit_r35_c240 bl_240 br_240 wl_35 vdd gnd cell_6t
Xbit_r36_c240 bl_240 br_240 wl_36 vdd gnd cell_6t
Xbit_r37_c240 bl_240 br_240 wl_37 vdd gnd cell_6t
Xbit_r38_c240 bl_240 br_240 wl_38 vdd gnd cell_6t
Xbit_r39_c240 bl_240 br_240 wl_39 vdd gnd cell_6t
Xbit_r40_c240 bl_240 br_240 wl_40 vdd gnd cell_6t
Xbit_r41_c240 bl_240 br_240 wl_41 vdd gnd cell_6t
Xbit_r42_c240 bl_240 br_240 wl_42 vdd gnd cell_6t
Xbit_r43_c240 bl_240 br_240 wl_43 vdd gnd cell_6t
Xbit_r44_c240 bl_240 br_240 wl_44 vdd gnd cell_6t
Xbit_r45_c240 bl_240 br_240 wl_45 vdd gnd cell_6t
Xbit_r46_c240 bl_240 br_240 wl_46 vdd gnd cell_6t
Xbit_r47_c240 bl_240 br_240 wl_47 vdd gnd cell_6t
Xbit_r48_c240 bl_240 br_240 wl_48 vdd gnd cell_6t
Xbit_r49_c240 bl_240 br_240 wl_49 vdd gnd cell_6t
Xbit_r50_c240 bl_240 br_240 wl_50 vdd gnd cell_6t
Xbit_r51_c240 bl_240 br_240 wl_51 vdd gnd cell_6t
Xbit_r52_c240 bl_240 br_240 wl_52 vdd gnd cell_6t
Xbit_r53_c240 bl_240 br_240 wl_53 vdd gnd cell_6t
Xbit_r54_c240 bl_240 br_240 wl_54 vdd gnd cell_6t
Xbit_r55_c240 bl_240 br_240 wl_55 vdd gnd cell_6t
Xbit_r56_c240 bl_240 br_240 wl_56 vdd gnd cell_6t
Xbit_r57_c240 bl_240 br_240 wl_57 vdd gnd cell_6t
Xbit_r58_c240 bl_240 br_240 wl_58 vdd gnd cell_6t
Xbit_r59_c240 bl_240 br_240 wl_59 vdd gnd cell_6t
Xbit_r60_c240 bl_240 br_240 wl_60 vdd gnd cell_6t
Xbit_r61_c240 bl_240 br_240 wl_61 vdd gnd cell_6t
Xbit_r62_c240 bl_240 br_240 wl_62 vdd gnd cell_6t
Xbit_r63_c240 bl_240 br_240 wl_63 vdd gnd cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd cell_6t
Xbit_r1_c241 bl_241 br_241 wl_1 vdd gnd cell_6t
Xbit_r2_c241 bl_241 br_241 wl_2 vdd gnd cell_6t
Xbit_r3_c241 bl_241 br_241 wl_3 vdd gnd cell_6t
Xbit_r4_c241 bl_241 br_241 wl_4 vdd gnd cell_6t
Xbit_r5_c241 bl_241 br_241 wl_5 vdd gnd cell_6t
Xbit_r6_c241 bl_241 br_241 wl_6 vdd gnd cell_6t
Xbit_r7_c241 bl_241 br_241 wl_7 vdd gnd cell_6t
Xbit_r8_c241 bl_241 br_241 wl_8 vdd gnd cell_6t
Xbit_r9_c241 bl_241 br_241 wl_9 vdd gnd cell_6t
Xbit_r10_c241 bl_241 br_241 wl_10 vdd gnd cell_6t
Xbit_r11_c241 bl_241 br_241 wl_11 vdd gnd cell_6t
Xbit_r12_c241 bl_241 br_241 wl_12 vdd gnd cell_6t
Xbit_r13_c241 bl_241 br_241 wl_13 vdd gnd cell_6t
Xbit_r14_c241 bl_241 br_241 wl_14 vdd gnd cell_6t
Xbit_r15_c241 bl_241 br_241 wl_15 vdd gnd cell_6t
Xbit_r16_c241 bl_241 br_241 wl_16 vdd gnd cell_6t
Xbit_r17_c241 bl_241 br_241 wl_17 vdd gnd cell_6t
Xbit_r18_c241 bl_241 br_241 wl_18 vdd gnd cell_6t
Xbit_r19_c241 bl_241 br_241 wl_19 vdd gnd cell_6t
Xbit_r20_c241 bl_241 br_241 wl_20 vdd gnd cell_6t
Xbit_r21_c241 bl_241 br_241 wl_21 vdd gnd cell_6t
Xbit_r22_c241 bl_241 br_241 wl_22 vdd gnd cell_6t
Xbit_r23_c241 bl_241 br_241 wl_23 vdd gnd cell_6t
Xbit_r24_c241 bl_241 br_241 wl_24 vdd gnd cell_6t
Xbit_r25_c241 bl_241 br_241 wl_25 vdd gnd cell_6t
Xbit_r26_c241 bl_241 br_241 wl_26 vdd gnd cell_6t
Xbit_r27_c241 bl_241 br_241 wl_27 vdd gnd cell_6t
Xbit_r28_c241 bl_241 br_241 wl_28 vdd gnd cell_6t
Xbit_r29_c241 bl_241 br_241 wl_29 vdd gnd cell_6t
Xbit_r30_c241 bl_241 br_241 wl_30 vdd gnd cell_6t
Xbit_r31_c241 bl_241 br_241 wl_31 vdd gnd cell_6t
Xbit_r32_c241 bl_241 br_241 wl_32 vdd gnd cell_6t
Xbit_r33_c241 bl_241 br_241 wl_33 vdd gnd cell_6t
Xbit_r34_c241 bl_241 br_241 wl_34 vdd gnd cell_6t
Xbit_r35_c241 bl_241 br_241 wl_35 vdd gnd cell_6t
Xbit_r36_c241 bl_241 br_241 wl_36 vdd gnd cell_6t
Xbit_r37_c241 bl_241 br_241 wl_37 vdd gnd cell_6t
Xbit_r38_c241 bl_241 br_241 wl_38 vdd gnd cell_6t
Xbit_r39_c241 bl_241 br_241 wl_39 vdd gnd cell_6t
Xbit_r40_c241 bl_241 br_241 wl_40 vdd gnd cell_6t
Xbit_r41_c241 bl_241 br_241 wl_41 vdd gnd cell_6t
Xbit_r42_c241 bl_241 br_241 wl_42 vdd gnd cell_6t
Xbit_r43_c241 bl_241 br_241 wl_43 vdd gnd cell_6t
Xbit_r44_c241 bl_241 br_241 wl_44 vdd gnd cell_6t
Xbit_r45_c241 bl_241 br_241 wl_45 vdd gnd cell_6t
Xbit_r46_c241 bl_241 br_241 wl_46 vdd gnd cell_6t
Xbit_r47_c241 bl_241 br_241 wl_47 vdd gnd cell_6t
Xbit_r48_c241 bl_241 br_241 wl_48 vdd gnd cell_6t
Xbit_r49_c241 bl_241 br_241 wl_49 vdd gnd cell_6t
Xbit_r50_c241 bl_241 br_241 wl_50 vdd gnd cell_6t
Xbit_r51_c241 bl_241 br_241 wl_51 vdd gnd cell_6t
Xbit_r52_c241 bl_241 br_241 wl_52 vdd gnd cell_6t
Xbit_r53_c241 bl_241 br_241 wl_53 vdd gnd cell_6t
Xbit_r54_c241 bl_241 br_241 wl_54 vdd gnd cell_6t
Xbit_r55_c241 bl_241 br_241 wl_55 vdd gnd cell_6t
Xbit_r56_c241 bl_241 br_241 wl_56 vdd gnd cell_6t
Xbit_r57_c241 bl_241 br_241 wl_57 vdd gnd cell_6t
Xbit_r58_c241 bl_241 br_241 wl_58 vdd gnd cell_6t
Xbit_r59_c241 bl_241 br_241 wl_59 vdd gnd cell_6t
Xbit_r60_c241 bl_241 br_241 wl_60 vdd gnd cell_6t
Xbit_r61_c241 bl_241 br_241 wl_61 vdd gnd cell_6t
Xbit_r62_c241 bl_241 br_241 wl_62 vdd gnd cell_6t
Xbit_r63_c241 bl_241 br_241 wl_63 vdd gnd cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd cell_6t
Xbit_r1_c242 bl_242 br_242 wl_1 vdd gnd cell_6t
Xbit_r2_c242 bl_242 br_242 wl_2 vdd gnd cell_6t
Xbit_r3_c242 bl_242 br_242 wl_3 vdd gnd cell_6t
Xbit_r4_c242 bl_242 br_242 wl_4 vdd gnd cell_6t
Xbit_r5_c242 bl_242 br_242 wl_5 vdd gnd cell_6t
Xbit_r6_c242 bl_242 br_242 wl_6 vdd gnd cell_6t
Xbit_r7_c242 bl_242 br_242 wl_7 vdd gnd cell_6t
Xbit_r8_c242 bl_242 br_242 wl_8 vdd gnd cell_6t
Xbit_r9_c242 bl_242 br_242 wl_9 vdd gnd cell_6t
Xbit_r10_c242 bl_242 br_242 wl_10 vdd gnd cell_6t
Xbit_r11_c242 bl_242 br_242 wl_11 vdd gnd cell_6t
Xbit_r12_c242 bl_242 br_242 wl_12 vdd gnd cell_6t
Xbit_r13_c242 bl_242 br_242 wl_13 vdd gnd cell_6t
Xbit_r14_c242 bl_242 br_242 wl_14 vdd gnd cell_6t
Xbit_r15_c242 bl_242 br_242 wl_15 vdd gnd cell_6t
Xbit_r16_c242 bl_242 br_242 wl_16 vdd gnd cell_6t
Xbit_r17_c242 bl_242 br_242 wl_17 vdd gnd cell_6t
Xbit_r18_c242 bl_242 br_242 wl_18 vdd gnd cell_6t
Xbit_r19_c242 bl_242 br_242 wl_19 vdd gnd cell_6t
Xbit_r20_c242 bl_242 br_242 wl_20 vdd gnd cell_6t
Xbit_r21_c242 bl_242 br_242 wl_21 vdd gnd cell_6t
Xbit_r22_c242 bl_242 br_242 wl_22 vdd gnd cell_6t
Xbit_r23_c242 bl_242 br_242 wl_23 vdd gnd cell_6t
Xbit_r24_c242 bl_242 br_242 wl_24 vdd gnd cell_6t
Xbit_r25_c242 bl_242 br_242 wl_25 vdd gnd cell_6t
Xbit_r26_c242 bl_242 br_242 wl_26 vdd gnd cell_6t
Xbit_r27_c242 bl_242 br_242 wl_27 vdd gnd cell_6t
Xbit_r28_c242 bl_242 br_242 wl_28 vdd gnd cell_6t
Xbit_r29_c242 bl_242 br_242 wl_29 vdd gnd cell_6t
Xbit_r30_c242 bl_242 br_242 wl_30 vdd gnd cell_6t
Xbit_r31_c242 bl_242 br_242 wl_31 vdd gnd cell_6t
Xbit_r32_c242 bl_242 br_242 wl_32 vdd gnd cell_6t
Xbit_r33_c242 bl_242 br_242 wl_33 vdd gnd cell_6t
Xbit_r34_c242 bl_242 br_242 wl_34 vdd gnd cell_6t
Xbit_r35_c242 bl_242 br_242 wl_35 vdd gnd cell_6t
Xbit_r36_c242 bl_242 br_242 wl_36 vdd gnd cell_6t
Xbit_r37_c242 bl_242 br_242 wl_37 vdd gnd cell_6t
Xbit_r38_c242 bl_242 br_242 wl_38 vdd gnd cell_6t
Xbit_r39_c242 bl_242 br_242 wl_39 vdd gnd cell_6t
Xbit_r40_c242 bl_242 br_242 wl_40 vdd gnd cell_6t
Xbit_r41_c242 bl_242 br_242 wl_41 vdd gnd cell_6t
Xbit_r42_c242 bl_242 br_242 wl_42 vdd gnd cell_6t
Xbit_r43_c242 bl_242 br_242 wl_43 vdd gnd cell_6t
Xbit_r44_c242 bl_242 br_242 wl_44 vdd gnd cell_6t
Xbit_r45_c242 bl_242 br_242 wl_45 vdd gnd cell_6t
Xbit_r46_c242 bl_242 br_242 wl_46 vdd gnd cell_6t
Xbit_r47_c242 bl_242 br_242 wl_47 vdd gnd cell_6t
Xbit_r48_c242 bl_242 br_242 wl_48 vdd gnd cell_6t
Xbit_r49_c242 bl_242 br_242 wl_49 vdd gnd cell_6t
Xbit_r50_c242 bl_242 br_242 wl_50 vdd gnd cell_6t
Xbit_r51_c242 bl_242 br_242 wl_51 vdd gnd cell_6t
Xbit_r52_c242 bl_242 br_242 wl_52 vdd gnd cell_6t
Xbit_r53_c242 bl_242 br_242 wl_53 vdd gnd cell_6t
Xbit_r54_c242 bl_242 br_242 wl_54 vdd gnd cell_6t
Xbit_r55_c242 bl_242 br_242 wl_55 vdd gnd cell_6t
Xbit_r56_c242 bl_242 br_242 wl_56 vdd gnd cell_6t
Xbit_r57_c242 bl_242 br_242 wl_57 vdd gnd cell_6t
Xbit_r58_c242 bl_242 br_242 wl_58 vdd gnd cell_6t
Xbit_r59_c242 bl_242 br_242 wl_59 vdd gnd cell_6t
Xbit_r60_c242 bl_242 br_242 wl_60 vdd gnd cell_6t
Xbit_r61_c242 bl_242 br_242 wl_61 vdd gnd cell_6t
Xbit_r62_c242 bl_242 br_242 wl_62 vdd gnd cell_6t
Xbit_r63_c242 bl_242 br_242 wl_63 vdd gnd cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd cell_6t
Xbit_r1_c243 bl_243 br_243 wl_1 vdd gnd cell_6t
Xbit_r2_c243 bl_243 br_243 wl_2 vdd gnd cell_6t
Xbit_r3_c243 bl_243 br_243 wl_3 vdd gnd cell_6t
Xbit_r4_c243 bl_243 br_243 wl_4 vdd gnd cell_6t
Xbit_r5_c243 bl_243 br_243 wl_5 vdd gnd cell_6t
Xbit_r6_c243 bl_243 br_243 wl_6 vdd gnd cell_6t
Xbit_r7_c243 bl_243 br_243 wl_7 vdd gnd cell_6t
Xbit_r8_c243 bl_243 br_243 wl_8 vdd gnd cell_6t
Xbit_r9_c243 bl_243 br_243 wl_9 vdd gnd cell_6t
Xbit_r10_c243 bl_243 br_243 wl_10 vdd gnd cell_6t
Xbit_r11_c243 bl_243 br_243 wl_11 vdd gnd cell_6t
Xbit_r12_c243 bl_243 br_243 wl_12 vdd gnd cell_6t
Xbit_r13_c243 bl_243 br_243 wl_13 vdd gnd cell_6t
Xbit_r14_c243 bl_243 br_243 wl_14 vdd gnd cell_6t
Xbit_r15_c243 bl_243 br_243 wl_15 vdd gnd cell_6t
Xbit_r16_c243 bl_243 br_243 wl_16 vdd gnd cell_6t
Xbit_r17_c243 bl_243 br_243 wl_17 vdd gnd cell_6t
Xbit_r18_c243 bl_243 br_243 wl_18 vdd gnd cell_6t
Xbit_r19_c243 bl_243 br_243 wl_19 vdd gnd cell_6t
Xbit_r20_c243 bl_243 br_243 wl_20 vdd gnd cell_6t
Xbit_r21_c243 bl_243 br_243 wl_21 vdd gnd cell_6t
Xbit_r22_c243 bl_243 br_243 wl_22 vdd gnd cell_6t
Xbit_r23_c243 bl_243 br_243 wl_23 vdd gnd cell_6t
Xbit_r24_c243 bl_243 br_243 wl_24 vdd gnd cell_6t
Xbit_r25_c243 bl_243 br_243 wl_25 vdd gnd cell_6t
Xbit_r26_c243 bl_243 br_243 wl_26 vdd gnd cell_6t
Xbit_r27_c243 bl_243 br_243 wl_27 vdd gnd cell_6t
Xbit_r28_c243 bl_243 br_243 wl_28 vdd gnd cell_6t
Xbit_r29_c243 bl_243 br_243 wl_29 vdd gnd cell_6t
Xbit_r30_c243 bl_243 br_243 wl_30 vdd gnd cell_6t
Xbit_r31_c243 bl_243 br_243 wl_31 vdd gnd cell_6t
Xbit_r32_c243 bl_243 br_243 wl_32 vdd gnd cell_6t
Xbit_r33_c243 bl_243 br_243 wl_33 vdd gnd cell_6t
Xbit_r34_c243 bl_243 br_243 wl_34 vdd gnd cell_6t
Xbit_r35_c243 bl_243 br_243 wl_35 vdd gnd cell_6t
Xbit_r36_c243 bl_243 br_243 wl_36 vdd gnd cell_6t
Xbit_r37_c243 bl_243 br_243 wl_37 vdd gnd cell_6t
Xbit_r38_c243 bl_243 br_243 wl_38 vdd gnd cell_6t
Xbit_r39_c243 bl_243 br_243 wl_39 vdd gnd cell_6t
Xbit_r40_c243 bl_243 br_243 wl_40 vdd gnd cell_6t
Xbit_r41_c243 bl_243 br_243 wl_41 vdd gnd cell_6t
Xbit_r42_c243 bl_243 br_243 wl_42 vdd gnd cell_6t
Xbit_r43_c243 bl_243 br_243 wl_43 vdd gnd cell_6t
Xbit_r44_c243 bl_243 br_243 wl_44 vdd gnd cell_6t
Xbit_r45_c243 bl_243 br_243 wl_45 vdd gnd cell_6t
Xbit_r46_c243 bl_243 br_243 wl_46 vdd gnd cell_6t
Xbit_r47_c243 bl_243 br_243 wl_47 vdd gnd cell_6t
Xbit_r48_c243 bl_243 br_243 wl_48 vdd gnd cell_6t
Xbit_r49_c243 bl_243 br_243 wl_49 vdd gnd cell_6t
Xbit_r50_c243 bl_243 br_243 wl_50 vdd gnd cell_6t
Xbit_r51_c243 bl_243 br_243 wl_51 vdd gnd cell_6t
Xbit_r52_c243 bl_243 br_243 wl_52 vdd gnd cell_6t
Xbit_r53_c243 bl_243 br_243 wl_53 vdd gnd cell_6t
Xbit_r54_c243 bl_243 br_243 wl_54 vdd gnd cell_6t
Xbit_r55_c243 bl_243 br_243 wl_55 vdd gnd cell_6t
Xbit_r56_c243 bl_243 br_243 wl_56 vdd gnd cell_6t
Xbit_r57_c243 bl_243 br_243 wl_57 vdd gnd cell_6t
Xbit_r58_c243 bl_243 br_243 wl_58 vdd gnd cell_6t
Xbit_r59_c243 bl_243 br_243 wl_59 vdd gnd cell_6t
Xbit_r60_c243 bl_243 br_243 wl_60 vdd gnd cell_6t
Xbit_r61_c243 bl_243 br_243 wl_61 vdd gnd cell_6t
Xbit_r62_c243 bl_243 br_243 wl_62 vdd gnd cell_6t
Xbit_r63_c243 bl_243 br_243 wl_63 vdd gnd cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd cell_6t
Xbit_r1_c244 bl_244 br_244 wl_1 vdd gnd cell_6t
Xbit_r2_c244 bl_244 br_244 wl_2 vdd gnd cell_6t
Xbit_r3_c244 bl_244 br_244 wl_3 vdd gnd cell_6t
Xbit_r4_c244 bl_244 br_244 wl_4 vdd gnd cell_6t
Xbit_r5_c244 bl_244 br_244 wl_5 vdd gnd cell_6t
Xbit_r6_c244 bl_244 br_244 wl_6 vdd gnd cell_6t
Xbit_r7_c244 bl_244 br_244 wl_7 vdd gnd cell_6t
Xbit_r8_c244 bl_244 br_244 wl_8 vdd gnd cell_6t
Xbit_r9_c244 bl_244 br_244 wl_9 vdd gnd cell_6t
Xbit_r10_c244 bl_244 br_244 wl_10 vdd gnd cell_6t
Xbit_r11_c244 bl_244 br_244 wl_11 vdd gnd cell_6t
Xbit_r12_c244 bl_244 br_244 wl_12 vdd gnd cell_6t
Xbit_r13_c244 bl_244 br_244 wl_13 vdd gnd cell_6t
Xbit_r14_c244 bl_244 br_244 wl_14 vdd gnd cell_6t
Xbit_r15_c244 bl_244 br_244 wl_15 vdd gnd cell_6t
Xbit_r16_c244 bl_244 br_244 wl_16 vdd gnd cell_6t
Xbit_r17_c244 bl_244 br_244 wl_17 vdd gnd cell_6t
Xbit_r18_c244 bl_244 br_244 wl_18 vdd gnd cell_6t
Xbit_r19_c244 bl_244 br_244 wl_19 vdd gnd cell_6t
Xbit_r20_c244 bl_244 br_244 wl_20 vdd gnd cell_6t
Xbit_r21_c244 bl_244 br_244 wl_21 vdd gnd cell_6t
Xbit_r22_c244 bl_244 br_244 wl_22 vdd gnd cell_6t
Xbit_r23_c244 bl_244 br_244 wl_23 vdd gnd cell_6t
Xbit_r24_c244 bl_244 br_244 wl_24 vdd gnd cell_6t
Xbit_r25_c244 bl_244 br_244 wl_25 vdd gnd cell_6t
Xbit_r26_c244 bl_244 br_244 wl_26 vdd gnd cell_6t
Xbit_r27_c244 bl_244 br_244 wl_27 vdd gnd cell_6t
Xbit_r28_c244 bl_244 br_244 wl_28 vdd gnd cell_6t
Xbit_r29_c244 bl_244 br_244 wl_29 vdd gnd cell_6t
Xbit_r30_c244 bl_244 br_244 wl_30 vdd gnd cell_6t
Xbit_r31_c244 bl_244 br_244 wl_31 vdd gnd cell_6t
Xbit_r32_c244 bl_244 br_244 wl_32 vdd gnd cell_6t
Xbit_r33_c244 bl_244 br_244 wl_33 vdd gnd cell_6t
Xbit_r34_c244 bl_244 br_244 wl_34 vdd gnd cell_6t
Xbit_r35_c244 bl_244 br_244 wl_35 vdd gnd cell_6t
Xbit_r36_c244 bl_244 br_244 wl_36 vdd gnd cell_6t
Xbit_r37_c244 bl_244 br_244 wl_37 vdd gnd cell_6t
Xbit_r38_c244 bl_244 br_244 wl_38 vdd gnd cell_6t
Xbit_r39_c244 bl_244 br_244 wl_39 vdd gnd cell_6t
Xbit_r40_c244 bl_244 br_244 wl_40 vdd gnd cell_6t
Xbit_r41_c244 bl_244 br_244 wl_41 vdd gnd cell_6t
Xbit_r42_c244 bl_244 br_244 wl_42 vdd gnd cell_6t
Xbit_r43_c244 bl_244 br_244 wl_43 vdd gnd cell_6t
Xbit_r44_c244 bl_244 br_244 wl_44 vdd gnd cell_6t
Xbit_r45_c244 bl_244 br_244 wl_45 vdd gnd cell_6t
Xbit_r46_c244 bl_244 br_244 wl_46 vdd gnd cell_6t
Xbit_r47_c244 bl_244 br_244 wl_47 vdd gnd cell_6t
Xbit_r48_c244 bl_244 br_244 wl_48 vdd gnd cell_6t
Xbit_r49_c244 bl_244 br_244 wl_49 vdd gnd cell_6t
Xbit_r50_c244 bl_244 br_244 wl_50 vdd gnd cell_6t
Xbit_r51_c244 bl_244 br_244 wl_51 vdd gnd cell_6t
Xbit_r52_c244 bl_244 br_244 wl_52 vdd gnd cell_6t
Xbit_r53_c244 bl_244 br_244 wl_53 vdd gnd cell_6t
Xbit_r54_c244 bl_244 br_244 wl_54 vdd gnd cell_6t
Xbit_r55_c244 bl_244 br_244 wl_55 vdd gnd cell_6t
Xbit_r56_c244 bl_244 br_244 wl_56 vdd gnd cell_6t
Xbit_r57_c244 bl_244 br_244 wl_57 vdd gnd cell_6t
Xbit_r58_c244 bl_244 br_244 wl_58 vdd gnd cell_6t
Xbit_r59_c244 bl_244 br_244 wl_59 vdd gnd cell_6t
Xbit_r60_c244 bl_244 br_244 wl_60 vdd gnd cell_6t
Xbit_r61_c244 bl_244 br_244 wl_61 vdd gnd cell_6t
Xbit_r62_c244 bl_244 br_244 wl_62 vdd gnd cell_6t
Xbit_r63_c244 bl_244 br_244 wl_63 vdd gnd cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd cell_6t
Xbit_r1_c245 bl_245 br_245 wl_1 vdd gnd cell_6t
Xbit_r2_c245 bl_245 br_245 wl_2 vdd gnd cell_6t
Xbit_r3_c245 bl_245 br_245 wl_3 vdd gnd cell_6t
Xbit_r4_c245 bl_245 br_245 wl_4 vdd gnd cell_6t
Xbit_r5_c245 bl_245 br_245 wl_5 vdd gnd cell_6t
Xbit_r6_c245 bl_245 br_245 wl_6 vdd gnd cell_6t
Xbit_r7_c245 bl_245 br_245 wl_7 vdd gnd cell_6t
Xbit_r8_c245 bl_245 br_245 wl_8 vdd gnd cell_6t
Xbit_r9_c245 bl_245 br_245 wl_9 vdd gnd cell_6t
Xbit_r10_c245 bl_245 br_245 wl_10 vdd gnd cell_6t
Xbit_r11_c245 bl_245 br_245 wl_11 vdd gnd cell_6t
Xbit_r12_c245 bl_245 br_245 wl_12 vdd gnd cell_6t
Xbit_r13_c245 bl_245 br_245 wl_13 vdd gnd cell_6t
Xbit_r14_c245 bl_245 br_245 wl_14 vdd gnd cell_6t
Xbit_r15_c245 bl_245 br_245 wl_15 vdd gnd cell_6t
Xbit_r16_c245 bl_245 br_245 wl_16 vdd gnd cell_6t
Xbit_r17_c245 bl_245 br_245 wl_17 vdd gnd cell_6t
Xbit_r18_c245 bl_245 br_245 wl_18 vdd gnd cell_6t
Xbit_r19_c245 bl_245 br_245 wl_19 vdd gnd cell_6t
Xbit_r20_c245 bl_245 br_245 wl_20 vdd gnd cell_6t
Xbit_r21_c245 bl_245 br_245 wl_21 vdd gnd cell_6t
Xbit_r22_c245 bl_245 br_245 wl_22 vdd gnd cell_6t
Xbit_r23_c245 bl_245 br_245 wl_23 vdd gnd cell_6t
Xbit_r24_c245 bl_245 br_245 wl_24 vdd gnd cell_6t
Xbit_r25_c245 bl_245 br_245 wl_25 vdd gnd cell_6t
Xbit_r26_c245 bl_245 br_245 wl_26 vdd gnd cell_6t
Xbit_r27_c245 bl_245 br_245 wl_27 vdd gnd cell_6t
Xbit_r28_c245 bl_245 br_245 wl_28 vdd gnd cell_6t
Xbit_r29_c245 bl_245 br_245 wl_29 vdd gnd cell_6t
Xbit_r30_c245 bl_245 br_245 wl_30 vdd gnd cell_6t
Xbit_r31_c245 bl_245 br_245 wl_31 vdd gnd cell_6t
Xbit_r32_c245 bl_245 br_245 wl_32 vdd gnd cell_6t
Xbit_r33_c245 bl_245 br_245 wl_33 vdd gnd cell_6t
Xbit_r34_c245 bl_245 br_245 wl_34 vdd gnd cell_6t
Xbit_r35_c245 bl_245 br_245 wl_35 vdd gnd cell_6t
Xbit_r36_c245 bl_245 br_245 wl_36 vdd gnd cell_6t
Xbit_r37_c245 bl_245 br_245 wl_37 vdd gnd cell_6t
Xbit_r38_c245 bl_245 br_245 wl_38 vdd gnd cell_6t
Xbit_r39_c245 bl_245 br_245 wl_39 vdd gnd cell_6t
Xbit_r40_c245 bl_245 br_245 wl_40 vdd gnd cell_6t
Xbit_r41_c245 bl_245 br_245 wl_41 vdd gnd cell_6t
Xbit_r42_c245 bl_245 br_245 wl_42 vdd gnd cell_6t
Xbit_r43_c245 bl_245 br_245 wl_43 vdd gnd cell_6t
Xbit_r44_c245 bl_245 br_245 wl_44 vdd gnd cell_6t
Xbit_r45_c245 bl_245 br_245 wl_45 vdd gnd cell_6t
Xbit_r46_c245 bl_245 br_245 wl_46 vdd gnd cell_6t
Xbit_r47_c245 bl_245 br_245 wl_47 vdd gnd cell_6t
Xbit_r48_c245 bl_245 br_245 wl_48 vdd gnd cell_6t
Xbit_r49_c245 bl_245 br_245 wl_49 vdd gnd cell_6t
Xbit_r50_c245 bl_245 br_245 wl_50 vdd gnd cell_6t
Xbit_r51_c245 bl_245 br_245 wl_51 vdd gnd cell_6t
Xbit_r52_c245 bl_245 br_245 wl_52 vdd gnd cell_6t
Xbit_r53_c245 bl_245 br_245 wl_53 vdd gnd cell_6t
Xbit_r54_c245 bl_245 br_245 wl_54 vdd gnd cell_6t
Xbit_r55_c245 bl_245 br_245 wl_55 vdd gnd cell_6t
Xbit_r56_c245 bl_245 br_245 wl_56 vdd gnd cell_6t
Xbit_r57_c245 bl_245 br_245 wl_57 vdd gnd cell_6t
Xbit_r58_c245 bl_245 br_245 wl_58 vdd gnd cell_6t
Xbit_r59_c245 bl_245 br_245 wl_59 vdd gnd cell_6t
Xbit_r60_c245 bl_245 br_245 wl_60 vdd gnd cell_6t
Xbit_r61_c245 bl_245 br_245 wl_61 vdd gnd cell_6t
Xbit_r62_c245 bl_245 br_245 wl_62 vdd gnd cell_6t
Xbit_r63_c245 bl_245 br_245 wl_63 vdd gnd cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd cell_6t
Xbit_r1_c246 bl_246 br_246 wl_1 vdd gnd cell_6t
Xbit_r2_c246 bl_246 br_246 wl_2 vdd gnd cell_6t
Xbit_r3_c246 bl_246 br_246 wl_3 vdd gnd cell_6t
Xbit_r4_c246 bl_246 br_246 wl_4 vdd gnd cell_6t
Xbit_r5_c246 bl_246 br_246 wl_5 vdd gnd cell_6t
Xbit_r6_c246 bl_246 br_246 wl_6 vdd gnd cell_6t
Xbit_r7_c246 bl_246 br_246 wl_7 vdd gnd cell_6t
Xbit_r8_c246 bl_246 br_246 wl_8 vdd gnd cell_6t
Xbit_r9_c246 bl_246 br_246 wl_9 vdd gnd cell_6t
Xbit_r10_c246 bl_246 br_246 wl_10 vdd gnd cell_6t
Xbit_r11_c246 bl_246 br_246 wl_11 vdd gnd cell_6t
Xbit_r12_c246 bl_246 br_246 wl_12 vdd gnd cell_6t
Xbit_r13_c246 bl_246 br_246 wl_13 vdd gnd cell_6t
Xbit_r14_c246 bl_246 br_246 wl_14 vdd gnd cell_6t
Xbit_r15_c246 bl_246 br_246 wl_15 vdd gnd cell_6t
Xbit_r16_c246 bl_246 br_246 wl_16 vdd gnd cell_6t
Xbit_r17_c246 bl_246 br_246 wl_17 vdd gnd cell_6t
Xbit_r18_c246 bl_246 br_246 wl_18 vdd gnd cell_6t
Xbit_r19_c246 bl_246 br_246 wl_19 vdd gnd cell_6t
Xbit_r20_c246 bl_246 br_246 wl_20 vdd gnd cell_6t
Xbit_r21_c246 bl_246 br_246 wl_21 vdd gnd cell_6t
Xbit_r22_c246 bl_246 br_246 wl_22 vdd gnd cell_6t
Xbit_r23_c246 bl_246 br_246 wl_23 vdd gnd cell_6t
Xbit_r24_c246 bl_246 br_246 wl_24 vdd gnd cell_6t
Xbit_r25_c246 bl_246 br_246 wl_25 vdd gnd cell_6t
Xbit_r26_c246 bl_246 br_246 wl_26 vdd gnd cell_6t
Xbit_r27_c246 bl_246 br_246 wl_27 vdd gnd cell_6t
Xbit_r28_c246 bl_246 br_246 wl_28 vdd gnd cell_6t
Xbit_r29_c246 bl_246 br_246 wl_29 vdd gnd cell_6t
Xbit_r30_c246 bl_246 br_246 wl_30 vdd gnd cell_6t
Xbit_r31_c246 bl_246 br_246 wl_31 vdd gnd cell_6t
Xbit_r32_c246 bl_246 br_246 wl_32 vdd gnd cell_6t
Xbit_r33_c246 bl_246 br_246 wl_33 vdd gnd cell_6t
Xbit_r34_c246 bl_246 br_246 wl_34 vdd gnd cell_6t
Xbit_r35_c246 bl_246 br_246 wl_35 vdd gnd cell_6t
Xbit_r36_c246 bl_246 br_246 wl_36 vdd gnd cell_6t
Xbit_r37_c246 bl_246 br_246 wl_37 vdd gnd cell_6t
Xbit_r38_c246 bl_246 br_246 wl_38 vdd gnd cell_6t
Xbit_r39_c246 bl_246 br_246 wl_39 vdd gnd cell_6t
Xbit_r40_c246 bl_246 br_246 wl_40 vdd gnd cell_6t
Xbit_r41_c246 bl_246 br_246 wl_41 vdd gnd cell_6t
Xbit_r42_c246 bl_246 br_246 wl_42 vdd gnd cell_6t
Xbit_r43_c246 bl_246 br_246 wl_43 vdd gnd cell_6t
Xbit_r44_c246 bl_246 br_246 wl_44 vdd gnd cell_6t
Xbit_r45_c246 bl_246 br_246 wl_45 vdd gnd cell_6t
Xbit_r46_c246 bl_246 br_246 wl_46 vdd gnd cell_6t
Xbit_r47_c246 bl_246 br_246 wl_47 vdd gnd cell_6t
Xbit_r48_c246 bl_246 br_246 wl_48 vdd gnd cell_6t
Xbit_r49_c246 bl_246 br_246 wl_49 vdd gnd cell_6t
Xbit_r50_c246 bl_246 br_246 wl_50 vdd gnd cell_6t
Xbit_r51_c246 bl_246 br_246 wl_51 vdd gnd cell_6t
Xbit_r52_c246 bl_246 br_246 wl_52 vdd gnd cell_6t
Xbit_r53_c246 bl_246 br_246 wl_53 vdd gnd cell_6t
Xbit_r54_c246 bl_246 br_246 wl_54 vdd gnd cell_6t
Xbit_r55_c246 bl_246 br_246 wl_55 vdd gnd cell_6t
Xbit_r56_c246 bl_246 br_246 wl_56 vdd gnd cell_6t
Xbit_r57_c246 bl_246 br_246 wl_57 vdd gnd cell_6t
Xbit_r58_c246 bl_246 br_246 wl_58 vdd gnd cell_6t
Xbit_r59_c246 bl_246 br_246 wl_59 vdd gnd cell_6t
Xbit_r60_c246 bl_246 br_246 wl_60 vdd gnd cell_6t
Xbit_r61_c246 bl_246 br_246 wl_61 vdd gnd cell_6t
Xbit_r62_c246 bl_246 br_246 wl_62 vdd gnd cell_6t
Xbit_r63_c246 bl_246 br_246 wl_63 vdd gnd cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd cell_6t
Xbit_r1_c247 bl_247 br_247 wl_1 vdd gnd cell_6t
Xbit_r2_c247 bl_247 br_247 wl_2 vdd gnd cell_6t
Xbit_r3_c247 bl_247 br_247 wl_3 vdd gnd cell_6t
Xbit_r4_c247 bl_247 br_247 wl_4 vdd gnd cell_6t
Xbit_r5_c247 bl_247 br_247 wl_5 vdd gnd cell_6t
Xbit_r6_c247 bl_247 br_247 wl_6 vdd gnd cell_6t
Xbit_r7_c247 bl_247 br_247 wl_7 vdd gnd cell_6t
Xbit_r8_c247 bl_247 br_247 wl_8 vdd gnd cell_6t
Xbit_r9_c247 bl_247 br_247 wl_9 vdd gnd cell_6t
Xbit_r10_c247 bl_247 br_247 wl_10 vdd gnd cell_6t
Xbit_r11_c247 bl_247 br_247 wl_11 vdd gnd cell_6t
Xbit_r12_c247 bl_247 br_247 wl_12 vdd gnd cell_6t
Xbit_r13_c247 bl_247 br_247 wl_13 vdd gnd cell_6t
Xbit_r14_c247 bl_247 br_247 wl_14 vdd gnd cell_6t
Xbit_r15_c247 bl_247 br_247 wl_15 vdd gnd cell_6t
Xbit_r16_c247 bl_247 br_247 wl_16 vdd gnd cell_6t
Xbit_r17_c247 bl_247 br_247 wl_17 vdd gnd cell_6t
Xbit_r18_c247 bl_247 br_247 wl_18 vdd gnd cell_6t
Xbit_r19_c247 bl_247 br_247 wl_19 vdd gnd cell_6t
Xbit_r20_c247 bl_247 br_247 wl_20 vdd gnd cell_6t
Xbit_r21_c247 bl_247 br_247 wl_21 vdd gnd cell_6t
Xbit_r22_c247 bl_247 br_247 wl_22 vdd gnd cell_6t
Xbit_r23_c247 bl_247 br_247 wl_23 vdd gnd cell_6t
Xbit_r24_c247 bl_247 br_247 wl_24 vdd gnd cell_6t
Xbit_r25_c247 bl_247 br_247 wl_25 vdd gnd cell_6t
Xbit_r26_c247 bl_247 br_247 wl_26 vdd gnd cell_6t
Xbit_r27_c247 bl_247 br_247 wl_27 vdd gnd cell_6t
Xbit_r28_c247 bl_247 br_247 wl_28 vdd gnd cell_6t
Xbit_r29_c247 bl_247 br_247 wl_29 vdd gnd cell_6t
Xbit_r30_c247 bl_247 br_247 wl_30 vdd gnd cell_6t
Xbit_r31_c247 bl_247 br_247 wl_31 vdd gnd cell_6t
Xbit_r32_c247 bl_247 br_247 wl_32 vdd gnd cell_6t
Xbit_r33_c247 bl_247 br_247 wl_33 vdd gnd cell_6t
Xbit_r34_c247 bl_247 br_247 wl_34 vdd gnd cell_6t
Xbit_r35_c247 bl_247 br_247 wl_35 vdd gnd cell_6t
Xbit_r36_c247 bl_247 br_247 wl_36 vdd gnd cell_6t
Xbit_r37_c247 bl_247 br_247 wl_37 vdd gnd cell_6t
Xbit_r38_c247 bl_247 br_247 wl_38 vdd gnd cell_6t
Xbit_r39_c247 bl_247 br_247 wl_39 vdd gnd cell_6t
Xbit_r40_c247 bl_247 br_247 wl_40 vdd gnd cell_6t
Xbit_r41_c247 bl_247 br_247 wl_41 vdd gnd cell_6t
Xbit_r42_c247 bl_247 br_247 wl_42 vdd gnd cell_6t
Xbit_r43_c247 bl_247 br_247 wl_43 vdd gnd cell_6t
Xbit_r44_c247 bl_247 br_247 wl_44 vdd gnd cell_6t
Xbit_r45_c247 bl_247 br_247 wl_45 vdd gnd cell_6t
Xbit_r46_c247 bl_247 br_247 wl_46 vdd gnd cell_6t
Xbit_r47_c247 bl_247 br_247 wl_47 vdd gnd cell_6t
Xbit_r48_c247 bl_247 br_247 wl_48 vdd gnd cell_6t
Xbit_r49_c247 bl_247 br_247 wl_49 vdd gnd cell_6t
Xbit_r50_c247 bl_247 br_247 wl_50 vdd gnd cell_6t
Xbit_r51_c247 bl_247 br_247 wl_51 vdd gnd cell_6t
Xbit_r52_c247 bl_247 br_247 wl_52 vdd gnd cell_6t
Xbit_r53_c247 bl_247 br_247 wl_53 vdd gnd cell_6t
Xbit_r54_c247 bl_247 br_247 wl_54 vdd gnd cell_6t
Xbit_r55_c247 bl_247 br_247 wl_55 vdd gnd cell_6t
Xbit_r56_c247 bl_247 br_247 wl_56 vdd gnd cell_6t
Xbit_r57_c247 bl_247 br_247 wl_57 vdd gnd cell_6t
Xbit_r58_c247 bl_247 br_247 wl_58 vdd gnd cell_6t
Xbit_r59_c247 bl_247 br_247 wl_59 vdd gnd cell_6t
Xbit_r60_c247 bl_247 br_247 wl_60 vdd gnd cell_6t
Xbit_r61_c247 bl_247 br_247 wl_61 vdd gnd cell_6t
Xbit_r62_c247 bl_247 br_247 wl_62 vdd gnd cell_6t
Xbit_r63_c247 bl_247 br_247 wl_63 vdd gnd cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd cell_6t
Xbit_r1_c248 bl_248 br_248 wl_1 vdd gnd cell_6t
Xbit_r2_c248 bl_248 br_248 wl_2 vdd gnd cell_6t
Xbit_r3_c248 bl_248 br_248 wl_3 vdd gnd cell_6t
Xbit_r4_c248 bl_248 br_248 wl_4 vdd gnd cell_6t
Xbit_r5_c248 bl_248 br_248 wl_5 vdd gnd cell_6t
Xbit_r6_c248 bl_248 br_248 wl_6 vdd gnd cell_6t
Xbit_r7_c248 bl_248 br_248 wl_7 vdd gnd cell_6t
Xbit_r8_c248 bl_248 br_248 wl_8 vdd gnd cell_6t
Xbit_r9_c248 bl_248 br_248 wl_9 vdd gnd cell_6t
Xbit_r10_c248 bl_248 br_248 wl_10 vdd gnd cell_6t
Xbit_r11_c248 bl_248 br_248 wl_11 vdd gnd cell_6t
Xbit_r12_c248 bl_248 br_248 wl_12 vdd gnd cell_6t
Xbit_r13_c248 bl_248 br_248 wl_13 vdd gnd cell_6t
Xbit_r14_c248 bl_248 br_248 wl_14 vdd gnd cell_6t
Xbit_r15_c248 bl_248 br_248 wl_15 vdd gnd cell_6t
Xbit_r16_c248 bl_248 br_248 wl_16 vdd gnd cell_6t
Xbit_r17_c248 bl_248 br_248 wl_17 vdd gnd cell_6t
Xbit_r18_c248 bl_248 br_248 wl_18 vdd gnd cell_6t
Xbit_r19_c248 bl_248 br_248 wl_19 vdd gnd cell_6t
Xbit_r20_c248 bl_248 br_248 wl_20 vdd gnd cell_6t
Xbit_r21_c248 bl_248 br_248 wl_21 vdd gnd cell_6t
Xbit_r22_c248 bl_248 br_248 wl_22 vdd gnd cell_6t
Xbit_r23_c248 bl_248 br_248 wl_23 vdd gnd cell_6t
Xbit_r24_c248 bl_248 br_248 wl_24 vdd gnd cell_6t
Xbit_r25_c248 bl_248 br_248 wl_25 vdd gnd cell_6t
Xbit_r26_c248 bl_248 br_248 wl_26 vdd gnd cell_6t
Xbit_r27_c248 bl_248 br_248 wl_27 vdd gnd cell_6t
Xbit_r28_c248 bl_248 br_248 wl_28 vdd gnd cell_6t
Xbit_r29_c248 bl_248 br_248 wl_29 vdd gnd cell_6t
Xbit_r30_c248 bl_248 br_248 wl_30 vdd gnd cell_6t
Xbit_r31_c248 bl_248 br_248 wl_31 vdd gnd cell_6t
Xbit_r32_c248 bl_248 br_248 wl_32 vdd gnd cell_6t
Xbit_r33_c248 bl_248 br_248 wl_33 vdd gnd cell_6t
Xbit_r34_c248 bl_248 br_248 wl_34 vdd gnd cell_6t
Xbit_r35_c248 bl_248 br_248 wl_35 vdd gnd cell_6t
Xbit_r36_c248 bl_248 br_248 wl_36 vdd gnd cell_6t
Xbit_r37_c248 bl_248 br_248 wl_37 vdd gnd cell_6t
Xbit_r38_c248 bl_248 br_248 wl_38 vdd gnd cell_6t
Xbit_r39_c248 bl_248 br_248 wl_39 vdd gnd cell_6t
Xbit_r40_c248 bl_248 br_248 wl_40 vdd gnd cell_6t
Xbit_r41_c248 bl_248 br_248 wl_41 vdd gnd cell_6t
Xbit_r42_c248 bl_248 br_248 wl_42 vdd gnd cell_6t
Xbit_r43_c248 bl_248 br_248 wl_43 vdd gnd cell_6t
Xbit_r44_c248 bl_248 br_248 wl_44 vdd gnd cell_6t
Xbit_r45_c248 bl_248 br_248 wl_45 vdd gnd cell_6t
Xbit_r46_c248 bl_248 br_248 wl_46 vdd gnd cell_6t
Xbit_r47_c248 bl_248 br_248 wl_47 vdd gnd cell_6t
Xbit_r48_c248 bl_248 br_248 wl_48 vdd gnd cell_6t
Xbit_r49_c248 bl_248 br_248 wl_49 vdd gnd cell_6t
Xbit_r50_c248 bl_248 br_248 wl_50 vdd gnd cell_6t
Xbit_r51_c248 bl_248 br_248 wl_51 vdd gnd cell_6t
Xbit_r52_c248 bl_248 br_248 wl_52 vdd gnd cell_6t
Xbit_r53_c248 bl_248 br_248 wl_53 vdd gnd cell_6t
Xbit_r54_c248 bl_248 br_248 wl_54 vdd gnd cell_6t
Xbit_r55_c248 bl_248 br_248 wl_55 vdd gnd cell_6t
Xbit_r56_c248 bl_248 br_248 wl_56 vdd gnd cell_6t
Xbit_r57_c248 bl_248 br_248 wl_57 vdd gnd cell_6t
Xbit_r58_c248 bl_248 br_248 wl_58 vdd gnd cell_6t
Xbit_r59_c248 bl_248 br_248 wl_59 vdd gnd cell_6t
Xbit_r60_c248 bl_248 br_248 wl_60 vdd gnd cell_6t
Xbit_r61_c248 bl_248 br_248 wl_61 vdd gnd cell_6t
Xbit_r62_c248 bl_248 br_248 wl_62 vdd gnd cell_6t
Xbit_r63_c248 bl_248 br_248 wl_63 vdd gnd cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd cell_6t
Xbit_r1_c249 bl_249 br_249 wl_1 vdd gnd cell_6t
Xbit_r2_c249 bl_249 br_249 wl_2 vdd gnd cell_6t
Xbit_r3_c249 bl_249 br_249 wl_3 vdd gnd cell_6t
Xbit_r4_c249 bl_249 br_249 wl_4 vdd gnd cell_6t
Xbit_r5_c249 bl_249 br_249 wl_5 vdd gnd cell_6t
Xbit_r6_c249 bl_249 br_249 wl_6 vdd gnd cell_6t
Xbit_r7_c249 bl_249 br_249 wl_7 vdd gnd cell_6t
Xbit_r8_c249 bl_249 br_249 wl_8 vdd gnd cell_6t
Xbit_r9_c249 bl_249 br_249 wl_9 vdd gnd cell_6t
Xbit_r10_c249 bl_249 br_249 wl_10 vdd gnd cell_6t
Xbit_r11_c249 bl_249 br_249 wl_11 vdd gnd cell_6t
Xbit_r12_c249 bl_249 br_249 wl_12 vdd gnd cell_6t
Xbit_r13_c249 bl_249 br_249 wl_13 vdd gnd cell_6t
Xbit_r14_c249 bl_249 br_249 wl_14 vdd gnd cell_6t
Xbit_r15_c249 bl_249 br_249 wl_15 vdd gnd cell_6t
Xbit_r16_c249 bl_249 br_249 wl_16 vdd gnd cell_6t
Xbit_r17_c249 bl_249 br_249 wl_17 vdd gnd cell_6t
Xbit_r18_c249 bl_249 br_249 wl_18 vdd gnd cell_6t
Xbit_r19_c249 bl_249 br_249 wl_19 vdd gnd cell_6t
Xbit_r20_c249 bl_249 br_249 wl_20 vdd gnd cell_6t
Xbit_r21_c249 bl_249 br_249 wl_21 vdd gnd cell_6t
Xbit_r22_c249 bl_249 br_249 wl_22 vdd gnd cell_6t
Xbit_r23_c249 bl_249 br_249 wl_23 vdd gnd cell_6t
Xbit_r24_c249 bl_249 br_249 wl_24 vdd gnd cell_6t
Xbit_r25_c249 bl_249 br_249 wl_25 vdd gnd cell_6t
Xbit_r26_c249 bl_249 br_249 wl_26 vdd gnd cell_6t
Xbit_r27_c249 bl_249 br_249 wl_27 vdd gnd cell_6t
Xbit_r28_c249 bl_249 br_249 wl_28 vdd gnd cell_6t
Xbit_r29_c249 bl_249 br_249 wl_29 vdd gnd cell_6t
Xbit_r30_c249 bl_249 br_249 wl_30 vdd gnd cell_6t
Xbit_r31_c249 bl_249 br_249 wl_31 vdd gnd cell_6t
Xbit_r32_c249 bl_249 br_249 wl_32 vdd gnd cell_6t
Xbit_r33_c249 bl_249 br_249 wl_33 vdd gnd cell_6t
Xbit_r34_c249 bl_249 br_249 wl_34 vdd gnd cell_6t
Xbit_r35_c249 bl_249 br_249 wl_35 vdd gnd cell_6t
Xbit_r36_c249 bl_249 br_249 wl_36 vdd gnd cell_6t
Xbit_r37_c249 bl_249 br_249 wl_37 vdd gnd cell_6t
Xbit_r38_c249 bl_249 br_249 wl_38 vdd gnd cell_6t
Xbit_r39_c249 bl_249 br_249 wl_39 vdd gnd cell_6t
Xbit_r40_c249 bl_249 br_249 wl_40 vdd gnd cell_6t
Xbit_r41_c249 bl_249 br_249 wl_41 vdd gnd cell_6t
Xbit_r42_c249 bl_249 br_249 wl_42 vdd gnd cell_6t
Xbit_r43_c249 bl_249 br_249 wl_43 vdd gnd cell_6t
Xbit_r44_c249 bl_249 br_249 wl_44 vdd gnd cell_6t
Xbit_r45_c249 bl_249 br_249 wl_45 vdd gnd cell_6t
Xbit_r46_c249 bl_249 br_249 wl_46 vdd gnd cell_6t
Xbit_r47_c249 bl_249 br_249 wl_47 vdd gnd cell_6t
Xbit_r48_c249 bl_249 br_249 wl_48 vdd gnd cell_6t
Xbit_r49_c249 bl_249 br_249 wl_49 vdd gnd cell_6t
Xbit_r50_c249 bl_249 br_249 wl_50 vdd gnd cell_6t
Xbit_r51_c249 bl_249 br_249 wl_51 vdd gnd cell_6t
Xbit_r52_c249 bl_249 br_249 wl_52 vdd gnd cell_6t
Xbit_r53_c249 bl_249 br_249 wl_53 vdd gnd cell_6t
Xbit_r54_c249 bl_249 br_249 wl_54 vdd gnd cell_6t
Xbit_r55_c249 bl_249 br_249 wl_55 vdd gnd cell_6t
Xbit_r56_c249 bl_249 br_249 wl_56 vdd gnd cell_6t
Xbit_r57_c249 bl_249 br_249 wl_57 vdd gnd cell_6t
Xbit_r58_c249 bl_249 br_249 wl_58 vdd gnd cell_6t
Xbit_r59_c249 bl_249 br_249 wl_59 vdd gnd cell_6t
Xbit_r60_c249 bl_249 br_249 wl_60 vdd gnd cell_6t
Xbit_r61_c249 bl_249 br_249 wl_61 vdd gnd cell_6t
Xbit_r62_c249 bl_249 br_249 wl_62 vdd gnd cell_6t
Xbit_r63_c249 bl_249 br_249 wl_63 vdd gnd cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd cell_6t
Xbit_r1_c250 bl_250 br_250 wl_1 vdd gnd cell_6t
Xbit_r2_c250 bl_250 br_250 wl_2 vdd gnd cell_6t
Xbit_r3_c250 bl_250 br_250 wl_3 vdd gnd cell_6t
Xbit_r4_c250 bl_250 br_250 wl_4 vdd gnd cell_6t
Xbit_r5_c250 bl_250 br_250 wl_5 vdd gnd cell_6t
Xbit_r6_c250 bl_250 br_250 wl_6 vdd gnd cell_6t
Xbit_r7_c250 bl_250 br_250 wl_7 vdd gnd cell_6t
Xbit_r8_c250 bl_250 br_250 wl_8 vdd gnd cell_6t
Xbit_r9_c250 bl_250 br_250 wl_9 vdd gnd cell_6t
Xbit_r10_c250 bl_250 br_250 wl_10 vdd gnd cell_6t
Xbit_r11_c250 bl_250 br_250 wl_11 vdd gnd cell_6t
Xbit_r12_c250 bl_250 br_250 wl_12 vdd gnd cell_6t
Xbit_r13_c250 bl_250 br_250 wl_13 vdd gnd cell_6t
Xbit_r14_c250 bl_250 br_250 wl_14 vdd gnd cell_6t
Xbit_r15_c250 bl_250 br_250 wl_15 vdd gnd cell_6t
Xbit_r16_c250 bl_250 br_250 wl_16 vdd gnd cell_6t
Xbit_r17_c250 bl_250 br_250 wl_17 vdd gnd cell_6t
Xbit_r18_c250 bl_250 br_250 wl_18 vdd gnd cell_6t
Xbit_r19_c250 bl_250 br_250 wl_19 vdd gnd cell_6t
Xbit_r20_c250 bl_250 br_250 wl_20 vdd gnd cell_6t
Xbit_r21_c250 bl_250 br_250 wl_21 vdd gnd cell_6t
Xbit_r22_c250 bl_250 br_250 wl_22 vdd gnd cell_6t
Xbit_r23_c250 bl_250 br_250 wl_23 vdd gnd cell_6t
Xbit_r24_c250 bl_250 br_250 wl_24 vdd gnd cell_6t
Xbit_r25_c250 bl_250 br_250 wl_25 vdd gnd cell_6t
Xbit_r26_c250 bl_250 br_250 wl_26 vdd gnd cell_6t
Xbit_r27_c250 bl_250 br_250 wl_27 vdd gnd cell_6t
Xbit_r28_c250 bl_250 br_250 wl_28 vdd gnd cell_6t
Xbit_r29_c250 bl_250 br_250 wl_29 vdd gnd cell_6t
Xbit_r30_c250 bl_250 br_250 wl_30 vdd gnd cell_6t
Xbit_r31_c250 bl_250 br_250 wl_31 vdd gnd cell_6t
Xbit_r32_c250 bl_250 br_250 wl_32 vdd gnd cell_6t
Xbit_r33_c250 bl_250 br_250 wl_33 vdd gnd cell_6t
Xbit_r34_c250 bl_250 br_250 wl_34 vdd gnd cell_6t
Xbit_r35_c250 bl_250 br_250 wl_35 vdd gnd cell_6t
Xbit_r36_c250 bl_250 br_250 wl_36 vdd gnd cell_6t
Xbit_r37_c250 bl_250 br_250 wl_37 vdd gnd cell_6t
Xbit_r38_c250 bl_250 br_250 wl_38 vdd gnd cell_6t
Xbit_r39_c250 bl_250 br_250 wl_39 vdd gnd cell_6t
Xbit_r40_c250 bl_250 br_250 wl_40 vdd gnd cell_6t
Xbit_r41_c250 bl_250 br_250 wl_41 vdd gnd cell_6t
Xbit_r42_c250 bl_250 br_250 wl_42 vdd gnd cell_6t
Xbit_r43_c250 bl_250 br_250 wl_43 vdd gnd cell_6t
Xbit_r44_c250 bl_250 br_250 wl_44 vdd gnd cell_6t
Xbit_r45_c250 bl_250 br_250 wl_45 vdd gnd cell_6t
Xbit_r46_c250 bl_250 br_250 wl_46 vdd gnd cell_6t
Xbit_r47_c250 bl_250 br_250 wl_47 vdd gnd cell_6t
Xbit_r48_c250 bl_250 br_250 wl_48 vdd gnd cell_6t
Xbit_r49_c250 bl_250 br_250 wl_49 vdd gnd cell_6t
Xbit_r50_c250 bl_250 br_250 wl_50 vdd gnd cell_6t
Xbit_r51_c250 bl_250 br_250 wl_51 vdd gnd cell_6t
Xbit_r52_c250 bl_250 br_250 wl_52 vdd gnd cell_6t
Xbit_r53_c250 bl_250 br_250 wl_53 vdd gnd cell_6t
Xbit_r54_c250 bl_250 br_250 wl_54 vdd gnd cell_6t
Xbit_r55_c250 bl_250 br_250 wl_55 vdd gnd cell_6t
Xbit_r56_c250 bl_250 br_250 wl_56 vdd gnd cell_6t
Xbit_r57_c250 bl_250 br_250 wl_57 vdd gnd cell_6t
Xbit_r58_c250 bl_250 br_250 wl_58 vdd gnd cell_6t
Xbit_r59_c250 bl_250 br_250 wl_59 vdd gnd cell_6t
Xbit_r60_c250 bl_250 br_250 wl_60 vdd gnd cell_6t
Xbit_r61_c250 bl_250 br_250 wl_61 vdd gnd cell_6t
Xbit_r62_c250 bl_250 br_250 wl_62 vdd gnd cell_6t
Xbit_r63_c250 bl_250 br_250 wl_63 vdd gnd cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd cell_6t
Xbit_r1_c251 bl_251 br_251 wl_1 vdd gnd cell_6t
Xbit_r2_c251 bl_251 br_251 wl_2 vdd gnd cell_6t
Xbit_r3_c251 bl_251 br_251 wl_3 vdd gnd cell_6t
Xbit_r4_c251 bl_251 br_251 wl_4 vdd gnd cell_6t
Xbit_r5_c251 bl_251 br_251 wl_5 vdd gnd cell_6t
Xbit_r6_c251 bl_251 br_251 wl_6 vdd gnd cell_6t
Xbit_r7_c251 bl_251 br_251 wl_7 vdd gnd cell_6t
Xbit_r8_c251 bl_251 br_251 wl_8 vdd gnd cell_6t
Xbit_r9_c251 bl_251 br_251 wl_9 vdd gnd cell_6t
Xbit_r10_c251 bl_251 br_251 wl_10 vdd gnd cell_6t
Xbit_r11_c251 bl_251 br_251 wl_11 vdd gnd cell_6t
Xbit_r12_c251 bl_251 br_251 wl_12 vdd gnd cell_6t
Xbit_r13_c251 bl_251 br_251 wl_13 vdd gnd cell_6t
Xbit_r14_c251 bl_251 br_251 wl_14 vdd gnd cell_6t
Xbit_r15_c251 bl_251 br_251 wl_15 vdd gnd cell_6t
Xbit_r16_c251 bl_251 br_251 wl_16 vdd gnd cell_6t
Xbit_r17_c251 bl_251 br_251 wl_17 vdd gnd cell_6t
Xbit_r18_c251 bl_251 br_251 wl_18 vdd gnd cell_6t
Xbit_r19_c251 bl_251 br_251 wl_19 vdd gnd cell_6t
Xbit_r20_c251 bl_251 br_251 wl_20 vdd gnd cell_6t
Xbit_r21_c251 bl_251 br_251 wl_21 vdd gnd cell_6t
Xbit_r22_c251 bl_251 br_251 wl_22 vdd gnd cell_6t
Xbit_r23_c251 bl_251 br_251 wl_23 vdd gnd cell_6t
Xbit_r24_c251 bl_251 br_251 wl_24 vdd gnd cell_6t
Xbit_r25_c251 bl_251 br_251 wl_25 vdd gnd cell_6t
Xbit_r26_c251 bl_251 br_251 wl_26 vdd gnd cell_6t
Xbit_r27_c251 bl_251 br_251 wl_27 vdd gnd cell_6t
Xbit_r28_c251 bl_251 br_251 wl_28 vdd gnd cell_6t
Xbit_r29_c251 bl_251 br_251 wl_29 vdd gnd cell_6t
Xbit_r30_c251 bl_251 br_251 wl_30 vdd gnd cell_6t
Xbit_r31_c251 bl_251 br_251 wl_31 vdd gnd cell_6t
Xbit_r32_c251 bl_251 br_251 wl_32 vdd gnd cell_6t
Xbit_r33_c251 bl_251 br_251 wl_33 vdd gnd cell_6t
Xbit_r34_c251 bl_251 br_251 wl_34 vdd gnd cell_6t
Xbit_r35_c251 bl_251 br_251 wl_35 vdd gnd cell_6t
Xbit_r36_c251 bl_251 br_251 wl_36 vdd gnd cell_6t
Xbit_r37_c251 bl_251 br_251 wl_37 vdd gnd cell_6t
Xbit_r38_c251 bl_251 br_251 wl_38 vdd gnd cell_6t
Xbit_r39_c251 bl_251 br_251 wl_39 vdd gnd cell_6t
Xbit_r40_c251 bl_251 br_251 wl_40 vdd gnd cell_6t
Xbit_r41_c251 bl_251 br_251 wl_41 vdd gnd cell_6t
Xbit_r42_c251 bl_251 br_251 wl_42 vdd gnd cell_6t
Xbit_r43_c251 bl_251 br_251 wl_43 vdd gnd cell_6t
Xbit_r44_c251 bl_251 br_251 wl_44 vdd gnd cell_6t
Xbit_r45_c251 bl_251 br_251 wl_45 vdd gnd cell_6t
Xbit_r46_c251 bl_251 br_251 wl_46 vdd gnd cell_6t
Xbit_r47_c251 bl_251 br_251 wl_47 vdd gnd cell_6t
Xbit_r48_c251 bl_251 br_251 wl_48 vdd gnd cell_6t
Xbit_r49_c251 bl_251 br_251 wl_49 vdd gnd cell_6t
Xbit_r50_c251 bl_251 br_251 wl_50 vdd gnd cell_6t
Xbit_r51_c251 bl_251 br_251 wl_51 vdd gnd cell_6t
Xbit_r52_c251 bl_251 br_251 wl_52 vdd gnd cell_6t
Xbit_r53_c251 bl_251 br_251 wl_53 vdd gnd cell_6t
Xbit_r54_c251 bl_251 br_251 wl_54 vdd gnd cell_6t
Xbit_r55_c251 bl_251 br_251 wl_55 vdd gnd cell_6t
Xbit_r56_c251 bl_251 br_251 wl_56 vdd gnd cell_6t
Xbit_r57_c251 bl_251 br_251 wl_57 vdd gnd cell_6t
Xbit_r58_c251 bl_251 br_251 wl_58 vdd gnd cell_6t
Xbit_r59_c251 bl_251 br_251 wl_59 vdd gnd cell_6t
Xbit_r60_c251 bl_251 br_251 wl_60 vdd gnd cell_6t
Xbit_r61_c251 bl_251 br_251 wl_61 vdd gnd cell_6t
Xbit_r62_c251 bl_251 br_251 wl_62 vdd gnd cell_6t
Xbit_r63_c251 bl_251 br_251 wl_63 vdd gnd cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd cell_6t
Xbit_r1_c252 bl_252 br_252 wl_1 vdd gnd cell_6t
Xbit_r2_c252 bl_252 br_252 wl_2 vdd gnd cell_6t
Xbit_r3_c252 bl_252 br_252 wl_3 vdd gnd cell_6t
Xbit_r4_c252 bl_252 br_252 wl_4 vdd gnd cell_6t
Xbit_r5_c252 bl_252 br_252 wl_5 vdd gnd cell_6t
Xbit_r6_c252 bl_252 br_252 wl_6 vdd gnd cell_6t
Xbit_r7_c252 bl_252 br_252 wl_7 vdd gnd cell_6t
Xbit_r8_c252 bl_252 br_252 wl_8 vdd gnd cell_6t
Xbit_r9_c252 bl_252 br_252 wl_9 vdd gnd cell_6t
Xbit_r10_c252 bl_252 br_252 wl_10 vdd gnd cell_6t
Xbit_r11_c252 bl_252 br_252 wl_11 vdd gnd cell_6t
Xbit_r12_c252 bl_252 br_252 wl_12 vdd gnd cell_6t
Xbit_r13_c252 bl_252 br_252 wl_13 vdd gnd cell_6t
Xbit_r14_c252 bl_252 br_252 wl_14 vdd gnd cell_6t
Xbit_r15_c252 bl_252 br_252 wl_15 vdd gnd cell_6t
Xbit_r16_c252 bl_252 br_252 wl_16 vdd gnd cell_6t
Xbit_r17_c252 bl_252 br_252 wl_17 vdd gnd cell_6t
Xbit_r18_c252 bl_252 br_252 wl_18 vdd gnd cell_6t
Xbit_r19_c252 bl_252 br_252 wl_19 vdd gnd cell_6t
Xbit_r20_c252 bl_252 br_252 wl_20 vdd gnd cell_6t
Xbit_r21_c252 bl_252 br_252 wl_21 vdd gnd cell_6t
Xbit_r22_c252 bl_252 br_252 wl_22 vdd gnd cell_6t
Xbit_r23_c252 bl_252 br_252 wl_23 vdd gnd cell_6t
Xbit_r24_c252 bl_252 br_252 wl_24 vdd gnd cell_6t
Xbit_r25_c252 bl_252 br_252 wl_25 vdd gnd cell_6t
Xbit_r26_c252 bl_252 br_252 wl_26 vdd gnd cell_6t
Xbit_r27_c252 bl_252 br_252 wl_27 vdd gnd cell_6t
Xbit_r28_c252 bl_252 br_252 wl_28 vdd gnd cell_6t
Xbit_r29_c252 bl_252 br_252 wl_29 vdd gnd cell_6t
Xbit_r30_c252 bl_252 br_252 wl_30 vdd gnd cell_6t
Xbit_r31_c252 bl_252 br_252 wl_31 vdd gnd cell_6t
Xbit_r32_c252 bl_252 br_252 wl_32 vdd gnd cell_6t
Xbit_r33_c252 bl_252 br_252 wl_33 vdd gnd cell_6t
Xbit_r34_c252 bl_252 br_252 wl_34 vdd gnd cell_6t
Xbit_r35_c252 bl_252 br_252 wl_35 vdd gnd cell_6t
Xbit_r36_c252 bl_252 br_252 wl_36 vdd gnd cell_6t
Xbit_r37_c252 bl_252 br_252 wl_37 vdd gnd cell_6t
Xbit_r38_c252 bl_252 br_252 wl_38 vdd gnd cell_6t
Xbit_r39_c252 bl_252 br_252 wl_39 vdd gnd cell_6t
Xbit_r40_c252 bl_252 br_252 wl_40 vdd gnd cell_6t
Xbit_r41_c252 bl_252 br_252 wl_41 vdd gnd cell_6t
Xbit_r42_c252 bl_252 br_252 wl_42 vdd gnd cell_6t
Xbit_r43_c252 bl_252 br_252 wl_43 vdd gnd cell_6t
Xbit_r44_c252 bl_252 br_252 wl_44 vdd gnd cell_6t
Xbit_r45_c252 bl_252 br_252 wl_45 vdd gnd cell_6t
Xbit_r46_c252 bl_252 br_252 wl_46 vdd gnd cell_6t
Xbit_r47_c252 bl_252 br_252 wl_47 vdd gnd cell_6t
Xbit_r48_c252 bl_252 br_252 wl_48 vdd gnd cell_6t
Xbit_r49_c252 bl_252 br_252 wl_49 vdd gnd cell_6t
Xbit_r50_c252 bl_252 br_252 wl_50 vdd gnd cell_6t
Xbit_r51_c252 bl_252 br_252 wl_51 vdd gnd cell_6t
Xbit_r52_c252 bl_252 br_252 wl_52 vdd gnd cell_6t
Xbit_r53_c252 bl_252 br_252 wl_53 vdd gnd cell_6t
Xbit_r54_c252 bl_252 br_252 wl_54 vdd gnd cell_6t
Xbit_r55_c252 bl_252 br_252 wl_55 vdd gnd cell_6t
Xbit_r56_c252 bl_252 br_252 wl_56 vdd gnd cell_6t
Xbit_r57_c252 bl_252 br_252 wl_57 vdd gnd cell_6t
Xbit_r58_c252 bl_252 br_252 wl_58 vdd gnd cell_6t
Xbit_r59_c252 bl_252 br_252 wl_59 vdd gnd cell_6t
Xbit_r60_c252 bl_252 br_252 wl_60 vdd gnd cell_6t
Xbit_r61_c252 bl_252 br_252 wl_61 vdd gnd cell_6t
Xbit_r62_c252 bl_252 br_252 wl_62 vdd gnd cell_6t
Xbit_r63_c252 bl_252 br_252 wl_63 vdd gnd cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd cell_6t
Xbit_r1_c253 bl_253 br_253 wl_1 vdd gnd cell_6t
Xbit_r2_c253 bl_253 br_253 wl_2 vdd gnd cell_6t
Xbit_r3_c253 bl_253 br_253 wl_3 vdd gnd cell_6t
Xbit_r4_c253 bl_253 br_253 wl_4 vdd gnd cell_6t
Xbit_r5_c253 bl_253 br_253 wl_5 vdd gnd cell_6t
Xbit_r6_c253 bl_253 br_253 wl_6 vdd gnd cell_6t
Xbit_r7_c253 bl_253 br_253 wl_7 vdd gnd cell_6t
Xbit_r8_c253 bl_253 br_253 wl_8 vdd gnd cell_6t
Xbit_r9_c253 bl_253 br_253 wl_9 vdd gnd cell_6t
Xbit_r10_c253 bl_253 br_253 wl_10 vdd gnd cell_6t
Xbit_r11_c253 bl_253 br_253 wl_11 vdd gnd cell_6t
Xbit_r12_c253 bl_253 br_253 wl_12 vdd gnd cell_6t
Xbit_r13_c253 bl_253 br_253 wl_13 vdd gnd cell_6t
Xbit_r14_c253 bl_253 br_253 wl_14 vdd gnd cell_6t
Xbit_r15_c253 bl_253 br_253 wl_15 vdd gnd cell_6t
Xbit_r16_c253 bl_253 br_253 wl_16 vdd gnd cell_6t
Xbit_r17_c253 bl_253 br_253 wl_17 vdd gnd cell_6t
Xbit_r18_c253 bl_253 br_253 wl_18 vdd gnd cell_6t
Xbit_r19_c253 bl_253 br_253 wl_19 vdd gnd cell_6t
Xbit_r20_c253 bl_253 br_253 wl_20 vdd gnd cell_6t
Xbit_r21_c253 bl_253 br_253 wl_21 vdd gnd cell_6t
Xbit_r22_c253 bl_253 br_253 wl_22 vdd gnd cell_6t
Xbit_r23_c253 bl_253 br_253 wl_23 vdd gnd cell_6t
Xbit_r24_c253 bl_253 br_253 wl_24 vdd gnd cell_6t
Xbit_r25_c253 bl_253 br_253 wl_25 vdd gnd cell_6t
Xbit_r26_c253 bl_253 br_253 wl_26 vdd gnd cell_6t
Xbit_r27_c253 bl_253 br_253 wl_27 vdd gnd cell_6t
Xbit_r28_c253 bl_253 br_253 wl_28 vdd gnd cell_6t
Xbit_r29_c253 bl_253 br_253 wl_29 vdd gnd cell_6t
Xbit_r30_c253 bl_253 br_253 wl_30 vdd gnd cell_6t
Xbit_r31_c253 bl_253 br_253 wl_31 vdd gnd cell_6t
Xbit_r32_c253 bl_253 br_253 wl_32 vdd gnd cell_6t
Xbit_r33_c253 bl_253 br_253 wl_33 vdd gnd cell_6t
Xbit_r34_c253 bl_253 br_253 wl_34 vdd gnd cell_6t
Xbit_r35_c253 bl_253 br_253 wl_35 vdd gnd cell_6t
Xbit_r36_c253 bl_253 br_253 wl_36 vdd gnd cell_6t
Xbit_r37_c253 bl_253 br_253 wl_37 vdd gnd cell_6t
Xbit_r38_c253 bl_253 br_253 wl_38 vdd gnd cell_6t
Xbit_r39_c253 bl_253 br_253 wl_39 vdd gnd cell_6t
Xbit_r40_c253 bl_253 br_253 wl_40 vdd gnd cell_6t
Xbit_r41_c253 bl_253 br_253 wl_41 vdd gnd cell_6t
Xbit_r42_c253 bl_253 br_253 wl_42 vdd gnd cell_6t
Xbit_r43_c253 bl_253 br_253 wl_43 vdd gnd cell_6t
Xbit_r44_c253 bl_253 br_253 wl_44 vdd gnd cell_6t
Xbit_r45_c253 bl_253 br_253 wl_45 vdd gnd cell_6t
Xbit_r46_c253 bl_253 br_253 wl_46 vdd gnd cell_6t
Xbit_r47_c253 bl_253 br_253 wl_47 vdd gnd cell_6t
Xbit_r48_c253 bl_253 br_253 wl_48 vdd gnd cell_6t
Xbit_r49_c253 bl_253 br_253 wl_49 vdd gnd cell_6t
Xbit_r50_c253 bl_253 br_253 wl_50 vdd gnd cell_6t
Xbit_r51_c253 bl_253 br_253 wl_51 vdd gnd cell_6t
Xbit_r52_c253 bl_253 br_253 wl_52 vdd gnd cell_6t
Xbit_r53_c253 bl_253 br_253 wl_53 vdd gnd cell_6t
Xbit_r54_c253 bl_253 br_253 wl_54 vdd gnd cell_6t
Xbit_r55_c253 bl_253 br_253 wl_55 vdd gnd cell_6t
Xbit_r56_c253 bl_253 br_253 wl_56 vdd gnd cell_6t
Xbit_r57_c253 bl_253 br_253 wl_57 vdd gnd cell_6t
Xbit_r58_c253 bl_253 br_253 wl_58 vdd gnd cell_6t
Xbit_r59_c253 bl_253 br_253 wl_59 vdd gnd cell_6t
Xbit_r60_c253 bl_253 br_253 wl_60 vdd gnd cell_6t
Xbit_r61_c253 bl_253 br_253 wl_61 vdd gnd cell_6t
Xbit_r62_c253 bl_253 br_253 wl_62 vdd gnd cell_6t
Xbit_r63_c253 bl_253 br_253 wl_63 vdd gnd cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd cell_6t
Xbit_r1_c254 bl_254 br_254 wl_1 vdd gnd cell_6t
Xbit_r2_c254 bl_254 br_254 wl_2 vdd gnd cell_6t
Xbit_r3_c254 bl_254 br_254 wl_3 vdd gnd cell_6t
Xbit_r4_c254 bl_254 br_254 wl_4 vdd gnd cell_6t
Xbit_r5_c254 bl_254 br_254 wl_5 vdd gnd cell_6t
Xbit_r6_c254 bl_254 br_254 wl_6 vdd gnd cell_6t
Xbit_r7_c254 bl_254 br_254 wl_7 vdd gnd cell_6t
Xbit_r8_c254 bl_254 br_254 wl_8 vdd gnd cell_6t
Xbit_r9_c254 bl_254 br_254 wl_9 vdd gnd cell_6t
Xbit_r10_c254 bl_254 br_254 wl_10 vdd gnd cell_6t
Xbit_r11_c254 bl_254 br_254 wl_11 vdd gnd cell_6t
Xbit_r12_c254 bl_254 br_254 wl_12 vdd gnd cell_6t
Xbit_r13_c254 bl_254 br_254 wl_13 vdd gnd cell_6t
Xbit_r14_c254 bl_254 br_254 wl_14 vdd gnd cell_6t
Xbit_r15_c254 bl_254 br_254 wl_15 vdd gnd cell_6t
Xbit_r16_c254 bl_254 br_254 wl_16 vdd gnd cell_6t
Xbit_r17_c254 bl_254 br_254 wl_17 vdd gnd cell_6t
Xbit_r18_c254 bl_254 br_254 wl_18 vdd gnd cell_6t
Xbit_r19_c254 bl_254 br_254 wl_19 vdd gnd cell_6t
Xbit_r20_c254 bl_254 br_254 wl_20 vdd gnd cell_6t
Xbit_r21_c254 bl_254 br_254 wl_21 vdd gnd cell_6t
Xbit_r22_c254 bl_254 br_254 wl_22 vdd gnd cell_6t
Xbit_r23_c254 bl_254 br_254 wl_23 vdd gnd cell_6t
Xbit_r24_c254 bl_254 br_254 wl_24 vdd gnd cell_6t
Xbit_r25_c254 bl_254 br_254 wl_25 vdd gnd cell_6t
Xbit_r26_c254 bl_254 br_254 wl_26 vdd gnd cell_6t
Xbit_r27_c254 bl_254 br_254 wl_27 vdd gnd cell_6t
Xbit_r28_c254 bl_254 br_254 wl_28 vdd gnd cell_6t
Xbit_r29_c254 bl_254 br_254 wl_29 vdd gnd cell_6t
Xbit_r30_c254 bl_254 br_254 wl_30 vdd gnd cell_6t
Xbit_r31_c254 bl_254 br_254 wl_31 vdd gnd cell_6t
Xbit_r32_c254 bl_254 br_254 wl_32 vdd gnd cell_6t
Xbit_r33_c254 bl_254 br_254 wl_33 vdd gnd cell_6t
Xbit_r34_c254 bl_254 br_254 wl_34 vdd gnd cell_6t
Xbit_r35_c254 bl_254 br_254 wl_35 vdd gnd cell_6t
Xbit_r36_c254 bl_254 br_254 wl_36 vdd gnd cell_6t
Xbit_r37_c254 bl_254 br_254 wl_37 vdd gnd cell_6t
Xbit_r38_c254 bl_254 br_254 wl_38 vdd gnd cell_6t
Xbit_r39_c254 bl_254 br_254 wl_39 vdd gnd cell_6t
Xbit_r40_c254 bl_254 br_254 wl_40 vdd gnd cell_6t
Xbit_r41_c254 bl_254 br_254 wl_41 vdd gnd cell_6t
Xbit_r42_c254 bl_254 br_254 wl_42 vdd gnd cell_6t
Xbit_r43_c254 bl_254 br_254 wl_43 vdd gnd cell_6t
Xbit_r44_c254 bl_254 br_254 wl_44 vdd gnd cell_6t
Xbit_r45_c254 bl_254 br_254 wl_45 vdd gnd cell_6t
Xbit_r46_c254 bl_254 br_254 wl_46 vdd gnd cell_6t
Xbit_r47_c254 bl_254 br_254 wl_47 vdd gnd cell_6t
Xbit_r48_c254 bl_254 br_254 wl_48 vdd gnd cell_6t
Xbit_r49_c254 bl_254 br_254 wl_49 vdd gnd cell_6t
Xbit_r50_c254 bl_254 br_254 wl_50 vdd gnd cell_6t
Xbit_r51_c254 bl_254 br_254 wl_51 vdd gnd cell_6t
Xbit_r52_c254 bl_254 br_254 wl_52 vdd gnd cell_6t
Xbit_r53_c254 bl_254 br_254 wl_53 vdd gnd cell_6t
Xbit_r54_c254 bl_254 br_254 wl_54 vdd gnd cell_6t
Xbit_r55_c254 bl_254 br_254 wl_55 vdd gnd cell_6t
Xbit_r56_c254 bl_254 br_254 wl_56 vdd gnd cell_6t
Xbit_r57_c254 bl_254 br_254 wl_57 vdd gnd cell_6t
Xbit_r58_c254 bl_254 br_254 wl_58 vdd gnd cell_6t
Xbit_r59_c254 bl_254 br_254 wl_59 vdd gnd cell_6t
Xbit_r60_c254 bl_254 br_254 wl_60 vdd gnd cell_6t
Xbit_r61_c254 bl_254 br_254 wl_61 vdd gnd cell_6t
Xbit_r62_c254 bl_254 br_254 wl_62 vdd gnd cell_6t
Xbit_r63_c254 bl_254 br_254 wl_63 vdd gnd cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd cell_6t
Xbit_r1_c255 bl_255 br_255 wl_1 vdd gnd cell_6t
Xbit_r2_c255 bl_255 br_255 wl_2 vdd gnd cell_6t
Xbit_r3_c255 bl_255 br_255 wl_3 vdd gnd cell_6t
Xbit_r4_c255 bl_255 br_255 wl_4 vdd gnd cell_6t
Xbit_r5_c255 bl_255 br_255 wl_5 vdd gnd cell_6t
Xbit_r6_c255 bl_255 br_255 wl_6 vdd gnd cell_6t
Xbit_r7_c255 bl_255 br_255 wl_7 vdd gnd cell_6t
Xbit_r8_c255 bl_255 br_255 wl_8 vdd gnd cell_6t
Xbit_r9_c255 bl_255 br_255 wl_9 vdd gnd cell_6t
Xbit_r10_c255 bl_255 br_255 wl_10 vdd gnd cell_6t
Xbit_r11_c255 bl_255 br_255 wl_11 vdd gnd cell_6t
Xbit_r12_c255 bl_255 br_255 wl_12 vdd gnd cell_6t
Xbit_r13_c255 bl_255 br_255 wl_13 vdd gnd cell_6t
Xbit_r14_c255 bl_255 br_255 wl_14 vdd gnd cell_6t
Xbit_r15_c255 bl_255 br_255 wl_15 vdd gnd cell_6t
Xbit_r16_c255 bl_255 br_255 wl_16 vdd gnd cell_6t
Xbit_r17_c255 bl_255 br_255 wl_17 vdd gnd cell_6t
Xbit_r18_c255 bl_255 br_255 wl_18 vdd gnd cell_6t
Xbit_r19_c255 bl_255 br_255 wl_19 vdd gnd cell_6t
Xbit_r20_c255 bl_255 br_255 wl_20 vdd gnd cell_6t
Xbit_r21_c255 bl_255 br_255 wl_21 vdd gnd cell_6t
Xbit_r22_c255 bl_255 br_255 wl_22 vdd gnd cell_6t
Xbit_r23_c255 bl_255 br_255 wl_23 vdd gnd cell_6t
Xbit_r24_c255 bl_255 br_255 wl_24 vdd gnd cell_6t
Xbit_r25_c255 bl_255 br_255 wl_25 vdd gnd cell_6t
Xbit_r26_c255 bl_255 br_255 wl_26 vdd gnd cell_6t
Xbit_r27_c255 bl_255 br_255 wl_27 vdd gnd cell_6t
Xbit_r28_c255 bl_255 br_255 wl_28 vdd gnd cell_6t
Xbit_r29_c255 bl_255 br_255 wl_29 vdd gnd cell_6t
Xbit_r30_c255 bl_255 br_255 wl_30 vdd gnd cell_6t
Xbit_r31_c255 bl_255 br_255 wl_31 vdd gnd cell_6t
Xbit_r32_c255 bl_255 br_255 wl_32 vdd gnd cell_6t
Xbit_r33_c255 bl_255 br_255 wl_33 vdd gnd cell_6t
Xbit_r34_c255 bl_255 br_255 wl_34 vdd gnd cell_6t
Xbit_r35_c255 bl_255 br_255 wl_35 vdd gnd cell_6t
Xbit_r36_c255 bl_255 br_255 wl_36 vdd gnd cell_6t
Xbit_r37_c255 bl_255 br_255 wl_37 vdd gnd cell_6t
Xbit_r38_c255 bl_255 br_255 wl_38 vdd gnd cell_6t
Xbit_r39_c255 bl_255 br_255 wl_39 vdd gnd cell_6t
Xbit_r40_c255 bl_255 br_255 wl_40 vdd gnd cell_6t
Xbit_r41_c255 bl_255 br_255 wl_41 vdd gnd cell_6t
Xbit_r42_c255 bl_255 br_255 wl_42 vdd gnd cell_6t
Xbit_r43_c255 bl_255 br_255 wl_43 vdd gnd cell_6t
Xbit_r44_c255 bl_255 br_255 wl_44 vdd gnd cell_6t
Xbit_r45_c255 bl_255 br_255 wl_45 vdd gnd cell_6t
Xbit_r46_c255 bl_255 br_255 wl_46 vdd gnd cell_6t
Xbit_r47_c255 bl_255 br_255 wl_47 vdd gnd cell_6t
Xbit_r48_c255 bl_255 br_255 wl_48 vdd gnd cell_6t
Xbit_r49_c255 bl_255 br_255 wl_49 vdd gnd cell_6t
Xbit_r50_c255 bl_255 br_255 wl_50 vdd gnd cell_6t
Xbit_r51_c255 bl_255 br_255 wl_51 vdd gnd cell_6t
Xbit_r52_c255 bl_255 br_255 wl_52 vdd gnd cell_6t
Xbit_r53_c255 bl_255 br_255 wl_53 vdd gnd cell_6t
Xbit_r54_c255 bl_255 br_255 wl_54 vdd gnd cell_6t
Xbit_r55_c255 bl_255 br_255 wl_55 vdd gnd cell_6t
Xbit_r56_c255 bl_255 br_255 wl_56 vdd gnd cell_6t
Xbit_r57_c255 bl_255 br_255 wl_57 vdd gnd cell_6t
Xbit_r58_c255 bl_255 br_255 wl_58 vdd gnd cell_6t
Xbit_r59_c255 bl_255 br_255 wl_59 vdd gnd cell_6t
Xbit_r60_c255 bl_255 br_255 wl_60 vdd gnd cell_6t
Xbit_r61_c255 bl_255 br_255 wl_61 vdd gnd cell_6t
Xbit_r62_c255 bl_255 br_255 wl_62 vdd gnd cell_6t
Xbit_r63_c255 bl_255 br_255 wl_63 vdd gnd cell_6t
.ENDS bitcell_array_0

.SUBCKT replica_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 vdd Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 vdd Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q vdd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q vdd vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl vdd gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT dummy_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl_noconn wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br_noconn wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT replica_column_0 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 vdd gnd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xrbc_1 bl_0 br_0 wl_1 vdd gnd replica_cell_6t
Xrbc_2 bl_0 br_0 wl_2 vdd gnd replica_cell_6t
Xrbc_3 bl_0 br_0 wl_3 vdd gnd replica_cell_6t
Xrbc_4 bl_0 br_0 wl_4 vdd gnd replica_cell_6t
Xrbc_5 bl_0 br_0 wl_5 vdd gnd replica_cell_6t
Xrbc_6 bl_0 br_0 wl_6 vdd gnd replica_cell_6t
Xrbc_7 bl_0 br_0 wl_7 vdd gnd replica_cell_6t
Xrbc_8 bl_0 br_0 wl_8 vdd gnd replica_cell_6t
Xrbc_9 bl_0 br_0 wl_9 vdd gnd replica_cell_6t
Xrbc_10 bl_0 br_0 wl_10 vdd gnd replica_cell_6t
Xrbc_11 bl_0 br_0 wl_11 vdd gnd replica_cell_6t
Xrbc_12 bl_0 br_0 wl_12 vdd gnd replica_cell_6t
Xrbc_13 bl_0 br_0 wl_13 vdd gnd replica_cell_6t
Xrbc_14 bl_0 br_0 wl_14 vdd gnd replica_cell_6t
Xrbc_15 bl_0 br_0 wl_15 vdd gnd replica_cell_6t
Xrbc_16 bl_0 br_0 wl_16 vdd gnd replica_cell_6t
Xrbc_17 bl_0 br_0 wl_17 vdd gnd replica_cell_6t
Xrbc_18 bl_0 br_0 wl_18 vdd gnd replica_cell_6t
Xrbc_19 bl_0 br_0 wl_19 vdd gnd replica_cell_6t
Xrbc_20 bl_0 br_0 wl_20 vdd gnd replica_cell_6t
Xrbc_21 bl_0 br_0 wl_21 vdd gnd replica_cell_6t
Xrbc_22 bl_0 br_0 wl_22 vdd gnd replica_cell_6t
Xrbc_23 bl_0 br_0 wl_23 vdd gnd replica_cell_6t
Xrbc_24 bl_0 br_0 wl_24 vdd gnd replica_cell_6t
Xrbc_25 bl_0 br_0 wl_25 vdd gnd replica_cell_6t
Xrbc_26 bl_0 br_0 wl_26 vdd gnd replica_cell_6t
Xrbc_27 bl_0 br_0 wl_27 vdd gnd replica_cell_6t
Xrbc_28 bl_0 br_0 wl_28 vdd gnd replica_cell_6t
Xrbc_29 bl_0 br_0 wl_29 vdd gnd replica_cell_6t
Xrbc_30 bl_0 br_0 wl_30 vdd gnd replica_cell_6t
Xrbc_31 bl_0 br_0 wl_31 vdd gnd replica_cell_6t
Xrbc_32 bl_0 br_0 wl_32 vdd gnd replica_cell_6t
Xrbc_33 bl_0 br_0 wl_33 vdd gnd replica_cell_6t
Xrbc_34 bl_0 br_0 wl_34 vdd gnd replica_cell_6t
Xrbc_35 bl_0 br_0 wl_35 vdd gnd replica_cell_6t
Xrbc_36 bl_0 br_0 wl_36 vdd gnd replica_cell_6t
Xrbc_37 bl_0 br_0 wl_37 vdd gnd replica_cell_6t
Xrbc_38 bl_0 br_0 wl_38 vdd gnd replica_cell_6t
Xrbc_39 bl_0 br_0 wl_39 vdd gnd replica_cell_6t
Xrbc_40 bl_0 br_0 wl_40 vdd gnd replica_cell_6t
Xrbc_41 bl_0 br_0 wl_41 vdd gnd replica_cell_6t
Xrbc_42 bl_0 br_0 wl_42 vdd gnd replica_cell_6t
Xrbc_43 bl_0 br_0 wl_43 vdd gnd replica_cell_6t
Xrbc_44 bl_0 br_0 wl_44 vdd gnd replica_cell_6t
Xrbc_45 bl_0 br_0 wl_45 vdd gnd replica_cell_6t
Xrbc_46 bl_0 br_0 wl_46 vdd gnd replica_cell_6t
Xrbc_47 bl_0 br_0 wl_47 vdd gnd replica_cell_6t
Xrbc_48 bl_0 br_0 wl_48 vdd gnd replica_cell_6t
Xrbc_49 bl_0 br_0 wl_49 vdd gnd replica_cell_6t
Xrbc_50 bl_0 br_0 wl_50 vdd gnd replica_cell_6t
Xrbc_51 bl_0 br_0 wl_51 vdd gnd replica_cell_6t
Xrbc_52 bl_0 br_0 wl_52 vdd gnd replica_cell_6t
Xrbc_53 bl_0 br_0 wl_53 vdd gnd replica_cell_6t
Xrbc_54 bl_0 br_0 wl_54 vdd gnd replica_cell_6t
Xrbc_55 bl_0 br_0 wl_55 vdd gnd replica_cell_6t
Xrbc_56 bl_0 br_0 wl_56 vdd gnd replica_cell_6t
Xrbc_57 bl_0 br_0 wl_57 vdd gnd replica_cell_6t
Xrbc_58 bl_0 br_0 wl_58 vdd gnd replica_cell_6t
Xrbc_59 bl_0 br_0 wl_59 vdd gnd replica_cell_6t
Xrbc_60 bl_0 br_0 wl_60 vdd gnd replica_cell_6t
Xrbc_61 bl_0 br_0 wl_61 vdd gnd replica_cell_6t
Xrbc_62 bl_0 br_0 wl_62 vdd gnd replica_cell_6t
Xrbc_63 bl_0 br_0 wl_63 vdd gnd replica_cell_6t
Xrbc_64 bl_0 br_0 wl_64 vdd gnd replica_cell_6t
Xrbc_65 bl_0 br_0 wl_65 vdd gnd replica_cell_6t
Xrbc_66 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
.ENDS replica_column_0

.SUBCKT dummy_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd dummy_cell_6t
.ENDS dummy_array_0

.SUBCKT dummy_array_1 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* POWER : vdd 
* GROUND: gnd 
* rows: 67 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
.ENDS dummy_array_1

.SUBCKT dummy_array_2 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* POWER : vdd 
* GROUND: gnd 
* rows: 67 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
.ENDS dummy_array_2

.SUBCKT replica_bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 rbl_wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: rbl_bl_0 
* OUTPUT: rbl_br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : rbl_wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 64 cols: 256
Xbitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 vdd gnd bitcell_array_0
Xreplica_col_0 rbl_bl_0 rbl_br_0 dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 dummy_wl_top vdd gnd replica_column_0
Xdummy_row_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_wl_0 vdd gnd dummy_array_0
Xdummy_row_bot bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_bot vdd gnd dummy_array_0
Xdummy_row_top bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_top vdd gnd dummy_array_0
Xdummy_col_left dummy_bl_left dummy_br_left dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 dummy_wl_top vdd gnd dummy_array_1
Xdummy_col_right dummy_bl_right dummy_br_right dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 dummy_wl_top vdd gnd dummy_array_2
.ENDS replica_bitcell_array_0

.SUBCKT bank dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 dout0_33 dout0_34 dout0_35 dout0_36 dout0_37 dout0_38 dout0_39 dout0_40 dout0_41 dout0_42 dout0_43 dout0_44 dout0_45 dout0_46 dout0_47 dout0_48 dout0_49 dout0_50 dout0_51 dout0_52 dout0_53 dout0_54 dout0_55 dout0_56 dout0_57 dout0_58 dout0_59 dout0_60 dout0_61 dout0_62 dout0_63 dout0_64 dout0_65 dout0_66 dout0_67 dout0_68 dout0_69 dout0_70 dout0_71 dout0_72 dout0_73 dout0_74 dout0_75 dout0_76 dout0_77 dout0_78 dout0_79 dout0_80 dout0_81 dout0_82 dout0_83 dout0_84 dout0_85 dout0_86 dout0_87 dout0_88 dout0_89 dout0_90 dout0_91 dout0_92 dout0_93 dout0_94 dout0_95 dout0_96 dout0_97 dout0_98 dout0_99 dout0_100 dout0_101 dout0_102 dout0_103 dout0_104 dout0_105 dout0_106 dout0_107 dout0_108 dout0_109 dout0_110 dout0_111 dout0_112 dout0_113 dout0_114 dout0_115 dout0_116 dout0_117 dout0_118 dout0_119 dout0_120 dout0_121 dout0_122 dout0_123 dout0_124 dout0_125 dout0_126 dout0_127 dout0_128 dout0_129 dout0_130 dout0_131 dout0_132 dout0_133 dout0_134 dout0_135 dout0_136 dout0_137 dout0_138 dout0_139 dout0_140 dout0_141 dout0_142 dout0_143 dout0_144 dout0_145 dout0_146 dout0_147 dout0_148 dout0_149 dout0_150 dout0_151 dout0_152 dout0_153 dout0_154 dout0_155 dout0_156 dout0_157 dout0_158 dout0_159 dout0_160 dout0_161 dout0_162 dout0_163 dout0_164 dout0_165 dout0_166 dout0_167 dout0_168 dout0_169 dout0_170 dout0_171 dout0_172 dout0_173 dout0_174 dout0_175 dout0_176 dout0_177 dout0_178 dout0_179 dout0_180 dout0_181 dout0_182 dout0_183 dout0_184 dout0_185 dout0_186 dout0_187 dout0_188 dout0_189 dout0_190 dout0_191 dout0_192 dout0_193 dout0_194 dout0_195 dout0_196 dout0_197 dout0_198 dout0_199 dout0_200 dout0_201 dout0_202 dout0_203 dout0_204 dout0_205 dout0_206 dout0_207 dout0_208 dout0_209 dout0_210 dout0_211 dout0_212 dout0_213 dout0_214 dout0_215 dout0_216 dout0_217 dout0_218 dout0_219 dout0_220 dout0_221 dout0_222 dout0_223 dout0_224 dout0_225 dout0_226 dout0_227 dout0_228 dout0_229 dout0_230 dout0_231 dout0_232 dout0_233 dout0_234 dout0_235 dout0_236 dout0_237 dout0_238 dout0_239 dout0_240 dout0_241 dout0_242 dout0_243 dout0_244 dout0_245 dout0_246 dout0_247 dout0_248 dout0_249 dout0_250 dout0_251 dout0_252 dout0_253 dout0_254 dout0_255 rbl_bl_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 din0_33 din0_34 din0_35 din0_36 din0_37 din0_38 din0_39 din0_40 din0_41 din0_42 din0_43 din0_44 din0_45 din0_46 din0_47 din0_48 din0_49 din0_50 din0_51 din0_52 din0_53 din0_54 din0_55 din0_56 din0_57 din0_58 din0_59 din0_60 din0_61 din0_62 din0_63 din0_64 din0_65 din0_66 din0_67 din0_68 din0_69 din0_70 din0_71 din0_72 din0_73 din0_74 din0_75 din0_76 din0_77 din0_78 din0_79 din0_80 din0_81 din0_82 din0_83 din0_84 din0_85 din0_86 din0_87 din0_88 din0_89 din0_90 din0_91 din0_92 din0_93 din0_94 din0_95 din0_96 din0_97 din0_98 din0_99 din0_100 din0_101 din0_102 din0_103 din0_104 din0_105 din0_106 din0_107 din0_108 din0_109 din0_110 din0_111 din0_112 din0_113 din0_114 din0_115 din0_116 din0_117 din0_118 din0_119 din0_120 din0_121 din0_122 din0_123 din0_124 din0_125 din0_126 din0_127 din0_128 din0_129 din0_130 din0_131 din0_132 din0_133 din0_134 din0_135 din0_136 din0_137 din0_138 din0_139 din0_140 din0_141 din0_142 din0_143 din0_144 din0_145 din0_146 din0_147 din0_148 din0_149 din0_150 din0_151 din0_152 din0_153 din0_154 din0_155 din0_156 din0_157 din0_158 din0_159 din0_160 din0_161 din0_162 din0_163 din0_164 din0_165 din0_166 din0_167 din0_168 din0_169 din0_170 din0_171 din0_172 din0_173 din0_174 din0_175 din0_176 din0_177 din0_178 din0_179 din0_180 din0_181 din0_182 din0_183 din0_184 din0_185 din0_186 din0_187 din0_188 din0_189 din0_190 din0_191 din0_192 din0_193 din0_194 din0_195 din0_196 din0_197 din0_198 din0_199 din0_200 din0_201 din0_202 din0_203 din0_204 din0_205 din0_206 din0_207 din0_208 din0_209 din0_210 din0_211 din0_212 din0_213 din0_214 din0_215 din0_216 din0_217 din0_218 din0_219 din0_220 din0_221 din0_222 din0_223 din0_224 din0_225 din0_226 din0_227 din0_228 din0_229 din0_230 din0_231 din0_232 din0_233 din0_234 din0_235 din0_236 din0_237 din0_238 din0_239 din0_240 din0_241 din0_242 din0_243 din0_244 din0_245 din0_246 din0_247 din0_248 din0_249 din0_250 din0_251 din0_252 din0_253 din0_254 din0_255 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout0_32 
* OUTPUT: dout0_33 
* OUTPUT: dout0_34 
* OUTPUT: dout0_35 
* OUTPUT: dout0_36 
* OUTPUT: dout0_37 
* OUTPUT: dout0_38 
* OUTPUT: dout0_39 
* OUTPUT: dout0_40 
* OUTPUT: dout0_41 
* OUTPUT: dout0_42 
* OUTPUT: dout0_43 
* OUTPUT: dout0_44 
* OUTPUT: dout0_45 
* OUTPUT: dout0_46 
* OUTPUT: dout0_47 
* OUTPUT: dout0_48 
* OUTPUT: dout0_49 
* OUTPUT: dout0_50 
* OUTPUT: dout0_51 
* OUTPUT: dout0_52 
* OUTPUT: dout0_53 
* OUTPUT: dout0_54 
* OUTPUT: dout0_55 
* OUTPUT: dout0_56 
* OUTPUT: dout0_57 
* OUTPUT: dout0_58 
* OUTPUT: dout0_59 
* OUTPUT: dout0_60 
* OUTPUT: dout0_61 
* OUTPUT: dout0_62 
* OUTPUT: dout0_63 
* OUTPUT: dout0_64 
* OUTPUT: dout0_65 
* OUTPUT: dout0_66 
* OUTPUT: dout0_67 
* OUTPUT: dout0_68 
* OUTPUT: dout0_69 
* OUTPUT: dout0_70 
* OUTPUT: dout0_71 
* OUTPUT: dout0_72 
* OUTPUT: dout0_73 
* OUTPUT: dout0_74 
* OUTPUT: dout0_75 
* OUTPUT: dout0_76 
* OUTPUT: dout0_77 
* OUTPUT: dout0_78 
* OUTPUT: dout0_79 
* OUTPUT: dout0_80 
* OUTPUT: dout0_81 
* OUTPUT: dout0_82 
* OUTPUT: dout0_83 
* OUTPUT: dout0_84 
* OUTPUT: dout0_85 
* OUTPUT: dout0_86 
* OUTPUT: dout0_87 
* OUTPUT: dout0_88 
* OUTPUT: dout0_89 
* OUTPUT: dout0_90 
* OUTPUT: dout0_91 
* OUTPUT: dout0_92 
* OUTPUT: dout0_93 
* OUTPUT: dout0_94 
* OUTPUT: dout0_95 
* OUTPUT: dout0_96 
* OUTPUT: dout0_97 
* OUTPUT: dout0_98 
* OUTPUT: dout0_99 
* OUTPUT: dout0_100 
* OUTPUT: dout0_101 
* OUTPUT: dout0_102 
* OUTPUT: dout0_103 
* OUTPUT: dout0_104 
* OUTPUT: dout0_105 
* OUTPUT: dout0_106 
* OUTPUT: dout0_107 
* OUTPUT: dout0_108 
* OUTPUT: dout0_109 
* OUTPUT: dout0_110 
* OUTPUT: dout0_111 
* OUTPUT: dout0_112 
* OUTPUT: dout0_113 
* OUTPUT: dout0_114 
* OUTPUT: dout0_115 
* OUTPUT: dout0_116 
* OUTPUT: dout0_117 
* OUTPUT: dout0_118 
* OUTPUT: dout0_119 
* OUTPUT: dout0_120 
* OUTPUT: dout0_121 
* OUTPUT: dout0_122 
* OUTPUT: dout0_123 
* OUTPUT: dout0_124 
* OUTPUT: dout0_125 
* OUTPUT: dout0_126 
* OUTPUT: dout0_127 
* OUTPUT: dout0_128 
* OUTPUT: dout0_129 
* OUTPUT: dout0_130 
* OUTPUT: dout0_131 
* OUTPUT: dout0_132 
* OUTPUT: dout0_133 
* OUTPUT: dout0_134 
* OUTPUT: dout0_135 
* OUTPUT: dout0_136 
* OUTPUT: dout0_137 
* OUTPUT: dout0_138 
* OUTPUT: dout0_139 
* OUTPUT: dout0_140 
* OUTPUT: dout0_141 
* OUTPUT: dout0_142 
* OUTPUT: dout0_143 
* OUTPUT: dout0_144 
* OUTPUT: dout0_145 
* OUTPUT: dout0_146 
* OUTPUT: dout0_147 
* OUTPUT: dout0_148 
* OUTPUT: dout0_149 
* OUTPUT: dout0_150 
* OUTPUT: dout0_151 
* OUTPUT: dout0_152 
* OUTPUT: dout0_153 
* OUTPUT: dout0_154 
* OUTPUT: dout0_155 
* OUTPUT: dout0_156 
* OUTPUT: dout0_157 
* OUTPUT: dout0_158 
* OUTPUT: dout0_159 
* OUTPUT: dout0_160 
* OUTPUT: dout0_161 
* OUTPUT: dout0_162 
* OUTPUT: dout0_163 
* OUTPUT: dout0_164 
* OUTPUT: dout0_165 
* OUTPUT: dout0_166 
* OUTPUT: dout0_167 
* OUTPUT: dout0_168 
* OUTPUT: dout0_169 
* OUTPUT: dout0_170 
* OUTPUT: dout0_171 
* OUTPUT: dout0_172 
* OUTPUT: dout0_173 
* OUTPUT: dout0_174 
* OUTPUT: dout0_175 
* OUTPUT: dout0_176 
* OUTPUT: dout0_177 
* OUTPUT: dout0_178 
* OUTPUT: dout0_179 
* OUTPUT: dout0_180 
* OUTPUT: dout0_181 
* OUTPUT: dout0_182 
* OUTPUT: dout0_183 
* OUTPUT: dout0_184 
* OUTPUT: dout0_185 
* OUTPUT: dout0_186 
* OUTPUT: dout0_187 
* OUTPUT: dout0_188 
* OUTPUT: dout0_189 
* OUTPUT: dout0_190 
* OUTPUT: dout0_191 
* OUTPUT: dout0_192 
* OUTPUT: dout0_193 
* OUTPUT: dout0_194 
* OUTPUT: dout0_195 
* OUTPUT: dout0_196 
* OUTPUT: dout0_197 
* OUTPUT: dout0_198 
* OUTPUT: dout0_199 
* OUTPUT: dout0_200 
* OUTPUT: dout0_201 
* OUTPUT: dout0_202 
* OUTPUT: dout0_203 
* OUTPUT: dout0_204 
* OUTPUT: dout0_205 
* OUTPUT: dout0_206 
* OUTPUT: dout0_207 
* OUTPUT: dout0_208 
* OUTPUT: dout0_209 
* OUTPUT: dout0_210 
* OUTPUT: dout0_211 
* OUTPUT: dout0_212 
* OUTPUT: dout0_213 
* OUTPUT: dout0_214 
* OUTPUT: dout0_215 
* OUTPUT: dout0_216 
* OUTPUT: dout0_217 
* OUTPUT: dout0_218 
* OUTPUT: dout0_219 
* OUTPUT: dout0_220 
* OUTPUT: dout0_221 
* OUTPUT: dout0_222 
* OUTPUT: dout0_223 
* OUTPUT: dout0_224 
* OUTPUT: dout0_225 
* OUTPUT: dout0_226 
* OUTPUT: dout0_227 
* OUTPUT: dout0_228 
* OUTPUT: dout0_229 
* OUTPUT: dout0_230 
* OUTPUT: dout0_231 
* OUTPUT: dout0_232 
* OUTPUT: dout0_233 
* OUTPUT: dout0_234 
* OUTPUT: dout0_235 
* OUTPUT: dout0_236 
* OUTPUT: dout0_237 
* OUTPUT: dout0_238 
* OUTPUT: dout0_239 
* OUTPUT: dout0_240 
* OUTPUT: dout0_241 
* OUTPUT: dout0_242 
* OUTPUT: dout0_243 
* OUTPUT: dout0_244 
* OUTPUT: dout0_245 
* OUTPUT: dout0_246 
* OUTPUT: dout0_247 
* OUTPUT: dout0_248 
* OUTPUT: dout0_249 
* OUTPUT: dout0_250 
* OUTPUT: dout0_251 
* OUTPUT: dout0_252 
* OUTPUT: dout0_253 
* OUTPUT: dout0_254 
* OUTPUT: dout0_255 
* OUTPUT: rbl_bl_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : din0_32 
* INPUT : din0_33 
* INPUT : din0_34 
* INPUT : din0_35 
* INPUT : din0_36 
* INPUT : din0_37 
* INPUT : din0_38 
* INPUT : din0_39 
* INPUT : din0_40 
* INPUT : din0_41 
* INPUT : din0_42 
* INPUT : din0_43 
* INPUT : din0_44 
* INPUT : din0_45 
* INPUT : din0_46 
* INPUT : din0_47 
* INPUT : din0_48 
* INPUT : din0_49 
* INPUT : din0_50 
* INPUT : din0_51 
* INPUT : din0_52 
* INPUT : din0_53 
* INPUT : din0_54 
* INPUT : din0_55 
* INPUT : din0_56 
* INPUT : din0_57 
* INPUT : din0_58 
* INPUT : din0_59 
* INPUT : din0_60 
* INPUT : din0_61 
* INPUT : din0_62 
* INPUT : din0_63 
* INPUT : din0_64 
* INPUT : din0_65 
* INPUT : din0_66 
* INPUT : din0_67 
* INPUT : din0_68 
* INPUT : din0_69 
* INPUT : din0_70 
* INPUT : din0_71 
* INPUT : din0_72 
* INPUT : din0_73 
* INPUT : din0_74 
* INPUT : din0_75 
* INPUT : din0_76 
* INPUT : din0_77 
* INPUT : din0_78 
* INPUT : din0_79 
* INPUT : din0_80 
* INPUT : din0_81 
* INPUT : din0_82 
* INPUT : din0_83 
* INPUT : din0_84 
* INPUT : din0_85 
* INPUT : din0_86 
* INPUT : din0_87 
* INPUT : din0_88 
* INPUT : din0_89 
* INPUT : din0_90 
* INPUT : din0_91 
* INPUT : din0_92 
* INPUT : din0_93 
* INPUT : din0_94 
* INPUT : din0_95 
* INPUT : din0_96 
* INPUT : din0_97 
* INPUT : din0_98 
* INPUT : din0_99 
* INPUT : din0_100 
* INPUT : din0_101 
* INPUT : din0_102 
* INPUT : din0_103 
* INPUT : din0_104 
* INPUT : din0_105 
* INPUT : din0_106 
* INPUT : din0_107 
* INPUT : din0_108 
* INPUT : din0_109 
* INPUT : din0_110 
* INPUT : din0_111 
* INPUT : din0_112 
* INPUT : din0_113 
* INPUT : din0_114 
* INPUT : din0_115 
* INPUT : din0_116 
* INPUT : din0_117 
* INPUT : din0_118 
* INPUT : din0_119 
* INPUT : din0_120 
* INPUT : din0_121 
* INPUT : din0_122 
* INPUT : din0_123 
* INPUT : din0_124 
* INPUT : din0_125 
* INPUT : din0_126 
* INPUT : din0_127 
* INPUT : din0_128 
* INPUT : din0_129 
* INPUT : din0_130 
* INPUT : din0_131 
* INPUT : din0_132 
* INPUT : din0_133 
* INPUT : din0_134 
* INPUT : din0_135 
* INPUT : din0_136 
* INPUT : din0_137 
* INPUT : din0_138 
* INPUT : din0_139 
* INPUT : din0_140 
* INPUT : din0_141 
* INPUT : din0_142 
* INPUT : din0_143 
* INPUT : din0_144 
* INPUT : din0_145 
* INPUT : din0_146 
* INPUT : din0_147 
* INPUT : din0_148 
* INPUT : din0_149 
* INPUT : din0_150 
* INPUT : din0_151 
* INPUT : din0_152 
* INPUT : din0_153 
* INPUT : din0_154 
* INPUT : din0_155 
* INPUT : din0_156 
* INPUT : din0_157 
* INPUT : din0_158 
* INPUT : din0_159 
* INPUT : din0_160 
* INPUT : din0_161 
* INPUT : din0_162 
* INPUT : din0_163 
* INPUT : din0_164 
* INPUT : din0_165 
* INPUT : din0_166 
* INPUT : din0_167 
* INPUT : din0_168 
* INPUT : din0_169 
* INPUT : din0_170 
* INPUT : din0_171 
* INPUT : din0_172 
* INPUT : din0_173 
* INPUT : din0_174 
* INPUT : din0_175 
* INPUT : din0_176 
* INPUT : din0_177 
* INPUT : din0_178 
* INPUT : din0_179 
* INPUT : din0_180 
* INPUT : din0_181 
* INPUT : din0_182 
* INPUT : din0_183 
* INPUT : din0_184 
* INPUT : din0_185 
* INPUT : din0_186 
* INPUT : din0_187 
* INPUT : din0_188 
* INPUT : din0_189 
* INPUT : din0_190 
* INPUT : din0_191 
* INPUT : din0_192 
* INPUT : din0_193 
* INPUT : din0_194 
* INPUT : din0_195 
* INPUT : din0_196 
* INPUT : din0_197 
* INPUT : din0_198 
* INPUT : din0_199 
* INPUT : din0_200 
* INPUT : din0_201 
* INPUT : din0_202 
* INPUT : din0_203 
* INPUT : din0_204 
* INPUT : din0_205 
* INPUT : din0_206 
* INPUT : din0_207 
* INPUT : din0_208 
* INPUT : din0_209 
* INPUT : din0_210 
* INPUT : din0_211 
* INPUT : din0_212 
* INPUT : din0_213 
* INPUT : din0_214 
* INPUT : din0_215 
* INPUT : din0_216 
* INPUT : din0_217 
* INPUT : din0_218 
* INPUT : din0_219 
* INPUT : din0_220 
* INPUT : din0_221 
* INPUT : din0_222 
* INPUT : din0_223 
* INPUT : din0_224 
* INPUT : din0_225 
* INPUT : din0_226 
* INPUT : din0_227 
* INPUT : din0_228 
* INPUT : din0_229 
* INPUT : din0_230 
* INPUT : din0_231 
* INPUT : din0_232 
* INPUT : din0_233 
* INPUT : din0_234 
* INPUT : din0_235 
* INPUT : din0_236 
* INPUT : din0_237 
* INPUT : din0_238 
* INPUT : din0_239 
* INPUT : din0_240 
* INPUT : din0_241 
* INPUT : din0_242 
* INPUT : din0_243 
* INPUT : din0_244 
* INPUT : din0_245 
* INPUT : din0_246 
* INPUT : din0_247 
* INPUT : din0_248 
* INPUT : din0_249 
* INPUT : din0_250 
* INPUT : din0_251 
* INPUT : din0_252 
* INPUT : din0_253 
* INPUT : din0_254 
* INPUT : din0_255 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xreplica_bitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_en0 vdd gnd replica_bitcell_array_0
Xport_data0 rbl_bl_0 rbl_br_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 dout0_33 dout0_34 dout0_35 dout0_36 dout0_37 dout0_38 dout0_39 dout0_40 dout0_41 dout0_42 dout0_43 dout0_44 dout0_45 dout0_46 dout0_47 dout0_48 dout0_49 dout0_50 dout0_51 dout0_52 dout0_53 dout0_54 dout0_55 dout0_56 dout0_57 dout0_58 dout0_59 dout0_60 dout0_61 dout0_62 dout0_63 dout0_64 dout0_65 dout0_66 dout0_67 dout0_68 dout0_69 dout0_70 dout0_71 dout0_72 dout0_73 dout0_74 dout0_75 dout0_76 dout0_77 dout0_78 dout0_79 dout0_80 dout0_81 dout0_82 dout0_83 dout0_84 dout0_85 dout0_86 dout0_87 dout0_88 dout0_89 dout0_90 dout0_91 dout0_92 dout0_93 dout0_94 dout0_95 dout0_96 dout0_97 dout0_98 dout0_99 dout0_100 dout0_101 dout0_102 dout0_103 dout0_104 dout0_105 dout0_106 dout0_107 dout0_108 dout0_109 dout0_110 dout0_111 dout0_112 dout0_113 dout0_114 dout0_115 dout0_116 dout0_117 dout0_118 dout0_119 dout0_120 dout0_121 dout0_122 dout0_123 dout0_124 dout0_125 dout0_126 dout0_127 dout0_128 dout0_129 dout0_130 dout0_131 dout0_132 dout0_133 dout0_134 dout0_135 dout0_136 dout0_137 dout0_138 dout0_139 dout0_140 dout0_141 dout0_142 dout0_143 dout0_144 dout0_145 dout0_146 dout0_147 dout0_148 dout0_149 dout0_150 dout0_151 dout0_152 dout0_153 dout0_154 dout0_155 dout0_156 dout0_157 dout0_158 dout0_159 dout0_160 dout0_161 dout0_162 dout0_163 dout0_164 dout0_165 dout0_166 dout0_167 dout0_168 dout0_169 dout0_170 dout0_171 dout0_172 dout0_173 dout0_174 dout0_175 dout0_176 dout0_177 dout0_178 dout0_179 dout0_180 dout0_181 dout0_182 dout0_183 dout0_184 dout0_185 dout0_186 dout0_187 dout0_188 dout0_189 dout0_190 dout0_191 dout0_192 dout0_193 dout0_194 dout0_195 dout0_196 dout0_197 dout0_198 dout0_199 dout0_200 dout0_201 dout0_202 dout0_203 dout0_204 dout0_205 dout0_206 dout0_207 dout0_208 dout0_209 dout0_210 dout0_211 dout0_212 dout0_213 dout0_214 dout0_215 dout0_216 dout0_217 dout0_218 dout0_219 dout0_220 dout0_221 dout0_222 dout0_223 dout0_224 dout0_225 dout0_226 dout0_227 dout0_228 dout0_229 dout0_230 dout0_231 dout0_232 dout0_233 dout0_234 dout0_235 dout0_236 dout0_237 dout0_238 dout0_239 dout0_240 dout0_241 dout0_242 dout0_243 dout0_244 dout0_245 dout0_246 dout0_247 dout0_248 dout0_249 dout0_250 dout0_251 dout0_252 dout0_253 dout0_254 dout0_255 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 din0_33 din0_34 din0_35 din0_36 din0_37 din0_38 din0_39 din0_40 din0_41 din0_42 din0_43 din0_44 din0_45 din0_46 din0_47 din0_48 din0_49 din0_50 din0_51 din0_52 din0_53 din0_54 din0_55 din0_56 din0_57 din0_58 din0_59 din0_60 din0_61 din0_62 din0_63 din0_64 din0_65 din0_66 din0_67 din0_68 din0_69 din0_70 din0_71 din0_72 din0_73 din0_74 din0_75 din0_76 din0_77 din0_78 din0_79 din0_80 din0_81 din0_82 din0_83 din0_84 din0_85 din0_86 din0_87 din0_88 din0_89 din0_90 din0_91 din0_92 din0_93 din0_94 din0_95 din0_96 din0_97 din0_98 din0_99 din0_100 din0_101 din0_102 din0_103 din0_104 din0_105 din0_106 din0_107 din0_108 din0_109 din0_110 din0_111 din0_112 din0_113 din0_114 din0_115 din0_116 din0_117 din0_118 din0_119 din0_120 din0_121 din0_122 din0_123 din0_124 din0_125 din0_126 din0_127 din0_128 din0_129 din0_130 din0_131 din0_132 din0_133 din0_134 din0_135 din0_136 din0_137 din0_138 din0_139 din0_140 din0_141 din0_142 din0_143 din0_144 din0_145 din0_146 din0_147 din0_148 din0_149 din0_150 din0_151 din0_152 din0_153 din0_154 din0_155 din0_156 din0_157 din0_158 din0_159 din0_160 din0_161 din0_162 din0_163 din0_164 din0_165 din0_166 din0_167 din0_168 din0_169 din0_170 din0_171 din0_172 din0_173 din0_174 din0_175 din0_176 din0_177 din0_178 din0_179 din0_180 din0_181 din0_182 din0_183 din0_184 din0_185 din0_186 din0_187 din0_188 din0_189 din0_190 din0_191 din0_192 din0_193 din0_194 din0_195 din0_196 din0_197 din0_198 din0_199 din0_200 din0_201 din0_202 din0_203 din0_204 din0_205 din0_206 din0_207 din0_208 din0_209 din0_210 din0_211 din0_212 din0_213 din0_214 din0_215 din0_216 din0_217 din0_218 din0_219 din0_220 din0_221 din0_222 din0_223 din0_224 din0_225 din0_226 din0_227 din0_228 din0_229 din0_230 din0_231 din0_232 din0_233 din0_234 din0_235 din0_236 din0_237 din0_238 din0_239 din0_240 din0_241 din0_242 din0_243 din0_244 din0_245 din0_246 din0_247 din0_248 din0_249 din0_250 din0_251 din0_252 din0_253 din0_254 din0_255 s_en0 p_en_bar0 w_en0 vdd gnd port_data_0
Xport_address0 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 wl_en0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 vdd gnd port_address_0
.ENDS bank

* ptx M{0} {1} pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_6 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_6

* ptx M{0} {1} nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* ptx M{0} {1} pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_7 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_7

.SUBCKT dff_buf_0 D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff D qint clk vdd gnd dff
Xdff_buf_inv1 qint Qb vdd gnd pinv_6
Xdff_buf_inv2 Qb Q vdd gnd pinv_7
.ENDS dff_buf_0

.SUBCKT dff_buf_array_0 din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
Xdff_r1_c0 din_1 dout_1 dout_bar_1 clk vdd gnd dff_buf_0
.ENDS dff_buf_array_0

.SUBCKT pnand2_1 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_1

.SUBCKT pinv_8 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_8

.SUBCKT pdriver_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 4]
Xbuf_inv1 A Zb1_int vdd gnd pinv_8
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_8
Xbuf_inv3 Zb2_int Z vdd gnd pinv_7
.ENDS pdriver_1

.SUBCKT pand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_1
Xpand2_inv zb_int Z vdd gnd pdriver_1
.ENDS pand2_0

* ptx M{0} {1} nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p

.SUBCKT pinv_9 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p
.ENDS pinv_9

* ptx M{0} {1} nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT pinv_10 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_10

.SUBCKT pbuf_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_9
Xbuf_inv2 zb_int Z vdd gnd pinv_10
.ENDS pbuf_0

* ptx M{0} {1} nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p

.SUBCKT pinv_11 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p
.ENDS pinv_11

* ptx M{0} {1} nmos_vtg m=6 w=0.24u l=0.05u pd=0.58u ps=0.58u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=6 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT pinv_12 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=6 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mpinv_nmos Z A gnd gnd nmos_vtg m=6 w=0.24u l=0.05u pd=0.58u ps=0.58u as=0.03p ad=0.03p
.ENDS pinv_12

* ptx M{0} {1} nmos_vtg m=16 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=16 w=0.8275u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p

.SUBCKT pinv_13 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=16 w=0.8275u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=16 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p
.ENDS pinv_13

* ptx M{0} {1} nmos_vtg m=47 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=47 w=0.845u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p

.SUBCKT pinv_14 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=47 w=0.845u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=47 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_14

* ptx M{0} {1} nmos_vtg m=140 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=140 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT pinv_15 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=140 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=140 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_15

.SUBCKT pdriver_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 1, 1, 1, 2, 5, 16, 49, 147, 442]
Xbuf_inv1 A Zb1_int vdd gnd pinv_8
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_8
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_8
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_8
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_8
Xbuf_inv6 Zb5_int Zb6_int vdd gnd pinv_8
Xbuf_inv7 Zb6_int Zb7_int vdd gnd pinv_6
Xbuf_inv8 Zb7_int Zb8_int vdd gnd pinv_11
Xbuf_inv9 Zb8_int Zb9_int vdd gnd pinv_12
Xbuf_inv10 Zb9_int Zb10_int vdd gnd pinv_13
Xbuf_inv11 Zb10_int Zb11_int vdd gnd pinv_14
Xbuf_inv12 Zb11_int Z vdd gnd pinv_15
.ENDS pdriver_2

* ptx M{0} {1} nmos_vtg m=3 w=0.21u l=0.05u pd=0.52u ps=0.52u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=3 w=0.63u l=0.05u pd=1.36u ps=1.36u as=0.08p ad=0.08p

.SUBCKT pinv_16 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.63u l=0.05u pd=1.36u ps=1.36u as=0.08p ad=0.08p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.21u l=0.05u pd=0.52u ps=0.52u as=0.03p ad=0.03p
.ENDS pinv_16

* ptx M{0} {1} nmos_vtg m=7 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=7 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_17 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=7 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=7 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_17

.SUBCKT pdriver_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 2, 7, 21]
Xbuf_inv1 A Zb1_int vdd gnd pinv_8
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_6
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_16
Xbuf_inv4 Zb3_int Z vdd gnd pinv_17
.ENDS pdriver_3

.SUBCKT pnand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_1

* ptx M{0} {1} nmos_vtg m=84 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=84 w=0.8475u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p

.SUBCKT pinv_18 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=84 w=0.8475u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=84 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_18

.SUBCKT pand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_18
.ENDS pand3_0

.SUBCKT pand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_10
.ENDS pand3_1

* ptx M{0} {1} nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_19 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_19

* ptx M{0} {1} nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_20 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_20

* ptx M{0} {1} nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p

.SUBCKT pinv_21 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS pinv_21

* ptx M{0} {1} nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p

.SUBCKT pinv_22 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_22

.SUBCKT pdriver_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_8
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_8
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_19
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_20
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_21
Xbuf_inv6 Zb5_int Z vdd gnd pinv_22
.ENDS pdriver_4

.SUBCKT pinv_23 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_23

.SUBCKT delay_chain_0 in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0 in dout_1 vdd gnd pinv_23
Xdload_0_0 dout_1 n_0_0 vdd gnd pinv_23
Xdload_0_1 dout_1 n_0_1 vdd gnd pinv_23
Xdload_0_2 dout_1 n_0_2 vdd gnd pinv_23
Xdload_0_3 dout_1 n_0_3 vdd gnd pinv_23
Xdinv1 dout_1 dout_2 vdd gnd pinv_23
Xdload_1_0 dout_2 n_1_0 vdd gnd pinv_23
Xdload_1_1 dout_2 n_1_1 vdd gnd pinv_23
Xdload_1_2 dout_2 n_1_2 vdd gnd pinv_23
Xdload_1_3 dout_2 n_1_3 vdd gnd pinv_23
Xdinv2 dout_2 dout_3 vdd gnd pinv_23
Xdload_2_0 dout_3 n_2_0 vdd gnd pinv_23
Xdload_2_1 dout_3 n_2_1 vdd gnd pinv_23
Xdload_2_2 dout_3 n_2_2 vdd gnd pinv_23
Xdload_2_3 dout_3 n_2_3 vdd gnd pinv_23
Xdinv3 dout_3 dout_4 vdd gnd pinv_23
Xdload_3_0 dout_4 n_3_0 vdd gnd pinv_23
Xdload_3_1 dout_4 n_3_1 vdd gnd pinv_23
Xdload_3_2 dout_4 n_3_2 vdd gnd pinv_23
Xdload_3_3 dout_4 n_3_3 vdd gnd pinv_23
Xdinv4 dout_4 dout_5 vdd gnd pinv_23
Xdload_4_0 dout_5 n_4_0 vdd gnd pinv_23
Xdload_4_1 dout_5 n_4_1 vdd gnd pinv_23
Xdload_4_2 dout_5 n_4_2 vdd gnd pinv_23
Xdload_4_3 dout_5 n_4_3 vdd gnd pinv_23
Xdinv5 dout_5 dout_6 vdd gnd pinv_23
Xdload_5_0 dout_6 n_5_0 vdd gnd pinv_23
Xdload_5_1 dout_6 n_5_1 vdd gnd pinv_23
Xdload_5_2 dout_6 n_5_2 vdd gnd pinv_23
Xdload_5_3 dout_6 n_5_3 vdd gnd pinv_23
Xdinv6 dout_6 dout_7 vdd gnd pinv_23
Xdload_6_0 dout_7 n_6_0 vdd gnd pinv_23
Xdload_6_1 dout_7 n_6_1 vdd gnd pinv_23
Xdload_6_2 dout_7 n_6_2 vdd gnd pinv_23
Xdload_6_3 dout_7 n_6_3 vdd gnd pinv_23
Xdinv7 dout_7 dout_8 vdd gnd pinv_23
Xdload_7_0 dout_8 n_7_0 vdd gnd pinv_23
Xdload_7_1 dout_8 n_7_1 vdd gnd pinv_23
Xdload_7_2 dout_8 n_7_2 vdd gnd pinv_23
Xdload_7_3 dout_8 n_7_3 vdd gnd pinv_23
Xdinv8 dout_8 out vdd gnd pinv_23
Xdload_8_0 out n_8_0 vdd gnd pinv_23
Xdload_8_1 out n_8_1 vdd gnd pinv_23
Xdload_8_2 out n_8_2 vdd gnd pinv_23
Xdload_8_3 out n_8_3 vdd gnd pinv_23
.ENDS delay_chain_0

.SUBCKT control_logic_rw csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 256
Xctrl_dffs csb web cs_bar cs we_bar we clk_buf vdd gnd dff_buf_array_0
Xclkbuf clk clk_buf vdd gnd pdriver_2
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_8
Xand2_gated_clk_bar cs clk_bar gated_clk_bar vdd gnd pand2_0
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_0
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_3
Xrbl_bl_delay_inv rbl_bl_delay rbl_bl_delay_bar vdd gnd pinv_8
Xw_en_and we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd pand3_0
Xbuf_s_en_and rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd pand3_1
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain_0
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_4
.ENDS control_logic_rw

.SUBCKT sram_64_256 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36] din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43] din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50] din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57] din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64] din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71] din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78] din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85] din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92] din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99] din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106] din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113] din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120] din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127] din0[128] din0[129] din0[130] din0[131] din0[132] din0[133] din0[134] din0[135] din0[136] din0[137] din0[138] din0[139] din0[140] din0[141] din0[142] din0[143] din0[144] din0[145] din0[146] din0[147] din0[148] din0[149] din0[150] din0[151] din0[152] din0[153] din0[154] din0[155] din0[156] din0[157] din0[158] din0[159] din0[160] din0[161] din0[162] din0[163] din0[164] din0[165] din0[166] din0[167] din0[168] din0[169] din0[170] din0[171] din0[172] din0[173] din0[174] din0[175] din0[176] din0[177] din0[178] din0[179] din0[180] din0[181] din0[182] din0[183] din0[184] din0[185] din0[186] din0[187] din0[188] din0[189] din0[190] din0[191] din0[192] din0[193] din0[194] din0[195] din0[196] din0[197] din0[198] din0[199] din0[200] din0[201] din0[202] din0[203] din0[204] din0[205] din0[206] din0[207] din0[208] din0[209] din0[210] din0[211] din0[212] din0[213] din0[214] din0[215] din0[216] din0[217] din0[218] din0[219] din0[220] din0[221] din0[222] din0[223] din0[224] din0[225] din0[226] din0[227] din0[228] din0[229] din0[230] din0[231] din0[232] din0[233] din0[234] din0[235] din0[236] din0[237] din0[238] din0[239] din0[240] din0[241] din0[242] din0[243] din0[244] din0[245] din0[246] din0[247] din0[248] din0[249] din0[250] din0[251] din0[252] din0[253] din0[254] din0[255] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] csb0 web0 clk0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35] dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41] dout0[42] dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62] dout0[63] dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69] dout0[70] dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76] dout0[77] dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83] dout0[84] dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90] dout0[91] dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97] dout0[98] dout0[99] dout0[100] dout0[101] dout0[102] dout0[103] dout0[104] dout0[105] dout0[106] dout0[107] dout0[108] dout0[109] dout0[110] dout0[111] dout0[112] dout0[113] dout0[114] dout0[115] dout0[116] dout0[117] dout0[118] dout0[119] dout0[120] dout0[121] dout0[122] dout0[123] dout0[124] dout0[125] dout0[126] dout0[127] dout0[128] dout0[129] dout0[130] dout0[131] dout0[132] dout0[133] dout0[134] dout0[135] dout0[136] dout0[137] dout0[138] dout0[139] dout0[140] dout0[141] dout0[142] dout0[143] dout0[144] dout0[145] dout0[146] dout0[147] dout0[148] dout0[149] dout0[150] dout0[151] dout0[152] dout0[153] dout0[154] dout0[155] dout0[156] dout0[157] dout0[158] dout0[159] dout0[160] dout0[161] dout0[162] dout0[163] dout0[164] dout0[165] dout0[166] dout0[167] dout0[168] dout0[169] dout0[170] dout0[171] dout0[172] dout0[173] dout0[174] dout0[175] dout0[176] dout0[177] dout0[178] dout0[179] dout0[180] dout0[181] dout0[182] dout0[183] dout0[184] dout0[185] dout0[186] dout0[187] dout0[188] dout0[189] dout0[190] dout0[191] dout0[192] dout0[193] dout0[194] dout0[195] dout0[196] dout0[197] dout0[198] dout0[199] dout0[200] dout0[201] dout0[202] dout0[203] dout0[204] dout0[205] dout0[206] dout0[207] dout0[208] dout0[209] dout0[210] dout0[211] dout0[212] dout0[213] dout0[214] dout0[215] dout0[216] dout0[217] dout0[218] dout0[219] dout0[220] dout0[221] dout0[222] dout0[223] dout0[224] dout0[225] dout0[226] dout0[227] dout0[228] dout0[229] dout0[230] dout0[231] dout0[232] dout0[233] dout0[234] dout0[235] dout0[236] dout0[237] dout0[238] dout0[239] dout0[240] dout0[241] dout0[242] dout0[243] dout0[244] dout0[245] dout0[246] dout0[247] dout0[248] dout0[249] dout0[250] dout0[251] dout0[252] dout0[253] dout0[254] dout0[255] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : din0[32] 
* INPUT : din0[33] 
* INPUT : din0[34] 
* INPUT : din0[35] 
* INPUT : din0[36] 
* INPUT : din0[37] 
* INPUT : din0[38] 
* INPUT : din0[39] 
* INPUT : din0[40] 
* INPUT : din0[41] 
* INPUT : din0[42] 
* INPUT : din0[43] 
* INPUT : din0[44] 
* INPUT : din0[45] 
* INPUT : din0[46] 
* INPUT : din0[47] 
* INPUT : din0[48] 
* INPUT : din0[49] 
* INPUT : din0[50] 
* INPUT : din0[51] 
* INPUT : din0[52] 
* INPUT : din0[53] 
* INPUT : din0[54] 
* INPUT : din0[55] 
* INPUT : din0[56] 
* INPUT : din0[57] 
* INPUT : din0[58] 
* INPUT : din0[59] 
* INPUT : din0[60] 
* INPUT : din0[61] 
* INPUT : din0[62] 
* INPUT : din0[63] 
* INPUT : din0[64] 
* INPUT : din0[65] 
* INPUT : din0[66] 
* INPUT : din0[67] 
* INPUT : din0[68] 
* INPUT : din0[69] 
* INPUT : din0[70] 
* INPUT : din0[71] 
* INPUT : din0[72] 
* INPUT : din0[73] 
* INPUT : din0[74] 
* INPUT : din0[75] 
* INPUT : din0[76] 
* INPUT : din0[77] 
* INPUT : din0[78] 
* INPUT : din0[79] 
* INPUT : din0[80] 
* INPUT : din0[81] 
* INPUT : din0[82] 
* INPUT : din0[83] 
* INPUT : din0[84] 
* INPUT : din0[85] 
* INPUT : din0[86] 
* INPUT : din0[87] 
* INPUT : din0[88] 
* INPUT : din0[89] 
* INPUT : din0[90] 
* INPUT : din0[91] 
* INPUT : din0[92] 
* INPUT : din0[93] 
* INPUT : din0[94] 
* INPUT : din0[95] 
* INPUT : din0[96] 
* INPUT : din0[97] 
* INPUT : din0[98] 
* INPUT : din0[99] 
* INPUT : din0[100] 
* INPUT : din0[101] 
* INPUT : din0[102] 
* INPUT : din0[103] 
* INPUT : din0[104] 
* INPUT : din0[105] 
* INPUT : din0[106] 
* INPUT : din0[107] 
* INPUT : din0[108] 
* INPUT : din0[109] 
* INPUT : din0[110] 
* INPUT : din0[111] 
* INPUT : din0[112] 
* INPUT : din0[113] 
* INPUT : din0[114] 
* INPUT : din0[115] 
* INPUT : din0[116] 
* INPUT : din0[117] 
* INPUT : din0[118] 
* INPUT : din0[119] 
* INPUT : din0[120] 
* INPUT : din0[121] 
* INPUT : din0[122] 
* INPUT : din0[123] 
* INPUT : din0[124] 
* INPUT : din0[125] 
* INPUT : din0[126] 
* INPUT : din0[127] 
* INPUT : din0[128] 
* INPUT : din0[129] 
* INPUT : din0[130] 
* INPUT : din0[131] 
* INPUT : din0[132] 
* INPUT : din0[133] 
* INPUT : din0[134] 
* INPUT : din0[135] 
* INPUT : din0[136] 
* INPUT : din0[137] 
* INPUT : din0[138] 
* INPUT : din0[139] 
* INPUT : din0[140] 
* INPUT : din0[141] 
* INPUT : din0[142] 
* INPUT : din0[143] 
* INPUT : din0[144] 
* INPUT : din0[145] 
* INPUT : din0[146] 
* INPUT : din0[147] 
* INPUT : din0[148] 
* INPUT : din0[149] 
* INPUT : din0[150] 
* INPUT : din0[151] 
* INPUT : din0[152] 
* INPUT : din0[153] 
* INPUT : din0[154] 
* INPUT : din0[155] 
* INPUT : din0[156] 
* INPUT : din0[157] 
* INPUT : din0[158] 
* INPUT : din0[159] 
* INPUT : din0[160] 
* INPUT : din0[161] 
* INPUT : din0[162] 
* INPUT : din0[163] 
* INPUT : din0[164] 
* INPUT : din0[165] 
* INPUT : din0[166] 
* INPUT : din0[167] 
* INPUT : din0[168] 
* INPUT : din0[169] 
* INPUT : din0[170] 
* INPUT : din0[171] 
* INPUT : din0[172] 
* INPUT : din0[173] 
* INPUT : din0[174] 
* INPUT : din0[175] 
* INPUT : din0[176] 
* INPUT : din0[177] 
* INPUT : din0[178] 
* INPUT : din0[179] 
* INPUT : din0[180] 
* INPUT : din0[181] 
* INPUT : din0[182] 
* INPUT : din0[183] 
* INPUT : din0[184] 
* INPUT : din0[185] 
* INPUT : din0[186] 
* INPUT : din0[187] 
* INPUT : din0[188] 
* INPUT : din0[189] 
* INPUT : din0[190] 
* INPUT : din0[191] 
* INPUT : din0[192] 
* INPUT : din0[193] 
* INPUT : din0[194] 
* INPUT : din0[195] 
* INPUT : din0[196] 
* INPUT : din0[197] 
* INPUT : din0[198] 
* INPUT : din0[199] 
* INPUT : din0[200] 
* INPUT : din0[201] 
* INPUT : din0[202] 
* INPUT : din0[203] 
* INPUT : din0[204] 
* INPUT : din0[205] 
* INPUT : din0[206] 
* INPUT : din0[207] 
* INPUT : din0[208] 
* INPUT : din0[209] 
* INPUT : din0[210] 
* INPUT : din0[211] 
* INPUT : din0[212] 
* INPUT : din0[213] 
* INPUT : din0[214] 
* INPUT : din0[215] 
* INPUT : din0[216] 
* INPUT : din0[217] 
* INPUT : din0[218] 
* INPUT : din0[219] 
* INPUT : din0[220] 
* INPUT : din0[221] 
* INPUT : din0[222] 
* INPUT : din0[223] 
* INPUT : din0[224] 
* INPUT : din0[225] 
* INPUT : din0[226] 
* INPUT : din0[227] 
* INPUT : din0[228] 
* INPUT : din0[229] 
* INPUT : din0[230] 
* INPUT : din0[231] 
* INPUT : din0[232] 
* INPUT : din0[233] 
* INPUT : din0[234] 
* INPUT : din0[235] 
* INPUT : din0[236] 
* INPUT : din0[237] 
* INPUT : din0[238] 
* INPUT : din0[239] 
* INPUT : din0[240] 
* INPUT : din0[241] 
* INPUT : din0[242] 
* INPUT : din0[243] 
* INPUT : din0[244] 
* INPUT : din0[245] 
* INPUT : din0[246] 
* INPUT : din0[247] 
* INPUT : din0[248] 
* INPUT : din0[249] 
* INPUT : din0[250] 
* INPUT : din0[251] 
* INPUT : din0[252] 
* INPUT : din0[253] 
* INPUT : din0[254] 
* INPUT : din0[255] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout0[32] 
* OUTPUT: dout0[33] 
* OUTPUT: dout0[34] 
* OUTPUT: dout0[35] 
* OUTPUT: dout0[36] 
* OUTPUT: dout0[37] 
* OUTPUT: dout0[38] 
* OUTPUT: dout0[39] 
* OUTPUT: dout0[40] 
* OUTPUT: dout0[41] 
* OUTPUT: dout0[42] 
* OUTPUT: dout0[43] 
* OUTPUT: dout0[44] 
* OUTPUT: dout0[45] 
* OUTPUT: dout0[46] 
* OUTPUT: dout0[47] 
* OUTPUT: dout0[48] 
* OUTPUT: dout0[49] 
* OUTPUT: dout0[50] 
* OUTPUT: dout0[51] 
* OUTPUT: dout0[52] 
* OUTPUT: dout0[53] 
* OUTPUT: dout0[54] 
* OUTPUT: dout0[55] 
* OUTPUT: dout0[56] 
* OUTPUT: dout0[57] 
* OUTPUT: dout0[58] 
* OUTPUT: dout0[59] 
* OUTPUT: dout0[60] 
* OUTPUT: dout0[61] 
* OUTPUT: dout0[62] 
* OUTPUT: dout0[63] 
* OUTPUT: dout0[64] 
* OUTPUT: dout0[65] 
* OUTPUT: dout0[66] 
* OUTPUT: dout0[67] 
* OUTPUT: dout0[68] 
* OUTPUT: dout0[69] 
* OUTPUT: dout0[70] 
* OUTPUT: dout0[71] 
* OUTPUT: dout0[72] 
* OUTPUT: dout0[73] 
* OUTPUT: dout0[74] 
* OUTPUT: dout0[75] 
* OUTPUT: dout0[76] 
* OUTPUT: dout0[77] 
* OUTPUT: dout0[78] 
* OUTPUT: dout0[79] 
* OUTPUT: dout0[80] 
* OUTPUT: dout0[81] 
* OUTPUT: dout0[82] 
* OUTPUT: dout0[83] 
* OUTPUT: dout0[84] 
* OUTPUT: dout0[85] 
* OUTPUT: dout0[86] 
* OUTPUT: dout0[87] 
* OUTPUT: dout0[88] 
* OUTPUT: dout0[89] 
* OUTPUT: dout0[90] 
* OUTPUT: dout0[91] 
* OUTPUT: dout0[92] 
* OUTPUT: dout0[93] 
* OUTPUT: dout0[94] 
* OUTPUT: dout0[95] 
* OUTPUT: dout0[96] 
* OUTPUT: dout0[97] 
* OUTPUT: dout0[98] 
* OUTPUT: dout0[99] 
* OUTPUT: dout0[100] 
* OUTPUT: dout0[101] 
* OUTPUT: dout0[102] 
* OUTPUT: dout0[103] 
* OUTPUT: dout0[104] 
* OUTPUT: dout0[105] 
* OUTPUT: dout0[106] 
* OUTPUT: dout0[107] 
* OUTPUT: dout0[108] 
* OUTPUT: dout0[109] 
* OUTPUT: dout0[110] 
* OUTPUT: dout0[111] 
* OUTPUT: dout0[112] 
* OUTPUT: dout0[113] 
* OUTPUT: dout0[114] 
* OUTPUT: dout0[115] 
* OUTPUT: dout0[116] 
* OUTPUT: dout0[117] 
* OUTPUT: dout0[118] 
* OUTPUT: dout0[119] 
* OUTPUT: dout0[120] 
* OUTPUT: dout0[121] 
* OUTPUT: dout0[122] 
* OUTPUT: dout0[123] 
* OUTPUT: dout0[124] 
* OUTPUT: dout0[125] 
* OUTPUT: dout0[126] 
* OUTPUT: dout0[127] 
* OUTPUT: dout0[128] 
* OUTPUT: dout0[129] 
* OUTPUT: dout0[130] 
* OUTPUT: dout0[131] 
* OUTPUT: dout0[132] 
* OUTPUT: dout0[133] 
* OUTPUT: dout0[134] 
* OUTPUT: dout0[135] 
* OUTPUT: dout0[136] 
* OUTPUT: dout0[137] 
* OUTPUT: dout0[138] 
* OUTPUT: dout0[139] 
* OUTPUT: dout0[140] 
* OUTPUT: dout0[141] 
* OUTPUT: dout0[142] 
* OUTPUT: dout0[143] 
* OUTPUT: dout0[144] 
* OUTPUT: dout0[145] 
* OUTPUT: dout0[146] 
* OUTPUT: dout0[147] 
* OUTPUT: dout0[148] 
* OUTPUT: dout0[149] 
* OUTPUT: dout0[150] 
* OUTPUT: dout0[151] 
* OUTPUT: dout0[152] 
* OUTPUT: dout0[153] 
* OUTPUT: dout0[154] 
* OUTPUT: dout0[155] 
* OUTPUT: dout0[156] 
* OUTPUT: dout0[157] 
* OUTPUT: dout0[158] 
* OUTPUT: dout0[159] 
* OUTPUT: dout0[160] 
* OUTPUT: dout0[161] 
* OUTPUT: dout0[162] 
* OUTPUT: dout0[163] 
* OUTPUT: dout0[164] 
* OUTPUT: dout0[165] 
* OUTPUT: dout0[166] 
* OUTPUT: dout0[167] 
* OUTPUT: dout0[168] 
* OUTPUT: dout0[169] 
* OUTPUT: dout0[170] 
* OUTPUT: dout0[171] 
* OUTPUT: dout0[172] 
* OUTPUT: dout0[173] 
* OUTPUT: dout0[174] 
* OUTPUT: dout0[175] 
* OUTPUT: dout0[176] 
* OUTPUT: dout0[177] 
* OUTPUT: dout0[178] 
* OUTPUT: dout0[179] 
* OUTPUT: dout0[180] 
* OUTPUT: dout0[181] 
* OUTPUT: dout0[182] 
* OUTPUT: dout0[183] 
* OUTPUT: dout0[184] 
* OUTPUT: dout0[185] 
* OUTPUT: dout0[186] 
* OUTPUT: dout0[187] 
* OUTPUT: dout0[188] 
* OUTPUT: dout0[189] 
* OUTPUT: dout0[190] 
* OUTPUT: dout0[191] 
* OUTPUT: dout0[192] 
* OUTPUT: dout0[193] 
* OUTPUT: dout0[194] 
* OUTPUT: dout0[195] 
* OUTPUT: dout0[196] 
* OUTPUT: dout0[197] 
* OUTPUT: dout0[198] 
* OUTPUT: dout0[199] 
* OUTPUT: dout0[200] 
* OUTPUT: dout0[201] 
* OUTPUT: dout0[202] 
* OUTPUT: dout0[203] 
* OUTPUT: dout0[204] 
* OUTPUT: dout0[205] 
* OUTPUT: dout0[206] 
* OUTPUT: dout0[207] 
* OUTPUT: dout0[208] 
* OUTPUT: dout0[209] 
* OUTPUT: dout0[210] 
* OUTPUT: dout0[211] 
* OUTPUT: dout0[212] 
* OUTPUT: dout0[213] 
* OUTPUT: dout0[214] 
* OUTPUT: dout0[215] 
* OUTPUT: dout0[216] 
* OUTPUT: dout0[217] 
* OUTPUT: dout0[218] 
* OUTPUT: dout0[219] 
* OUTPUT: dout0[220] 
* OUTPUT: dout0[221] 
* OUTPUT: dout0[222] 
* OUTPUT: dout0[223] 
* OUTPUT: dout0[224] 
* OUTPUT: dout0[225] 
* OUTPUT: dout0[226] 
* OUTPUT: dout0[227] 
* OUTPUT: dout0[228] 
* OUTPUT: dout0[229] 
* OUTPUT: dout0[230] 
* OUTPUT: dout0[231] 
* OUTPUT: dout0[232] 
* OUTPUT: dout0[233] 
* OUTPUT: dout0[234] 
* OUTPUT: dout0[235] 
* OUTPUT: dout0[236] 
* OUTPUT: dout0[237] 
* OUTPUT: dout0[238] 
* OUTPUT: dout0[239] 
* OUTPUT: dout0[240] 
* OUTPUT: dout0[241] 
* OUTPUT: dout0[242] 
* OUTPUT: dout0[243] 
* OUTPUT: dout0[244] 
* OUTPUT: dout0[245] 
* OUTPUT: dout0[246] 
* OUTPUT: dout0[247] 
* OUTPUT: dout0[248] 
* OUTPUT: dout0[249] 
* OUTPUT: dout0[250] 
* OUTPUT: dout0[251] 
* OUTPUT: dout0[252] 
* OUTPUT: dout0[253] 
* OUTPUT: dout0[254] 
* OUTPUT: dout0[255] 
* POWER : vdd 
* GROUND: gnd 
Xbank0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35] dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41] dout0[42] dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62] dout0[63] dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69] dout0[70] dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76] dout0[77] dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83] dout0[84] dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90] dout0[91] dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97] dout0[98] dout0[99] dout0[100] dout0[101] dout0[102] dout0[103] dout0[104] dout0[105] dout0[106] dout0[107] dout0[108] dout0[109] dout0[110] dout0[111] dout0[112] dout0[113] dout0[114] dout0[115] dout0[116] dout0[117] dout0[118] dout0[119] dout0[120] dout0[121] dout0[122] dout0[123] dout0[124] dout0[125] dout0[126] dout0[127] dout0[128] dout0[129] dout0[130] dout0[131] dout0[132] dout0[133] dout0[134] dout0[135] dout0[136] dout0[137] dout0[138] dout0[139] dout0[140] dout0[141] dout0[142] dout0[143] dout0[144] dout0[145] dout0[146] dout0[147] dout0[148] dout0[149] dout0[150] dout0[151] dout0[152] dout0[153] dout0[154] dout0[155] dout0[156] dout0[157] dout0[158] dout0[159] dout0[160] dout0[161] dout0[162] dout0[163] dout0[164] dout0[165] dout0[166] dout0[167] dout0[168] dout0[169] dout0[170] dout0[171] dout0[172] dout0[173] dout0[174] dout0[175] dout0[176] dout0[177] dout0[178] dout0[179] dout0[180] dout0[181] dout0[182] dout0[183] dout0[184] dout0[185] dout0[186] dout0[187] dout0[188] dout0[189] dout0[190] dout0[191] dout0[192] dout0[193] dout0[194] dout0[195] dout0[196] dout0[197] dout0[198] dout0[199] dout0[200] dout0[201] dout0[202] dout0[203] dout0[204] dout0[205] dout0[206] dout0[207] dout0[208] dout0[209] dout0[210] dout0[211] dout0[212] dout0[213] dout0[214] dout0[215] dout0[216] dout0[217] dout0[218] dout0[219] dout0[220] dout0[221] dout0[222] dout0[223] dout0[224] dout0[225] dout0[226] dout0[227] dout0[228] dout0[229] dout0[230] dout0[231] dout0[232] dout0[233] dout0[234] dout0[235] dout0[236] dout0[237] dout0[238] dout0[239] dout0[240] dout0[241] dout0[242] dout0[243] dout0[244] dout0[245] dout0[246] dout0[247] dout0[248] dout0[249] dout0[250] dout0[251] dout0[252] dout0[253] dout0[254] dout0[255] rbl_bl0 bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] bank_din0[32] bank_din0[33] bank_din0[34] bank_din0[35] bank_din0[36] bank_din0[37] bank_din0[38] bank_din0[39] bank_din0[40] bank_din0[41] bank_din0[42] bank_din0[43] bank_din0[44] bank_din0[45] bank_din0[46] bank_din0[47] bank_din0[48] bank_din0[49] bank_din0[50] bank_din0[51] bank_din0[52] bank_din0[53] bank_din0[54] bank_din0[55] bank_din0[56] bank_din0[57] bank_din0[58] bank_din0[59] bank_din0[60] bank_din0[61] bank_din0[62] bank_din0[63] bank_din0[64] bank_din0[65] bank_din0[66] bank_din0[67] bank_din0[68] bank_din0[69] bank_din0[70] bank_din0[71] bank_din0[72] bank_din0[73] bank_din0[74] bank_din0[75] bank_din0[76] bank_din0[77] bank_din0[78] bank_din0[79] bank_din0[80] bank_din0[81] bank_din0[82] bank_din0[83] bank_din0[84] bank_din0[85] bank_din0[86] bank_din0[87] bank_din0[88] bank_din0[89] bank_din0[90] bank_din0[91] bank_din0[92] bank_din0[93] bank_din0[94] bank_din0[95] bank_din0[96] bank_din0[97] bank_din0[98] bank_din0[99] bank_din0[100] bank_din0[101] bank_din0[102] bank_din0[103] bank_din0[104] bank_din0[105] bank_din0[106] bank_din0[107] bank_din0[108] bank_din0[109] bank_din0[110] bank_din0[111] bank_din0[112] bank_din0[113] bank_din0[114] bank_din0[115] bank_din0[116] bank_din0[117] bank_din0[118] bank_din0[119] bank_din0[120] bank_din0[121] bank_din0[122] bank_din0[123] bank_din0[124] bank_din0[125] bank_din0[126] bank_din0[127] bank_din0[128] bank_din0[129] bank_din0[130] bank_din0[131] bank_din0[132] bank_din0[133] bank_din0[134] bank_din0[135] bank_din0[136] bank_din0[137] bank_din0[138] bank_din0[139] bank_din0[140] bank_din0[141] bank_din0[142] bank_din0[143] bank_din0[144] bank_din0[145] bank_din0[146] bank_din0[147] bank_din0[148] bank_din0[149] bank_din0[150] bank_din0[151] bank_din0[152] bank_din0[153] bank_din0[154] bank_din0[155] bank_din0[156] bank_din0[157] bank_din0[158] bank_din0[159] bank_din0[160] bank_din0[161] bank_din0[162] bank_din0[163] bank_din0[164] bank_din0[165] bank_din0[166] bank_din0[167] bank_din0[168] bank_din0[169] bank_din0[170] bank_din0[171] bank_din0[172] bank_din0[173] bank_din0[174] bank_din0[175] bank_din0[176] bank_din0[177] bank_din0[178] bank_din0[179] bank_din0[180] bank_din0[181] bank_din0[182] bank_din0[183] bank_din0[184] bank_din0[185] bank_din0[186] bank_din0[187] bank_din0[188] bank_din0[189] bank_din0[190] bank_din0[191] bank_din0[192] bank_din0[193] bank_din0[194] bank_din0[195] bank_din0[196] bank_din0[197] bank_din0[198] bank_din0[199] bank_din0[200] bank_din0[201] bank_din0[202] bank_din0[203] bank_din0[204] bank_din0[205] bank_din0[206] bank_din0[207] bank_din0[208] bank_din0[209] bank_din0[210] bank_din0[211] bank_din0[212] bank_din0[213] bank_din0[214] bank_din0[215] bank_din0[216] bank_din0[217] bank_din0[218] bank_din0[219] bank_din0[220] bank_din0[221] bank_din0[222] bank_din0[223] bank_din0[224] bank_din0[225] bank_din0[226] bank_din0[227] bank_din0[228] bank_din0[229] bank_din0[230] bank_din0[231] bank_din0[232] bank_din0[233] bank_din0[234] bank_din0[235] bank_din0[236] bank_din0[237] bank_din0[238] bank_din0[239] bank_din0[240] bank_din0[241] bank_din0[242] bank_din0[243] bank_din0[244] bank_din0[245] bank_din0[246] bank_din0[247] bank_din0[248] bank_din0[249] bank_din0[250] bank_din0[251] bank_din0[252] bank_din0[253] bank_din0[254] bank_din0[255] a0[0] a0[1] a0[2] a0[3] a0[4] a0[5] s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd bank
Xcontrol0 csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd control_logic_rw
Xrow_address0 addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] a0[0] a0[1] a0[2] a0[3] a0[4] a0[5] clk_buf0 vdd gnd row_addr_dff
Xdata_dff0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36] din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43] din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50] din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57] din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64] din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71] din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78] din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85] din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92] din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99] din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106] din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113] din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120] din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127] din0[128] din0[129] din0[130] din0[131] din0[132] din0[133] din0[134] din0[135] din0[136] din0[137] din0[138] din0[139] din0[140] din0[141] din0[142] din0[143] din0[144] din0[145] din0[146] din0[147] din0[148] din0[149] din0[150] din0[151] din0[152] din0[153] din0[154] din0[155] din0[156] din0[157] din0[158] din0[159] din0[160] din0[161] din0[162] din0[163] din0[164] din0[165] din0[166] din0[167] din0[168] din0[169] din0[170] din0[171] din0[172] din0[173] din0[174] din0[175] din0[176] din0[177] din0[178] din0[179] din0[180] din0[181] din0[182] din0[183] din0[184] din0[185] din0[186] din0[187] din0[188] din0[189] din0[190] din0[191] din0[192] din0[193] din0[194] din0[195] din0[196] din0[197] din0[198] din0[199] din0[200] din0[201] din0[202] din0[203] din0[204] din0[205] din0[206] din0[207] din0[208] din0[209] din0[210] din0[211] din0[212] din0[213] din0[214] din0[215] din0[216] din0[217] din0[218] din0[219] din0[220] din0[221] din0[222] din0[223] din0[224] din0[225] din0[226] din0[227] din0[228] din0[229] din0[230] din0[231] din0[232] din0[233] din0[234] din0[235] din0[236] din0[237] din0[238] din0[239] din0[240] din0[241] din0[242] din0[243] din0[244] din0[245] din0[246] din0[247] din0[248] din0[249] din0[250] din0[251] din0[252] din0[253] din0[254] din0[255] bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] bank_din0[32] bank_din0[33] bank_din0[34] bank_din0[35] bank_din0[36] bank_din0[37] bank_din0[38] bank_din0[39] bank_din0[40] bank_din0[41] bank_din0[42] bank_din0[43] bank_din0[44] bank_din0[45] bank_din0[46] bank_din0[47] bank_din0[48] bank_din0[49] bank_din0[50] bank_din0[51] bank_din0[52] bank_din0[53] bank_din0[54] bank_din0[55] bank_din0[56] bank_din0[57] bank_din0[58] bank_din0[59] bank_din0[60] bank_din0[61] bank_din0[62] bank_din0[63] bank_din0[64] bank_din0[65] bank_din0[66] bank_din0[67] bank_din0[68] bank_din0[69] bank_din0[70] bank_din0[71] bank_din0[72] bank_din0[73] bank_din0[74] bank_din0[75] bank_din0[76] bank_din0[77] bank_din0[78] bank_din0[79] bank_din0[80] bank_din0[81] bank_din0[82] bank_din0[83] bank_din0[84] bank_din0[85] bank_din0[86] bank_din0[87] bank_din0[88] bank_din0[89] bank_din0[90] bank_din0[91] bank_din0[92] bank_din0[93] bank_din0[94] bank_din0[95] bank_din0[96] bank_din0[97] bank_din0[98] bank_din0[99] bank_din0[100] bank_din0[101] bank_din0[102] bank_din0[103] bank_din0[104] bank_din0[105] bank_din0[106] bank_din0[107] bank_din0[108] bank_din0[109] bank_din0[110] bank_din0[111] bank_din0[112] bank_din0[113] bank_din0[114] bank_din0[115] bank_din0[116] bank_din0[117] bank_din0[118] bank_din0[119] bank_din0[120] bank_din0[121] bank_din0[122] bank_din0[123] bank_din0[124] bank_din0[125] bank_din0[126] bank_din0[127] bank_din0[128] bank_din0[129] bank_din0[130] bank_din0[131] bank_din0[132] bank_din0[133] bank_din0[134] bank_din0[135] bank_din0[136] bank_din0[137] bank_din0[138] bank_din0[139] bank_din0[140] bank_din0[141] bank_din0[142] bank_din0[143] bank_din0[144] bank_din0[145] bank_din0[146] bank_din0[147] bank_din0[148] bank_din0[149] bank_din0[150] bank_din0[151] bank_din0[152] bank_din0[153] bank_din0[154] bank_din0[155] bank_din0[156] bank_din0[157] bank_din0[158] bank_din0[159] bank_din0[160] bank_din0[161] bank_din0[162] bank_din0[163] bank_din0[164] bank_din0[165] bank_din0[166] bank_din0[167] bank_din0[168] bank_din0[169] bank_din0[170] bank_din0[171] bank_din0[172] bank_din0[173] bank_din0[174] bank_din0[175] bank_din0[176] bank_din0[177] bank_din0[178] bank_din0[179] bank_din0[180] bank_din0[181] bank_din0[182] bank_din0[183] bank_din0[184] bank_din0[185] bank_din0[186] bank_din0[187] bank_din0[188] bank_din0[189] bank_din0[190] bank_din0[191] bank_din0[192] bank_din0[193] bank_din0[194] bank_din0[195] bank_din0[196] bank_din0[197] bank_din0[198] bank_din0[199] bank_din0[200] bank_din0[201] bank_din0[202] bank_din0[203] bank_din0[204] bank_din0[205] bank_din0[206] bank_din0[207] bank_din0[208] bank_din0[209] bank_din0[210] bank_din0[211] bank_din0[212] bank_din0[213] bank_din0[214] bank_din0[215] bank_din0[216] bank_din0[217] bank_din0[218] bank_din0[219] bank_din0[220] bank_din0[221] bank_din0[222] bank_din0[223] bank_din0[224] bank_din0[225] bank_din0[226] bank_din0[227] bank_din0[228] bank_din0[229] bank_din0[230] bank_din0[231] bank_din0[232] bank_din0[233] bank_din0[234] bank_din0[235] bank_din0[236] bank_din0[237] bank_din0[238] bank_din0[239] bank_din0[240] bank_din0[241] bank_din0[242] bank_din0[243] bank_din0[244] bank_din0[245] bank_din0[246] bank_din0[247] bank_din0[248] bank_din0[249] bank_din0[250] bank_din0[251] bank_din0[252] bank_din0[253] bank_din0[254] bank_din0[255] clk_buf0 vdd gnd data_dff
.ENDS sram_64_256
