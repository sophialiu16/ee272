
//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/Fifo_ODTYPE_16__b082e045ab0825c90c856c0668d6e3347c56_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:12 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_16_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_16_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;
  reg [15:0] regs_13_sva_dfm;
  reg [15:0] regs_14_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd97),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd98),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd117),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_14_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_14_sva_dfm <= 16'b0000000000000000;
      regs_13_sva_dfm <= 16'b0000000000000000;
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_14_sva_dfm <= regs_13_sva_dfm;
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_16
// ------------------------------------------------------------------


module Fifo_ODTYPE_16 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_16_run Fifo_ODTYPE_16_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_15__30ad9192d0464f2c737edb11c85d93b679f7_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:20 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_15_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_15_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;
  reg [15:0] regs_13_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd94),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd95),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd118),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_13_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_13_sva_dfm <= 16'b0000000000000000;
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_15
// ------------------------------------------------------------------


module Fifo_ODTYPE_15 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_15_run Fifo_ODTYPE_15_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_14__9ee6c6d92769a02e65b3e79b2bfd82597798_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:27 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_14_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_14_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd91),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd92),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd119),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_12_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_14
// ------------------------------------------------------------------


module Fifo_ODTYPE_14 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_14_run Fifo_ODTYPE_14_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_13__2e906883fcda2ed1d8b8dfd8b0b4a2be7539_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:35 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_13_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_13_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd88),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd89),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd120),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_11_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_13
// ------------------------------------------------------------------


module Fifo_ODTYPE_13 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_13_run Fifo_ODTYPE_13_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_12__9e26134eb7d12b3f93ee918d40b1533b72da_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:43 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_12_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_12_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd85),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd86),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd121),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_10_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_12
// ------------------------------------------------------------------


module Fifo_ODTYPE_12 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_12_run Fifo_ODTYPE_12_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_11__31bade9fd05fb924a7bedeeff0d44833707b_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:51:51 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_11_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_11_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd82),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd83),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd122),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_9_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_11
// ------------------------------------------------------------------


module Fifo_ODTYPE_11 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_11_run Fifo_ODTYPE_11_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_10__f200e82bf6c1ead98f116d1648e23cec6e1d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:01 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_10_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_10_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd79),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd80),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd123),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_8_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_10
// ------------------------------------------------------------------


module Fifo_ODTYPE_10 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_10_run Fifo_ODTYPE_10_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_9__e738e5f75f1907c347b631a57f9915616bb3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:09 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_9_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_9_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd76),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd77),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd124),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_7_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_9
// ------------------------------------------------------------------


module Fifo_ODTYPE_9 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_9_run Fifo_ODTYPE_9_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_8__1fc8233da49ef9875c5241d4c5f4759f6955_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:17 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_8_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_8_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd73),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd74),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd125),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_6_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_8
// ------------------------------------------------------------------


module Fifo_ODTYPE_8 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_8_run Fifo_ODTYPE_8_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_7__044ac23b573abf031bfbf74b6c3218c666f7_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:25 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_7_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_7_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd70),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd71),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd126),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_5_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_7
// ------------------------------------------------------------------


module Fifo_ODTYPE_7 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_7_run Fifo_ODTYPE_7_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_6__ac9d9dc3ef096245180b91b761fa49fc6499_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:32 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_6_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_6_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd67),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd68),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd127),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_4_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_6
// ------------------------------------------------------------------


module Fifo_ODTYPE_6 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_6_run Fifo_ODTYPE_6_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_5__672f25d54775cea8cbecbd56d50e496a623b_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:40 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_5_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_5_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd64),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd65),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd128),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_3_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_5
// ------------------------------------------------------------------


module Fifo_ODTYPE_5 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_5_run Fifo_ODTYPE_5_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_4__cd2b76537cb81c7e66b90a768c8e6be75fdd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:48 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_4_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_4_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd61),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd62),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd129),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_2_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_4
// ------------------------------------------------------------------


module Fifo_ODTYPE_4 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_4_run Fifo_ODTYPE_4_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_3__02d3e5a754710daba473b818f4f831bf5d7f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:52:56 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_3_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_3_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd58),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd59),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd130),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_1_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_3
// ------------------------------------------------------------------


module Fifo_ODTYPE_3 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_3_run Fifo_ODTYPE_3_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_2__ac03de2b4e2534734bb0faf2dd2257465b21_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:04 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_2_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_2_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [15:0] regs_0_sva;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd55),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd56),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd131),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_0_sva;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_2
// ------------------------------------------------------------------


module Fifo_ODTYPE_2 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_2_run Fifo_ODTYPE_2_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_16__95124708f0678fb3fc12f90f4757ba9d7c29_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:20 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_16_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_16_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;
  reg [7:0] regs_13_sva_dfm;
  reg [7:0] regs_14_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd50),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd51),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd133),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_14_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_14_sva_dfm <= 8'b00000000;
      regs_13_sva_dfm <= 8'b00000000;
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_14_sva_dfm <= regs_13_sva_dfm;
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_16
// ------------------------------------------------------------------


module Fifo_IDTYPE_16 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_16_run Fifo_IDTYPE_16_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_15__f960108503a4c5f8415ed5adc9a9911579cb_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:28 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_15_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_15_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;
  reg [7:0] regs_13_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd47),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd48),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd134),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_13_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_13_sva_dfm <= 8'b00000000;
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_15
// ------------------------------------------------------------------


module Fifo_IDTYPE_15 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_15_run Fifo_IDTYPE_15_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_14__5498672fc186849f1a453e7578913ba4776d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:37 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_14_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_14_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd45),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd135),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_12_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_14
// ------------------------------------------------------------------


module Fifo_IDTYPE_14 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_14_run Fifo_IDTYPE_14_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_13__140c58040441cb68db13d83a1b3529a3750f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:45 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_13_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_13_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd41),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd42),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd136),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_11_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_13
// ------------------------------------------------------------------


module Fifo_IDTYPE_13 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_13_run Fifo_IDTYPE_13_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_12__97b113b64506d203c951f30f24019f9672b1_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:54 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_12_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_12_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd38),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd39),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd137),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_10_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_12
// ------------------------------------------------------------------


module Fifo_IDTYPE_12 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_12_run Fifo_IDTYPE_12_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_11__a50a5e9a32c085bccf8cadd9828ced0c7053_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:02 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_11_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_11_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd35),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd36),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd138),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_9_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_11
// ------------------------------------------------------------------


module Fifo_IDTYPE_11 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_11_run Fifo_IDTYPE_11_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_10__306a33ab3b28e00f5fee43b67cdfb4566df6_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:11 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_10_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_10_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd32),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd33),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd139),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_8_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_10
// ------------------------------------------------------------------


module Fifo_IDTYPE_10 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_10_run Fifo_IDTYPE_10_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_9__2cd80038408356854038769ee7a34b1b6b8d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:19 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_9_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_9_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd29),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd30),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd140),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_7_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_9
// ------------------------------------------------------------------


module Fifo_IDTYPE_9 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_9_run Fifo_IDTYPE_9_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_8__05bd72a244f928e63128b6b19625769c6930_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:28 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_8_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_8_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd26),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd27),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd141),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_6_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_8
// ------------------------------------------------------------------


module Fifo_IDTYPE_8 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_8_run Fifo_IDTYPE_8_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_7__d852beaa1f4c8fd838fbd9904419990066d3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:36 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_7_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_7_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd23),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd24),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd142),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_5_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_7
// ------------------------------------------------------------------


module Fifo_IDTYPE_7 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_7_run Fifo_IDTYPE_7_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_6__da4fb178783bbcbec6c48145d90a717b6476_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:45 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_6_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_6_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd20),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd21),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd143),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_4_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_6
// ------------------------------------------------------------------


module Fifo_IDTYPE_6 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_6_run Fifo_IDTYPE_6_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_5__ba9d0340e9908208b9fe8dbb6bf986706219_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:54:53 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_5_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_5_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd17),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd18),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd144),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_3_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_5
// ------------------------------------------------------------------


module Fifo_IDTYPE_5 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_5_run Fifo_IDTYPE_5_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_4__95ce258b6624ba5b1bc2748b6d950f545fbc_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:55:02 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_4_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_4_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd14),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd15),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd145),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_2_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_4
// ------------------------------------------------------------------


module Fifo_IDTYPE_4 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_4_run Fifo_IDTYPE_4_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_3__dbe2c0b9a0576493f3e2da2d3c31e1ff5d5f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:55:10 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_3_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_3_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd12),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd146),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_1_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_3
// ------------------------------------------------------------------


module Fifo_IDTYPE_3 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_3_run Fifo_IDTYPE_3_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_2__62c8d9056024328273aec1a1afbe23285b00_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:55:18 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_2_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_2_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [7:0] regs_0_sva;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd147),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_0_sva;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_0_sva <= 8'b00000000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_2
// ------------------------------------------------------------------


module Fifo_IDTYPE_2 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_2_run Fifo_IDTYPE_2_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../ProcessingElementless_IDTYPEcomma_ODTYPEgreater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy07
//  Generated date: Sun Feb 23 19:23:19 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ProcessingElement_IDTYPE_ODTYPE_run
// ------------------------------------------------------------------


module ProcessingElement_IDTYPE_ODTYPE_run (
  clk, arst_n, input_in_rsc_dat, psum_in_rsc_dat, weight_rsc_dat, input_out_rsc_z,
      psum_out_rsc_z, ccs_ccore_en
);
  input clk;
  input arst_n;
  input [7:0] input_in_rsc_dat;
  input [15:0] psum_in_rsc_dat;
  input [7:0] weight_rsc_dat;
  output [7:0] input_out_rsc_z;
  output [15:0] psum_out_rsc_z;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_in_rsci_idat;
  wire [15:0] psum_in_rsci_idat;
  wire [7:0] weight_rsci_idat;
  reg [7:0] input_out_rsci_d;
  reg [15:0] psum_out_rsci_d;
  wire [16:0] nl_psum_out_rsci_d;

  wire[15:0] mul_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd8)) input_in_rsci (
      .dat(input_in_rsc_dat),
      .idat(input_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) psum_in_rsci (
      .dat(psum_in_rsc_dat),
      .idat(psum_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd8)) weight_rsci (
      .dat(weight_rsc_dat),
      .idat(weight_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd8)) input_out_rsci (
      .d(input_out_rsci_d),
      .z(input_out_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd5),
  .width(32'sd16)) psum_out_rsci (
      .d(psum_out_rsci_d),
      .z(psum_out_rsc_z)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_out_rsci_d <= 8'b00000000;
      psum_out_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      input_out_rsci_d <= input_in_rsci_idat;
      psum_out_rsci_d <= nl_psum_out_rsci_d[15:0];
    end
  end
  assign mul_nl = conv_s2u_16_16($signed((input_in_rsci_idat)) * $signed((weight_rsci_idat)));
  assign nl_psum_out_rsci_d  = (mul_nl) + psum_in_rsci_idat;

  function automatic [15:0] conv_s2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_16 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ProcessingElement_IDTYPE_ODTYPE
// ------------------------------------------------------------------


module ProcessingElement_IDTYPE_ODTYPE (
  clk, arst_n, input_in_rsc_dat, psum_in_rsc_dat, weight_rsc_dat, input_out_rsc_z,
      psum_out_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_en
);
  input clk;
  input arst_n;
  input [7:0] input_in_rsc_dat;
  input [15:0] psum_in_rsc_dat;
  input [7:0] weight_rsc_dat;
  output [7:0] input_out_rsc_z;
  output [15:0] psum_out_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  ProcessingElement_IDTYPE_ODTYPE_run ProcessingElement_IDTYPE_ODTYPE_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .input_in_rsc_dat(input_in_rsc_dat),
      .psum_in_rsc_dat(psum_in_rsc_dat),
      .weight_rsc_dat(weight_rsc_dat),
      .input_out_rsc_z(input_out_rsc_z),
      .psum_out_rsc_z(psum_out_rsc_z),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_1__e8724e5d64a0158fc7643301a5bd75415451_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:53:12 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_1_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_1_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_clk, ccs_ccore_arst, ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd53),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd54),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_1
// ------------------------------------------------------------------


module Fifo_ODTYPE_1 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_1_run Fifo_ODTYPE_1_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_1__4010773ccc4167191cf2f733a2c976455432_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy16
//  Generated date: Sun Feb 23 16:55:27 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_1_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_1_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_clk, ccs_ccore_arst, ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_1
// ------------------------------------------------------------------


module Fifo_IDTYPE_1 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_1_run Fifo_IDTYPE_1_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../../../ee272-hw5/temp/sram_512_128.v 
// macro alternative to $clog2, which isn't supported by some tools
`define CLOG2(x) \
((x <= 1) || (x > 16384)) ? 0 : \
(x <= 2) ? 1 : \
(x <= 4) ? 2 : \
(x <= 8) ? 3 : \
(x <= 16) ? 4 : \
(x <= 32) ? 5 : \
(x <= 64) ? 6 : \
(x <= 128) ? 7: \
(x <= 256) ? 8: \
(x <= 512) ? 9 : \
(x <= 1024) ? 10: \
(x <= 2048) ? 11 : \
(x <= 4096) ? 12 : \
(x <= 8192) ? 13 : \
(x <= 16384) ? 14 : 0

// Wrapper module to create larger memories from smaller generated memories
module sram_512_128(
    clk, csb, web, addr, din, dout
);
    // set these values 
    parameter WRAPPER_DEPTH = 512;
    parameter WRAPPER_WIDTH = 128;
    parameter WRAPPER_ADDR_BITS = 9;

    input clk;
    input csb;
    input web;
    input [WRAPPER_ADDR_BITS-1:0] addr;
    input [WRAPPER_WIDTH-1:0] din;
    output [WRAPPER_WIDTH-1:0] dout;


    // Change these SRAM values:
    parameter SRAM_DEPTH = 128;
    parameter SRAM_WIDTH = 128;
    parameter SRAM_ADDR_BITS = 7;
    parameter num_inst_depth = WRAPPER_DEPTH / SRAM_DEPTH;
    parameter num_inst_width = WRAPPER_WIDTH / SRAM_WIDTH;
    genvar i,j;

    wire [num_inst_depth-1:0] sram_csb;
    wire [num_inst_depth-1:0] sram_web;
    wire [SRAM_ADDR_BITS-1:0] sram_address;
    wire [SRAM_WIDTH-1:0] sram_din [num_inst_width-1:0];
    wire [SRAM_WIDTH-1:0] sram_dout [num_inst_depth-1:0][num_inst_width-1:0];

    // upper bits of address are used as mem_select
    wire [WRAPPER_ADDR_BITS-SRAM_ADDR_BITS-1:0] mem_select;
    assign mem_select = addr[WRAPPER_ADDR_BITS-1:SRAM_ADDR_BITS];
    reg [WRAPPER_ADDR_BITS-SRAM_ADDR_BITS-1:0] output_mem_select;

    assign sram_csb = ~(csb) ? ~(1 << mem_select) : ~0;
    assign sram_web = ~(web) ? ~(1 << mem_select) : ~0;

    always @(posedge clk) begin
        if(csb == 0 & web == 0) begin
            output_mem_select <= mem_select;
        end
    end

    generate
    for(j = 0; j < num_inst_width; j=j+1) begin
        assign dout[(j+1)*SRAM_WIDTH-1:j*SRAM_WIDTH] = sram_dout[output_mem_select][j];
    end
    endgenerate

    generate
    for(i = 0; i < num_inst_depth; i=i+1) begin
        for(j = 0; j < num_inst_width; j=j+1) begin
            sram_128_128 #(.DELAY(1)) memory (
                .clk0(clk),
                .csb0(sram_csb[i]),
                .web0(sram_web[i]),
                .addr0(addr[SRAM_ADDR_BITS-1:0]),
                .din0(din[(j+1)*SRAM_WIDTH-1:j*SRAM_WIDTH]),
                .dout0(sram_dout[i][j])
            );
        end
    end
    endgenerate
endmodule



// synopsys translate_off
`include "/afs/ir.stanford.edu/class/ee272/OpenRAM/generated_memories/1RW/sram_128_128/sram_128_128.v"
// synopsys translate_on

//------> /afs/ir.stanford.edu/class/ee272/OpenRAM/generated_memories/1RW/sram_128_128/sram_128_128.v 
// OpenRAM SRAM model
// Words: 128
// Word size: 128

module sram_128_128(
// Port 0: RW
    clk0,csb0,web0,addr0,din0,dout0
  );

  parameter DATA_WIDTH = 128 ;
  parameter ADDR_WIDTH = 7 ;
  parameter RAM_DEPTH = 1 << ADDR_WIDTH;
  // FIXME: This delay is arbitrary.
  parameter DELAY = 3 ;

  input  clk0; // clock
  input   csb0; // active low chip select
  input  web0; // active low write control
  input [ADDR_WIDTH-1:0]  addr0;
  input [DATA_WIDTH-1:0]  din0;
  output [DATA_WIDTH-1:0] dout0;

  reg  csb0_reg;
  reg  web0_reg;
  reg [ADDR_WIDTH-1:0]  addr0_reg;
  reg [DATA_WIDTH-1:0]  din0_reg;
  reg [DATA_WIDTH-1:0]  dout0;

reg [DATA_WIDTH-1:0]    mem [0:RAM_DEPTH-1];

  // All inputs are registers
  always @(posedge clk0)
  begin
    csb0_reg = csb0;
    web0_reg = web0;
    addr0_reg = addr0;
    din0_reg = din0;
    dout0 = 128'bx;
    if ( !csb0_reg && web0_reg ) 
      $display($time," Reading %m addr0=%b dout0=%b",addr0_reg,mem[addr0_reg]);
    if ( !csb0_reg && !web0_reg )
      $display($time," Writing %m addr0=%b din0=%b",addr0_reg,din0_reg);
  end


  // Memory Write Block Port 0
  // Write Operation : When web0 = 0, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_WRITE0
    if ( !csb0_reg && !web0_reg )
        mem[addr0_reg] = din0_reg;
  end

  // Memory Read Block Port 0
  // Read Operation : When web0 = 1, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_READ0
    if (!csb0_reg && web0_reg)
       dout0 <= #(DELAY) mem[addr0_reg];
  end

endmodule

//------> ../SystolicArrayCoreless_IDTYPEcomma_WDTYPEcomma_ODTYPEcomma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy07
//  Generated date: Sun Feb 23 19:43:21 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_164_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_164_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_163_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_163_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_162_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_162_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_161_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_161_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_160_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_160_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_159_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_159_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_158_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_158_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_157_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_157_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_156_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_156_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_155_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_155_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_154_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_154_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_153_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_153_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_152_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_152_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_151_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_151_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_150_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_150_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_149_16_12_256_16_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_149_16_12_256_16_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [15:0] dout;
  output [15:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [15:0] din_d;
  output [15:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire accumulation_buffer_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign accumulation_buffer_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) &
      (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (accumulation_buffer_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, step_C_0_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input step_C_0_tr0;


  // FSM State Type Declaration for SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 9'd0,
    main_C_0 = 9'd1,
    step_C_0 = 9'd2,
    step_C_1 = 9'd3,
    step_C_2 = 9'd4,
    step_C_3 = 9'd5,
    step_C_4 = 9'd6,
    step_C_5 = 9'd7,
    step_C_6 = 9'd8,
    step_C_7 = 9'd9,
    step_C_8 = 9'd10,
    step_C_9 = 9'd11,
    step_C_10 = 9'd12,
    step_C_11 = 9'd13,
    step_C_12 = 9'd14,
    step_C_13 = 9'd15,
    step_C_14 = 9'd16,
    step_C_15 = 9'd17,
    step_C_16 = 9'd18,
    step_C_17 = 9'd19,
    step_C_18 = 9'd20,
    step_C_19 = 9'd21,
    step_C_20 = 9'd22,
    step_C_21 = 9'd23,
    step_C_22 = 9'd24,
    step_C_23 = 9'd25,
    step_C_24 = 9'd26,
    step_C_25 = 9'd27,
    step_C_26 = 9'd28,
    step_C_27 = 9'd29,
    step_C_28 = 9'd30,
    step_C_29 = 9'd31,
    step_C_30 = 9'd32,
    step_C_31 = 9'd33,
    step_C_32 = 9'd34,
    step_C_33 = 9'd35,
    step_C_34 = 9'd36,
    step_C_35 = 9'd37,
    step_C_36 = 9'd38,
    step_C_37 = 9'd39,
    step_C_38 = 9'd40,
    step_C_39 = 9'd41,
    step_C_40 = 9'd42,
    step_C_41 = 9'd43,
    step_C_42 = 9'd44,
    step_C_43 = 9'd45,
    step_C_44 = 9'd46,
    step_C_45 = 9'd47,
    step_C_46 = 9'd48,
    step_C_47 = 9'd49,
    step_C_48 = 9'd50,
    step_C_49 = 9'd51,
    step_C_50 = 9'd52,
    step_C_51 = 9'd53,
    step_C_52 = 9'd54,
    step_C_53 = 9'd55,
    step_C_54 = 9'd56,
    step_C_55 = 9'd57,
    step_C_56 = 9'd58,
    step_C_57 = 9'd59,
    step_C_58 = 9'd60,
    step_C_59 = 9'd61,
    step_C_60 = 9'd62,
    step_C_61 = 9'd63,
    step_C_62 = 9'd64,
    step_C_63 = 9'd65,
    step_C_64 = 9'd66,
    step_C_65 = 9'd67,
    step_C_66 = 9'd68,
    step_C_67 = 9'd69,
    step_C_68 = 9'd70,
    step_C_69 = 9'd71,
    step_C_70 = 9'd72,
    step_C_71 = 9'd73,
    step_C_72 = 9'd74,
    step_C_73 = 9'd75,
    step_C_74 = 9'd76,
    step_C_75 = 9'd77,
    step_C_76 = 9'd78,
    step_C_77 = 9'd79,
    step_C_78 = 9'd80,
    step_C_79 = 9'd81,
    step_C_80 = 9'd82,
    step_C_81 = 9'd83,
    step_C_82 = 9'd84,
    step_C_83 = 9'd85,
    step_C_84 = 9'd86,
    step_C_85 = 9'd87,
    step_C_86 = 9'd88,
    step_C_87 = 9'd89,
    step_C_88 = 9'd90,
    step_C_89 = 9'd91,
    step_C_90 = 9'd92,
    step_C_91 = 9'd93,
    step_C_92 = 9'd94,
    step_C_93 = 9'd95,
    step_C_94 = 9'd96,
    step_C_95 = 9'd97,
    step_C_96 = 9'd98,
    step_C_97 = 9'd99,
    step_C_98 = 9'd100,
    step_C_99 = 9'd101,
    step_C_100 = 9'd102,
    step_C_101 = 9'd103,
    step_C_102 = 9'd104,
    step_C_103 = 9'd105,
    step_C_104 = 9'd106,
    step_C_105 = 9'd107,
    step_C_106 = 9'd108,
    step_C_107 = 9'd109,
    step_C_108 = 9'd110,
    step_C_109 = 9'd111,
    step_C_110 = 9'd112,
    step_C_111 = 9'd113,
    step_C_112 = 9'd114,
    step_C_113 = 9'd115,
    step_C_114 = 9'd116,
    step_C_115 = 9'd117,
    step_C_116 = 9'd118,
    step_C_117 = 9'd119,
    step_C_118 = 9'd120,
    step_C_119 = 9'd121,
    step_C_120 = 9'd122,
    step_C_121 = 9'd123,
    step_C_122 = 9'd124,
    step_C_123 = 9'd125,
    step_C_124 = 9'd126,
    step_C_125 = 9'd127,
    step_C_126 = 9'd128,
    step_C_127 = 9'd129,
    step_C_128 = 9'd130,
    step_C_129 = 9'd131,
    step_C_130 = 9'd132,
    step_C_131 = 9'd133,
    step_C_132 = 9'd134,
    step_C_133 = 9'd135,
    step_C_134 = 9'd136,
    step_C_135 = 9'd137,
    step_C_136 = 9'd138,
    step_C_137 = 9'd139,
    step_C_138 = 9'd140,
    step_C_139 = 9'd141,
    step_C_140 = 9'd142,
    step_C_141 = 9'd143,
    step_C_142 = 9'd144,
    step_C_143 = 9'd145,
    step_C_144 = 9'd146,
    step_C_145 = 9'd147,
    step_C_146 = 9'd148,
    step_C_147 = 9'd149,
    step_C_148 = 9'd150,
    step_C_149 = 9'd151,
    step_C_150 = 9'd152,
    step_C_151 = 9'd153,
    step_C_152 = 9'd154,
    step_C_153 = 9'd155,
    step_C_154 = 9'd156,
    step_C_155 = 9'd157,
    step_C_156 = 9'd158,
    step_C_157 = 9'd159,
    step_C_158 = 9'd160,
    step_C_159 = 9'd161,
    step_C_160 = 9'd162,
    step_C_161 = 9'd163,
    step_C_162 = 9'd164,
    step_C_163 = 9'd165,
    step_C_164 = 9'd166,
    step_C_165 = 9'd167,
    step_C_166 = 9'd168,
    step_C_167 = 9'd169,
    step_C_168 = 9'd170,
    step_C_169 = 9'd171,
    step_C_170 = 9'd172,
    step_C_171 = 9'd173,
    step_C_172 = 9'd174,
    step_C_173 = 9'd175,
    step_C_174 = 9'd176,
    step_C_175 = 9'd177,
    step_C_176 = 9'd178,
    step_C_177 = 9'd179,
    step_C_178 = 9'd180,
    step_C_179 = 9'd181,
    step_C_180 = 9'd182,
    step_C_181 = 9'd183,
    step_C_182 = 9'd184,
    step_C_183 = 9'd185,
    step_C_184 = 9'd186,
    step_C_185 = 9'd187,
    step_C_186 = 9'd188,
    step_C_187 = 9'd189,
    step_C_188 = 9'd190,
    step_C_189 = 9'd191,
    step_C_190 = 9'd192,
    step_C_191 = 9'd193,
    step_C_192 = 9'd194,
    step_C_193 = 9'd195,
    step_C_194 = 9'd196,
    step_C_195 = 9'd197,
    step_C_196 = 9'd198,
    step_C_197 = 9'd199,
    step_C_198 = 9'd200,
    step_C_199 = 9'd201,
    step_C_200 = 9'd202,
    step_C_201 = 9'd203,
    step_C_202 = 9'd204,
    step_C_203 = 9'd205,
    step_C_204 = 9'd206,
    step_C_205 = 9'd207,
    step_C_206 = 9'd208,
    step_C_207 = 9'd209,
    step_C_208 = 9'd210,
    step_C_209 = 9'd211,
    step_C_210 = 9'd212,
    step_C_211 = 9'd213,
    step_C_212 = 9'd214,
    step_C_213 = 9'd215,
    step_C_214 = 9'd216,
    step_C_215 = 9'd217,
    step_C_216 = 9'd218,
    step_C_217 = 9'd219,
    step_C_218 = 9'd220,
    step_C_219 = 9'd221,
    step_C_220 = 9'd222,
    step_C_221 = 9'd223,
    step_C_222 = 9'd224,
    step_C_223 = 9'd225,
    step_C_224 = 9'd226,
    step_C_225 = 9'd227,
    step_C_226 = 9'd228,
    step_C_227 = 9'd229,
    step_C_228 = 9'd230,
    step_C_229 = 9'd231,
    step_C_230 = 9'd232,
    step_C_231 = 9'd233,
    step_C_232 = 9'd234,
    step_C_233 = 9'd235,
    step_C_234 = 9'd236,
    step_C_235 = 9'd237,
    step_C_236 = 9'd238,
    step_C_237 = 9'd239,
    step_C_238 = 9'd240,
    step_C_239 = 9'd241,
    step_C_240 = 9'd242,
    step_C_241 = 9'd243,
    step_C_242 = 9'd244,
    step_C_243 = 9'd245,
    step_C_244 = 9'd246,
    step_C_245 = 9'd247,
    step_C_246 = 9'd248,
    step_C_247 = 9'd249,
    step_C_248 = 9'd250,
    step_C_249 = 9'd251,
    step_C_250 = 9'd252,
    step_C_251 = 9'd253,
    step_C_252 = 9'd254,
    step_C_253 = 9'd255,
    step_C_254 = 9'd256,
    step_C_255 = 9'd257,
    step_C_256 = 9'd258,
    step_C_257 = 9'd259;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000001;
        state_var_NS = step_C_0;
      end
      step_C_0 : begin
        fsm_output = 9'b000000010;
        if ( step_C_0_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = step_C_1;
        end
      end
      step_C_1 : begin
        fsm_output = 9'b000000011;
        state_var_NS = step_C_2;
      end
      step_C_2 : begin
        fsm_output = 9'b000000100;
        state_var_NS = step_C_3;
      end
      step_C_3 : begin
        fsm_output = 9'b000000101;
        state_var_NS = step_C_4;
      end
      step_C_4 : begin
        fsm_output = 9'b000000110;
        state_var_NS = step_C_5;
      end
      step_C_5 : begin
        fsm_output = 9'b000000111;
        state_var_NS = step_C_6;
      end
      step_C_6 : begin
        fsm_output = 9'b000001000;
        state_var_NS = step_C_7;
      end
      step_C_7 : begin
        fsm_output = 9'b000001001;
        state_var_NS = step_C_8;
      end
      step_C_8 : begin
        fsm_output = 9'b000001010;
        state_var_NS = step_C_9;
      end
      step_C_9 : begin
        fsm_output = 9'b000001011;
        state_var_NS = step_C_10;
      end
      step_C_10 : begin
        fsm_output = 9'b000001100;
        state_var_NS = step_C_11;
      end
      step_C_11 : begin
        fsm_output = 9'b000001101;
        state_var_NS = step_C_12;
      end
      step_C_12 : begin
        fsm_output = 9'b000001110;
        state_var_NS = step_C_13;
      end
      step_C_13 : begin
        fsm_output = 9'b000001111;
        state_var_NS = step_C_14;
      end
      step_C_14 : begin
        fsm_output = 9'b000010000;
        state_var_NS = step_C_15;
      end
      step_C_15 : begin
        fsm_output = 9'b000010001;
        state_var_NS = step_C_16;
      end
      step_C_16 : begin
        fsm_output = 9'b000010010;
        state_var_NS = step_C_17;
      end
      step_C_17 : begin
        fsm_output = 9'b000010011;
        state_var_NS = step_C_18;
      end
      step_C_18 : begin
        fsm_output = 9'b000010100;
        state_var_NS = step_C_19;
      end
      step_C_19 : begin
        fsm_output = 9'b000010101;
        state_var_NS = step_C_20;
      end
      step_C_20 : begin
        fsm_output = 9'b000010110;
        state_var_NS = step_C_21;
      end
      step_C_21 : begin
        fsm_output = 9'b000010111;
        state_var_NS = step_C_22;
      end
      step_C_22 : begin
        fsm_output = 9'b000011000;
        state_var_NS = step_C_23;
      end
      step_C_23 : begin
        fsm_output = 9'b000011001;
        state_var_NS = step_C_24;
      end
      step_C_24 : begin
        fsm_output = 9'b000011010;
        state_var_NS = step_C_25;
      end
      step_C_25 : begin
        fsm_output = 9'b000011011;
        state_var_NS = step_C_26;
      end
      step_C_26 : begin
        fsm_output = 9'b000011100;
        state_var_NS = step_C_27;
      end
      step_C_27 : begin
        fsm_output = 9'b000011101;
        state_var_NS = step_C_28;
      end
      step_C_28 : begin
        fsm_output = 9'b000011110;
        state_var_NS = step_C_29;
      end
      step_C_29 : begin
        fsm_output = 9'b000011111;
        state_var_NS = step_C_30;
      end
      step_C_30 : begin
        fsm_output = 9'b000100000;
        state_var_NS = step_C_31;
      end
      step_C_31 : begin
        fsm_output = 9'b000100001;
        state_var_NS = step_C_32;
      end
      step_C_32 : begin
        fsm_output = 9'b000100010;
        state_var_NS = step_C_33;
      end
      step_C_33 : begin
        fsm_output = 9'b000100011;
        state_var_NS = step_C_34;
      end
      step_C_34 : begin
        fsm_output = 9'b000100100;
        state_var_NS = step_C_35;
      end
      step_C_35 : begin
        fsm_output = 9'b000100101;
        state_var_NS = step_C_36;
      end
      step_C_36 : begin
        fsm_output = 9'b000100110;
        state_var_NS = step_C_37;
      end
      step_C_37 : begin
        fsm_output = 9'b000100111;
        state_var_NS = step_C_38;
      end
      step_C_38 : begin
        fsm_output = 9'b000101000;
        state_var_NS = step_C_39;
      end
      step_C_39 : begin
        fsm_output = 9'b000101001;
        state_var_NS = step_C_40;
      end
      step_C_40 : begin
        fsm_output = 9'b000101010;
        state_var_NS = step_C_41;
      end
      step_C_41 : begin
        fsm_output = 9'b000101011;
        state_var_NS = step_C_42;
      end
      step_C_42 : begin
        fsm_output = 9'b000101100;
        state_var_NS = step_C_43;
      end
      step_C_43 : begin
        fsm_output = 9'b000101101;
        state_var_NS = step_C_44;
      end
      step_C_44 : begin
        fsm_output = 9'b000101110;
        state_var_NS = step_C_45;
      end
      step_C_45 : begin
        fsm_output = 9'b000101111;
        state_var_NS = step_C_46;
      end
      step_C_46 : begin
        fsm_output = 9'b000110000;
        state_var_NS = step_C_47;
      end
      step_C_47 : begin
        fsm_output = 9'b000110001;
        state_var_NS = step_C_48;
      end
      step_C_48 : begin
        fsm_output = 9'b000110010;
        state_var_NS = step_C_49;
      end
      step_C_49 : begin
        fsm_output = 9'b000110011;
        state_var_NS = step_C_50;
      end
      step_C_50 : begin
        fsm_output = 9'b000110100;
        state_var_NS = step_C_51;
      end
      step_C_51 : begin
        fsm_output = 9'b000110101;
        state_var_NS = step_C_52;
      end
      step_C_52 : begin
        fsm_output = 9'b000110110;
        state_var_NS = step_C_53;
      end
      step_C_53 : begin
        fsm_output = 9'b000110111;
        state_var_NS = step_C_54;
      end
      step_C_54 : begin
        fsm_output = 9'b000111000;
        state_var_NS = step_C_55;
      end
      step_C_55 : begin
        fsm_output = 9'b000111001;
        state_var_NS = step_C_56;
      end
      step_C_56 : begin
        fsm_output = 9'b000111010;
        state_var_NS = step_C_57;
      end
      step_C_57 : begin
        fsm_output = 9'b000111011;
        state_var_NS = step_C_58;
      end
      step_C_58 : begin
        fsm_output = 9'b000111100;
        state_var_NS = step_C_59;
      end
      step_C_59 : begin
        fsm_output = 9'b000111101;
        state_var_NS = step_C_60;
      end
      step_C_60 : begin
        fsm_output = 9'b000111110;
        state_var_NS = step_C_61;
      end
      step_C_61 : begin
        fsm_output = 9'b000111111;
        state_var_NS = step_C_62;
      end
      step_C_62 : begin
        fsm_output = 9'b001000000;
        state_var_NS = step_C_63;
      end
      step_C_63 : begin
        fsm_output = 9'b001000001;
        state_var_NS = step_C_64;
      end
      step_C_64 : begin
        fsm_output = 9'b001000010;
        state_var_NS = step_C_65;
      end
      step_C_65 : begin
        fsm_output = 9'b001000011;
        state_var_NS = step_C_66;
      end
      step_C_66 : begin
        fsm_output = 9'b001000100;
        state_var_NS = step_C_67;
      end
      step_C_67 : begin
        fsm_output = 9'b001000101;
        state_var_NS = step_C_68;
      end
      step_C_68 : begin
        fsm_output = 9'b001000110;
        state_var_NS = step_C_69;
      end
      step_C_69 : begin
        fsm_output = 9'b001000111;
        state_var_NS = step_C_70;
      end
      step_C_70 : begin
        fsm_output = 9'b001001000;
        state_var_NS = step_C_71;
      end
      step_C_71 : begin
        fsm_output = 9'b001001001;
        state_var_NS = step_C_72;
      end
      step_C_72 : begin
        fsm_output = 9'b001001010;
        state_var_NS = step_C_73;
      end
      step_C_73 : begin
        fsm_output = 9'b001001011;
        state_var_NS = step_C_74;
      end
      step_C_74 : begin
        fsm_output = 9'b001001100;
        state_var_NS = step_C_75;
      end
      step_C_75 : begin
        fsm_output = 9'b001001101;
        state_var_NS = step_C_76;
      end
      step_C_76 : begin
        fsm_output = 9'b001001110;
        state_var_NS = step_C_77;
      end
      step_C_77 : begin
        fsm_output = 9'b001001111;
        state_var_NS = step_C_78;
      end
      step_C_78 : begin
        fsm_output = 9'b001010000;
        state_var_NS = step_C_79;
      end
      step_C_79 : begin
        fsm_output = 9'b001010001;
        state_var_NS = step_C_80;
      end
      step_C_80 : begin
        fsm_output = 9'b001010010;
        state_var_NS = step_C_81;
      end
      step_C_81 : begin
        fsm_output = 9'b001010011;
        state_var_NS = step_C_82;
      end
      step_C_82 : begin
        fsm_output = 9'b001010100;
        state_var_NS = step_C_83;
      end
      step_C_83 : begin
        fsm_output = 9'b001010101;
        state_var_NS = step_C_84;
      end
      step_C_84 : begin
        fsm_output = 9'b001010110;
        state_var_NS = step_C_85;
      end
      step_C_85 : begin
        fsm_output = 9'b001010111;
        state_var_NS = step_C_86;
      end
      step_C_86 : begin
        fsm_output = 9'b001011000;
        state_var_NS = step_C_87;
      end
      step_C_87 : begin
        fsm_output = 9'b001011001;
        state_var_NS = step_C_88;
      end
      step_C_88 : begin
        fsm_output = 9'b001011010;
        state_var_NS = step_C_89;
      end
      step_C_89 : begin
        fsm_output = 9'b001011011;
        state_var_NS = step_C_90;
      end
      step_C_90 : begin
        fsm_output = 9'b001011100;
        state_var_NS = step_C_91;
      end
      step_C_91 : begin
        fsm_output = 9'b001011101;
        state_var_NS = step_C_92;
      end
      step_C_92 : begin
        fsm_output = 9'b001011110;
        state_var_NS = step_C_93;
      end
      step_C_93 : begin
        fsm_output = 9'b001011111;
        state_var_NS = step_C_94;
      end
      step_C_94 : begin
        fsm_output = 9'b001100000;
        state_var_NS = step_C_95;
      end
      step_C_95 : begin
        fsm_output = 9'b001100001;
        state_var_NS = step_C_96;
      end
      step_C_96 : begin
        fsm_output = 9'b001100010;
        state_var_NS = step_C_97;
      end
      step_C_97 : begin
        fsm_output = 9'b001100011;
        state_var_NS = step_C_98;
      end
      step_C_98 : begin
        fsm_output = 9'b001100100;
        state_var_NS = step_C_99;
      end
      step_C_99 : begin
        fsm_output = 9'b001100101;
        state_var_NS = step_C_100;
      end
      step_C_100 : begin
        fsm_output = 9'b001100110;
        state_var_NS = step_C_101;
      end
      step_C_101 : begin
        fsm_output = 9'b001100111;
        state_var_NS = step_C_102;
      end
      step_C_102 : begin
        fsm_output = 9'b001101000;
        state_var_NS = step_C_103;
      end
      step_C_103 : begin
        fsm_output = 9'b001101001;
        state_var_NS = step_C_104;
      end
      step_C_104 : begin
        fsm_output = 9'b001101010;
        state_var_NS = step_C_105;
      end
      step_C_105 : begin
        fsm_output = 9'b001101011;
        state_var_NS = step_C_106;
      end
      step_C_106 : begin
        fsm_output = 9'b001101100;
        state_var_NS = step_C_107;
      end
      step_C_107 : begin
        fsm_output = 9'b001101101;
        state_var_NS = step_C_108;
      end
      step_C_108 : begin
        fsm_output = 9'b001101110;
        state_var_NS = step_C_109;
      end
      step_C_109 : begin
        fsm_output = 9'b001101111;
        state_var_NS = step_C_110;
      end
      step_C_110 : begin
        fsm_output = 9'b001110000;
        state_var_NS = step_C_111;
      end
      step_C_111 : begin
        fsm_output = 9'b001110001;
        state_var_NS = step_C_112;
      end
      step_C_112 : begin
        fsm_output = 9'b001110010;
        state_var_NS = step_C_113;
      end
      step_C_113 : begin
        fsm_output = 9'b001110011;
        state_var_NS = step_C_114;
      end
      step_C_114 : begin
        fsm_output = 9'b001110100;
        state_var_NS = step_C_115;
      end
      step_C_115 : begin
        fsm_output = 9'b001110101;
        state_var_NS = step_C_116;
      end
      step_C_116 : begin
        fsm_output = 9'b001110110;
        state_var_NS = step_C_117;
      end
      step_C_117 : begin
        fsm_output = 9'b001110111;
        state_var_NS = step_C_118;
      end
      step_C_118 : begin
        fsm_output = 9'b001111000;
        state_var_NS = step_C_119;
      end
      step_C_119 : begin
        fsm_output = 9'b001111001;
        state_var_NS = step_C_120;
      end
      step_C_120 : begin
        fsm_output = 9'b001111010;
        state_var_NS = step_C_121;
      end
      step_C_121 : begin
        fsm_output = 9'b001111011;
        state_var_NS = step_C_122;
      end
      step_C_122 : begin
        fsm_output = 9'b001111100;
        state_var_NS = step_C_123;
      end
      step_C_123 : begin
        fsm_output = 9'b001111101;
        state_var_NS = step_C_124;
      end
      step_C_124 : begin
        fsm_output = 9'b001111110;
        state_var_NS = step_C_125;
      end
      step_C_125 : begin
        fsm_output = 9'b001111111;
        state_var_NS = step_C_126;
      end
      step_C_126 : begin
        fsm_output = 9'b010000000;
        state_var_NS = step_C_127;
      end
      step_C_127 : begin
        fsm_output = 9'b010000001;
        state_var_NS = step_C_128;
      end
      step_C_128 : begin
        fsm_output = 9'b010000010;
        state_var_NS = step_C_129;
      end
      step_C_129 : begin
        fsm_output = 9'b010000011;
        state_var_NS = step_C_130;
      end
      step_C_130 : begin
        fsm_output = 9'b010000100;
        state_var_NS = step_C_131;
      end
      step_C_131 : begin
        fsm_output = 9'b010000101;
        state_var_NS = step_C_132;
      end
      step_C_132 : begin
        fsm_output = 9'b010000110;
        state_var_NS = step_C_133;
      end
      step_C_133 : begin
        fsm_output = 9'b010000111;
        state_var_NS = step_C_134;
      end
      step_C_134 : begin
        fsm_output = 9'b010001000;
        state_var_NS = step_C_135;
      end
      step_C_135 : begin
        fsm_output = 9'b010001001;
        state_var_NS = step_C_136;
      end
      step_C_136 : begin
        fsm_output = 9'b010001010;
        state_var_NS = step_C_137;
      end
      step_C_137 : begin
        fsm_output = 9'b010001011;
        state_var_NS = step_C_138;
      end
      step_C_138 : begin
        fsm_output = 9'b010001100;
        state_var_NS = step_C_139;
      end
      step_C_139 : begin
        fsm_output = 9'b010001101;
        state_var_NS = step_C_140;
      end
      step_C_140 : begin
        fsm_output = 9'b010001110;
        state_var_NS = step_C_141;
      end
      step_C_141 : begin
        fsm_output = 9'b010001111;
        state_var_NS = step_C_142;
      end
      step_C_142 : begin
        fsm_output = 9'b010010000;
        state_var_NS = step_C_143;
      end
      step_C_143 : begin
        fsm_output = 9'b010010001;
        state_var_NS = step_C_144;
      end
      step_C_144 : begin
        fsm_output = 9'b010010010;
        state_var_NS = step_C_145;
      end
      step_C_145 : begin
        fsm_output = 9'b010010011;
        state_var_NS = step_C_146;
      end
      step_C_146 : begin
        fsm_output = 9'b010010100;
        state_var_NS = step_C_147;
      end
      step_C_147 : begin
        fsm_output = 9'b010010101;
        state_var_NS = step_C_148;
      end
      step_C_148 : begin
        fsm_output = 9'b010010110;
        state_var_NS = step_C_149;
      end
      step_C_149 : begin
        fsm_output = 9'b010010111;
        state_var_NS = step_C_150;
      end
      step_C_150 : begin
        fsm_output = 9'b010011000;
        state_var_NS = step_C_151;
      end
      step_C_151 : begin
        fsm_output = 9'b010011001;
        state_var_NS = step_C_152;
      end
      step_C_152 : begin
        fsm_output = 9'b010011010;
        state_var_NS = step_C_153;
      end
      step_C_153 : begin
        fsm_output = 9'b010011011;
        state_var_NS = step_C_154;
      end
      step_C_154 : begin
        fsm_output = 9'b010011100;
        state_var_NS = step_C_155;
      end
      step_C_155 : begin
        fsm_output = 9'b010011101;
        state_var_NS = step_C_156;
      end
      step_C_156 : begin
        fsm_output = 9'b010011110;
        state_var_NS = step_C_157;
      end
      step_C_157 : begin
        fsm_output = 9'b010011111;
        state_var_NS = step_C_158;
      end
      step_C_158 : begin
        fsm_output = 9'b010100000;
        state_var_NS = step_C_159;
      end
      step_C_159 : begin
        fsm_output = 9'b010100001;
        state_var_NS = step_C_160;
      end
      step_C_160 : begin
        fsm_output = 9'b010100010;
        state_var_NS = step_C_161;
      end
      step_C_161 : begin
        fsm_output = 9'b010100011;
        state_var_NS = step_C_162;
      end
      step_C_162 : begin
        fsm_output = 9'b010100100;
        state_var_NS = step_C_163;
      end
      step_C_163 : begin
        fsm_output = 9'b010100101;
        state_var_NS = step_C_164;
      end
      step_C_164 : begin
        fsm_output = 9'b010100110;
        state_var_NS = step_C_165;
      end
      step_C_165 : begin
        fsm_output = 9'b010100111;
        state_var_NS = step_C_166;
      end
      step_C_166 : begin
        fsm_output = 9'b010101000;
        state_var_NS = step_C_167;
      end
      step_C_167 : begin
        fsm_output = 9'b010101001;
        state_var_NS = step_C_168;
      end
      step_C_168 : begin
        fsm_output = 9'b010101010;
        state_var_NS = step_C_169;
      end
      step_C_169 : begin
        fsm_output = 9'b010101011;
        state_var_NS = step_C_170;
      end
      step_C_170 : begin
        fsm_output = 9'b010101100;
        state_var_NS = step_C_171;
      end
      step_C_171 : begin
        fsm_output = 9'b010101101;
        state_var_NS = step_C_172;
      end
      step_C_172 : begin
        fsm_output = 9'b010101110;
        state_var_NS = step_C_173;
      end
      step_C_173 : begin
        fsm_output = 9'b010101111;
        state_var_NS = step_C_174;
      end
      step_C_174 : begin
        fsm_output = 9'b010110000;
        state_var_NS = step_C_175;
      end
      step_C_175 : begin
        fsm_output = 9'b010110001;
        state_var_NS = step_C_176;
      end
      step_C_176 : begin
        fsm_output = 9'b010110010;
        state_var_NS = step_C_177;
      end
      step_C_177 : begin
        fsm_output = 9'b010110011;
        state_var_NS = step_C_178;
      end
      step_C_178 : begin
        fsm_output = 9'b010110100;
        state_var_NS = step_C_179;
      end
      step_C_179 : begin
        fsm_output = 9'b010110101;
        state_var_NS = step_C_180;
      end
      step_C_180 : begin
        fsm_output = 9'b010110110;
        state_var_NS = step_C_181;
      end
      step_C_181 : begin
        fsm_output = 9'b010110111;
        state_var_NS = step_C_182;
      end
      step_C_182 : begin
        fsm_output = 9'b010111000;
        state_var_NS = step_C_183;
      end
      step_C_183 : begin
        fsm_output = 9'b010111001;
        state_var_NS = step_C_184;
      end
      step_C_184 : begin
        fsm_output = 9'b010111010;
        state_var_NS = step_C_185;
      end
      step_C_185 : begin
        fsm_output = 9'b010111011;
        state_var_NS = step_C_186;
      end
      step_C_186 : begin
        fsm_output = 9'b010111100;
        state_var_NS = step_C_187;
      end
      step_C_187 : begin
        fsm_output = 9'b010111101;
        state_var_NS = step_C_188;
      end
      step_C_188 : begin
        fsm_output = 9'b010111110;
        state_var_NS = step_C_189;
      end
      step_C_189 : begin
        fsm_output = 9'b010111111;
        state_var_NS = step_C_190;
      end
      step_C_190 : begin
        fsm_output = 9'b011000000;
        state_var_NS = step_C_191;
      end
      step_C_191 : begin
        fsm_output = 9'b011000001;
        state_var_NS = step_C_192;
      end
      step_C_192 : begin
        fsm_output = 9'b011000010;
        state_var_NS = step_C_193;
      end
      step_C_193 : begin
        fsm_output = 9'b011000011;
        state_var_NS = step_C_194;
      end
      step_C_194 : begin
        fsm_output = 9'b011000100;
        state_var_NS = step_C_195;
      end
      step_C_195 : begin
        fsm_output = 9'b011000101;
        state_var_NS = step_C_196;
      end
      step_C_196 : begin
        fsm_output = 9'b011000110;
        state_var_NS = step_C_197;
      end
      step_C_197 : begin
        fsm_output = 9'b011000111;
        state_var_NS = step_C_198;
      end
      step_C_198 : begin
        fsm_output = 9'b011001000;
        state_var_NS = step_C_199;
      end
      step_C_199 : begin
        fsm_output = 9'b011001001;
        state_var_NS = step_C_200;
      end
      step_C_200 : begin
        fsm_output = 9'b011001010;
        state_var_NS = step_C_201;
      end
      step_C_201 : begin
        fsm_output = 9'b011001011;
        state_var_NS = step_C_202;
      end
      step_C_202 : begin
        fsm_output = 9'b011001100;
        state_var_NS = step_C_203;
      end
      step_C_203 : begin
        fsm_output = 9'b011001101;
        state_var_NS = step_C_204;
      end
      step_C_204 : begin
        fsm_output = 9'b011001110;
        state_var_NS = step_C_205;
      end
      step_C_205 : begin
        fsm_output = 9'b011001111;
        state_var_NS = step_C_206;
      end
      step_C_206 : begin
        fsm_output = 9'b011010000;
        state_var_NS = step_C_207;
      end
      step_C_207 : begin
        fsm_output = 9'b011010001;
        state_var_NS = step_C_208;
      end
      step_C_208 : begin
        fsm_output = 9'b011010010;
        state_var_NS = step_C_209;
      end
      step_C_209 : begin
        fsm_output = 9'b011010011;
        state_var_NS = step_C_210;
      end
      step_C_210 : begin
        fsm_output = 9'b011010100;
        state_var_NS = step_C_211;
      end
      step_C_211 : begin
        fsm_output = 9'b011010101;
        state_var_NS = step_C_212;
      end
      step_C_212 : begin
        fsm_output = 9'b011010110;
        state_var_NS = step_C_213;
      end
      step_C_213 : begin
        fsm_output = 9'b011010111;
        state_var_NS = step_C_214;
      end
      step_C_214 : begin
        fsm_output = 9'b011011000;
        state_var_NS = step_C_215;
      end
      step_C_215 : begin
        fsm_output = 9'b011011001;
        state_var_NS = step_C_216;
      end
      step_C_216 : begin
        fsm_output = 9'b011011010;
        state_var_NS = step_C_217;
      end
      step_C_217 : begin
        fsm_output = 9'b011011011;
        state_var_NS = step_C_218;
      end
      step_C_218 : begin
        fsm_output = 9'b011011100;
        state_var_NS = step_C_219;
      end
      step_C_219 : begin
        fsm_output = 9'b011011101;
        state_var_NS = step_C_220;
      end
      step_C_220 : begin
        fsm_output = 9'b011011110;
        state_var_NS = step_C_221;
      end
      step_C_221 : begin
        fsm_output = 9'b011011111;
        state_var_NS = step_C_222;
      end
      step_C_222 : begin
        fsm_output = 9'b011100000;
        state_var_NS = step_C_223;
      end
      step_C_223 : begin
        fsm_output = 9'b011100001;
        state_var_NS = step_C_224;
      end
      step_C_224 : begin
        fsm_output = 9'b011100010;
        state_var_NS = step_C_225;
      end
      step_C_225 : begin
        fsm_output = 9'b011100011;
        state_var_NS = step_C_226;
      end
      step_C_226 : begin
        fsm_output = 9'b011100100;
        state_var_NS = step_C_227;
      end
      step_C_227 : begin
        fsm_output = 9'b011100101;
        state_var_NS = step_C_228;
      end
      step_C_228 : begin
        fsm_output = 9'b011100110;
        state_var_NS = step_C_229;
      end
      step_C_229 : begin
        fsm_output = 9'b011100111;
        state_var_NS = step_C_230;
      end
      step_C_230 : begin
        fsm_output = 9'b011101000;
        state_var_NS = step_C_231;
      end
      step_C_231 : begin
        fsm_output = 9'b011101001;
        state_var_NS = step_C_232;
      end
      step_C_232 : begin
        fsm_output = 9'b011101010;
        state_var_NS = step_C_233;
      end
      step_C_233 : begin
        fsm_output = 9'b011101011;
        state_var_NS = step_C_234;
      end
      step_C_234 : begin
        fsm_output = 9'b011101100;
        state_var_NS = step_C_235;
      end
      step_C_235 : begin
        fsm_output = 9'b011101101;
        state_var_NS = step_C_236;
      end
      step_C_236 : begin
        fsm_output = 9'b011101110;
        state_var_NS = step_C_237;
      end
      step_C_237 : begin
        fsm_output = 9'b011101111;
        state_var_NS = step_C_238;
      end
      step_C_238 : begin
        fsm_output = 9'b011110000;
        state_var_NS = step_C_239;
      end
      step_C_239 : begin
        fsm_output = 9'b011110001;
        state_var_NS = step_C_240;
      end
      step_C_240 : begin
        fsm_output = 9'b011110010;
        state_var_NS = step_C_241;
      end
      step_C_241 : begin
        fsm_output = 9'b011110011;
        state_var_NS = step_C_242;
      end
      step_C_242 : begin
        fsm_output = 9'b011110100;
        state_var_NS = step_C_243;
      end
      step_C_243 : begin
        fsm_output = 9'b011110101;
        state_var_NS = step_C_244;
      end
      step_C_244 : begin
        fsm_output = 9'b011110110;
        state_var_NS = step_C_245;
      end
      step_C_245 : begin
        fsm_output = 9'b011110111;
        state_var_NS = step_C_246;
      end
      step_C_246 : begin
        fsm_output = 9'b011111000;
        state_var_NS = step_C_247;
      end
      step_C_247 : begin
        fsm_output = 9'b011111001;
        state_var_NS = step_C_248;
      end
      step_C_248 : begin
        fsm_output = 9'b011111010;
        state_var_NS = step_C_249;
      end
      step_C_249 : begin
        fsm_output = 9'b011111011;
        state_var_NS = step_C_250;
      end
      step_C_250 : begin
        fsm_output = 9'b011111100;
        state_var_NS = step_C_251;
      end
      step_C_251 : begin
        fsm_output = 9'b011111101;
        state_var_NS = step_C_252;
      end
      step_C_252 : begin
        fsm_output = 9'b011111110;
        state_var_NS = step_C_253;
      end
      step_C_253 : begin
        fsm_output = 9'b011111111;
        state_var_NS = step_C_254;
      end
      step_C_254 : begin
        fsm_output = 9'b100000000;
        state_var_NS = step_C_255;
      end
      step_C_255 : begin
        fsm_output = 9'b100000001;
        state_var_NS = step_C_256;
      end
      step_C_256 : begin
        fsm_output = 9'b100000010;
        state_var_NS = step_C_257;
      end
      step_C_257 : begin
        fsm_output = 9'b100000011;
        state_var_NS = step_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, input_rsci_wen_comp, weight_rsci_wen_comp, output_rsci_wen_comp,
      paramsIn_rsci_wen_comp, loopIndicesIn_rsci_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input input_rsci_wen_comp;
  input weight_rsci_wen_comp;
  input output_rsci_wen_comp;
  input paramsIn_rsci_wen_comp;
  input loopIndicesIn_rsci_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_rsci_wen_comp & weight_rsci_wen_comp & output_rsci_wen_comp
      & paramsIn_rsci_wen_comp & loopIndicesIn_rsci_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp (
  ensig_cgo_iro, ensig_cgo_iro_1, ensig_cgo_iro_30, ensig_cgo_iro_45, ensig_cgo_iro_46,
      run_wen, ensig_cgo, accum_fifo_15_rsci_ccs_ccore_en, ensig_cgo_1, output_fifo_0_rsci_ccs_ccore_en,
      ensig_cgo_30, input_fifo_15_rsci_ccs_ccore_en, ensig_cgo_45, pe_0_0_run_cmp_ccs_ccore_en,
      ensig_cgo_46, accum_fifo_0_run_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo_iro_1;
  input ensig_cgo_iro_30;
  input ensig_cgo_iro_45;
  input ensig_cgo_iro_46;
  input run_wen;
  input ensig_cgo;
  output accum_fifo_15_rsci_ccs_ccore_en;
  input ensig_cgo_1;
  output output_fifo_0_rsci_ccs_ccore_en;
  input ensig_cgo_30;
  output input_fifo_15_rsci_ccs_ccore_en;
  input ensig_cgo_45;
  output pe_0_0_run_cmp_ccs_ccore_en;
  input ensig_cgo_46;
  output accum_fifo_0_run_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign accum_fifo_15_rsci_ccs_ccore_en = run_wen & (ensig_cgo | ensig_cgo_iro);
  assign output_fifo_0_rsci_ccs_ccore_en = run_wen & (ensig_cgo_1 | ensig_cgo_iro_1);
  assign input_fifo_15_rsci_ccs_ccore_en = run_wen & (ensig_cgo_30 | ensig_cgo_iro_30);
  assign pe_0_0_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_45 | ensig_cgo_iro_45);
  assign accum_fifo_0_run_cmp_ccs_ccore_en = run_wen & (ensig_cgo_46 | ensig_cgo_iro_46);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CGHpart
// ------------------------------------------------------------------


module CGHpart (
  CGHpart_isig
);
  input CGHpart_isig;



  // Interconnect Declarations for Component Instantiations 
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_15_i_web_d, accumulation_buffer_rsc_0_15_i_addr_d,
      accumulation_buffer_rsc_0_15_i_dout_d, accumulation_buffer_rsc_0_15_i_addr_d_run,
      accumulation_buffer_rsc_0_15_i_dout_d_mxwt, accumulation_buffer_rsc_0_15_i_biwt,
      accumulation_buffer_rsc_0_15_i_bdwt, accumulation_buffer_rsc_0_15_i_web_d_run_sct,
      accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_15_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_15_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_15_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_15_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_15_i_biwt;
  input accumulation_buffer_rsc_0_15_i_bdwt;
  input accumulation_buffer_rsc_0_15_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_15_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_15_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_15_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_15_i_dout_d,
      accumulation_buffer_rsc_0_15_i_dout_d_bfwt, accumulation_buffer_rsc_0_15_i_bcwt);
  assign accumulation_buffer_rsc_0_15_i_web_d = ~ accumulation_buffer_rsc_0_15_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_15_i_addr_d = {(~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_15_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_15_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_15_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_15_i_bcwt <= ~((~(accumulation_buffer_rsc_0_15_i_bcwt
          | accumulation_buffer_rsc_0_15_i_biwt)) | accumulation_buffer_rsc_0_15_i_bdwt);
      accumulation_buffer_rsc_0_15_i_dout_d_bfwt <= accumulation_buffer_rsc_0_15_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_15_i_oswt, accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_15_i_biwt, accumulation_buffer_rsc_0_15_i_bdwt, accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_15_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_15_i_oswt_pff, accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_15_i_oswt;
  input accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_15_i_biwt;
  output accumulation_buffer_rsc_0_15_i_bdwt;
  output accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_15_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_15_i_oswt_pff;
  output accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_15_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_15_i_bdwt = accumulation_buffer_rsc_0_15_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_15_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_15_i_oswt;
  assign accumulation_buffer_rsc_0_15_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_15_i_dswt_pff;
  assign accumulation_buffer_rsc_0_15_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_15_i_oswt_pff;
  assign accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_15_i_dswt_pff;
  assign accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_15_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_14_i_web_d, accumulation_buffer_rsc_0_14_i_addr_d,
      accumulation_buffer_rsc_0_14_i_dout_d, accumulation_buffer_rsc_0_14_i_addr_d_run,
      accumulation_buffer_rsc_0_14_i_dout_d_mxwt, accumulation_buffer_rsc_0_14_i_biwt,
      accumulation_buffer_rsc_0_14_i_bdwt, accumulation_buffer_rsc_0_14_i_web_d_run_sct,
      accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_14_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_14_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_14_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_14_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_14_i_biwt;
  input accumulation_buffer_rsc_0_14_i_bdwt;
  input accumulation_buffer_rsc_0_14_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_14_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_14_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_14_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_14_i_dout_d,
      accumulation_buffer_rsc_0_14_i_dout_d_bfwt, accumulation_buffer_rsc_0_14_i_bcwt);
  assign accumulation_buffer_rsc_0_14_i_web_d = ~ accumulation_buffer_rsc_0_14_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_14_i_addr_d = {(~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_14_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_14_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_14_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_14_i_bcwt <= ~((~(accumulation_buffer_rsc_0_14_i_bcwt
          | accumulation_buffer_rsc_0_14_i_biwt)) | accumulation_buffer_rsc_0_14_i_bdwt);
      accumulation_buffer_rsc_0_14_i_dout_d_bfwt <= accumulation_buffer_rsc_0_14_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_14_i_oswt, accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_14_i_biwt, accumulation_buffer_rsc_0_14_i_bdwt, accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_14_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_14_i_oswt_pff, accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_14_i_oswt;
  input accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_14_i_biwt;
  output accumulation_buffer_rsc_0_14_i_bdwt;
  output accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_14_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_14_i_oswt_pff;
  output accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_14_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_14_i_bdwt = accumulation_buffer_rsc_0_14_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_14_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_14_i_oswt;
  assign accumulation_buffer_rsc_0_14_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_14_i_dswt_pff;
  assign accumulation_buffer_rsc_0_14_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_14_i_oswt_pff;
  assign accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_14_i_dswt_pff;
  assign accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_14_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_13_i_web_d, accumulation_buffer_rsc_0_13_i_addr_d,
      accumulation_buffer_rsc_0_13_i_dout_d, accumulation_buffer_rsc_0_13_i_addr_d_run,
      accumulation_buffer_rsc_0_13_i_dout_d_mxwt, accumulation_buffer_rsc_0_13_i_biwt,
      accumulation_buffer_rsc_0_13_i_bdwt, accumulation_buffer_rsc_0_13_i_web_d_run_sct,
      accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_13_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_13_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_13_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_13_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_13_i_biwt;
  input accumulation_buffer_rsc_0_13_i_bdwt;
  input accumulation_buffer_rsc_0_13_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_13_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_13_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_13_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_13_i_dout_d,
      accumulation_buffer_rsc_0_13_i_dout_d_bfwt, accumulation_buffer_rsc_0_13_i_bcwt);
  assign accumulation_buffer_rsc_0_13_i_web_d = ~ accumulation_buffer_rsc_0_13_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_13_i_addr_d = {(~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_13_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_13_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_13_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_13_i_bcwt <= ~((~(accumulation_buffer_rsc_0_13_i_bcwt
          | accumulation_buffer_rsc_0_13_i_biwt)) | accumulation_buffer_rsc_0_13_i_bdwt);
      accumulation_buffer_rsc_0_13_i_dout_d_bfwt <= accumulation_buffer_rsc_0_13_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_13_i_oswt, accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_13_i_biwt, accumulation_buffer_rsc_0_13_i_bdwt, accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_13_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_13_i_oswt_pff, accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_13_i_oswt;
  input accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_13_i_biwt;
  output accumulation_buffer_rsc_0_13_i_bdwt;
  output accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_13_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_13_i_oswt_pff;
  output accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_13_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_13_i_bdwt = accumulation_buffer_rsc_0_13_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_13_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_13_i_oswt;
  assign accumulation_buffer_rsc_0_13_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_13_i_dswt_pff;
  assign accumulation_buffer_rsc_0_13_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_13_i_oswt_pff;
  assign accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_13_i_dswt_pff;
  assign accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_13_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_12_i_web_d, accumulation_buffer_rsc_0_12_i_addr_d,
      accumulation_buffer_rsc_0_12_i_dout_d, accumulation_buffer_rsc_0_12_i_addr_d_run,
      accumulation_buffer_rsc_0_12_i_dout_d_mxwt, accumulation_buffer_rsc_0_12_i_biwt,
      accumulation_buffer_rsc_0_12_i_bdwt, accumulation_buffer_rsc_0_12_i_web_d_run_sct,
      accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_12_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_12_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_12_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_12_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_12_i_biwt;
  input accumulation_buffer_rsc_0_12_i_bdwt;
  input accumulation_buffer_rsc_0_12_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_12_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_12_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_12_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_12_i_dout_d,
      accumulation_buffer_rsc_0_12_i_dout_d_bfwt, accumulation_buffer_rsc_0_12_i_bcwt);
  assign accumulation_buffer_rsc_0_12_i_web_d = ~ accumulation_buffer_rsc_0_12_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_12_i_addr_d = {(~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_12_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_12_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_12_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_12_i_bcwt <= ~((~(accumulation_buffer_rsc_0_12_i_bcwt
          | accumulation_buffer_rsc_0_12_i_biwt)) | accumulation_buffer_rsc_0_12_i_bdwt);
      accumulation_buffer_rsc_0_12_i_dout_d_bfwt <= accumulation_buffer_rsc_0_12_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_12_i_oswt, accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_12_i_biwt, accumulation_buffer_rsc_0_12_i_bdwt, accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_12_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_12_i_oswt_pff, accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_12_i_oswt;
  input accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_12_i_biwt;
  output accumulation_buffer_rsc_0_12_i_bdwt;
  output accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_12_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_12_i_oswt_pff;
  output accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_12_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_12_i_bdwt = accumulation_buffer_rsc_0_12_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_12_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_12_i_oswt;
  assign accumulation_buffer_rsc_0_12_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_12_i_dswt_pff;
  assign accumulation_buffer_rsc_0_12_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_12_i_oswt_pff;
  assign accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_12_i_dswt_pff;
  assign accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_12_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_11_i_web_d, accumulation_buffer_rsc_0_11_i_addr_d,
      accumulation_buffer_rsc_0_11_i_dout_d, accumulation_buffer_rsc_0_11_i_addr_d_run,
      accumulation_buffer_rsc_0_11_i_dout_d_mxwt, accumulation_buffer_rsc_0_11_i_biwt,
      accumulation_buffer_rsc_0_11_i_bdwt, accumulation_buffer_rsc_0_11_i_web_d_run_sct,
      accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_11_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_11_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_11_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_11_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_11_i_biwt;
  input accumulation_buffer_rsc_0_11_i_bdwt;
  input accumulation_buffer_rsc_0_11_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_11_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_11_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_11_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_11_i_dout_d,
      accumulation_buffer_rsc_0_11_i_dout_d_bfwt, accumulation_buffer_rsc_0_11_i_bcwt);
  assign accumulation_buffer_rsc_0_11_i_web_d = ~ accumulation_buffer_rsc_0_11_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_11_i_addr_d = {(~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_11_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_11_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_11_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_11_i_bcwt <= ~((~(accumulation_buffer_rsc_0_11_i_bcwt
          | accumulation_buffer_rsc_0_11_i_biwt)) | accumulation_buffer_rsc_0_11_i_bdwt);
      accumulation_buffer_rsc_0_11_i_dout_d_bfwt <= accumulation_buffer_rsc_0_11_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_11_i_oswt, accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_11_i_biwt, accumulation_buffer_rsc_0_11_i_bdwt, accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_11_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_11_i_oswt_pff, accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_11_i_oswt;
  input accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_11_i_biwt;
  output accumulation_buffer_rsc_0_11_i_bdwt;
  output accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_11_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_11_i_oswt_pff;
  output accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_11_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_11_i_bdwt = accumulation_buffer_rsc_0_11_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_11_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_11_i_oswt;
  assign accumulation_buffer_rsc_0_11_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_11_i_dswt_pff;
  assign accumulation_buffer_rsc_0_11_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_11_i_oswt_pff;
  assign accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_11_i_dswt_pff;
  assign accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_11_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_10_i_web_d, accumulation_buffer_rsc_0_10_i_addr_d,
      accumulation_buffer_rsc_0_10_i_dout_d, accumulation_buffer_rsc_0_10_i_addr_d_run,
      accumulation_buffer_rsc_0_10_i_dout_d_mxwt, accumulation_buffer_rsc_0_10_i_biwt,
      accumulation_buffer_rsc_0_10_i_bdwt, accumulation_buffer_rsc_0_10_i_web_d_run_sct,
      accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_10_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_10_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_10_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_10_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_10_i_biwt;
  input accumulation_buffer_rsc_0_10_i_bdwt;
  input accumulation_buffer_rsc_0_10_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_10_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_10_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_10_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_10_i_dout_d,
      accumulation_buffer_rsc_0_10_i_dout_d_bfwt, accumulation_buffer_rsc_0_10_i_bcwt);
  assign accumulation_buffer_rsc_0_10_i_web_d = ~ accumulation_buffer_rsc_0_10_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_10_i_addr_d = {(~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_10_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_10_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_10_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_10_i_bcwt <= ~((~(accumulation_buffer_rsc_0_10_i_bcwt
          | accumulation_buffer_rsc_0_10_i_biwt)) | accumulation_buffer_rsc_0_10_i_bdwt);
      accumulation_buffer_rsc_0_10_i_dout_d_bfwt <= accumulation_buffer_rsc_0_10_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_10_i_oswt, accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_10_i_biwt, accumulation_buffer_rsc_0_10_i_bdwt, accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_10_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_10_i_oswt_pff, accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_10_i_oswt;
  input accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_10_i_biwt;
  output accumulation_buffer_rsc_0_10_i_bdwt;
  output accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_10_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_10_i_oswt_pff;
  output accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_10_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_10_i_bdwt = accumulation_buffer_rsc_0_10_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_10_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_10_i_oswt;
  assign accumulation_buffer_rsc_0_10_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_10_i_dswt_pff;
  assign accumulation_buffer_rsc_0_10_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_10_i_oswt_pff;
  assign accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_10_i_dswt_pff;
  assign accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_10_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_9_i_web_d, accumulation_buffer_rsc_0_9_i_addr_d,
      accumulation_buffer_rsc_0_9_i_dout_d, accumulation_buffer_rsc_0_9_i_addr_d_run,
      accumulation_buffer_rsc_0_9_i_dout_d_mxwt, accumulation_buffer_rsc_0_9_i_biwt,
      accumulation_buffer_rsc_0_9_i_bdwt, accumulation_buffer_rsc_0_9_i_web_d_run_sct,
      accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_9_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_9_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_9_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_9_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_9_i_biwt;
  input accumulation_buffer_rsc_0_9_i_bdwt;
  input accumulation_buffer_rsc_0_9_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_9_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_9_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_9_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_9_i_dout_d,
      accumulation_buffer_rsc_0_9_i_dout_d_bfwt, accumulation_buffer_rsc_0_9_i_bcwt);
  assign accumulation_buffer_rsc_0_9_i_web_d = ~ accumulation_buffer_rsc_0_9_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_9_i_addr_d = {(~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_9_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_9_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_9_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_9_i_bcwt <= ~((~(accumulation_buffer_rsc_0_9_i_bcwt
          | accumulation_buffer_rsc_0_9_i_biwt)) | accumulation_buffer_rsc_0_9_i_bdwt);
      accumulation_buffer_rsc_0_9_i_dout_d_bfwt <= accumulation_buffer_rsc_0_9_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_9_i_oswt, accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_9_i_biwt, accumulation_buffer_rsc_0_9_i_bdwt, accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_9_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_9_i_oswt_pff, accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_9_i_oswt;
  input accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_9_i_biwt;
  output accumulation_buffer_rsc_0_9_i_bdwt;
  output accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_9_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_9_i_oswt_pff;
  output accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_9_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_9_i_bdwt = accumulation_buffer_rsc_0_9_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_9_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_9_i_oswt;
  assign accumulation_buffer_rsc_0_9_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_9_i_dswt_pff;
  assign accumulation_buffer_rsc_0_9_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_9_i_oswt_pff;
  assign accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_9_i_dswt_pff;
  assign accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_9_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_8_i_web_d, accumulation_buffer_rsc_0_8_i_addr_d,
      accumulation_buffer_rsc_0_8_i_dout_d, accumulation_buffer_rsc_0_8_i_addr_d_run,
      accumulation_buffer_rsc_0_8_i_dout_d_mxwt, accumulation_buffer_rsc_0_8_i_biwt,
      accumulation_buffer_rsc_0_8_i_bdwt, accumulation_buffer_rsc_0_8_i_web_d_run_sct,
      accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_8_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_8_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_8_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_8_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_8_i_biwt;
  input accumulation_buffer_rsc_0_8_i_bdwt;
  input accumulation_buffer_rsc_0_8_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_8_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_8_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_8_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_8_i_dout_d,
      accumulation_buffer_rsc_0_8_i_dout_d_bfwt, accumulation_buffer_rsc_0_8_i_bcwt);
  assign accumulation_buffer_rsc_0_8_i_web_d = ~ accumulation_buffer_rsc_0_8_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_8_i_addr_d = {(~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_8_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_8_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_8_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_8_i_bcwt <= ~((~(accumulation_buffer_rsc_0_8_i_bcwt
          | accumulation_buffer_rsc_0_8_i_biwt)) | accumulation_buffer_rsc_0_8_i_bdwt);
      accumulation_buffer_rsc_0_8_i_dout_d_bfwt <= accumulation_buffer_rsc_0_8_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_8_i_oswt, accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_8_i_biwt, accumulation_buffer_rsc_0_8_i_bdwt, accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_8_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_8_i_oswt_pff, accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_8_i_oswt;
  input accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_8_i_biwt;
  output accumulation_buffer_rsc_0_8_i_bdwt;
  output accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_8_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_8_i_oswt_pff;
  output accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_8_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_8_i_bdwt = accumulation_buffer_rsc_0_8_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_8_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_8_i_oswt;
  assign accumulation_buffer_rsc_0_8_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_8_i_dswt_pff;
  assign accumulation_buffer_rsc_0_8_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_8_i_oswt_pff;
  assign accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_8_i_dswt_pff;
  assign accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_8_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_7_i_web_d, accumulation_buffer_rsc_0_7_i_addr_d,
      accumulation_buffer_rsc_0_7_i_dout_d, accumulation_buffer_rsc_0_7_i_addr_d_run,
      accumulation_buffer_rsc_0_7_i_dout_d_mxwt, accumulation_buffer_rsc_0_7_i_biwt,
      accumulation_buffer_rsc_0_7_i_bdwt, accumulation_buffer_rsc_0_7_i_web_d_run_sct,
      accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_7_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_7_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_7_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_7_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_7_i_biwt;
  input accumulation_buffer_rsc_0_7_i_bdwt;
  input accumulation_buffer_rsc_0_7_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_7_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_7_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_7_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_7_i_dout_d,
      accumulation_buffer_rsc_0_7_i_dout_d_bfwt, accumulation_buffer_rsc_0_7_i_bcwt);
  assign accumulation_buffer_rsc_0_7_i_web_d = ~ accumulation_buffer_rsc_0_7_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_7_i_addr_d = {(~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_7_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_7_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_7_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_7_i_bcwt <= ~((~(accumulation_buffer_rsc_0_7_i_bcwt
          | accumulation_buffer_rsc_0_7_i_biwt)) | accumulation_buffer_rsc_0_7_i_bdwt);
      accumulation_buffer_rsc_0_7_i_dout_d_bfwt <= accumulation_buffer_rsc_0_7_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_7_i_oswt, accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_7_i_biwt, accumulation_buffer_rsc_0_7_i_bdwt, accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_7_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_7_i_oswt_pff, accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_7_i_oswt;
  input accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_7_i_biwt;
  output accumulation_buffer_rsc_0_7_i_bdwt;
  output accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_7_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_7_i_oswt_pff;
  output accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_7_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_7_i_bdwt = accumulation_buffer_rsc_0_7_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_7_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_7_i_oswt;
  assign accumulation_buffer_rsc_0_7_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_7_i_dswt_pff;
  assign accumulation_buffer_rsc_0_7_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_7_i_oswt_pff;
  assign accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_7_i_dswt_pff;
  assign accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_7_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_6_i_web_d, accumulation_buffer_rsc_0_6_i_addr_d,
      accumulation_buffer_rsc_0_6_i_dout_d, accumulation_buffer_rsc_0_6_i_addr_d_run,
      accumulation_buffer_rsc_0_6_i_dout_d_mxwt, accumulation_buffer_rsc_0_6_i_biwt,
      accumulation_buffer_rsc_0_6_i_bdwt, accumulation_buffer_rsc_0_6_i_web_d_run_sct,
      accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_6_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_6_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_6_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_6_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_6_i_biwt;
  input accumulation_buffer_rsc_0_6_i_bdwt;
  input accumulation_buffer_rsc_0_6_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_6_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_6_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_6_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_6_i_dout_d,
      accumulation_buffer_rsc_0_6_i_dout_d_bfwt, accumulation_buffer_rsc_0_6_i_bcwt);
  assign accumulation_buffer_rsc_0_6_i_web_d = ~ accumulation_buffer_rsc_0_6_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_6_i_addr_d = {(~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_6_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_6_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_6_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_6_i_bcwt <= ~((~(accumulation_buffer_rsc_0_6_i_bcwt
          | accumulation_buffer_rsc_0_6_i_biwt)) | accumulation_buffer_rsc_0_6_i_bdwt);
      accumulation_buffer_rsc_0_6_i_dout_d_bfwt <= accumulation_buffer_rsc_0_6_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_6_i_oswt, accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_6_i_biwt, accumulation_buffer_rsc_0_6_i_bdwt, accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_6_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_6_i_oswt_pff, accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_6_i_oswt;
  input accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_6_i_biwt;
  output accumulation_buffer_rsc_0_6_i_bdwt;
  output accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_6_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_6_i_oswt_pff;
  output accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_6_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_6_i_bdwt = accumulation_buffer_rsc_0_6_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_6_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_6_i_oswt;
  assign accumulation_buffer_rsc_0_6_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_6_i_dswt_pff;
  assign accumulation_buffer_rsc_0_6_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_6_i_oswt_pff;
  assign accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_6_i_dswt_pff;
  assign accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_6_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_5_i_web_d, accumulation_buffer_rsc_0_5_i_addr_d,
      accumulation_buffer_rsc_0_5_i_dout_d, accumulation_buffer_rsc_0_5_i_addr_d_run,
      accumulation_buffer_rsc_0_5_i_dout_d_mxwt, accumulation_buffer_rsc_0_5_i_biwt,
      accumulation_buffer_rsc_0_5_i_bdwt, accumulation_buffer_rsc_0_5_i_web_d_run_sct,
      accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_5_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_5_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_5_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_5_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_5_i_biwt;
  input accumulation_buffer_rsc_0_5_i_bdwt;
  input accumulation_buffer_rsc_0_5_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_5_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_5_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_5_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_5_i_dout_d,
      accumulation_buffer_rsc_0_5_i_dout_d_bfwt, accumulation_buffer_rsc_0_5_i_bcwt);
  assign accumulation_buffer_rsc_0_5_i_web_d = ~ accumulation_buffer_rsc_0_5_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_5_i_addr_d = {(~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_5_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_5_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_5_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_5_i_bcwt <= ~((~(accumulation_buffer_rsc_0_5_i_bcwt
          | accumulation_buffer_rsc_0_5_i_biwt)) | accumulation_buffer_rsc_0_5_i_bdwt);
      accumulation_buffer_rsc_0_5_i_dout_d_bfwt <= accumulation_buffer_rsc_0_5_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_5_i_oswt, accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_5_i_biwt, accumulation_buffer_rsc_0_5_i_bdwt, accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_5_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_5_i_oswt_pff, accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_5_i_oswt;
  input accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_5_i_biwt;
  output accumulation_buffer_rsc_0_5_i_bdwt;
  output accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_5_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_5_i_oswt_pff;
  output accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_5_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_5_i_bdwt = accumulation_buffer_rsc_0_5_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_5_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_5_i_oswt;
  assign accumulation_buffer_rsc_0_5_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_5_i_dswt_pff;
  assign accumulation_buffer_rsc_0_5_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_5_i_oswt_pff;
  assign accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_5_i_dswt_pff;
  assign accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_5_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_4_i_web_d, accumulation_buffer_rsc_0_4_i_addr_d,
      accumulation_buffer_rsc_0_4_i_dout_d, accumulation_buffer_rsc_0_4_i_addr_d_run,
      accumulation_buffer_rsc_0_4_i_dout_d_mxwt, accumulation_buffer_rsc_0_4_i_biwt,
      accumulation_buffer_rsc_0_4_i_bdwt, accumulation_buffer_rsc_0_4_i_web_d_run_sct,
      accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_4_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_4_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_4_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_4_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_4_i_biwt;
  input accumulation_buffer_rsc_0_4_i_bdwt;
  input accumulation_buffer_rsc_0_4_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_4_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_4_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_4_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_4_i_dout_d,
      accumulation_buffer_rsc_0_4_i_dout_d_bfwt, accumulation_buffer_rsc_0_4_i_bcwt);
  assign accumulation_buffer_rsc_0_4_i_web_d = ~ accumulation_buffer_rsc_0_4_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_4_i_addr_d = {(~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_4_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_4_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_4_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_4_i_bcwt <= ~((~(accumulation_buffer_rsc_0_4_i_bcwt
          | accumulation_buffer_rsc_0_4_i_biwt)) | accumulation_buffer_rsc_0_4_i_bdwt);
      accumulation_buffer_rsc_0_4_i_dout_d_bfwt <= accumulation_buffer_rsc_0_4_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_4_i_oswt, accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_4_i_biwt, accumulation_buffer_rsc_0_4_i_bdwt, accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_4_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_4_i_oswt_pff, accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_4_i_oswt;
  input accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_4_i_biwt;
  output accumulation_buffer_rsc_0_4_i_bdwt;
  output accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_4_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_4_i_oswt_pff;
  output accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_4_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_4_i_bdwt = accumulation_buffer_rsc_0_4_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_4_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_4_i_oswt;
  assign accumulation_buffer_rsc_0_4_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_4_i_dswt_pff;
  assign accumulation_buffer_rsc_0_4_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_4_i_oswt_pff;
  assign accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_4_i_dswt_pff;
  assign accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_4_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_3_i_web_d, accumulation_buffer_rsc_0_3_i_addr_d,
      accumulation_buffer_rsc_0_3_i_dout_d, accumulation_buffer_rsc_0_3_i_addr_d_run,
      accumulation_buffer_rsc_0_3_i_dout_d_mxwt, accumulation_buffer_rsc_0_3_i_biwt,
      accumulation_buffer_rsc_0_3_i_bdwt, accumulation_buffer_rsc_0_3_i_web_d_run_sct,
      accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_3_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_3_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_3_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_3_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_3_i_biwt;
  input accumulation_buffer_rsc_0_3_i_bdwt;
  input accumulation_buffer_rsc_0_3_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_3_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_3_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_3_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_3_i_dout_d,
      accumulation_buffer_rsc_0_3_i_dout_d_bfwt, accumulation_buffer_rsc_0_3_i_bcwt);
  assign accumulation_buffer_rsc_0_3_i_web_d = ~ accumulation_buffer_rsc_0_3_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_3_i_addr_d = {(~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_3_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_3_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_3_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_3_i_bcwt <= ~((~(accumulation_buffer_rsc_0_3_i_bcwt
          | accumulation_buffer_rsc_0_3_i_biwt)) | accumulation_buffer_rsc_0_3_i_bdwt);
      accumulation_buffer_rsc_0_3_i_dout_d_bfwt <= accumulation_buffer_rsc_0_3_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_3_i_oswt, accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_3_i_biwt, accumulation_buffer_rsc_0_3_i_bdwt, accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_3_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_3_i_oswt_pff, accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_3_i_oswt;
  input accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_3_i_biwt;
  output accumulation_buffer_rsc_0_3_i_bdwt;
  output accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_3_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_3_i_oswt_pff;
  output accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_3_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_3_i_bdwt = accumulation_buffer_rsc_0_3_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_3_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_3_i_oswt;
  assign accumulation_buffer_rsc_0_3_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_3_i_dswt_pff;
  assign accumulation_buffer_rsc_0_3_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_3_i_oswt_pff;
  assign accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_3_i_dswt_pff;
  assign accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_3_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_2_i_web_d, accumulation_buffer_rsc_0_2_i_addr_d,
      accumulation_buffer_rsc_0_2_i_dout_d, accumulation_buffer_rsc_0_2_i_addr_d_run,
      accumulation_buffer_rsc_0_2_i_dout_d_mxwt, accumulation_buffer_rsc_0_2_i_biwt,
      accumulation_buffer_rsc_0_2_i_bdwt, accumulation_buffer_rsc_0_2_i_web_d_run_sct,
      accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_2_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_2_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_2_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_2_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_2_i_biwt;
  input accumulation_buffer_rsc_0_2_i_bdwt;
  input accumulation_buffer_rsc_0_2_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_2_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_2_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_2_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_2_i_dout_d,
      accumulation_buffer_rsc_0_2_i_dout_d_bfwt, accumulation_buffer_rsc_0_2_i_bcwt);
  assign accumulation_buffer_rsc_0_2_i_web_d = ~ accumulation_buffer_rsc_0_2_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_2_i_addr_d = {(~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_2_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_2_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_2_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_2_i_bcwt <= ~((~(accumulation_buffer_rsc_0_2_i_bcwt
          | accumulation_buffer_rsc_0_2_i_biwt)) | accumulation_buffer_rsc_0_2_i_bdwt);
      accumulation_buffer_rsc_0_2_i_dout_d_bfwt <= accumulation_buffer_rsc_0_2_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_2_i_oswt, accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_2_i_biwt, accumulation_buffer_rsc_0_2_i_bdwt, accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_2_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_2_i_oswt_pff, accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_2_i_oswt;
  input accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_2_i_biwt;
  output accumulation_buffer_rsc_0_2_i_bdwt;
  output accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_2_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_2_i_oswt_pff;
  output accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_2_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_2_i_bdwt = accumulation_buffer_rsc_0_2_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_2_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_2_i_oswt;
  assign accumulation_buffer_rsc_0_2_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_2_i_dswt_pff;
  assign accumulation_buffer_rsc_0_2_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_2_i_oswt_pff;
  assign accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_2_i_dswt_pff;
  assign accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_2_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_1_i_web_d, accumulation_buffer_rsc_0_1_i_addr_d,
      accumulation_buffer_rsc_0_1_i_dout_d, accumulation_buffer_rsc_0_1_i_addr_d_run,
      accumulation_buffer_rsc_0_1_i_dout_d_mxwt, accumulation_buffer_rsc_0_1_i_biwt,
      accumulation_buffer_rsc_0_1_i_bdwt, accumulation_buffer_rsc_0_1_i_web_d_run_sct,
      accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_1_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_1_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_1_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_1_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_1_i_biwt;
  input accumulation_buffer_rsc_0_1_i_bdwt;
  input accumulation_buffer_rsc_0_1_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_1_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_1_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_1_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_1_i_dout_d,
      accumulation_buffer_rsc_0_1_i_dout_d_bfwt, accumulation_buffer_rsc_0_1_i_bcwt);
  assign accumulation_buffer_rsc_0_1_i_web_d = ~ accumulation_buffer_rsc_0_1_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_1_i_addr_d = {(~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_1_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_1_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_1_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_1_i_bcwt <= ~((~(accumulation_buffer_rsc_0_1_i_bcwt
          | accumulation_buffer_rsc_0_1_i_biwt)) | accumulation_buffer_rsc_0_1_i_bdwt);
      accumulation_buffer_rsc_0_1_i_dout_d_bfwt <= accumulation_buffer_rsc_0_1_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_1_i_oswt, accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_1_i_biwt, accumulation_buffer_rsc_0_1_i_bdwt, accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_1_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_1_i_oswt_pff, accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_1_i_oswt;
  input accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_1_i_biwt;
  output accumulation_buffer_rsc_0_1_i_bdwt;
  output accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_1_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_1_i_oswt_pff;
  output accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_1_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_1_i_bdwt = accumulation_buffer_rsc_0_1_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_1_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_1_i_oswt;
  assign accumulation_buffer_rsc_0_1_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_1_i_dswt_pff;
  assign accumulation_buffer_rsc_0_1_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_1_i_oswt_pff;
  assign accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_1_i_dswt_pff;
  assign accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_1_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_0_i_web_d, accumulation_buffer_rsc_0_0_i_addr_d,
      accumulation_buffer_rsc_0_0_i_dout_d, accumulation_buffer_rsc_0_0_i_addr_d_run,
      accumulation_buffer_rsc_0_0_i_dout_d_mxwt, accumulation_buffer_rsc_0_0_i_biwt,
      accumulation_buffer_rsc_0_0_i_bdwt, accumulation_buffer_rsc_0_0_i_web_d_run_sct,
      accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_0_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_0_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_dout_d;
  input [11:0] accumulation_buffer_rsc_0_0_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_0_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_0_i_biwt;
  input accumulation_buffer_rsc_0_0_i_bdwt;
  input accumulation_buffer_rsc_0_0_i_web_d_run_sct;
  input accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_0_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_0_i_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_0_i_dout_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_0_i_dout_d,
      accumulation_buffer_rsc_0_0_i_dout_d_bfwt, accumulation_buffer_rsc_0_0_i_bcwt);
  assign accumulation_buffer_rsc_0_0_i_web_d = ~ accumulation_buffer_rsc_0_0_i_web_d_run_sct;
  assign accumulation_buffer_rsc_0_0_i_addr_d = {(~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff) , (~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff) , (accumulation_buffer_rsc_0_0_i_addr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_0_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_0_i_dout_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_0_i_bcwt <= ~((~(accumulation_buffer_rsc_0_0_i_bcwt
          | accumulation_buffer_rsc_0_0_i_biwt)) | accumulation_buffer_rsc_0_0_i_bdwt);
      accumulation_buffer_rsc_0_0_i_dout_d_bfwt <= accumulation_buffer_rsc_0_0_i_dout_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_0_i_oswt, accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_0_i_biwt, accumulation_buffer_rsc_0_0_i_bdwt, accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct,
      accumulation_buffer_rsc_0_0_i_web_d_run_sct_pff, accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff,
      accumulation_buffer_rsc_0_0_i_oswt_pff, accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_0_i_oswt;
  input accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  output accumulation_buffer_rsc_0_0_i_biwt;
  output accumulation_buffer_rsc_0_0_i_bdwt;
  output accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  output accumulation_buffer_rsc_0_0_i_web_d_run_sct_pff;
  input accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_0_i_oswt_pff;
  output accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_0_i_dswt_pff;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_0_i_bdwt = accumulation_buffer_rsc_0_0_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_0_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_0_i_oswt;
  assign accumulation_buffer_rsc_0_0_i_web_d_run_sct_pff = accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff
      & accumulation_buffer_rsc_0_0_i_dswt_pff;
  assign accumulation_buffer_rsc_0_0_i_dswt_pff = run_wen & accumulation_buffer_rsc_0_0_i_oswt_pff;
  assign accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff = accumulation_buffer_rsc_0_0_i_dswt_pff;
  assign accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct
      = accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct
      & accumulation_buffer_rsc_0_0_i_dswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
    (
  clk, arst_n, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt,
      loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt, loopIndicesIn_rsci_bcwt,
      loopIndicesIn_rsci_idat
);
  input clk;
  input arst_n;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [47:0] loopIndicesIn_rsci_idat_mxwt;
  input loopIndicesIn_rsci_biwt;
  input loopIndicesIn_rsci_bdwt;
  output loopIndicesIn_rsci_bcwt;
  reg loopIndicesIn_rsci_bcwt;
  input [47:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations
  reg [47:0] loopIndicesIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_wen_comp = (~ loopIndicesIn_rsci_oswt) | loopIndicesIn_rsci_biwt
      | loopIndicesIn_rsci_bcwt;
  assign loopIndicesIn_rsci_idat_mxwt = MUX_v_48_2_2(loopIndicesIn_rsci_idat, loopIndicesIn_rsci_idat_bfwt,
      loopIndicesIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_rsci_bcwt <= 1'b0;
    end
    else begin
      loopIndicesIn_rsci_bcwt <= ~((~(loopIndicesIn_rsci_bcwt | loopIndicesIn_rsci_biwt))
          | loopIndicesIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_rsci_idat_bfwt <= 48'b000000000000000000000000000000000000000000000000;
    end
    else if ( ~ loopIndicesIn_rsci_bcwt ) begin
      loopIndicesIn_rsci_idat_bfwt <= loopIndicesIn_rsci_idat_mxwt;
    end
  end

  function automatic [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
    (
  run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt,
      loopIndicesIn_rsci_bcwt, loopIndicesIn_rsci_irdy_run_sct, loopIndicesIn_rsci_ivld
);
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_biwt;
  output loopIndicesIn_rsci_bdwt;
  input loopIndicesIn_rsci_bcwt;
  output loopIndicesIn_rsci_irdy_run_sct;
  input loopIndicesIn_rsci_ivld;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_bdwt = loopIndicesIn_rsci_oswt & run_wen;
  assign loopIndicesIn_rsci_biwt = loopIndicesIn_rsci_ogwt & loopIndicesIn_rsci_ivld;
  assign loopIndicesIn_rsci_ogwt = loopIndicesIn_rsci_oswt & (~ loopIndicesIn_rsci_bcwt);
  assign loopIndicesIn_rsci_irdy_run_sct = loopIndicesIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
    (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [95:0] paramsIn_rsci_idat_bfwt_127_32;
  wire [95:0] paramsIn_rsci_idat_mxwt_opt_127_32;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_127_32 = MUX_v_96_2_2((paramsIn_rsci_idat[127:32]),
      paramsIn_rsci_idat_bfwt_127_32, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_opt_127_32;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt_127_32 <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt_127_32 <= paramsIn_rsci_idat_mxwt_opt_127_32;
    end
  end

  function automatic [95:0] MUX_v_96_2_2;
    input [95:0] input_0;
    input [95:0] input_1;
    input [0:0] sel;
    reg [95:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_96_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
    (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp
    (
  clk, arst_n, output_rsci_oswt, output_rsci_wen_comp, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_bcwt
);
  input clk;
  input arst_n;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input output_rsci_biwt;
  input output_rsci_bdwt;
  output output_rsci_bcwt;
  reg output_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt | output_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_rsci_bcwt <= 1'b0;
    end
    else begin
      output_rsci_bcwt <= ~((~(output_rsci_bcwt | output_rsci_biwt)) | output_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl
    (
  run_wen, output_rsci_oswt, output_rsci_irdy, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_bcwt, output_rsci_ivld_run_sct
);
  input run_wen;
  input output_rsci_oswt;
  input output_rsci_irdy;
  output output_rsci_biwt;
  output output_rsci_bdwt;
  input output_rsci_bcwt;
  output output_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire output_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_bdwt = output_rsci_oswt & run_wen;
  assign output_rsci_biwt = output_rsci_ogwt & output_rsci_irdy;
  assign output_rsci_ogwt = output_rsci_oswt & (~ output_rsci_bcwt);
  assign output_rsci_ivld_run_sct = output_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp
    (
  clk, arst_n, weight_rsci_oswt, weight_rsci_wen_comp, weight_rsci_idat_mxwt, weight_rsci_biwt,
      weight_rsci_bdwt, weight_rsci_bcwt, weight_rsci_idat
);
  input clk;
  input arst_n;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [127:0] weight_rsci_idat_mxwt;
  input weight_rsci_biwt;
  input weight_rsci_bdwt;
  output weight_rsci_bcwt;
  reg weight_rsci_bcwt;
  input [127:0] weight_rsci_idat;


  // Interconnect Declarations
  reg [127:0] weight_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_wen_comp = (~ weight_rsci_oswt) | weight_rsci_biwt | weight_rsci_bcwt;
  assign weight_rsci_idat_mxwt = MUX_v_128_2_2(weight_rsci_idat, weight_rsci_idat_bfwt,
      weight_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_rsci_bcwt <= 1'b0;
      weight_rsci_idat_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      weight_rsci_bcwt <= ~((~(weight_rsci_bcwt | weight_rsci_biwt)) | weight_rsci_bdwt);
      weight_rsci_idat_bfwt <= weight_rsci_idat_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl
    (
  run_wen, weight_rsci_oswt, weight_rsci_biwt, weight_rsci_bdwt, weight_rsci_bcwt,
      weight_rsci_irdy_run_sct, weight_rsci_ivld
);
  input run_wen;
  input weight_rsci_oswt;
  output weight_rsci_biwt;
  output weight_rsci_bdwt;
  input weight_rsci_bcwt;
  output weight_rsci_irdy_run_sct;
  input weight_rsci_ivld;


  // Interconnect Declarations
  wire weight_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_bdwt = weight_rsci_oswt & run_wen;
  assign weight_rsci_biwt = weight_rsci_ogwt & weight_rsci_ivld;
  assign weight_rsci_ogwt = weight_rsci_oswt & (~ weight_rsci_bcwt);
  assign weight_rsci_irdy_run_sct = weight_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp
    (
  clk, arst_n, input_rsci_oswt, input_rsci_wen_comp, input_rsci_idat_mxwt, input_rsci_biwt,
      input_rsci_bdwt, input_rsci_bcwt, input_rsci_idat
);
  input clk;
  input arst_n;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [127:0] input_rsci_idat_mxwt;
  input input_rsci_biwt;
  input input_rsci_bdwt;
  output input_rsci_bcwt;
  reg input_rsci_bcwt;
  input [127:0] input_rsci_idat;


  // Interconnect Declarations
  reg [127:0] input_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_wen_comp = (~ input_rsci_oswt) | input_rsci_biwt | input_rsci_bcwt;
  assign input_rsci_idat_mxwt = MUX_v_128_2_2(input_rsci_idat, input_rsci_idat_bfwt,
      input_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_rsci_bcwt <= 1'b0;
      input_rsci_idat_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      input_rsci_bcwt <= ~((~(input_rsci_bcwt | input_rsci_biwt)) | input_rsci_bdwt);
      input_rsci_idat_bfwt <= input_rsci_idat_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl
    (
  run_wen, input_rsci_oswt, input_rsci_biwt, input_rsci_bdwt, input_rsci_bcwt, input_rsci_irdy_run_sct,
      input_rsci_ivld
);
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_biwt;
  output input_rsci_bdwt;
  input input_rsci_bcwt;
  output input_rsci_irdy_run_sct;
  input input_rsci_ivld;


  // Interconnect Declarations
  wire input_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_bdwt = input_rsci_oswt & run_wen;
  assign input_rsci_biwt = input_rsci_ogwt & input_rsci_ivld;
  assign input_rsci_ogwt = input_rsci_oswt & (~ input_rsci_bcwt);
  assign input_rsci_irdy_run_sct = input_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_15_i_web_d, accumulation_buffer_rsc_0_15_i_addr_d,
      accumulation_buffer_rsc_0_15_i_dout_d, accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_15_i_oswt, accumulation_buffer_rsc_0_15_i_addr_d_run,
      accumulation_buffer_rsc_0_15_i_dout_d_mxwt, accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_15_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_15_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_15_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_dout_d;
  output accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_15_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_15_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_15_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_15_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_15_i_biwt;
  wire accumulation_buffer_rsc_0_15_i_bdwt;
  wire accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_15_i_web_d_reg;
  wire accumulation_buffer_rsc_0_15_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_15_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_15_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_15_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_15_i_oswt(accumulation_buffer_rsc_0_15_i_oswt),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_15_i_biwt(accumulation_buffer_rsc_0_15_i_biwt),
      .accumulation_buffer_rsc_0_15_i_bdwt(accumulation_buffer_rsc_0_15_i_bdwt),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_15_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_15_i_oswt_pff(accumulation_buffer_rsc_0_15_i_oswt_pff),
      .accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_15_i_web_d(accumulation_buffer_rsc_0_15_i_web_d_reg),
      .accumulation_buffer_rsc_0_15_i_addr_d(accumulation_buffer_rsc_0_15_i_addr_d_reg),
      .accumulation_buffer_rsc_0_15_i_dout_d(accumulation_buffer_rsc_0_15_i_dout_d),
      .accumulation_buffer_rsc_0_15_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_15_i_dout_d_mxwt(accumulation_buffer_rsc_0_15_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_15_i_biwt(accumulation_buffer_rsc_0_15_i_biwt),
      .accumulation_buffer_rsc_0_15_i_bdwt(accumulation_buffer_rsc_0_15_i_bdwt),
      .accumulation_buffer_rsc_0_15_i_web_d_run_sct(accumulation_buffer_rsc_0_15_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_15_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_15_i_web_d = accumulation_buffer_rsc_0_15_i_web_d_reg;
  assign accumulation_buffer_rsc_0_15_i_addr_d = accumulation_buffer_rsc_0_15_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_15_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_14_i_web_d, accumulation_buffer_rsc_0_14_i_addr_d,
      accumulation_buffer_rsc_0_14_i_dout_d, accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_14_i_oswt, accumulation_buffer_rsc_0_14_i_addr_d_run,
      accumulation_buffer_rsc_0_14_i_dout_d_mxwt, accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_14_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_14_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_14_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_dout_d;
  output accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_14_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_14_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_14_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_14_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_14_i_biwt;
  wire accumulation_buffer_rsc_0_14_i_bdwt;
  wire accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_14_i_web_d_reg;
  wire accumulation_buffer_rsc_0_14_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_14_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_14_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_14_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_14_i_oswt(accumulation_buffer_rsc_0_14_i_oswt),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_14_i_biwt(accumulation_buffer_rsc_0_14_i_biwt),
      .accumulation_buffer_rsc_0_14_i_bdwt(accumulation_buffer_rsc_0_14_i_bdwt),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_14_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_14_i_oswt_pff(accumulation_buffer_rsc_0_14_i_oswt_pff),
      .accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_14_i_web_d(accumulation_buffer_rsc_0_14_i_web_d_reg),
      .accumulation_buffer_rsc_0_14_i_addr_d(accumulation_buffer_rsc_0_14_i_addr_d_reg),
      .accumulation_buffer_rsc_0_14_i_dout_d(accumulation_buffer_rsc_0_14_i_dout_d),
      .accumulation_buffer_rsc_0_14_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_14_i_dout_d_mxwt(accumulation_buffer_rsc_0_14_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_14_i_biwt(accumulation_buffer_rsc_0_14_i_biwt),
      .accumulation_buffer_rsc_0_14_i_bdwt(accumulation_buffer_rsc_0_14_i_bdwt),
      .accumulation_buffer_rsc_0_14_i_web_d_run_sct(accumulation_buffer_rsc_0_14_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_14_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_14_i_web_d = accumulation_buffer_rsc_0_14_i_web_d_reg;
  assign accumulation_buffer_rsc_0_14_i_addr_d = accumulation_buffer_rsc_0_14_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_14_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_13_i_web_d, accumulation_buffer_rsc_0_13_i_addr_d,
      accumulation_buffer_rsc_0_13_i_dout_d, accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_13_i_oswt, accumulation_buffer_rsc_0_13_i_addr_d_run,
      accumulation_buffer_rsc_0_13_i_dout_d_mxwt, accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_13_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_13_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_13_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_dout_d;
  output accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_13_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_13_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_13_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_13_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_13_i_biwt;
  wire accumulation_buffer_rsc_0_13_i_bdwt;
  wire accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_13_i_web_d_reg;
  wire accumulation_buffer_rsc_0_13_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_13_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_13_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_13_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_13_i_oswt(accumulation_buffer_rsc_0_13_i_oswt),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_13_i_biwt(accumulation_buffer_rsc_0_13_i_biwt),
      .accumulation_buffer_rsc_0_13_i_bdwt(accumulation_buffer_rsc_0_13_i_bdwt),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_13_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_13_i_oswt_pff(accumulation_buffer_rsc_0_13_i_oswt_pff),
      .accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_13_i_web_d(accumulation_buffer_rsc_0_13_i_web_d_reg),
      .accumulation_buffer_rsc_0_13_i_addr_d(accumulation_buffer_rsc_0_13_i_addr_d_reg),
      .accumulation_buffer_rsc_0_13_i_dout_d(accumulation_buffer_rsc_0_13_i_dout_d),
      .accumulation_buffer_rsc_0_13_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_13_i_dout_d_mxwt(accumulation_buffer_rsc_0_13_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_13_i_biwt(accumulation_buffer_rsc_0_13_i_biwt),
      .accumulation_buffer_rsc_0_13_i_bdwt(accumulation_buffer_rsc_0_13_i_bdwt),
      .accumulation_buffer_rsc_0_13_i_web_d_run_sct(accumulation_buffer_rsc_0_13_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_13_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_13_i_web_d = accumulation_buffer_rsc_0_13_i_web_d_reg;
  assign accumulation_buffer_rsc_0_13_i_addr_d = accumulation_buffer_rsc_0_13_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_13_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_12_i_web_d, accumulation_buffer_rsc_0_12_i_addr_d,
      accumulation_buffer_rsc_0_12_i_dout_d, accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_12_i_oswt, accumulation_buffer_rsc_0_12_i_addr_d_run,
      accumulation_buffer_rsc_0_12_i_dout_d_mxwt, accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_12_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_12_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_12_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_dout_d;
  output accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_12_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_12_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_12_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_12_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_12_i_biwt;
  wire accumulation_buffer_rsc_0_12_i_bdwt;
  wire accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_12_i_web_d_reg;
  wire accumulation_buffer_rsc_0_12_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_12_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_12_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_12_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_12_i_oswt(accumulation_buffer_rsc_0_12_i_oswt),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_12_i_biwt(accumulation_buffer_rsc_0_12_i_biwt),
      .accumulation_buffer_rsc_0_12_i_bdwt(accumulation_buffer_rsc_0_12_i_bdwt),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_12_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_12_i_oswt_pff(accumulation_buffer_rsc_0_12_i_oswt_pff),
      .accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_12_i_web_d(accumulation_buffer_rsc_0_12_i_web_d_reg),
      .accumulation_buffer_rsc_0_12_i_addr_d(accumulation_buffer_rsc_0_12_i_addr_d_reg),
      .accumulation_buffer_rsc_0_12_i_dout_d(accumulation_buffer_rsc_0_12_i_dout_d),
      .accumulation_buffer_rsc_0_12_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_12_i_dout_d_mxwt(accumulation_buffer_rsc_0_12_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_12_i_biwt(accumulation_buffer_rsc_0_12_i_biwt),
      .accumulation_buffer_rsc_0_12_i_bdwt(accumulation_buffer_rsc_0_12_i_bdwt),
      .accumulation_buffer_rsc_0_12_i_web_d_run_sct(accumulation_buffer_rsc_0_12_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_12_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_12_i_web_d = accumulation_buffer_rsc_0_12_i_web_d_reg;
  assign accumulation_buffer_rsc_0_12_i_addr_d = accumulation_buffer_rsc_0_12_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_12_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_11_i_web_d, accumulation_buffer_rsc_0_11_i_addr_d,
      accumulation_buffer_rsc_0_11_i_dout_d, accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_11_i_oswt, accumulation_buffer_rsc_0_11_i_addr_d_run,
      accumulation_buffer_rsc_0_11_i_dout_d_mxwt, accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_11_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_11_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_11_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_dout_d;
  output accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_11_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_11_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_11_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_11_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_11_i_biwt;
  wire accumulation_buffer_rsc_0_11_i_bdwt;
  wire accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_11_i_web_d_reg;
  wire accumulation_buffer_rsc_0_11_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_11_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_11_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_11_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_11_i_oswt(accumulation_buffer_rsc_0_11_i_oswt),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_11_i_biwt(accumulation_buffer_rsc_0_11_i_biwt),
      .accumulation_buffer_rsc_0_11_i_bdwt(accumulation_buffer_rsc_0_11_i_bdwt),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_11_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_11_i_oswt_pff(accumulation_buffer_rsc_0_11_i_oswt_pff),
      .accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_11_i_web_d(accumulation_buffer_rsc_0_11_i_web_d_reg),
      .accumulation_buffer_rsc_0_11_i_addr_d(accumulation_buffer_rsc_0_11_i_addr_d_reg),
      .accumulation_buffer_rsc_0_11_i_dout_d(accumulation_buffer_rsc_0_11_i_dout_d),
      .accumulation_buffer_rsc_0_11_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_11_i_dout_d_mxwt(accumulation_buffer_rsc_0_11_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_11_i_biwt(accumulation_buffer_rsc_0_11_i_biwt),
      .accumulation_buffer_rsc_0_11_i_bdwt(accumulation_buffer_rsc_0_11_i_bdwt),
      .accumulation_buffer_rsc_0_11_i_web_d_run_sct(accumulation_buffer_rsc_0_11_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_11_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_11_i_web_d = accumulation_buffer_rsc_0_11_i_web_d_reg;
  assign accumulation_buffer_rsc_0_11_i_addr_d = accumulation_buffer_rsc_0_11_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_11_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_10_i_web_d, accumulation_buffer_rsc_0_10_i_addr_d,
      accumulation_buffer_rsc_0_10_i_dout_d, accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_10_i_oswt, accumulation_buffer_rsc_0_10_i_addr_d_run,
      accumulation_buffer_rsc_0_10_i_dout_d_mxwt, accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_10_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_10_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_10_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_dout_d;
  output accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_10_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_10_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_10_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_10_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_10_i_biwt;
  wire accumulation_buffer_rsc_0_10_i_bdwt;
  wire accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_10_i_web_d_reg;
  wire accumulation_buffer_rsc_0_10_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_10_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_10_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_10_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_10_i_oswt(accumulation_buffer_rsc_0_10_i_oswt),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_10_i_biwt(accumulation_buffer_rsc_0_10_i_biwt),
      .accumulation_buffer_rsc_0_10_i_bdwt(accumulation_buffer_rsc_0_10_i_bdwt),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_10_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_10_i_oswt_pff(accumulation_buffer_rsc_0_10_i_oswt_pff),
      .accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_10_i_web_d(accumulation_buffer_rsc_0_10_i_web_d_reg),
      .accumulation_buffer_rsc_0_10_i_addr_d(accumulation_buffer_rsc_0_10_i_addr_d_reg),
      .accumulation_buffer_rsc_0_10_i_dout_d(accumulation_buffer_rsc_0_10_i_dout_d),
      .accumulation_buffer_rsc_0_10_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_10_i_dout_d_mxwt(accumulation_buffer_rsc_0_10_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_10_i_biwt(accumulation_buffer_rsc_0_10_i_biwt),
      .accumulation_buffer_rsc_0_10_i_bdwt(accumulation_buffer_rsc_0_10_i_bdwt),
      .accumulation_buffer_rsc_0_10_i_web_d_run_sct(accumulation_buffer_rsc_0_10_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_10_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_10_i_web_d = accumulation_buffer_rsc_0_10_i_web_d_reg;
  assign accumulation_buffer_rsc_0_10_i_addr_d = accumulation_buffer_rsc_0_10_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_10_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_9_i_web_d, accumulation_buffer_rsc_0_9_i_addr_d,
      accumulation_buffer_rsc_0_9_i_dout_d, accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_9_i_oswt, accumulation_buffer_rsc_0_9_i_addr_d_run,
      accumulation_buffer_rsc_0_9_i_dout_d_mxwt, accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_9_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_9_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_9_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_dout_d;
  output accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_9_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_9_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_9_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_9_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_9_i_biwt;
  wire accumulation_buffer_rsc_0_9_i_bdwt;
  wire accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_9_i_web_d_reg;
  wire accumulation_buffer_rsc_0_9_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_9_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_9_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_9_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_9_i_oswt(accumulation_buffer_rsc_0_9_i_oswt),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_9_i_biwt(accumulation_buffer_rsc_0_9_i_biwt),
      .accumulation_buffer_rsc_0_9_i_bdwt(accumulation_buffer_rsc_0_9_i_bdwt),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_9_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_9_i_oswt_pff(accumulation_buffer_rsc_0_9_i_oswt_pff),
      .accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_9_i_web_d(accumulation_buffer_rsc_0_9_i_web_d_reg),
      .accumulation_buffer_rsc_0_9_i_addr_d(accumulation_buffer_rsc_0_9_i_addr_d_reg),
      .accumulation_buffer_rsc_0_9_i_dout_d(accumulation_buffer_rsc_0_9_i_dout_d),
      .accumulation_buffer_rsc_0_9_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_9_i_dout_d_mxwt(accumulation_buffer_rsc_0_9_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_9_i_biwt(accumulation_buffer_rsc_0_9_i_biwt),
      .accumulation_buffer_rsc_0_9_i_bdwt(accumulation_buffer_rsc_0_9_i_bdwt),
      .accumulation_buffer_rsc_0_9_i_web_d_run_sct(accumulation_buffer_rsc_0_9_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_9_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_9_i_web_d = accumulation_buffer_rsc_0_9_i_web_d_reg;
  assign accumulation_buffer_rsc_0_9_i_addr_d = accumulation_buffer_rsc_0_9_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_9_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_8_i_web_d, accumulation_buffer_rsc_0_8_i_addr_d,
      accumulation_buffer_rsc_0_8_i_dout_d, accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_8_i_oswt, accumulation_buffer_rsc_0_8_i_addr_d_run,
      accumulation_buffer_rsc_0_8_i_dout_d_mxwt, accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_8_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_8_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_8_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_dout_d;
  output accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_8_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_8_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_8_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_8_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_8_i_biwt;
  wire accumulation_buffer_rsc_0_8_i_bdwt;
  wire accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_8_i_web_d_reg;
  wire accumulation_buffer_rsc_0_8_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_8_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_8_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_8_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_8_i_oswt(accumulation_buffer_rsc_0_8_i_oswt),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_8_i_biwt(accumulation_buffer_rsc_0_8_i_biwt),
      .accumulation_buffer_rsc_0_8_i_bdwt(accumulation_buffer_rsc_0_8_i_bdwt),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_8_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_8_i_oswt_pff(accumulation_buffer_rsc_0_8_i_oswt_pff),
      .accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_8_i_web_d(accumulation_buffer_rsc_0_8_i_web_d_reg),
      .accumulation_buffer_rsc_0_8_i_addr_d(accumulation_buffer_rsc_0_8_i_addr_d_reg),
      .accumulation_buffer_rsc_0_8_i_dout_d(accumulation_buffer_rsc_0_8_i_dout_d),
      .accumulation_buffer_rsc_0_8_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_8_i_dout_d_mxwt(accumulation_buffer_rsc_0_8_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_8_i_biwt(accumulation_buffer_rsc_0_8_i_biwt),
      .accumulation_buffer_rsc_0_8_i_bdwt(accumulation_buffer_rsc_0_8_i_bdwt),
      .accumulation_buffer_rsc_0_8_i_web_d_run_sct(accumulation_buffer_rsc_0_8_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_8_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_8_i_web_d = accumulation_buffer_rsc_0_8_i_web_d_reg;
  assign accumulation_buffer_rsc_0_8_i_addr_d = accumulation_buffer_rsc_0_8_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_8_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_7_i_web_d, accumulation_buffer_rsc_0_7_i_addr_d,
      accumulation_buffer_rsc_0_7_i_dout_d, accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_7_i_oswt, accumulation_buffer_rsc_0_7_i_addr_d_run,
      accumulation_buffer_rsc_0_7_i_dout_d_mxwt, accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_7_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_7_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_7_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_dout_d;
  output accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_7_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_7_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_7_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_7_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_7_i_biwt;
  wire accumulation_buffer_rsc_0_7_i_bdwt;
  wire accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_7_i_web_d_reg;
  wire accumulation_buffer_rsc_0_7_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_7_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_7_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_7_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_7_i_oswt(accumulation_buffer_rsc_0_7_i_oswt),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_7_i_biwt(accumulation_buffer_rsc_0_7_i_biwt),
      .accumulation_buffer_rsc_0_7_i_bdwt(accumulation_buffer_rsc_0_7_i_bdwt),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_7_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_7_i_oswt_pff(accumulation_buffer_rsc_0_7_i_oswt_pff),
      .accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_7_i_web_d(accumulation_buffer_rsc_0_7_i_web_d_reg),
      .accumulation_buffer_rsc_0_7_i_addr_d(accumulation_buffer_rsc_0_7_i_addr_d_reg),
      .accumulation_buffer_rsc_0_7_i_dout_d(accumulation_buffer_rsc_0_7_i_dout_d),
      .accumulation_buffer_rsc_0_7_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_7_i_dout_d_mxwt(accumulation_buffer_rsc_0_7_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_7_i_biwt(accumulation_buffer_rsc_0_7_i_biwt),
      .accumulation_buffer_rsc_0_7_i_bdwt(accumulation_buffer_rsc_0_7_i_bdwt),
      .accumulation_buffer_rsc_0_7_i_web_d_run_sct(accumulation_buffer_rsc_0_7_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_7_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_7_i_web_d = accumulation_buffer_rsc_0_7_i_web_d_reg;
  assign accumulation_buffer_rsc_0_7_i_addr_d = accumulation_buffer_rsc_0_7_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_7_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_6_i_web_d, accumulation_buffer_rsc_0_6_i_addr_d,
      accumulation_buffer_rsc_0_6_i_dout_d, accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_6_i_oswt, accumulation_buffer_rsc_0_6_i_addr_d_run,
      accumulation_buffer_rsc_0_6_i_dout_d_mxwt, accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_6_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_6_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_6_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_dout_d;
  output accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_6_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_6_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_6_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_6_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_6_i_biwt;
  wire accumulation_buffer_rsc_0_6_i_bdwt;
  wire accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_6_i_web_d_reg;
  wire accumulation_buffer_rsc_0_6_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_6_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_6_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_6_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_6_i_oswt(accumulation_buffer_rsc_0_6_i_oswt),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_6_i_biwt(accumulation_buffer_rsc_0_6_i_biwt),
      .accumulation_buffer_rsc_0_6_i_bdwt(accumulation_buffer_rsc_0_6_i_bdwt),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_6_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_6_i_oswt_pff(accumulation_buffer_rsc_0_6_i_oswt_pff),
      .accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_6_i_web_d(accumulation_buffer_rsc_0_6_i_web_d_reg),
      .accumulation_buffer_rsc_0_6_i_addr_d(accumulation_buffer_rsc_0_6_i_addr_d_reg),
      .accumulation_buffer_rsc_0_6_i_dout_d(accumulation_buffer_rsc_0_6_i_dout_d),
      .accumulation_buffer_rsc_0_6_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_6_i_dout_d_mxwt(accumulation_buffer_rsc_0_6_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_6_i_biwt(accumulation_buffer_rsc_0_6_i_biwt),
      .accumulation_buffer_rsc_0_6_i_bdwt(accumulation_buffer_rsc_0_6_i_bdwt),
      .accumulation_buffer_rsc_0_6_i_web_d_run_sct(accumulation_buffer_rsc_0_6_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_6_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_6_i_web_d = accumulation_buffer_rsc_0_6_i_web_d_reg;
  assign accumulation_buffer_rsc_0_6_i_addr_d = accumulation_buffer_rsc_0_6_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_6_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_5_i_web_d, accumulation_buffer_rsc_0_5_i_addr_d,
      accumulation_buffer_rsc_0_5_i_dout_d, accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_5_i_oswt, accumulation_buffer_rsc_0_5_i_addr_d_run,
      accumulation_buffer_rsc_0_5_i_dout_d_mxwt, accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_5_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_5_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_5_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_dout_d;
  output accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_5_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_5_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_5_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_5_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_5_i_biwt;
  wire accumulation_buffer_rsc_0_5_i_bdwt;
  wire accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_5_i_web_d_reg;
  wire accumulation_buffer_rsc_0_5_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_5_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_5_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_5_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_5_i_oswt(accumulation_buffer_rsc_0_5_i_oswt),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_5_i_biwt(accumulation_buffer_rsc_0_5_i_biwt),
      .accumulation_buffer_rsc_0_5_i_bdwt(accumulation_buffer_rsc_0_5_i_bdwt),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_5_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_5_i_oswt_pff(accumulation_buffer_rsc_0_5_i_oswt_pff),
      .accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_5_i_web_d(accumulation_buffer_rsc_0_5_i_web_d_reg),
      .accumulation_buffer_rsc_0_5_i_addr_d(accumulation_buffer_rsc_0_5_i_addr_d_reg),
      .accumulation_buffer_rsc_0_5_i_dout_d(accumulation_buffer_rsc_0_5_i_dout_d),
      .accumulation_buffer_rsc_0_5_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_5_i_dout_d_mxwt(accumulation_buffer_rsc_0_5_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_5_i_biwt(accumulation_buffer_rsc_0_5_i_biwt),
      .accumulation_buffer_rsc_0_5_i_bdwt(accumulation_buffer_rsc_0_5_i_bdwt),
      .accumulation_buffer_rsc_0_5_i_web_d_run_sct(accumulation_buffer_rsc_0_5_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_5_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_5_i_web_d = accumulation_buffer_rsc_0_5_i_web_d_reg;
  assign accumulation_buffer_rsc_0_5_i_addr_d = accumulation_buffer_rsc_0_5_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_5_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_4_i_web_d, accumulation_buffer_rsc_0_4_i_addr_d,
      accumulation_buffer_rsc_0_4_i_dout_d, accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_4_i_oswt, accumulation_buffer_rsc_0_4_i_addr_d_run,
      accumulation_buffer_rsc_0_4_i_dout_d_mxwt, accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_4_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_4_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_4_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_dout_d;
  output accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_4_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_4_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_4_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_4_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_4_i_biwt;
  wire accumulation_buffer_rsc_0_4_i_bdwt;
  wire accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_4_i_web_d_reg;
  wire accumulation_buffer_rsc_0_4_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_4_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_4_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_4_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_4_i_oswt(accumulation_buffer_rsc_0_4_i_oswt),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_4_i_biwt(accumulation_buffer_rsc_0_4_i_biwt),
      .accumulation_buffer_rsc_0_4_i_bdwt(accumulation_buffer_rsc_0_4_i_bdwt),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_4_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_4_i_oswt_pff(accumulation_buffer_rsc_0_4_i_oswt_pff),
      .accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_4_i_web_d(accumulation_buffer_rsc_0_4_i_web_d_reg),
      .accumulation_buffer_rsc_0_4_i_addr_d(accumulation_buffer_rsc_0_4_i_addr_d_reg),
      .accumulation_buffer_rsc_0_4_i_dout_d(accumulation_buffer_rsc_0_4_i_dout_d),
      .accumulation_buffer_rsc_0_4_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_4_i_dout_d_mxwt(accumulation_buffer_rsc_0_4_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_4_i_biwt(accumulation_buffer_rsc_0_4_i_biwt),
      .accumulation_buffer_rsc_0_4_i_bdwt(accumulation_buffer_rsc_0_4_i_bdwt),
      .accumulation_buffer_rsc_0_4_i_web_d_run_sct(accumulation_buffer_rsc_0_4_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_4_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_4_i_web_d = accumulation_buffer_rsc_0_4_i_web_d_reg;
  assign accumulation_buffer_rsc_0_4_i_addr_d = accumulation_buffer_rsc_0_4_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_4_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_3_i_web_d, accumulation_buffer_rsc_0_3_i_addr_d,
      accumulation_buffer_rsc_0_3_i_dout_d, accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_3_i_oswt, accumulation_buffer_rsc_0_3_i_addr_d_run,
      accumulation_buffer_rsc_0_3_i_dout_d_mxwt, accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_3_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_3_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_3_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_dout_d;
  output accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_3_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_3_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_3_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_3_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_3_i_biwt;
  wire accumulation_buffer_rsc_0_3_i_bdwt;
  wire accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_3_i_web_d_reg;
  wire accumulation_buffer_rsc_0_3_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_3_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_3_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_3_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_3_i_oswt(accumulation_buffer_rsc_0_3_i_oswt),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_3_i_biwt(accumulation_buffer_rsc_0_3_i_biwt),
      .accumulation_buffer_rsc_0_3_i_bdwt(accumulation_buffer_rsc_0_3_i_bdwt),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_3_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_3_i_oswt_pff(accumulation_buffer_rsc_0_3_i_oswt_pff),
      .accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_3_i_web_d(accumulation_buffer_rsc_0_3_i_web_d_reg),
      .accumulation_buffer_rsc_0_3_i_addr_d(accumulation_buffer_rsc_0_3_i_addr_d_reg),
      .accumulation_buffer_rsc_0_3_i_dout_d(accumulation_buffer_rsc_0_3_i_dout_d),
      .accumulation_buffer_rsc_0_3_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_3_i_dout_d_mxwt(accumulation_buffer_rsc_0_3_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_3_i_biwt(accumulation_buffer_rsc_0_3_i_biwt),
      .accumulation_buffer_rsc_0_3_i_bdwt(accumulation_buffer_rsc_0_3_i_bdwt),
      .accumulation_buffer_rsc_0_3_i_web_d_run_sct(accumulation_buffer_rsc_0_3_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_3_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_3_i_web_d = accumulation_buffer_rsc_0_3_i_web_d_reg;
  assign accumulation_buffer_rsc_0_3_i_addr_d = accumulation_buffer_rsc_0_3_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_3_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_2_i_web_d, accumulation_buffer_rsc_0_2_i_addr_d,
      accumulation_buffer_rsc_0_2_i_dout_d, accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_2_i_oswt, accumulation_buffer_rsc_0_2_i_addr_d_run,
      accumulation_buffer_rsc_0_2_i_dout_d_mxwt, accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_2_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_2_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_2_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_dout_d;
  output accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_2_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_2_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_2_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_2_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_2_i_biwt;
  wire accumulation_buffer_rsc_0_2_i_bdwt;
  wire accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_2_i_web_d_reg;
  wire accumulation_buffer_rsc_0_2_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_2_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_2_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_2_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_2_i_oswt(accumulation_buffer_rsc_0_2_i_oswt),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_2_i_biwt(accumulation_buffer_rsc_0_2_i_biwt),
      .accumulation_buffer_rsc_0_2_i_bdwt(accumulation_buffer_rsc_0_2_i_bdwt),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_2_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_2_i_oswt_pff(accumulation_buffer_rsc_0_2_i_oswt_pff),
      .accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_2_i_web_d(accumulation_buffer_rsc_0_2_i_web_d_reg),
      .accumulation_buffer_rsc_0_2_i_addr_d(accumulation_buffer_rsc_0_2_i_addr_d_reg),
      .accumulation_buffer_rsc_0_2_i_dout_d(accumulation_buffer_rsc_0_2_i_dout_d),
      .accumulation_buffer_rsc_0_2_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_2_i_dout_d_mxwt(accumulation_buffer_rsc_0_2_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_2_i_biwt(accumulation_buffer_rsc_0_2_i_biwt),
      .accumulation_buffer_rsc_0_2_i_bdwt(accumulation_buffer_rsc_0_2_i_bdwt),
      .accumulation_buffer_rsc_0_2_i_web_d_run_sct(accumulation_buffer_rsc_0_2_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_2_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_2_i_web_d = accumulation_buffer_rsc_0_2_i_web_d_reg;
  assign accumulation_buffer_rsc_0_2_i_addr_d = accumulation_buffer_rsc_0_2_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_2_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_1_i_web_d, accumulation_buffer_rsc_0_1_i_addr_d,
      accumulation_buffer_rsc_0_1_i_dout_d, accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_1_i_oswt, accumulation_buffer_rsc_0_1_i_addr_d_run,
      accumulation_buffer_rsc_0_1_i_dout_d_mxwt, accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_1_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_1_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_1_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_dout_d;
  output accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_1_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_1_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_1_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_1_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_1_i_biwt;
  wire accumulation_buffer_rsc_0_1_i_bdwt;
  wire accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_1_i_web_d_reg;
  wire accumulation_buffer_rsc_0_1_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_1_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_1_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_1_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_1_i_oswt(accumulation_buffer_rsc_0_1_i_oswt),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_1_i_biwt(accumulation_buffer_rsc_0_1_i_biwt),
      .accumulation_buffer_rsc_0_1_i_bdwt(accumulation_buffer_rsc_0_1_i_bdwt),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_1_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_1_i_oswt_pff(accumulation_buffer_rsc_0_1_i_oswt_pff),
      .accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_1_i_web_d(accumulation_buffer_rsc_0_1_i_web_d_reg),
      .accumulation_buffer_rsc_0_1_i_addr_d(accumulation_buffer_rsc_0_1_i_addr_d_reg),
      .accumulation_buffer_rsc_0_1_i_dout_d(accumulation_buffer_rsc_0_1_i_dout_d),
      .accumulation_buffer_rsc_0_1_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_1_i_dout_d_mxwt(accumulation_buffer_rsc_0_1_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_1_i_biwt(accumulation_buffer_rsc_0_1_i_biwt),
      .accumulation_buffer_rsc_0_1_i_bdwt(accumulation_buffer_rsc_0_1_i_bdwt),
      .accumulation_buffer_rsc_0_1_i_web_d_run_sct(accumulation_buffer_rsc_0_1_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_1_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_1_i_web_d = accumulation_buffer_rsc_0_1_i_web_d_reg;
  assign accumulation_buffer_rsc_0_1_i_addr_d = accumulation_buffer_rsc_0_1_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_1_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_0_i_web_d, accumulation_buffer_rsc_0_0_i_addr_d,
      accumulation_buffer_rsc_0_0_i_dout_d, accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d,
      accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d, run_wen,
      run_wten, accumulation_buffer_rsc_0_0_i_oswt, accumulation_buffer_rsc_0_0_i_addr_d_run,
      accumulation_buffer_rsc_0_0_i_dout_d_mxwt, accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct,
      accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff, accumulation_buffer_rsc_0_0_i_oswt_pff
);
  input clk;
  input arst_n;
  output accumulation_buffer_rsc_0_0_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_0_i_addr_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_dout_d;
  output accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_0_i_oswt;
  input [11:0] accumulation_buffer_rsc_0_0_i_addr_d_run;
  output [15:0] accumulation_buffer_rsc_0_0_i_dout_d_mxwt;
  input accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct;
  input accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff;
  input accumulation_buffer_rsc_0_0_i_oswt_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_0_i_biwt;
  wire accumulation_buffer_rsc_0_0_i_bdwt;
  wire accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  wire accumulation_buffer_rsc_0_0_i_web_d_reg;
  wire accumulation_buffer_rsc_0_0_i_web_d_run_sct_iff;
  wire [11:0] accumulation_buffer_rsc_0_0_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_0_i_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_addr_d_run
      = {6'b000000 , (accumulation_buffer_rsc_0_0_i_addr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_0_i_oswt(accumulation_buffer_rsc_0_0_i_oswt),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct),
      .accumulation_buffer_rsc_0_0_i_biwt(accumulation_buffer_rsc_0_0_i_biwt),
      .accumulation_buffer_rsc_0_0_i_bdwt(accumulation_buffer_rsc_0_0_i_bdwt),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct),
      .accumulation_buffer_rsc_0_0_i_web_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff(accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff),
      .accumulation_buffer_rsc_0_0_i_oswt_pff(accumulation_buffer_rsc_0_0_i_oswt_pff),
      .accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_addr_d_run_sct_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_0_i_web_d(accumulation_buffer_rsc_0_0_i_web_d_reg),
      .accumulation_buffer_rsc_0_0_i_addr_d(accumulation_buffer_rsc_0_0_i_addr_d_reg),
      .accumulation_buffer_rsc_0_0_i_dout_d(accumulation_buffer_rsc_0_0_i_dout_d),
      .accumulation_buffer_rsc_0_0_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_0_i_dout_d_mxwt(accumulation_buffer_rsc_0_0_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_0_i_biwt(accumulation_buffer_rsc_0_0_i_biwt),
      .accumulation_buffer_rsc_0_0_i_bdwt(accumulation_buffer_rsc_0_0_i_bdwt),
      .accumulation_buffer_rsc_0_0_i_web_d_run_sct(accumulation_buffer_rsc_0_0_i_web_d_run_sct_iff),
      .accumulation_buffer_rsc_0_0_i_addr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_addr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_0_i_web_d = accumulation_buffer_rsc_0_0_i_web_d_reg;
  assign accumulation_buffer_rsc_0_0_i_addr_d = accumulation_buffer_rsc_0_0_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_sct;
  assign accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_0_i_web_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci (
  clk, arst_n, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld, loopIndicesIn_rsc_rdy,
      run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [47:0] loopIndicesIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_biwt;
  wire loopIndicesIn_rsci_bdwt;
  wire loopIndicesIn_rsci_bcwt;
  wire loopIndicesIn_rsci_irdy_run_sct;
  wire loopIndicesIn_rsci_ivld;
  wire [47:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd104),
  .width(32'sd48)) loopIndicesIn_rsci (
      .rdy(loopIndicesIn_rsc_rdy),
      .vld(loopIndicesIn_rsc_vld),
      .dat(loopIndicesIn_rsc_dat),
      .irdy(loopIndicesIn_rsci_irdy_run_sct),
      .ivld(loopIndicesIn_rsci_ivld),
      .idat(loopIndicesIn_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_irdy_run_sct(loopIndicesIn_rsci_irdy_run_sct),
      .loopIndicesIn_rsci_ivld(loopIndicesIn_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_idat(loopIndicesIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [95:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd103),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci (
  clk, arst_n, output_rsc_dat, output_rsc_vld, output_rsc_rdy, run_wen, output_rsci_oswt,
      output_rsci_wen_comp, output_rsci_idat
);
  input clk;
  input arst_n;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input run_wen;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [255:0] output_rsci_idat;


  // Interconnect Declarations
  wire output_rsci_irdy;
  wire output_rsci_biwt;
  wire output_rsci_bdwt;
  wire output_rsci_bcwt;
  wire output_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd102),
  .width(32'sd256)) output_rsci (
      .irdy(output_rsci_irdy),
      .ivld(output_rsci_ivld_run_sct),
      .idat(output_rsci_idat),
      .rdy(output_rsc_rdy),
      .vld(output_rsc_vld),
      .dat(output_rsc_dat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_irdy(output_rsci_irdy),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt),
      .output_rsci_ivld_run_sct(output_rsci_ivld_run_sct)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci (
  clk, arst_n, weight_rsc_dat, weight_rsc_vld, weight_rsc_rdy, run_wen, weight_rsci_oswt,
      weight_rsci_wen_comp, weight_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  input run_wen;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [127:0] weight_rsci_idat_mxwt;


  // Interconnect Declarations
  wire weight_rsci_biwt;
  wire weight_rsci_bdwt;
  wire weight_rsci_bcwt;
  wire weight_rsci_irdy_run_sct;
  wire weight_rsci_ivld;
  wire [127:0] weight_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd101),
  .width(32'sd128)) weight_rsci (
      .rdy(weight_rsc_rdy),
      .vld(weight_rsc_vld),
      .dat(weight_rsc_dat),
      .irdy(weight_rsci_irdy_run_sct),
      .ivld(weight_rsci_ivld),
      .idat(weight_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_bcwt(weight_rsci_bcwt),
      .weight_rsci_irdy_run_sct(weight_rsci_irdy_run_sct),
      .weight_rsci_ivld(weight_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_idat_mxwt(weight_rsci_idat_mxwt),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_bcwt(weight_rsci_bcwt),
      .weight_rsci_idat(weight_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, run_wen, input_rsci_oswt,
      input_rsci_wen_comp, input_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [127:0] input_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_rsci_biwt;
  wire input_rsci_bdwt;
  wire input_rsci_bcwt;
  wire input_rsci_irdy_run_sct;
  wire input_rsci_ivld;
  wire [127:0] input_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd100),
  .width(32'sd128)) input_rsci (
      .rdy(input_rsc_rdy),
      .vld(input_rsc_vld),
      .dat(input_rsc_dat),
      .irdy(input_rsci_irdy_run_sct),
      .ivld(input_rsci_ivld),
      .idat(input_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_irdy_run_sct(input_rsci_irdy_run_sct),
      .input_rsci_ivld(input_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_idat(input_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy, accumulation_buffer_rsc_0_0_i_web_d, accumulation_buffer_rsc_0_0_i_addr_d,
      accumulation_buffer_rsc_0_0_i_din_d, accumulation_buffer_rsc_0_0_i_dout_d,
      accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_1_i_web_d, accumulation_buffer_rsc_0_1_i_addr_d,
      accumulation_buffer_rsc_0_1_i_din_d, accumulation_buffer_rsc_0_1_i_dout_d,
      accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_2_i_web_d, accumulation_buffer_rsc_0_2_i_addr_d,
      accumulation_buffer_rsc_0_2_i_din_d, accumulation_buffer_rsc_0_2_i_dout_d,
      accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_3_i_web_d, accumulation_buffer_rsc_0_3_i_addr_d,
      accumulation_buffer_rsc_0_3_i_din_d, accumulation_buffer_rsc_0_3_i_dout_d,
      accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_4_i_web_d, accumulation_buffer_rsc_0_4_i_addr_d,
      accumulation_buffer_rsc_0_4_i_din_d, accumulation_buffer_rsc_0_4_i_dout_d,
      accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_5_i_web_d, accumulation_buffer_rsc_0_5_i_addr_d,
      accumulation_buffer_rsc_0_5_i_din_d, accumulation_buffer_rsc_0_5_i_dout_d,
      accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_6_i_web_d, accumulation_buffer_rsc_0_6_i_addr_d,
      accumulation_buffer_rsc_0_6_i_din_d, accumulation_buffer_rsc_0_6_i_dout_d,
      accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_7_i_web_d, accumulation_buffer_rsc_0_7_i_addr_d,
      accumulation_buffer_rsc_0_7_i_din_d, accumulation_buffer_rsc_0_7_i_dout_d,
      accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_8_i_web_d, accumulation_buffer_rsc_0_8_i_addr_d,
      accumulation_buffer_rsc_0_8_i_din_d, accumulation_buffer_rsc_0_8_i_dout_d,
      accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_9_i_web_d, accumulation_buffer_rsc_0_9_i_addr_d,
      accumulation_buffer_rsc_0_9_i_din_d, accumulation_buffer_rsc_0_9_i_dout_d,
      accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_10_i_web_d, accumulation_buffer_rsc_0_10_i_addr_d,
      accumulation_buffer_rsc_0_10_i_din_d, accumulation_buffer_rsc_0_10_i_dout_d,
      accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_11_i_web_d, accumulation_buffer_rsc_0_11_i_addr_d,
      accumulation_buffer_rsc_0_11_i_din_d, accumulation_buffer_rsc_0_11_i_dout_d,
      accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_12_i_web_d, accumulation_buffer_rsc_0_12_i_addr_d,
      accumulation_buffer_rsc_0_12_i_din_d, accumulation_buffer_rsc_0_12_i_dout_d,
      accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_13_i_web_d, accumulation_buffer_rsc_0_13_i_addr_d,
      accumulation_buffer_rsc_0_13_i_din_d, accumulation_buffer_rsc_0_13_i_dout_d,
      accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_14_i_web_d, accumulation_buffer_rsc_0_14_i_addr_d,
      accumulation_buffer_rsc_0_14_i_din_d, accumulation_buffer_rsc_0_14_i_dout_d,
      accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d,
      accumulation_buffer_rsc_0_15_i_web_d, accumulation_buffer_rsc_0_15_i_addr_d,
      accumulation_buffer_rsc_0_15_i_din_d, accumulation_buffer_rsc_0_15_i_dout_d,
      accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d, accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  output accumulation_buffer_rsc_0_0_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_0_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_0_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_dout_d;
  output accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_1_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_1_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_1_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_dout_d;
  output accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_2_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_2_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_2_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_dout_d;
  output accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_3_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_3_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_3_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_dout_d;
  output accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_4_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_4_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_4_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_dout_d;
  output accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_5_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_5_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_5_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_dout_d;
  output accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_6_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_6_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_6_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_dout_d;
  output accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_7_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_7_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_7_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_dout_d;
  output accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_8_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_8_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_8_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_dout_d;
  output accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_9_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_9_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_9_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_dout_d;
  output accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_10_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_10_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_10_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_dout_d;
  output accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_11_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_11_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_11_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_dout_d;
  output accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_12_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_12_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_12_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_dout_d;
  output accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_13_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_13_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_13_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_dout_d;
  output accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_14_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_14_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_14_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_dout_d;
  output accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  output accumulation_buffer_rsc_0_15_i_web_d;
  output [11:0] accumulation_buffer_rsc_0_15_i_addr_d;
  output [15:0] accumulation_buffer_rsc_0_15_i_din_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_dout_d;
  output accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  output accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire input_rsci_wen_comp;
  wire [127:0] input_rsci_idat_mxwt;
  wire weight_rsci_wen_comp;
  wire [127:0] weight_rsci_idat_mxwt;
  wire output_rsci_wen_comp;
  wire paramsIn_rsci_wen_comp;
  wire [95:0] paramsIn_rsci_idat_mxwt;
  wire loopIndicesIn_rsci_wen_comp;
  wire [47:0] loopIndicesIn_rsci_idat_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_0_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_1_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_2_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_3_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_4_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_5_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_6_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_7_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_8_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_9_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_10_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_11_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_12_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_13_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_14_i_dout_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_15_i_dout_d_mxwt;
  wire [15:0] accum_fifo_15_rsci_output_rsc_z;
  wire accum_fifo_15_rsci_ccs_ccore_en;
  wire [15:0] output_fifo_0_rsci_output_rsc_z;
  wire output_fifo_0_rsci_ccs_ccore_en;
  wire [15:0] accum_fifo_14_rsci_output_rsc_z;
  wire [15:0] output_fifo_1_rsci_output_rsc_z;
  wire [15:0] accum_fifo_13_rsci_output_rsc_z;
  wire [15:0] output_fifo_2_rsci_output_rsc_z;
  wire [15:0] accum_fifo_12_rsci_output_rsc_z;
  wire [15:0] output_fifo_3_rsci_output_rsc_z;
  wire [15:0] accum_fifo_11_rsci_output_rsc_z;
  wire [15:0] output_fifo_4_rsci_output_rsc_z;
  wire [15:0] accum_fifo_10_rsci_output_rsc_z;
  wire [15:0] output_fifo_5_rsci_output_rsc_z;
  wire [15:0] accum_fifo_9_rsci_output_rsc_z;
  wire [15:0] output_fifo_6_rsci_output_rsc_z;
  wire [15:0] accum_fifo_8_rsci_output_rsc_z;
  wire [15:0] output_fifo_7_rsci_output_rsc_z;
  wire [15:0] accum_fifo_7_rsci_output_rsc_z;
  wire [15:0] output_fifo_8_rsci_output_rsc_z;
  wire [15:0] accum_fifo_6_rsci_output_rsc_z;
  wire [15:0] output_fifo_9_rsci_output_rsc_z;
  wire [15:0] accum_fifo_5_rsci_output_rsc_z;
  wire [15:0] output_fifo_10_rsci_output_rsc_z;
  wire [15:0] accum_fifo_4_rsci_output_rsc_z;
  wire [15:0] output_fifo_11_rsci_output_rsc_z;
  wire [15:0] accum_fifo_3_rsci_output_rsc_z;
  wire [15:0] output_fifo_12_rsci_output_rsc_z;
  wire [15:0] accum_fifo_2_rsci_output_rsc_z;
  wire [15:0] output_fifo_13_rsci_output_rsc_z;
  wire [15:0] accum_fifo_1_rsci_output_rsc_z;
  wire [15:0] output_fifo_14_rsci_output_rsc_z;
  wire [7:0] input_fifo_15_rsci_output_rsc_z;
  wire input_fifo_15_rsci_ccs_ccore_en;
  wire [7:0] input_fifo_14_rsci_output_rsc_z;
  wire [7:0] input_fifo_13_rsci_output_rsc_z;
  wire [7:0] input_fifo_12_rsci_output_rsc_z;
  wire [7:0] input_fifo_11_rsci_output_rsc_z;
  wire [7:0] input_fifo_10_rsci_output_rsc_z;
  wire [7:0] input_fifo_9_rsci_output_rsc_z;
  wire [7:0] input_fifo_8_rsci_output_rsc_z;
  wire [7:0] input_fifo_7_rsci_output_rsc_z;
  wire [7:0] input_fifo_6_rsci_output_rsc_z;
  wire [7:0] input_fifo_5_rsci_output_rsc_z;
  wire [7:0] input_fifo_4_rsci_output_rsc_z;
  wire [7:0] input_fifo_3_rsci_output_rsc_z;
  wire [7:0] input_fifo_2_rsci_output_rsc_z;
  wire [7:0] input_fifo_1_rsci_output_rsc_z;
  wire [7:0] pe_0_0_run_cmp_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_psum_out_rsc_z;
  wire pe_0_0_run_cmp_ccs_ccore_en;
  wire [15:0] accum_fifo_0_run_cmp_output_rsc_z;
  wire accum_fifo_0_run_cmp_ccs_ccore_en;
  wire [7:0] input_fifo_0_run_cmp_output_rsc_z;
  reg [15:0] output_rsci_idat_255_240;
  reg [15:0] output_rsci_idat_239_224;
  reg [15:0] output_rsci_idat_223_208;
  reg [15:0] output_rsci_idat_207_192;
  reg [15:0] output_rsci_idat_191_176;
  reg [15:0] output_rsci_idat_175_160;
  reg [15:0] output_rsci_idat_159_144;
  reg [15:0] output_rsci_idat_143_128;
  reg [15:0] output_rsci_idat_127_112;
  reg [15:0] output_rsci_idat_111_96;
  reg [15:0] output_rsci_idat_95_80;
  reg [15:0] output_rsci_idat_79_64;
  reg [15:0] output_rsci_idat_63_48;
  reg [15:0] output_rsci_idat_47_32;
  reg [15:0] output_rsci_idat_31_16;
  reg [15:0] output_rsci_idat_15_0;
  wire [8:0] fsm_output;
  wire step_if_3_aif_1_step_if_3_aelse_1_step_if_3_aelse_1_nor_tmp;
  wire step_if_3_aif_step_if_3_aelse_step_if_3_aelse_nor_tmp;
  wire step_if_3_step_if_3_if_step_if_3_if_nor_tmp;
  wire step_if_2_if_step_if_2_if_and_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire or_dcpl_4;
  wire or_dcpl_10;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_12;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire mux_tmp_80;
  wire or_tmp_121;
  wire or_tmp_122;
  wire and_dcpl_20;
  wire or_dcpl_14;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_27;
  wire and_dcpl_29;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_121;
  wire and_dcpl_122;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_132;
  wire and_dcpl_133;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_145;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_148;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_195;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_213;
  wire and_dcpl_214;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire and_dcpl_222;
  wire and_dcpl_223;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_226;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_229;
  wire and_dcpl_230;
  wire and_dcpl_231;
  wire and_dcpl_232;
  wire and_dcpl_233;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_236;
  wire and_dcpl_237;
  wire and_dcpl_238;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_243;
  wire and_dcpl_244;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_248;
  wire and_dcpl_249;
  wire and_dcpl_250;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_253;
  wire and_dcpl_254;
  wire and_dcpl_255;
  wire and_dcpl_256;
  wire and_dcpl_257;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire and_dcpl_266;
  wire and_dcpl_267;
  wire and_dcpl_268;
  wire and_dcpl_269;
  wire and_dcpl_270;
  wire and_dcpl_271;
  wire and_dcpl_272;
  wire and_dcpl_273;
  wire and_dcpl_274;
  wire and_dcpl_275;
  wire and_dcpl_276;
  wire and_dcpl_277;
  wire and_dcpl_278;
  wire and_dcpl_279;
  wire and_dcpl_280;
  wire and_dcpl_281;
  wire and_dcpl_282;
  wire and_dcpl_283;
  wire and_dcpl_284;
  wire and_dcpl_285;
  wire and_dcpl_286;
  wire and_dcpl_287;
  wire and_dcpl_288;
  wire and_dcpl_289;
  wire and_dcpl_290;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_297;
  wire and_dcpl_298;
  wire and_dcpl_299;
  wire and_dcpl_300;
  wire and_dcpl_301;
  wire and_dcpl_302;
  wire and_dcpl_303;
  wire and_dcpl_304;
  wire and_dcpl_305;
  wire and_dcpl_306;
  wire and_dcpl_307;
  wire and_dcpl_308;
  wire and_dcpl_309;
  wire and_dcpl_310;
  wire and_dcpl_311;
  wire and_dcpl_312;
  wire and_dcpl_313;
  wire and_dcpl_314;
  wire and_dcpl_315;
  wire and_dcpl_316;
  wire and_dcpl_317;
  wire and_dcpl_318;
  wire and_dcpl_319;
  wire and_dcpl_320;
  wire and_dcpl_321;
  wire and_dcpl_322;
  wire and_dcpl_323;
  wire and_dcpl_324;
  wire and_dcpl_325;
  wire and_dcpl_326;
  wire and_dcpl_327;
  wire and_dcpl_328;
  wire and_dcpl_329;
  wire and_dcpl_330;
  wire and_dcpl_333;
  wire and_dcpl_334;
  wire and_dcpl_335;
  wire and_dcpl_336;
  wire and_dcpl_341;
  wire or_tmp_126;
  wire or_tmp_127;
  wire or_tmp_129;
  wire or_tmp_130;
  wire mux_tmp_91;
  wire or_tmp_133;
  wire mux_tmp_93;
  wire mux_tmp_103;
  wire nand_tmp_5;
  wire nor_tmp_20;
  wire mux_tmp_118;
  wire mux_tmp_153;
  wire nand_tmp_14;
  wire nor_tmp_41;
  wire or_tmp_213;
  wire mux_tmp_205;
  wire mux_tmp_206;
  wire or_tmp_219;
  wire or_tmp_225;
  wire mux_tmp_217;
  wire or_tmp_239;
  wire mux_tmp_231;
  wire mux_tmp_232;
  wire or_tmp_262;
  wire or_tmp_264;
  wire or_tmp_268;
  wire or_tmp_270;
  wire mux_tmp_253;
  wire or_tmp_282;
  wire or_tmp_292;
  wire mux_tmp_275;
  wire mux_tmp_280;
  wire mux_tmp_282;
  wire and_dcpl_360;
  wire and_dcpl_362;
  wire and_dcpl_376;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire and_dcpl_388;
  wire and_dcpl_394;
  wire and_dcpl_395;
  wire and_dcpl_397;
  wire and_dcpl_399;
  wire and_dcpl_401;
  wire and_dcpl_405;
  wire and_dcpl_406;
  wire and_dcpl_408;
  wire and_dcpl_410;
  wire and_dcpl_411;
  wire and_dcpl_412;
  wire and_dcpl_414;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_419;
  wire and_dcpl_421;
  wire and_dcpl_422;
  wire and_dcpl_424;
  wire and_dcpl_426;
  wire and_dcpl_427;
  wire and_dcpl_429;
  wire and_dcpl_431;
  wire and_dcpl_432;
  wire and_dcpl_434;
  wire and_dcpl_436;
  wire and_dcpl_438;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_35;
  wire or_dcpl_37;
  wire or_dcpl_38;
  wire or_dcpl_40;
  wire or_dcpl_41;
  wire or_dcpl_43;
  wire or_dcpl_44;
  wire or_dcpl_45;
  wire or_dcpl_46;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_50;
  wire or_dcpl_52;
  wire or_dcpl_54;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_59;
  wire or_dcpl_61;
  wire or_dcpl_63;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire or_dcpl_75;
  wire or_dcpl_76;
  wire or_dcpl_85;
  wire or_dcpl_94;
  wire or_dcpl_95;
  wire or_dcpl_97;
  wire or_dcpl_99;
  wire or_dcpl_101;
  wire or_dcpl_103;
  wire or_dcpl_132;
  wire or_dcpl_133;
  wire or_dcpl_142;
  wire or_dcpl_151;
  wire or_dcpl_159;
  wire or_dcpl_200;
  wire or_dcpl_201;
  wire or_dcpl_210;
  wire or_dcpl_219;
  wire or_dcpl_228;
  wire or_dcpl_269;
  wire or_dcpl_278;
  wire or_dcpl_287;
  wire and_dcpl_445;
  wire mux_tmp_337;
  wire mux_tmp_345;
  reg [15:0] step_step_sva;
  reg operator_16_false_slc_operator_16_false_acc_16_itm;
  reg operator_16_false_slc_operator_16_false_acc_12_svs;
  reg step_if_1_acc_cse_32;
  reg [47:0] loopIndicesIn_crt_sva;
  wire [16:0] operator_16_false_1_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_1_acc_psp_sva_1;
  wire output_and_cse;
  wire or_170_cse;
  wire nand_111_cse;
  wire or_186_cse;
  wire or_169_cse;
  wire or_201_cse;
  wire or_187_cse;
  wire or_220_cse;
  reg reg_ensig_cgo_47_cse;
  reg reg_ensig_cgo_29_cse;
  reg reg_ensig_cgo_28_cse;
  reg reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse;
  reg reg_loopIndicesIn_rsci_irdy_run_psct_cse;
  reg reg_output_rsci_ivld_run_psct_cse;
  reg reg_weight_rsci_irdy_run_psct_cse;
  reg reg_input_rsci_irdy_run_psct_cse;
  reg reg_ensig_cgo_46_cse;
  reg reg_ensig_cgo_45_cse;
  wire input_reg_and_1_cse;
  wire input_reg_and_2_cse;
  wire input_reg_and_3_cse;
  wire input_reg_and_4_cse;
  wire input_reg_and_5_cse;
  wire input_reg_and_6_cse;
  wire input_reg_and_7_cse;
  wire input_reg_and_8_cse;
  wire input_reg_and_9_cse;
  wire input_reg_and_10_cse;
  wire input_reg_and_11_cse;
  wire input_reg_and_12_cse;
  wire input_reg_and_13_cse;
  wire input_reg_and_14_cse;
  wire input_reg_and_16_cse;
  wire input_reg_and_17_cse;
  wire input_reg_and_18_cse;
  wire input_reg_and_19_cse;
  wire input_reg_and_20_cse;
  wire input_reg_and_21_cse;
  wire input_reg_and_22_cse;
  wire input_reg_and_23_cse;
  wire input_reg_and_24_cse;
  wire input_reg_and_25_cse;
  wire input_reg_and_26_cse;
  wire input_reg_and_27_cse;
  wire input_reg_and_28_cse;
  wire input_reg_and_29_cse;
  wire input_reg_and_31_cse;
  wire input_reg_and_32_cse;
  wire input_reg_and_33_cse;
  wire input_reg_and_34_cse;
  wire input_reg_and_35_cse;
  wire input_reg_and_36_cse;
  wire input_reg_and_37_cse;
  wire input_reg_and_38_cse;
  wire input_reg_and_39_cse;
  wire input_reg_and_40_cse;
  wire input_reg_and_41_cse;
  wire input_reg_and_42_cse;
  wire input_reg_and_43_cse;
  wire input_reg_and_44_cse;
  wire input_reg_and_46_cse;
  wire input_reg_and_47_cse;
  wire input_reg_and_48_cse;
  wire input_reg_and_49_cse;
  wire input_reg_and_50_cse;
  wire input_reg_and_51_cse;
  wire input_reg_and_52_cse;
  wire input_reg_and_53_cse;
  wire input_reg_and_54_cse;
  wire input_reg_and_55_cse;
  wire input_reg_and_56_cse;
  wire input_reg_and_57_cse;
  wire input_reg_and_58_cse;
  wire input_reg_and_59_cse;
  wire input_reg_and_61_cse;
  wire input_reg_and_62_cse;
  wire input_reg_and_63_cse;
  wire input_reg_and_64_cse;
  wire input_reg_and_65_cse;
  wire input_reg_and_66_cse;
  wire input_reg_and_67_cse;
  wire input_reg_and_68_cse;
  wire input_reg_and_69_cse;
  wire input_reg_and_70_cse;
  wire input_reg_and_71_cse;
  wire input_reg_and_72_cse;
  wire input_reg_and_73_cse;
  wire input_reg_and_74_cse;
  wire input_reg_and_75_cse;
  wire input_reg_and_76_cse;
  wire input_reg_and_77_cse;
  wire input_reg_and_78_cse;
  wire input_reg_and_79_cse;
  wire input_reg_and_80_cse;
  wire input_reg_and_81_cse;
  wire input_reg_and_82_cse;
  wire input_reg_and_83_cse;
  wire input_reg_and_84_cse;
  wire input_reg_and_85_cse;
  wire input_reg_and_86_cse;
  wire input_reg_and_87_cse;
  wire input_reg_and_88_cse;
  wire input_reg_and_89_cse;
  wire input_reg_and_91_cse;
  wire input_reg_and_92_cse;
  wire input_reg_and_93_cse;
  wire input_reg_and_94_cse;
  wire input_reg_and_95_cse;
  wire input_reg_and_96_cse;
  wire input_reg_and_97_cse;
  wire input_reg_and_98_cse;
  wire input_reg_and_99_cse;
  wire input_reg_and_100_cse;
  wire input_reg_and_101_cse;
  wire input_reg_and_102_cse;
  wire input_reg_and_103_cse;
  wire input_reg_and_104_cse;
  wire input_reg_and_105_cse;
  wire input_reg_and_107_cse;
  wire input_reg_and_108_cse;
  wire input_reg_and_109_cse;
  wire input_reg_and_110_cse;
  wire input_reg_and_111_cse;
  wire input_reg_and_112_cse;
  wire input_reg_and_113_cse;
  wire input_reg_and_114_cse;
  wire input_reg_and_115_cse;
  wire input_reg_and_116_cse;
  wire input_reg_and_117_cse;
  wire input_reg_and_118_cse;
  wire input_reg_and_119_cse;
  wire input_reg_and_120_cse;
  wire input_reg_and_121_cse;
  wire input_reg_and_123_cse;
  wire input_reg_and_124_cse;
  wire input_reg_and_125_cse;
  wire input_reg_and_126_cse;
  wire input_reg_and_127_cse;
  wire input_reg_and_128_cse;
  wire input_reg_and_129_cse;
  wire input_reg_and_130_cse;
  wire input_reg_and_131_cse;
  wire input_reg_and_132_cse;
  wire input_reg_and_133_cse;
  wire input_reg_and_134_cse;
  wire input_reg_and_135_cse;
  wire input_reg_and_136_cse;
  wire input_reg_and_137_cse;
  wire input_reg_and_139_cse;
  wire input_reg_and_140_cse;
  wire input_reg_and_141_cse;
  wire input_reg_and_142_cse;
  wire input_reg_and_143_cse;
  wire input_reg_and_144_cse;
  wire input_reg_and_145_cse;
  wire input_reg_and_146_cse;
  wire input_reg_and_147_cse;
  wire input_reg_and_148_cse;
  wire input_reg_and_149_cse;
  wire input_reg_and_150_cse;
  wire input_reg_and_151_cse;
  wire input_reg_and_152_cse;
  wire input_reg_and_153_cse;
  wire input_reg_and_155_cse;
  wire input_reg_and_156_cse;
  wire input_reg_and_157_cse;
  wire input_reg_and_158_cse;
  wire input_reg_and_159_cse;
  wire input_reg_and_160_cse;
  wire input_reg_and_161_cse;
  wire input_reg_and_162_cse;
  wire input_reg_and_163_cse;
  wire input_reg_and_164_cse;
  wire input_reg_and_165_cse;
  wire input_reg_and_166_cse;
  wire input_reg_and_167_cse;
  wire input_reg_and_168_cse;
  wire input_reg_and_169_cse;
  wire input_reg_and_171_cse;
  wire input_reg_and_172_cse;
  wire input_reg_and_173_cse;
  wire input_reg_and_174_cse;
  wire input_reg_and_175_cse;
  wire input_reg_and_176_cse;
  wire input_reg_and_177_cse;
  wire input_reg_and_178_cse;
  wire input_reg_and_179_cse;
  wire input_reg_and_180_cse;
  wire input_reg_and_181_cse;
  wire input_reg_and_182_cse;
  wire input_reg_and_183_cse;
  wire input_reg_and_184_cse;
  wire input_reg_and_185_cse;
  wire input_reg_and_187_cse;
  wire input_reg_and_188_cse;
  wire input_reg_and_189_cse;
  wire input_reg_and_190_cse;
  wire input_reg_and_191_cse;
  wire input_reg_and_192_cse;
  wire input_reg_and_193_cse;
  wire input_reg_and_194_cse;
  wire input_reg_and_195_cse;
  wire input_reg_and_196_cse;
  wire input_reg_and_197_cse;
  wire input_reg_and_198_cse;
  wire input_reg_and_199_cse;
  wire input_reg_and_200_cse;
  wire input_reg_and_201_cse;
  wire input_reg_and_203_cse;
  wire input_reg_and_204_cse;
  wire input_reg_and_205_cse;
  wire input_reg_and_206_cse;
  wire input_reg_and_207_cse;
  wire input_reg_and_208_cse;
  wire input_reg_and_209_cse;
  wire input_reg_and_210_cse;
  wire input_reg_and_211_cse;
  wire input_reg_and_212_cse;
  wire input_reg_and_213_cse;
  wire input_reg_and_214_cse;
  wire input_reg_and_215_cse;
  wire input_reg_and_216_cse;
  wire input_reg_and_217_cse;
  wire input_reg_and_219_cse;
  wire input_reg_and_220_cse;
  wire input_reg_and_221_cse;
  wire input_reg_and_222_cse;
  wire input_reg_and_223_cse;
  wire input_reg_and_224_cse;
  wire input_reg_and_225_cse;
  wire input_reg_and_226_cse;
  wire input_reg_and_227_cse;
  wire input_reg_and_228_cse;
  wire input_reg_and_229_cse;
  wire input_reg_and_230_cse;
  wire input_reg_and_231_cse;
  wire input_reg_and_232_cse;
  wire input_reg_and_233_cse;
  wire input_reg_and_30_cse;
  wire input_reg_and_45_cse;
  wire input_reg_and_60_cse;
  wire or_338_cse;
  wire nor_133_cse;
  wire nor_150_cse;
  wire or_645_cse;
  wire or_52_cse;
  wire or_58_cse;
  wire or_55_cse;
  wire nor_174_cse;
  wire or_94_cse;
  wire or_827_cse;
  wire nand_62_cse;
  wire nand_94_cse;
  wire input_reg_and_239_cse;
  wire and_463_cse;
  wire or_47_cse;
  wire and_cse;
  wire or_228_cse;
  wire mux_434_cse;
  wire or_765_cse;
  wire nand_100_cse;
  wire or_322_cse;
  wire mux_130_cse;
  wire mux_111_cse;
  wire mux_109_cse;
  wire mux_239_cse;
  wire mux_234_cse;
  wire mux_306_cse;
  wire mux_322_cse;
  wire mux_245_cse;
  wire mux_377_cse;
  wire or_176_cse;
  wire or_743_cse;
  wire or_177_cse;
  wire nand_10_cse;
  wire mux_142_cse;
  wire mux_210_cse;
  wire or_178_cse;
  wire mux_156_cse;
  wire mux_207_cse;
  wire mux_199_cse;
  wire or_222_cse;
  wire accumulation_buffer_rsc_0_0_i_web_d_reg;
  wire and_372_rmff;
  wire and_380_rmff;
  wire [11:0] accumulation_buffer_rsc_0_0_i_addr_d_reg;
  wire [5:0] operator_16_false_mux_rmff;
  wire accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire and_377_rmff;
  wire accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_1_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_1_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_2_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_2_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_3_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_3_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_4_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_4_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_5_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_5_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_6_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_6_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_7_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_7_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_8_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_8_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_9_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_9_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_10_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_10_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_11_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_11_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_12_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_12_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_13_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_13_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_14_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_14_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_15_i_web_d_reg;
  wire [11:0] accumulation_buffer_rsc_0_15_i_addr_d_reg;
  wire accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  wire and_368_rmff;
  wire and_364_rmff;
  wire and_17_rmff;
  wire and_23_rmff;
  reg [15:0] step_output_buf_value_0_sva;
  reg [15:0] psum_reg_16_8_lpi_2;
  reg [15:0] psum_reg_15_16_lpi_2;
  reg [15:0] psum_reg_16_15_lpi_2;
  reg [15:0] psum_reg_16_16_lpi_2;
  reg [15:0] psum_reg_16_2_lpi_2;
  reg [15:0] psum_reg_16_3_lpi_2;
  reg [15:0] psum_reg_16_4_lpi_2;
  reg [15:0] psum_reg_16_5_lpi_2;
  reg [15:0] psum_reg_16_6_lpi_2;
  reg [15:0] psum_reg_16_7_lpi_2;
  reg [15:0] psum_reg_16_1_lpi_2;
  reg [15:0] psum_reg_16_10_lpi_2;
  reg [15:0] psum_reg_16_11_lpi_2;
  reg [15:0] psum_reg_16_12_lpi_2;
  reg [15:0] psum_reg_16_14_lpi_2;
  reg [15:0] psum_reg_16_9_lpi_2;
  wire [127:0] step_in_col_value_lpi_2_dfm_mx0;
  reg [7:0] input_reg_16_15_lpi_2;
  reg [7:0] input_reg_16_14_lpi_2;
  reg [7:0] input_reg_16_13_lpi_2;
  reg [7:0] input_reg_16_10_lpi_2;
  reg [7:0] input_reg_16_11_lpi_2;
  reg [7:0] input_reg_16_12_lpi_2;
  reg [7:0] ROW_asn_142_itm;
  reg [7:0] ROW_asn_143_itm;
  reg [7:0] ROW_asn_145_itm;
  reg [7:0] ROW_asn_147_itm;
  reg [7:0] ROW_asn_149_itm;
  reg [7:0] ROW_asn_151_itm;
  reg [7:0] ROW_asn_153_itm;
  reg [7:0] ROW_asn_155_itm;
  reg [7:0] ROW_asn_157_itm;
  reg [7:0] ROW_asn_159_itm;
  reg [7:0] ROW_asn_161_itm;
  reg [7:0] ROW_asn_163_itm;
  reg [7:0] ROW_asn_165_itm;
  reg [7:0] ROW_asn_167_itm;
  reg [7:0] ROW_asn_169_itm;
  reg [15:0] psum_reg_15_15_lpi_2;
  reg [15:0] psum_reg_15_14_lpi_2;
  reg [15:0] psum_reg_15_11_lpi_2;
  reg [15:0] psum_reg_15_12_lpi_2;
  reg [15:0] psum_reg_15_13_lpi_2;
  reg [15:0] psum_reg_1_1_lpi_2;
  reg [15:0] psum_reg_2_1_lpi_2;
  reg [15:0] psum_reg_3_1_lpi_2;
  reg [15:0] psum_reg_4_1_lpi_2;
  reg [15:0] psum_reg_5_1_lpi_2;
  reg [15:0] psum_reg_6_1_lpi_2;
  reg [15:0] psum_reg_7_1_lpi_2;
  reg [15:0] psum_reg_8_1_lpi_2;
  reg [15:0] psum_reg_9_1_lpi_2;
  reg [15:0] psum_reg_10_1_lpi_2;
  reg [15:0] psum_reg_11_1_lpi_2;
  reg [15:0] psum_reg_12_1_lpi_2;
  reg [15:0] psum_reg_13_1_lpi_2;
  reg [15:0] psum_reg_14_1_lpi_2;
  reg [15:0] psum_reg_15_1_lpi_2;
  reg [15:0] psum_reg_1_2_lpi_2;
  reg [15:0] psum_reg_2_2_lpi_2;
  reg [15:0] psum_reg_3_2_lpi_2;
  reg [15:0] psum_reg_4_2_lpi_2;
  reg [15:0] psum_reg_5_2_lpi_2;
  reg [15:0] psum_reg_6_2_lpi_2;
  reg [15:0] psum_reg_7_2_lpi_2;
  reg [15:0] psum_reg_8_2_lpi_2;
  reg [15:0] psum_reg_9_2_lpi_2;
  reg [15:0] psum_reg_10_2_lpi_2;
  reg [15:0] psum_reg_11_2_lpi_2;
  reg [15:0] psum_reg_12_2_lpi_2;
  reg [15:0] psum_reg_13_2_lpi_2;
  reg [15:0] psum_reg_14_2_lpi_2;
  reg [15:0] psum_reg_15_2_lpi_2;
  reg [15:0] psum_reg_1_3_lpi_2;
  reg [15:0] psum_reg_2_3_lpi_2;
  reg [15:0] psum_reg_3_3_lpi_2;
  reg [15:0] psum_reg_4_3_lpi_2;
  reg [15:0] psum_reg_5_3_lpi_2;
  reg [15:0] psum_reg_6_3_lpi_2;
  reg [15:0] psum_reg_7_3_lpi_2;
  reg [15:0] psum_reg_8_3_lpi_2;
  reg [15:0] psum_reg_9_3_lpi_2;
  reg [15:0] psum_reg_10_3_lpi_2;
  reg [15:0] psum_reg_11_3_lpi_2;
  reg [15:0] psum_reg_12_3_lpi_2;
  reg [15:0] psum_reg_13_3_lpi_2;
  reg [15:0] psum_reg_14_3_lpi_2;
  reg [15:0] psum_reg_15_3_lpi_2;
  reg [15:0] psum_reg_1_4_lpi_2;
  reg [15:0] psum_reg_2_4_lpi_2;
  reg [15:0] psum_reg_3_4_lpi_2;
  reg [15:0] psum_reg_4_4_lpi_2;
  reg [15:0] psum_reg_5_4_lpi_2;
  reg [15:0] psum_reg_6_4_lpi_2;
  reg [15:0] psum_reg_7_4_lpi_2;
  reg [15:0] psum_reg_8_4_lpi_2;
  reg [15:0] psum_reg_9_4_lpi_2;
  reg [15:0] psum_reg_10_4_lpi_2;
  reg [15:0] psum_reg_11_4_lpi_2;
  reg [15:0] psum_reg_12_4_lpi_2;
  reg [15:0] psum_reg_13_4_lpi_2;
  reg [15:0] psum_reg_14_4_lpi_2;
  reg [15:0] psum_reg_15_4_lpi_2;
  reg [15:0] psum_reg_1_5_lpi_2;
  reg [15:0] psum_reg_2_5_lpi_2;
  reg [15:0] psum_reg_3_5_lpi_2;
  reg [15:0] psum_reg_4_5_lpi_2;
  reg [15:0] psum_reg_5_5_lpi_2;
  reg [15:0] psum_reg_6_5_lpi_2;
  reg [15:0] psum_reg_7_5_lpi_2;
  reg [15:0] psum_reg_8_5_lpi_2;
  reg [15:0] psum_reg_9_5_lpi_2;
  reg [15:0] psum_reg_10_5_lpi_2;
  reg [15:0] psum_reg_11_5_lpi_2;
  reg [15:0] psum_reg_12_5_lpi_2;
  reg [15:0] psum_reg_13_5_lpi_2;
  reg [15:0] psum_reg_14_5_lpi_2;
  reg [15:0] psum_reg_15_5_lpi_2;
  reg [15:0] psum_reg_1_6_lpi_2;
  reg [15:0] psum_reg_2_6_lpi_2;
  reg [15:0] psum_reg_3_6_lpi_2;
  reg [15:0] psum_reg_4_6_lpi_2;
  reg [15:0] psum_reg_5_6_lpi_2;
  reg [15:0] psum_reg_6_6_lpi_2;
  reg [15:0] psum_reg_7_6_lpi_2;
  reg [15:0] psum_reg_8_6_lpi_2;
  reg [15:0] psum_reg_9_6_lpi_2;
  reg [15:0] psum_reg_10_6_lpi_2;
  reg [15:0] psum_reg_11_6_lpi_2;
  reg [15:0] psum_reg_12_6_lpi_2;
  reg [15:0] psum_reg_13_6_lpi_2;
  reg [15:0] psum_reg_14_6_lpi_2;
  reg [15:0] psum_reg_15_6_lpi_2;
  reg [15:0] psum_reg_1_7_lpi_2;
  reg [15:0] psum_reg_2_7_lpi_2;
  reg [15:0] psum_reg_3_7_lpi_2;
  reg [15:0] psum_reg_4_7_lpi_2;
  reg [15:0] psum_reg_5_7_lpi_2;
  reg [15:0] psum_reg_6_7_lpi_2;
  reg [15:0] psum_reg_7_7_lpi_2;
  reg [15:0] psum_reg_8_7_lpi_2;
  reg [15:0] psum_reg_9_7_lpi_2;
  reg [15:0] psum_reg_10_7_lpi_2;
  reg [15:0] psum_reg_11_7_lpi_2;
  reg [15:0] psum_reg_12_7_lpi_2;
  reg [15:0] psum_reg_13_7_lpi_2;
  reg [15:0] psum_reg_14_7_lpi_2;
  reg [15:0] psum_reg_15_7_lpi_2;
  reg [15:0] psum_reg_1_8_lpi_2;
  reg [15:0] psum_reg_2_8_lpi_2;
  reg [15:0] psum_reg_3_8_lpi_2;
  reg [15:0] psum_reg_4_8_lpi_2;
  reg [15:0] psum_reg_5_8_lpi_2;
  reg [15:0] psum_reg_6_8_lpi_2;
  reg [15:0] psum_reg_7_8_lpi_2;
  reg [15:0] psum_reg_8_8_lpi_2;
  reg [15:0] psum_reg_9_8_lpi_2;
  reg [15:0] psum_reg_10_8_lpi_2;
  reg [15:0] psum_reg_11_8_lpi_2;
  reg [15:0] psum_reg_12_8_lpi_2;
  reg [15:0] psum_reg_13_8_lpi_2;
  reg [15:0] psum_reg_14_8_lpi_2;
  reg [15:0] psum_reg_15_8_lpi_2;
  reg [15:0] psum_reg_1_9_lpi_2;
  reg [15:0] psum_reg_2_9_lpi_2;
  reg [15:0] psum_reg_3_9_lpi_2;
  reg [15:0] psum_reg_4_9_lpi_2;
  reg [15:0] psum_reg_5_9_lpi_2;
  reg [15:0] psum_reg_6_9_lpi_2;
  reg [15:0] psum_reg_7_9_lpi_2;
  reg [15:0] psum_reg_8_9_lpi_2;
  reg [15:0] psum_reg_9_9_lpi_2;
  reg [15:0] psum_reg_10_9_lpi_2;
  reg [15:0] psum_reg_11_9_lpi_2;
  reg [15:0] psum_reg_12_9_lpi_2;
  reg [15:0] psum_reg_13_9_lpi_2;
  reg [15:0] psum_reg_14_9_lpi_2;
  reg [15:0] psum_reg_15_9_lpi_2;
  reg [15:0] psum_reg_1_10_lpi_2;
  reg [15:0] psum_reg_2_10_lpi_2;
  reg [15:0] psum_reg_3_10_lpi_2;
  reg [15:0] psum_reg_4_10_lpi_2;
  reg [15:0] psum_reg_5_10_lpi_2;
  reg [15:0] psum_reg_6_10_lpi_2;
  reg [15:0] psum_reg_7_10_lpi_2;
  reg [15:0] psum_reg_8_10_lpi_2;
  reg [15:0] psum_reg_9_10_lpi_2;
  reg [15:0] psum_reg_10_10_lpi_2;
  reg [15:0] psum_reg_11_10_lpi_2;
  reg [15:0] psum_reg_12_10_lpi_2;
  reg [15:0] psum_reg_13_10_lpi_2;
  reg [15:0] psum_reg_14_10_lpi_2;
  reg [15:0] psum_reg_15_10_lpi_2;
  reg [15:0] step_accum_fifo_input_15_asn_9_ncse_sva;
  reg [15:0] psum_reg_1_11_lpi_2;
  reg [15:0] psum_reg_2_11_lpi_2;
  reg [15:0] psum_reg_3_11_lpi_2;
  reg [15:0] psum_reg_4_11_lpi_2;
  reg [15:0] psum_reg_5_11_lpi_2;
  reg [15:0] psum_reg_6_11_lpi_2;
  reg [15:0] psum_reg_7_11_lpi_2;
  reg [15:0] psum_reg_8_11_lpi_2;
  reg [15:0] psum_reg_9_11_lpi_2;
  reg [15:0] psum_reg_10_11_lpi_2;
  reg [15:0] psum_reg_11_11_lpi_2;
  reg [15:0] psum_reg_12_11_lpi_2;
  reg [15:0] psum_reg_13_11_lpi_2;
  reg [15:0] psum_reg_14_11_lpi_2;
  reg [15:0] psum_reg_1_12_lpi_2;
  reg [15:0] psum_reg_2_12_lpi_2;
  reg [15:0] psum_reg_3_12_lpi_2;
  reg [15:0] psum_reg_4_12_lpi_2;
  reg [15:0] psum_reg_5_12_lpi_2;
  reg [15:0] psum_reg_6_12_lpi_2;
  reg [15:0] psum_reg_7_12_lpi_2;
  reg [15:0] psum_reg_8_12_lpi_2;
  reg [15:0] psum_reg_9_12_lpi_2;
  reg [15:0] psum_reg_10_12_lpi_2;
  reg [15:0] psum_reg_11_12_lpi_2;
  reg [15:0] psum_reg_12_12_lpi_2;
  reg [15:0] psum_reg_13_12_lpi_2;
  reg [15:0] psum_reg_14_12_lpi_2;
  reg [15:0] psum_reg_1_13_lpi_2;
  reg [15:0] psum_reg_2_13_lpi_2;
  reg [15:0] psum_reg_3_13_lpi_2;
  reg [15:0] psum_reg_4_13_lpi_2;
  reg [15:0] psum_reg_5_13_lpi_2;
  reg [15:0] psum_reg_6_13_lpi_2;
  reg [15:0] psum_reg_7_13_lpi_2;
  reg [15:0] psum_reg_8_13_lpi_2;
  reg [15:0] psum_reg_9_13_lpi_2;
  reg [15:0] psum_reg_10_13_lpi_2;
  reg [15:0] psum_reg_11_13_lpi_2;
  reg [15:0] psum_reg_12_13_lpi_2;
  reg [15:0] psum_reg_13_13_lpi_2;
  reg [15:0] psum_reg_14_13_lpi_2;
  reg [15:0] step_accum_fifo_input_15_asn_12_ncse_sva;
  reg [15:0] psum_reg_1_14_lpi_2;
  reg [15:0] psum_reg_2_14_lpi_2;
  reg [15:0] psum_reg_3_14_lpi_2;
  reg [15:0] psum_reg_4_14_lpi_2;
  reg [15:0] psum_reg_5_14_lpi_2;
  reg [15:0] psum_reg_6_14_lpi_2;
  reg [15:0] psum_reg_7_14_lpi_2;
  reg [15:0] psum_reg_8_14_lpi_2;
  reg [15:0] psum_reg_9_14_lpi_2;
  reg [15:0] psum_reg_10_14_lpi_2;
  reg [15:0] psum_reg_11_14_lpi_2;
  reg [15:0] psum_reg_12_14_lpi_2;
  reg [15:0] psum_reg_13_14_lpi_2;
  reg [15:0] psum_reg_14_14_lpi_2;
  reg [15:0] step_accum_fifo_input_15_asn_13_ncse_sva;
  reg [15:0] psum_reg_1_15_lpi_2;
  reg [15:0] psum_reg_2_15_lpi_2;
  reg [15:0] psum_reg_3_15_lpi_2;
  reg [15:0] psum_reg_4_15_lpi_2;
  reg [15:0] psum_reg_5_15_lpi_2;
  reg [15:0] psum_reg_6_15_lpi_2;
  reg [15:0] psum_reg_7_15_lpi_2;
  reg [15:0] psum_reg_8_15_lpi_2;
  reg [15:0] psum_reg_9_15_lpi_2;
  reg [15:0] psum_reg_10_15_lpi_2;
  reg [15:0] psum_reg_11_15_lpi_2;
  reg [15:0] psum_reg_12_15_lpi_2;
  reg [15:0] psum_reg_13_15_lpi_2;
  reg [15:0] psum_reg_14_15_lpi_2;
  reg [15:0] step_accum_fifo_input_15_asn_14_ncse_sva;
  reg [15:0] psum_reg_1_16_lpi_2;
  reg [15:0] psum_reg_2_16_lpi_2;
  reg [15:0] psum_reg_3_16_lpi_2;
  reg [15:0] psum_reg_4_16_lpi_2;
  reg [15:0] psum_reg_5_16_lpi_2;
  reg [15:0] psum_reg_6_16_lpi_2;
  reg [15:0] psum_reg_7_16_lpi_2;
  reg [15:0] psum_reg_8_16_lpi_2;
  reg [15:0] psum_reg_9_16_lpi_2;
  reg [15:0] psum_reg_10_16_lpi_2;
  reg [15:0] psum_reg_11_16_lpi_2;
  reg [15:0] psum_reg_12_16_lpi_2;
  reg [15:0] psum_reg_13_16_lpi_2;
  reg [15:0] psum_reg_14_16_lpi_2;
  reg [7:0] weight_reg_15_15_lpi_2;
  reg [7:0] weight_reg_15_14_lpi_2;
  reg [7:0] weight_reg_15_13_lpi_2;
  reg [7:0] weight_reg_15_10_lpi_2;
  reg [7:0] weight_reg_15_11_lpi_2;
  reg [7:0] weight_reg_15_12_lpi_2;
  reg [7:0] weight_reg_0_0_lpi_2;
  reg [7:0] weight_reg_1_0_lpi_2;
  reg [7:0] weight_reg_2_0_lpi_2;
  reg [7:0] weight_reg_3_0_lpi_2;
  reg [7:0] weight_reg_4_0_lpi_2;
  reg [7:0] weight_reg_5_0_lpi_2;
  reg [7:0] weight_reg_6_0_lpi_2;
  reg [7:0] weight_reg_7_0_lpi_2;
  reg [7:0] weight_reg_8_0_lpi_2;
  reg [7:0] weight_reg_9_0_lpi_2;
  reg [7:0] weight_reg_10_0_lpi_2;
  reg [7:0] weight_reg_11_0_lpi_2;
  reg [7:0] weight_reg_12_0_lpi_2;
  reg [7:0] weight_reg_13_0_lpi_2;
  reg [7:0] weight_reg_14_0_lpi_2;
  reg [7:0] weight_reg_15_0_lpi_2;
  reg [7:0] weight_reg_0_1_lpi_2;
  reg [7:0] weight_reg_1_1_lpi_2;
  reg [7:0] weight_reg_2_1_lpi_2;
  reg [7:0] weight_reg_3_1_lpi_2;
  reg [7:0] weight_reg_4_1_lpi_2;
  reg [7:0] weight_reg_5_1_lpi_2;
  reg [7:0] weight_reg_6_1_lpi_2;
  reg [7:0] weight_reg_7_1_lpi_2;
  reg [7:0] weight_reg_8_1_lpi_2;
  reg [7:0] weight_reg_9_1_lpi_2;
  reg [7:0] weight_reg_10_1_lpi_2;
  reg [7:0] weight_reg_11_1_lpi_2;
  reg [7:0] weight_reg_12_1_lpi_2;
  reg [7:0] weight_reg_13_1_lpi_2;
  reg [7:0] weight_reg_14_1_lpi_2;
  reg [7:0] weight_reg_15_1_lpi_2;
  reg [7:0] weight_reg_0_2_lpi_2;
  reg [7:0] weight_reg_1_2_lpi_2;
  reg [7:0] weight_reg_2_2_lpi_2;
  reg [7:0] weight_reg_3_2_lpi_2;
  reg [7:0] weight_reg_4_2_lpi_2;
  reg [7:0] weight_reg_5_2_lpi_2;
  reg [7:0] weight_reg_6_2_lpi_2;
  reg [7:0] weight_reg_7_2_lpi_2;
  reg [7:0] weight_reg_8_2_lpi_2;
  reg [7:0] weight_reg_9_2_lpi_2;
  reg [7:0] weight_reg_10_2_lpi_2;
  reg [7:0] weight_reg_11_2_lpi_2;
  reg [7:0] weight_reg_12_2_lpi_2;
  reg [7:0] weight_reg_13_2_lpi_2;
  reg [7:0] weight_reg_14_2_lpi_2;
  reg [7:0] weight_reg_15_2_lpi_2;
  reg [7:0] weight_reg_0_3_lpi_2;
  reg [7:0] weight_reg_1_3_lpi_2;
  reg [7:0] weight_reg_2_3_lpi_2;
  reg [7:0] weight_reg_3_3_lpi_2;
  reg [7:0] weight_reg_4_3_lpi_2;
  reg [7:0] weight_reg_5_3_lpi_2;
  reg [7:0] weight_reg_6_3_lpi_2;
  reg [7:0] weight_reg_7_3_lpi_2;
  reg [7:0] weight_reg_8_3_lpi_2;
  reg [7:0] weight_reg_9_3_lpi_2;
  reg [7:0] weight_reg_10_3_lpi_2;
  reg [7:0] weight_reg_11_3_lpi_2;
  reg [7:0] weight_reg_12_3_lpi_2;
  reg [7:0] weight_reg_13_3_lpi_2;
  reg [7:0] weight_reg_14_3_lpi_2;
  reg [7:0] weight_reg_15_3_lpi_2;
  reg [7:0] weight_reg_0_4_lpi_2;
  reg [7:0] weight_reg_1_4_lpi_2;
  reg [7:0] weight_reg_2_4_lpi_2;
  reg [7:0] weight_reg_3_4_lpi_2;
  reg [7:0] weight_reg_4_4_lpi_2;
  reg [7:0] weight_reg_5_4_lpi_2;
  reg [7:0] weight_reg_6_4_lpi_2;
  reg [7:0] weight_reg_7_4_lpi_2;
  reg [7:0] weight_reg_8_4_lpi_2;
  reg [7:0] weight_reg_9_4_lpi_2;
  reg [7:0] weight_reg_10_4_lpi_2;
  reg [7:0] weight_reg_11_4_lpi_2;
  reg [7:0] weight_reg_12_4_lpi_2;
  reg [7:0] weight_reg_13_4_lpi_2;
  reg [7:0] weight_reg_14_4_lpi_2;
  reg [7:0] weight_reg_15_4_lpi_2;
  reg [7:0] weight_reg_0_5_lpi_2;
  reg [7:0] weight_reg_1_5_lpi_2;
  reg [7:0] weight_reg_2_5_lpi_2;
  reg [7:0] weight_reg_3_5_lpi_2;
  reg [7:0] weight_reg_4_5_lpi_2;
  reg [7:0] weight_reg_5_5_lpi_2;
  reg [7:0] weight_reg_6_5_lpi_2;
  reg [7:0] weight_reg_7_5_lpi_2;
  reg [7:0] weight_reg_8_5_lpi_2;
  reg [7:0] weight_reg_9_5_lpi_2;
  reg [7:0] weight_reg_10_5_lpi_2;
  reg [7:0] weight_reg_11_5_lpi_2;
  reg [7:0] weight_reg_12_5_lpi_2;
  reg [7:0] weight_reg_13_5_lpi_2;
  reg [7:0] weight_reg_14_5_lpi_2;
  reg [7:0] weight_reg_15_5_lpi_2;
  reg [7:0] weight_reg_0_6_lpi_2;
  reg [7:0] weight_reg_1_6_lpi_2;
  reg [7:0] weight_reg_2_6_lpi_2;
  reg [7:0] weight_reg_3_6_lpi_2;
  reg [7:0] weight_reg_4_6_lpi_2;
  reg [7:0] weight_reg_5_6_lpi_2;
  reg [7:0] weight_reg_6_6_lpi_2;
  reg [7:0] weight_reg_7_6_lpi_2;
  reg [7:0] weight_reg_8_6_lpi_2;
  reg [7:0] weight_reg_9_6_lpi_2;
  reg [7:0] weight_reg_10_6_lpi_2;
  reg [7:0] weight_reg_11_6_lpi_2;
  reg [7:0] weight_reg_12_6_lpi_2;
  reg [7:0] weight_reg_13_6_lpi_2;
  reg [7:0] weight_reg_14_6_lpi_2;
  reg [7:0] weight_reg_15_6_lpi_2;
  reg [7:0] weight_reg_0_7_lpi_2;
  reg [7:0] weight_reg_1_7_lpi_2;
  reg [7:0] weight_reg_2_7_lpi_2;
  reg [7:0] weight_reg_3_7_lpi_2;
  reg [7:0] weight_reg_4_7_lpi_2;
  reg [7:0] weight_reg_5_7_lpi_2;
  reg [7:0] weight_reg_6_7_lpi_2;
  reg [7:0] weight_reg_7_7_lpi_2;
  reg [7:0] weight_reg_8_7_lpi_2;
  reg [7:0] weight_reg_9_7_lpi_2;
  reg [7:0] weight_reg_10_7_lpi_2;
  reg [7:0] weight_reg_11_7_lpi_2;
  reg [7:0] weight_reg_12_7_lpi_2;
  reg [7:0] weight_reg_13_7_lpi_2;
  reg [7:0] weight_reg_14_7_lpi_2;
  reg [7:0] weight_reg_15_7_lpi_2;
  reg [7:0] weight_reg_0_8_lpi_2;
  reg [7:0] weight_reg_1_8_lpi_2;
  reg [7:0] weight_reg_2_8_lpi_2;
  reg [7:0] weight_reg_3_8_lpi_2;
  reg [7:0] weight_reg_4_8_lpi_2;
  reg [7:0] weight_reg_5_8_lpi_2;
  reg [7:0] weight_reg_6_8_lpi_2;
  reg [7:0] weight_reg_7_8_lpi_2;
  reg [7:0] weight_reg_8_8_lpi_2;
  reg [7:0] weight_reg_9_8_lpi_2;
  reg [7:0] weight_reg_10_8_lpi_2;
  reg [7:0] weight_reg_11_8_lpi_2;
  reg [7:0] weight_reg_12_8_lpi_2;
  reg [7:0] weight_reg_13_8_lpi_2;
  reg [7:0] weight_reg_14_8_lpi_2;
  reg [7:0] weight_reg_15_8_lpi_2;
  reg [7:0] weight_reg_0_9_lpi_2;
  reg [7:0] weight_reg_1_9_lpi_2;
  reg [7:0] weight_reg_2_9_lpi_2;
  reg [7:0] weight_reg_3_9_lpi_2;
  reg [7:0] weight_reg_4_9_lpi_2;
  reg [7:0] weight_reg_5_9_lpi_2;
  reg [7:0] weight_reg_6_9_lpi_2;
  reg [7:0] weight_reg_7_9_lpi_2;
  reg [7:0] weight_reg_8_9_lpi_2;
  reg [7:0] weight_reg_9_9_lpi_2;
  reg [7:0] weight_reg_10_9_lpi_2;
  reg [7:0] weight_reg_11_9_lpi_2;
  reg [7:0] weight_reg_12_9_lpi_2;
  reg [7:0] weight_reg_13_9_lpi_2;
  reg [7:0] weight_reg_14_9_lpi_2;
  reg [7:0] weight_reg_15_9_lpi_2;
  reg [7:0] weight_reg_0_10_lpi_2;
  reg [7:0] weight_reg_1_10_lpi_2;
  reg [7:0] weight_reg_2_10_lpi_2;
  reg [7:0] weight_reg_3_10_lpi_2;
  reg [7:0] weight_reg_4_10_lpi_2;
  reg [7:0] weight_reg_5_10_lpi_2;
  reg [7:0] weight_reg_6_10_lpi_2;
  reg [7:0] weight_reg_7_10_lpi_2;
  reg [7:0] weight_reg_8_10_lpi_2;
  reg [7:0] weight_reg_9_10_lpi_2;
  reg [7:0] weight_reg_10_10_lpi_2;
  reg [7:0] weight_reg_11_10_lpi_2;
  reg [7:0] weight_reg_12_10_lpi_2;
  reg [7:0] weight_reg_13_10_lpi_2;
  reg [7:0] weight_reg_14_10_lpi_2;
  reg [7:0] weight_reg_0_11_lpi_2;
  reg [7:0] weight_reg_1_11_lpi_2;
  reg [7:0] weight_reg_2_11_lpi_2;
  reg [7:0] weight_reg_3_11_lpi_2;
  reg [7:0] weight_reg_4_11_lpi_2;
  reg [7:0] weight_reg_5_11_lpi_2;
  reg [7:0] weight_reg_6_11_lpi_2;
  reg [7:0] weight_reg_7_11_lpi_2;
  reg [7:0] weight_reg_8_11_lpi_2;
  reg [7:0] weight_reg_9_11_lpi_2;
  reg [7:0] weight_reg_10_11_lpi_2;
  reg [7:0] weight_reg_11_11_lpi_2;
  reg [7:0] weight_reg_12_11_lpi_2;
  reg [7:0] weight_reg_13_11_lpi_2;
  reg [7:0] weight_reg_14_11_lpi_2;
  reg [7:0] weight_reg_0_12_lpi_2;
  reg [7:0] weight_reg_1_12_lpi_2;
  reg [7:0] weight_reg_2_12_lpi_2;
  reg [7:0] weight_reg_3_12_lpi_2;
  reg [7:0] weight_reg_4_12_lpi_2;
  reg [7:0] weight_reg_5_12_lpi_2;
  reg [7:0] weight_reg_6_12_lpi_2;
  reg [7:0] weight_reg_7_12_lpi_2;
  reg [7:0] weight_reg_8_12_lpi_2;
  reg [7:0] weight_reg_9_12_lpi_2;
  reg [7:0] weight_reg_10_12_lpi_2;
  reg [7:0] weight_reg_11_12_lpi_2;
  reg [7:0] weight_reg_12_12_lpi_2;
  reg [7:0] weight_reg_13_12_lpi_2;
  reg [7:0] weight_reg_14_12_lpi_2;
  reg [7:0] weight_reg_0_13_lpi_2;
  reg [7:0] weight_reg_1_13_lpi_2;
  reg [7:0] weight_reg_2_13_lpi_2;
  reg [7:0] weight_reg_3_13_lpi_2;
  reg [7:0] weight_reg_4_13_lpi_2;
  reg [7:0] weight_reg_5_13_lpi_2;
  reg [7:0] weight_reg_6_13_lpi_2;
  reg [7:0] weight_reg_7_13_lpi_2;
  reg [7:0] weight_reg_8_13_lpi_2;
  reg [7:0] weight_reg_9_13_lpi_2;
  reg [7:0] weight_reg_10_13_lpi_2;
  reg [7:0] weight_reg_11_13_lpi_2;
  reg [7:0] weight_reg_12_13_lpi_2;
  reg [7:0] weight_reg_13_13_lpi_2;
  reg [7:0] weight_reg_14_13_lpi_2;
  reg [7:0] weight_reg_0_14_lpi_2;
  reg [7:0] weight_reg_1_14_lpi_2;
  reg [7:0] weight_reg_2_14_lpi_2;
  reg [7:0] weight_reg_3_14_lpi_2;
  reg [7:0] weight_reg_4_14_lpi_2;
  reg [7:0] weight_reg_5_14_lpi_2;
  reg [7:0] weight_reg_6_14_lpi_2;
  reg [7:0] weight_reg_7_14_lpi_2;
  reg [7:0] weight_reg_8_14_lpi_2;
  reg [7:0] weight_reg_9_14_lpi_2;
  reg [7:0] weight_reg_10_14_lpi_2;
  reg [7:0] weight_reg_11_14_lpi_2;
  reg [7:0] weight_reg_12_14_lpi_2;
  reg [7:0] weight_reg_13_14_lpi_2;
  reg [7:0] weight_reg_14_14_lpi_2;
  reg [7:0] weight_reg_0_15_lpi_2;
  reg [7:0] weight_reg_1_15_lpi_2;
  reg [7:0] weight_reg_2_15_lpi_2;
  reg [7:0] weight_reg_3_15_lpi_2;
  reg [7:0] weight_reg_4_15_lpi_2;
  reg [7:0] weight_reg_5_15_lpi_2;
  reg [7:0] weight_reg_6_15_lpi_2;
  reg [7:0] weight_reg_7_15_lpi_2;
  reg [7:0] weight_reg_8_15_lpi_2;
  reg [7:0] weight_reg_9_15_lpi_2;
  reg [7:0] weight_reg_10_15_lpi_2;
  reg [7:0] weight_reg_11_15_lpi_2;
  reg [7:0] weight_reg_12_15_lpi_2;
  reg [7:0] weight_reg_13_15_lpi_2;
  reg [7:0] weight_reg_14_15_lpi_2;
  wire mux_302_itm;
  reg [127:0] step_in_col_value_lpi_2;
  reg [7:0] input_reg_1_1_lpi_2;
  reg [7:0] input_reg_2_1_lpi_2;
  reg [7:0] input_reg_3_1_lpi_2;
  reg [7:0] input_reg_4_1_lpi_2;
  reg [7:0] input_reg_5_1_lpi_2;
  reg [7:0] input_reg_6_1_lpi_2;
  reg [7:0] input_reg_7_1_lpi_2;
  reg [7:0] input_reg_8_1_lpi_2;
  reg [7:0] input_reg_9_1_lpi_2;
  reg [7:0] input_reg_10_1_lpi_2;
  reg [7:0] input_reg_11_1_lpi_2;
  reg [7:0] input_reg_12_1_lpi_2;
  reg [7:0] input_reg_13_1_lpi_2;
  reg [7:0] input_reg_14_1_lpi_2;
  reg [7:0] input_reg_15_1_lpi_2;
  reg [7:0] input_reg_16_1_lpi_2;
  reg [7:0] input_reg_1_2_lpi_2;
  reg [7:0] input_reg_2_2_lpi_2;
  reg [7:0] input_reg_3_2_lpi_2;
  reg [7:0] input_reg_4_2_lpi_2;
  reg [7:0] input_reg_5_2_lpi_2;
  reg [7:0] input_reg_6_2_lpi_2;
  reg [7:0] input_reg_7_2_lpi_2;
  reg [7:0] input_reg_8_2_lpi_2;
  reg [7:0] input_reg_9_2_lpi_2;
  reg [7:0] input_reg_10_2_lpi_2;
  reg [7:0] input_reg_11_2_lpi_2;
  reg [7:0] input_reg_12_2_lpi_2;
  reg [7:0] input_reg_13_2_lpi_2;
  reg [7:0] input_reg_14_2_lpi_2;
  reg [7:0] input_reg_15_2_lpi_2;
  reg [7:0] input_reg_16_2_lpi_2;
  reg [7:0] input_reg_1_3_lpi_2;
  reg [7:0] input_reg_2_3_lpi_2;
  reg [7:0] input_reg_3_3_lpi_2;
  reg [7:0] input_reg_4_3_lpi_2;
  reg [7:0] input_reg_5_3_lpi_2;
  reg [7:0] input_reg_6_3_lpi_2;
  reg [7:0] input_reg_7_3_lpi_2;
  reg [7:0] input_reg_8_3_lpi_2;
  reg [7:0] input_reg_9_3_lpi_2;
  reg [7:0] input_reg_10_3_lpi_2;
  reg [7:0] input_reg_11_3_lpi_2;
  reg [7:0] input_reg_12_3_lpi_2;
  reg [7:0] input_reg_13_3_lpi_2;
  reg [7:0] input_reg_14_3_lpi_2;
  reg [7:0] input_reg_15_3_lpi_2;
  reg [7:0] input_reg_16_3_lpi_2;
  reg [7:0] input_reg_1_4_lpi_2;
  reg [7:0] input_reg_2_4_lpi_2;
  reg [7:0] input_reg_3_4_lpi_2;
  reg [7:0] input_reg_4_4_lpi_2;
  reg [7:0] input_reg_5_4_lpi_2;
  reg [7:0] input_reg_6_4_lpi_2;
  reg [7:0] input_reg_7_4_lpi_2;
  reg [7:0] input_reg_8_4_lpi_2;
  reg [7:0] input_reg_9_4_lpi_2;
  reg [7:0] input_reg_10_4_lpi_2;
  reg [7:0] input_reg_11_4_lpi_2;
  reg [7:0] input_reg_12_4_lpi_2;
  reg [7:0] input_reg_13_4_lpi_2;
  reg [7:0] input_reg_14_4_lpi_2;
  reg [7:0] input_reg_15_4_lpi_2;
  reg [7:0] input_reg_16_4_lpi_2;
  reg [7:0] input_reg_1_5_lpi_2;
  reg [7:0] input_reg_2_5_lpi_2;
  reg [7:0] input_reg_3_5_lpi_2;
  reg [7:0] input_reg_4_5_lpi_2;
  reg [7:0] input_reg_5_5_lpi_2;
  reg [7:0] input_reg_6_5_lpi_2;
  reg [7:0] input_reg_7_5_lpi_2;
  reg [7:0] input_reg_8_5_lpi_2;
  reg [7:0] input_reg_9_5_lpi_2;
  reg [7:0] input_reg_10_5_lpi_2;
  reg [7:0] input_reg_11_5_lpi_2;
  reg [7:0] input_reg_12_5_lpi_2;
  reg [7:0] input_reg_13_5_lpi_2;
  reg [7:0] input_reg_14_5_lpi_2;
  reg [7:0] input_reg_15_5_lpi_2;
  reg [7:0] input_reg_16_5_lpi_2;
  reg [7:0] input_reg_1_6_lpi_2;
  reg [7:0] input_reg_2_6_lpi_2;
  reg [7:0] input_reg_3_6_lpi_2;
  reg [7:0] input_reg_4_6_lpi_2;
  reg [7:0] input_reg_5_6_lpi_2;
  reg [7:0] input_reg_6_6_lpi_2;
  reg [7:0] input_reg_7_6_lpi_2;
  reg [7:0] input_reg_8_6_lpi_2;
  reg [7:0] input_reg_9_6_lpi_2;
  reg [7:0] input_reg_10_6_lpi_2;
  reg [7:0] input_reg_11_6_lpi_2;
  reg [7:0] input_reg_12_6_lpi_2;
  reg [7:0] input_reg_13_6_lpi_2;
  reg [7:0] input_reg_14_6_lpi_2;
  reg [7:0] input_reg_15_6_lpi_2;
  reg [7:0] input_reg_16_6_lpi_2;
  reg [7:0] input_reg_1_7_lpi_2;
  reg [7:0] input_reg_2_7_lpi_2;
  reg [7:0] input_reg_3_7_lpi_2;
  reg [7:0] input_reg_4_7_lpi_2;
  reg [7:0] input_reg_5_7_lpi_2;
  reg [7:0] input_reg_6_7_lpi_2;
  reg [7:0] input_reg_7_7_lpi_2;
  reg [7:0] input_reg_8_7_lpi_2;
  reg [7:0] input_reg_9_7_lpi_2;
  reg [7:0] input_reg_10_7_lpi_2;
  reg [7:0] input_reg_11_7_lpi_2;
  reg [7:0] input_reg_12_7_lpi_2;
  reg [7:0] input_reg_13_7_lpi_2;
  reg [7:0] input_reg_14_7_lpi_2;
  reg [7:0] input_reg_15_7_lpi_2;
  reg [7:0] input_reg_16_7_lpi_2;
  reg [7:0] input_reg_1_8_lpi_2;
  reg [7:0] input_reg_2_8_lpi_2;
  reg [7:0] input_reg_3_8_lpi_2;
  reg [7:0] input_reg_4_8_lpi_2;
  reg [7:0] input_reg_5_8_lpi_2;
  reg [7:0] input_reg_6_8_lpi_2;
  reg [7:0] input_reg_7_8_lpi_2;
  reg [7:0] input_reg_8_8_lpi_2;
  reg [7:0] input_reg_9_8_lpi_2;
  reg [7:0] input_reg_10_8_lpi_2;
  reg [7:0] input_reg_11_8_lpi_2;
  reg [7:0] input_reg_12_8_lpi_2;
  reg [7:0] input_reg_13_8_lpi_2;
  reg [7:0] input_reg_14_8_lpi_2;
  reg [7:0] input_reg_15_8_lpi_2;
  reg [7:0] input_reg_16_8_lpi_2;
  reg [7:0] input_reg_1_9_lpi_2;
  reg [7:0] input_reg_2_9_lpi_2;
  reg [7:0] input_reg_3_9_lpi_2;
  reg [7:0] input_reg_4_9_lpi_2;
  reg [7:0] input_reg_5_9_lpi_2;
  reg [7:0] input_reg_6_9_lpi_2;
  reg [7:0] input_reg_7_9_lpi_2;
  reg [7:0] input_reg_8_9_lpi_2;
  reg [7:0] input_reg_9_9_lpi_2;
  reg [7:0] input_reg_10_9_lpi_2;
  reg [7:0] input_reg_11_9_lpi_2;
  reg [7:0] input_reg_12_9_lpi_2;
  reg [7:0] input_reg_13_9_lpi_2;
  reg [7:0] input_reg_14_9_lpi_2;
  reg [7:0] input_reg_15_9_lpi_2;
  reg [7:0] input_reg_16_9_lpi_2;
  reg [7:0] input_reg_1_10_lpi_2;
  reg [7:0] input_reg_2_10_lpi_2;
  reg [7:0] input_reg_3_10_lpi_2;
  reg [7:0] input_reg_4_10_lpi_2;
  reg [7:0] input_reg_5_10_lpi_2;
  reg [7:0] input_reg_6_10_lpi_2;
  reg [7:0] input_reg_7_10_lpi_2;
  reg [7:0] input_reg_8_10_lpi_2;
  reg [7:0] input_reg_9_10_lpi_2;
  reg [7:0] input_reg_10_10_lpi_2;
  reg [7:0] input_reg_11_10_lpi_2;
  reg [7:0] input_reg_12_10_lpi_2;
  reg [7:0] input_reg_13_10_lpi_2;
  reg [7:0] input_reg_14_10_lpi_2;
  reg [7:0] input_reg_15_10_lpi_2;
  reg [7:0] input_reg_1_11_lpi_2;
  reg [7:0] input_reg_2_11_lpi_2;
  reg [7:0] input_reg_3_11_lpi_2;
  reg [7:0] input_reg_4_11_lpi_2;
  reg [7:0] input_reg_5_11_lpi_2;
  reg [7:0] input_reg_6_11_lpi_2;
  reg [7:0] input_reg_7_11_lpi_2;
  reg [7:0] input_reg_8_11_lpi_2;
  reg [7:0] input_reg_9_11_lpi_2;
  reg [7:0] input_reg_10_11_lpi_2;
  reg [7:0] input_reg_11_11_lpi_2;
  reg [7:0] input_reg_12_11_lpi_2;
  reg [7:0] input_reg_13_11_lpi_2;
  reg [7:0] input_reg_14_11_lpi_2;
  reg [7:0] input_reg_15_11_lpi_2;
  reg [7:0] input_reg_1_12_lpi_2;
  reg [7:0] input_reg_2_12_lpi_2;
  reg [7:0] input_reg_3_12_lpi_2;
  reg [7:0] input_reg_4_12_lpi_2;
  reg [7:0] input_reg_5_12_lpi_2;
  reg [7:0] input_reg_6_12_lpi_2;
  reg [7:0] input_reg_7_12_lpi_2;
  reg [7:0] input_reg_8_12_lpi_2;
  reg [7:0] input_reg_9_12_lpi_2;
  reg [7:0] input_reg_10_12_lpi_2;
  reg [7:0] input_reg_11_12_lpi_2;
  reg [7:0] input_reg_12_12_lpi_2;
  reg [7:0] input_reg_13_12_lpi_2;
  reg [7:0] input_reg_14_12_lpi_2;
  reg [7:0] input_reg_15_12_lpi_2;
  reg [7:0] input_reg_1_13_lpi_2;
  reg [7:0] input_reg_2_13_lpi_2;
  reg [7:0] input_reg_3_13_lpi_2;
  reg [7:0] input_reg_4_13_lpi_2;
  reg [7:0] input_reg_5_13_lpi_2;
  reg [7:0] input_reg_6_13_lpi_2;
  reg [7:0] input_reg_7_13_lpi_2;
  reg [7:0] input_reg_8_13_lpi_2;
  reg [7:0] input_reg_9_13_lpi_2;
  reg [7:0] input_reg_10_13_lpi_2;
  reg [7:0] input_reg_11_13_lpi_2;
  reg [7:0] input_reg_12_13_lpi_2;
  reg [7:0] input_reg_13_13_lpi_2;
  reg [7:0] input_reg_14_13_lpi_2;
  reg [7:0] input_reg_15_13_lpi_2;
  reg [7:0] input_reg_1_14_lpi_2;
  reg [7:0] input_reg_2_14_lpi_2;
  reg [7:0] input_reg_3_14_lpi_2;
  reg [7:0] input_reg_4_14_lpi_2;
  reg [7:0] input_reg_5_14_lpi_2;
  reg [7:0] input_reg_6_14_lpi_2;
  reg [7:0] input_reg_7_14_lpi_2;
  reg [7:0] input_reg_8_14_lpi_2;
  reg [7:0] input_reg_9_14_lpi_2;
  reg [7:0] input_reg_10_14_lpi_2;
  reg [7:0] input_reg_11_14_lpi_2;
  reg [7:0] input_reg_12_14_lpi_2;
  reg [7:0] input_reg_13_14_lpi_2;
  reg [7:0] input_reg_14_14_lpi_2;
  reg [7:0] input_reg_15_14_lpi_2;
  reg [7:0] input_reg_1_15_lpi_2;
  reg [7:0] input_reg_2_15_lpi_2;
  reg [7:0] input_reg_3_15_lpi_2;
  reg [7:0] input_reg_4_15_lpi_2;
  reg [7:0] input_reg_5_15_lpi_2;
  reg [7:0] input_reg_6_15_lpi_2;
  reg [7:0] input_reg_7_15_lpi_2;
  reg [7:0] input_reg_8_15_lpi_2;
  reg [7:0] input_reg_9_15_lpi_2;
  reg [7:0] input_reg_10_15_lpi_2;
  reg [7:0] input_reg_11_15_lpi_2;
  reg [7:0] input_reg_12_15_lpi_2;
  reg [7:0] input_reg_13_15_lpi_2;
  reg [7:0] input_reg_14_15_lpi_2;
  reg [7:0] input_reg_15_15_lpi_2;
  reg [95:0] paramsIn_crt_sva_127_32;
  wire psum_reg_15_16_lpi_2_mx0c2;
  wire ROW_asn_142_itm_mx0c0;
  wire [16:0] operator_16_false_3_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_3_acc_psp_sva_1;
  wire [16:0] operator_16_false_2_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_2_acc_psp_sva_1;
  wire and_443_m1c;
  wire operator_16_false_and_1_cse;
  wire [31:0] step_mul_itm;
  wire step_if_1_acc_itm_32_1;
  wire operator_16_false_acc_itm_12_1;
  wire operator_32_false_acc_itm_31_1;

  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] or_137_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] or_250_nl;
  wire[0:0] or_258_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] or_225_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] or_223_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_329_nl;
  wire[0:0] nand_84_nl;
  wire[0:0] or_326_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] or_337_nl;
  wire[0:0] and_441_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] or_35_nl;
  wire[0:0] psum_reg_or_4_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] or_924_nl;
  wire[0:0] or_920_nl;
  wire[0:0] psum_reg_and_242_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] or_664_nl;
  wire[0:0] or_662_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] or_669_nl;
  wire[0:0] or_674_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] or_676_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] or_51_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_57_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] or_685_nl;
  wire[0:0] or_67_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] or_918_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] nand_28_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] and_461_nl;
  wire[0:0] nor_117_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] or_76_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] or_83_nl;
  wire[0:0] or_82_nl;
  wire[0:0] or_80_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] or_706_nl;
  wire[0:0] or_92_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] or_714_nl;
  wire[0:0] nand_2_nl;
  wire[7:0] step_input_fifo_input_15_mux_nl;
  wire[0:0] and_451_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] or_720_nl;
  wire[0:0] or_104_nl;
  wire[0:0] or_103_nl;
  wire[0:0] or_102_nl;
  wire[0:0] and_447_nl;
  wire[15:0] step_acc_3_nl;
  wire[16:0] nl_step_acc_3_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] and_460_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_168_nl;
  wire[0:0] or_729_nl;
  wire[0:0] or_727_nl;
  wire[15:0] step_step_mux_nl;
  wire[0:0] step_step_not_nl;
  wire[16:0] operator_16_false_acc_nl;
  wire[17:0] nl_operator_16_false_acc_nl;
  wire[5:0] operator_16_false_mux_1_nl;
  wire[5:0] step_if_3_for_1_operator_16_false_acc_nl;
  wire[6:0] nl_step_if_3_for_1_operator_16_false_acc_nl;
  wire[32:0] step_if_1_acc_nl;
  wire[34:0] nl_step_if_1_acc_nl;
  wire[12:0] operator_16_false_acc_nl_1;
  wire[13:0] nl_operator_16_false_acc_nl_1;
  wire[0:0] or_133_nl;
  wire[0:0] or_132_nl;
  wire[0:0] or_848_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] or_240_nl;
  wire[0:0] or_254_nl;
  wire[0:0] nand_121_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] or_264_nl;
  wire[0:0] or_270_nl;
  wire[0:0] or_269_nl;
  wire[0:0] or_297_nl;
  wire[0:0] or_318_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] or_906_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] and_472_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] mux_355_nl;
  wire[31:0] operator_32_false_acc_nl;
  wire[32:0] nl_operator_32_false_acc_nl;
  wire[32:0] operator_32_false_acc_1_nl;
  wire[33:0] nl_operator_32_false_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[0:0] step_if_2_aelse_1_not_33_nl;
  wire [15:0] nl_accum_fifo_15_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_33_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_15_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_15_i_dout_d_mxwt, (step_if_2_aelse_1_not_33_nl));
  wire [15:0] nl_output_fifo_0_rsci_input_rsc_dat;
  assign nl_output_fifo_0_rsci_input_rsc_dat = psum_reg_16_1_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_34_nl;
  wire [15:0] nl_accum_fifo_14_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_34_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_14_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_14_i_dout_d_mxwt, (step_if_2_aelse_1_not_34_nl));
  wire [15:0] nl_output_fifo_1_rsci_input_rsc_dat;
  assign nl_output_fifo_1_rsci_input_rsc_dat = psum_reg_16_2_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_35_nl;
  wire [15:0] nl_accum_fifo_13_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_35_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_13_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_13_i_dout_d_mxwt, (step_if_2_aelse_1_not_35_nl));
  wire [15:0] nl_output_fifo_2_rsci_input_rsc_dat;
  assign nl_output_fifo_2_rsci_input_rsc_dat = psum_reg_16_3_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_36_nl;
  wire [15:0] nl_accum_fifo_12_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_36_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_12_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_12_i_dout_d_mxwt, (step_if_2_aelse_1_not_36_nl));
  wire [15:0] nl_output_fifo_3_rsci_input_rsc_dat;
  assign nl_output_fifo_3_rsci_input_rsc_dat = psum_reg_16_4_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_37_nl;
  wire [15:0] nl_accum_fifo_11_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_37_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_11_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_11_i_dout_d_mxwt, (step_if_2_aelse_1_not_37_nl));
  wire [15:0] nl_output_fifo_4_rsci_input_rsc_dat;
  assign nl_output_fifo_4_rsci_input_rsc_dat = psum_reg_16_5_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_38_nl;
  wire [15:0] nl_accum_fifo_10_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_38_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_10_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_10_i_dout_d_mxwt, (step_if_2_aelse_1_not_38_nl));
  wire [15:0] nl_output_fifo_5_rsci_input_rsc_dat;
  assign nl_output_fifo_5_rsci_input_rsc_dat = psum_reg_16_6_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_39_nl;
  wire [15:0] nl_accum_fifo_9_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_39_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_9_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_9_i_dout_d_mxwt, (step_if_2_aelse_1_not_39_nl));
  wire [15:0] nl_output_fifo_6_rsci_input_rsc_dat;
  assign nl_output_fifo_6_rsci_input_rsc_dat = psum_reg_16_7_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_40_nl;
  wire [15:0] nl_accum_fifo_8_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_40_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_8_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_8_i_dout_d_mxwt, (step_if_2_aelse_1_not_40_nl));
  wire [15:0] nl_output_fifo_7_rsci_input_rsc_dat;
  assign nl_output_fifo_7_rsci_input_rsc_dat = psum_reg_16_8_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_41_nl;
  wire [15:0] nl_accum_fifo_7_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_41_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_7_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_7_i_dout_d_mxwt, (step_if_2_aelse_1_not_41_nl));
  wire [15:0] nl_output_fifo_8_rsci_input_rsc_dat;
  assign nl_output_fifo_8_rsci_input_rsc_dat = psum_reg_16_9_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_42_nl;
  wire [15:0] nl_accum_fifo_6_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_42_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_6_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_6_i_dout_d_mxwt, (step_if_2_aelse_1_not_42_nl));
  wire [15:0] nl_output_fifo_9_rsci_input_rsc_dat;
  assign nl_output_fifo_9_rsci_input_rsc_dat = psum_reg_16_10_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_43_nl;
  wire [15:0] nl_accum_fifo_5_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_43_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_5_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_5_i_dout_d_mxwt, (step_if_2_aelse_1_not_43_nl));
  wire [15:0] nl_output_fifo_10_rsci_input_rsc_dat;
  assign nl_output_fifo_10_rsci_input_rsc_dat = psum_reg_16_11_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_44_nl;
  wire [15:0] nl_accum_fifo_4_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_44_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_4_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_4_i_dout_d_mxwt, (step_if_2_aelse_1_not_44_nl));
  wire [15:0] nl_output_fifo_11_rsci_input_rsc_dat;
  assign nl_output_fifo_11_rsci_input_rsc_dat = psum_reg_16_12_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_45_nl;
  wire [15:0] nl_accum_fifo_3_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_45_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_3_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_3_i_dout_d_mxwt, (step_if_2_aelse_1_not_45_nl));
  wire [15:0] nl_output_fifo_12_rsci_input_rsc_dat;
  assign nl_output_fifo_12_rsci_input_rsc_dat = step_output_buf_value_0_sva;
  wire[0:0] step_if_2_aelse_1_not_46_nl;
  wire [15:0] nl_accum_fifo_2_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_46_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_2_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_2_i_dout_d_mxwt, (step_if_2_aelse_1_not_46_nl));
  wire [15:0] nl_output_fifo_13_rsci_input_rsc_dat;
  assign nl_output_fifo_13_rsci_input_rsc_dat = psum_reg_16_14_lpi_2;
  wire[0:0] step_if_2_aelse_1_not_47_nl;
  wire [15:0] nl_accum_fifo_1_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_47_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign nl_accum_fifo_1_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_1_i_dout_d_mxwt, (step_if_2_aelse_1_not_47_nl));
  wire [15:0] nl_output_fifo_14_rsci_input_rsc_dat;
  assign nl_output_fifo_14_rsci_input_rsc_dat = psum_reg_16_15_lpi_2;
  wire [7:0] nl_input_fifo_15_rsci_input_rsc_dat;
  assign nl_input_fifo_15_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[127:120];
  wire [7:0] nl_input_fifo_14_rsci_input_rsc_dat;
  assign nl_input_fifo_14_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[119:112];
  wire [7:0] nl_input_fifo_13_rsci_input_rsc_dat;
  assign nl_input_fifo_13_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[111:104];
  wire [7:0] nl_input_fifo_12_rsci_input_rsc_dat;
  assign nl_input_fifo_12_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[103:96];
  wire [7:0] nl_input_fifo_11_rsci_input_rsc_dat;
  assign nl_input_fifo_11_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[95:88];
  wire [7:0] nl_input_fifo_10_rsci_input_rsc_dat;
  assign nl_input_fifo_10_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[87:80];
  wire [7:0] nl_input_fifo_9_rsci_input_rsc_dat;
  assign nl_input_fifo_9_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[79:72];
  wire [7:0] nl_input_fifo_8_rsci_input_rsc_dat;
  assign nl_input_fifo_8_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[71:64];
  wire [7:0] nl_input_fifo_7_rsci_input_rsc_dat;
  assign nl_input_fifo_7_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[63:56];
  wire [7:0] nl_input_fifo_6_rsci_input_rsc_dat;
  assign nl_input_fifo_6_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[55:48];
  wire [7:0] nl_input_fifo_5_rsci_input_rsc_dat;
  assign nl_input_fifo_5_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[47:40];
  wire [7:0] nl_input_fifo_4_rsci_input_rsc_dat;
  assign nl_input_fifo_4_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[39:32];
  wire [7:0] nl_input_fifo_3_rsci_input_rsc_dat;
  assign nl_input_fifo_3_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[31:24];
  wire [7:0] nl_input_fifo_2_rsci_input_rsc_dat;
  assign nl_input_fifo_2_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[23:16];
  wire [7:0] nl_input_fifo_1_rsci_input_rsc_dat;
  assign nl_input_fifo_1_rsci_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[15:8];
  wire[0:0] nor_206_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] or_163_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] or_162_nl;
  wire[0:0] or_161_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] or_159_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] or_155_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] nor_144_nl;
  wire[0:0] or_167_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] or_166_nl;
  wire[0:0] nor_204_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] nor_202_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] or_194_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] nor_201_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] or_199_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] or_198_nl;
  wire[0:0] nor_200_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] or_214_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] or_213_nl;
  wire[0:0] or_212_nl;
  wire[0:0] or_921_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] or_922_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_186_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] or_207_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] nor_199_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] or_219_nl;
  wire[0:0] nor_198_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] nand_16_nl;
  wire[0:0] nor_197_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] or_248_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] nand_132_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] or_245_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] or_241_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] or_238_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] nor_196_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] or_938_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] or_261_nl;
  wire[0:0] nand_124_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] or_256_nl;
  wire[0:0] nand_18_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] or_939_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] or_283_nl;
  wire[0:0] or_282_nl;
  wire[0:0] or_280_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] nor_138_nl;
  wire[0:0] nor_139_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] or_274_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] or_272_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] or_271_nl;
  wire[0:0] or_267_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] or_300_nl;
  wire[0:0] nand_21_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] or_298_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] or_296_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] or_295_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] or_293_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] or_290_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] or_289_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] or_285_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] or_313_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] or_312_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] or_308_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] or_304_nl;
  wire[0:0] or_301_nl;
  wire[0:0] nor_195_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] nand_122_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] nand_123_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] or_936_nl;
  wire[0:0] or_937_nl;
  wire [7:0] nl_pe_0_0_run_cmp_input_in_rsc_dat;
  assign or_162_nl = (fsm_output[6]) | (fsm_output[7]) | (fsm_output[2]);
  assign mux_119_nl = MUX_s_1_2_2(mux_tmp_93, (or_162_nl), fsm_output[3]);
  assign nand_4_nl = ~((fsm_output[5]) & (~ (mux_119_nl)));
  assign or_161_nl = (fsm_output[5]) | (fsm_output[3]) | mux_tmp_93;
  assign mux_120_nl = MUX_s_1_2_2((nand_4_nl), (or_161_nl), fsm_output[1]);
  assign or_163_nl = (fsm_output[4]) | (mux_120_nl);
  assign or_159_nl = (fsm_output[5]) | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[2]);
  assign nand_113_nl = ~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]) & (~
      (fsm_output[2])));
  assign mux_116_nl = MUX_s_1_2_2((nand_113_nl), mux_tmp_91, fsm_output[5]);
  assign mux_117_nl = MUX_s_1_2_2((or_159_nl), (mux_116_nl), fsm_output[1]);
  assign mux_113_nl = MUX_s_1_2_2(mux_tmp_93, mux_111_cse, fsm_output[3]);
  assign mux_114_nl = MUX_s_1_2_2((mux_113_nl), mux_tmp_91, fsm_output[5]);
  assign or_155_nl = (~ (fsm_output[5])) | (fsm_output[3]) | mux_109_cse;
  assign mux_115_nl = MUX_s_1_2_2((mux_114_nl), (or_155_nl), fsm_output[1]);
  assign mux_118_nl = MUX_s_1_2_2((mux_117_nl), (mux_115_nl), fsm_output[4]);
  assign mux_121_nl = MUX_s_1_2_2((or_163_nl), (mux_118_nl), fsm_output[0]);
  assign nor_206_nl = ~((mux_121_nl) | (fsm_output[8]));
  assign mux_126_nl = MUX_s_1_2_2(mux_tmp_103, (~ nor_tmp_20), fsm_output[6]);
  assign mux_127_nl = MUX_s_1_2_2((mux_126_nl), or_187_cse, fsm_output[2]);
  assign nor_144_nl = ~((~ (fsm_output[7])) | (fsm_output[3]));
  assign mux_125_nl = MUX_s_1_2_2(nor_tmp_20, (nor_144_nl), fsm_output[6]);
  assign nand_6_nl = ~((fsm_output[2]) & (mux_125_nl));
  assign mux_128_nl = MUX_s_1_2_2((mux_127_nl), (nand_6_nl), fsm_output[5]);
  assign mux_129_nl = MUX_s_1_2_2(nand_tmp_5, (mux_128_nl), fsm_output[1]);
  assign mux_131_nl = MUX_s_1_2_2(or_170_cse, (mux_129_nl), fsm_output[4]);
  assign or_166_nl = (fsm_output[5]) | mux_377_cse;
  assign mux_124_nl = MUX_s_1_2_2(nand_tmp_5, (or_166_nl), fsm_output[1]);
  assign or_167_nl = (fsm_output[4]) | (mux_124_nl);
  assign mux_132_nl = MUX_s_1_2_2((mux_131_nl), (or_167_nl), fsm_output[0]);
  assign nor_205_nl = ~((mux_132_nl) | (fsm_output[8]));
  assign mux_134_nl = MUX_s_1_2_2(or_827_cse, (~ mux_434_cse), fsm_output[7]);
  assign mux_135_nl = MUX_s_1_2_2((mux_134_nl), or_187_cse, fsm_output[2]);
  assign nand_7_nl = ~((fsm_output[2]) & (fsm_output[7]) & (~ mux_434_cse));
  assign mux_136_nl = MUX_s_1_2_2((mux_135_nl), (nand_7_nl), fsm_output[5]);
  assign mux_139_nl = MUX_s_1_2_2(nand_10_cse, (mux_136_nl), fsm_output[1]);
  assign mux_141_nl = MUX_s_1_2_2(or_170_cse, (mux_139_nl), fsm_output[4]);
  assign mux_144_nl = MUX_s_1_2_2(or_178_cse, (mux_141_nl), fsm_output[0]);
  assign nor_204_nl = ~((mux_144_nl) | (fsm_output[8]));
  assign mux_157_nl = MUX_s_1_2_2(mux_156_cse, or_178_cse, fsm_output[0]);
  assign nor_203_nl = ~((mux_157_nl) | (fsm_output[8]));
  assign nand_11_nl = ~((fsm_output[5]) & (~ mux_142_cse));
  assign mux_169_nl = MUX_s_1_2_2((nand_11_nl), or_177_cse, fsm_output[1]);
  assign or_194_nl = (fsm_output[4]) | (mux_169_nl);
  assign mux_170_nl = MUX_s_1_2_2((or_194_nl), mux_156_cse, fsm_output[0]);
  assign nor_202_nl = ~((mux_170_nl) | (fsm_output[8]));
  assign nand_99_nl = ~((fsm_output[5]) & (fsm_output[2]) & (fsm_output[6]) & (fsm_output[7])
      & (fsm_output[3]));
  assign mux_179_nl = MUX_s_1_2_2((nand_99_nl), or_186_cse, fsm_output[1]);
  assign mux_177_nl = MUX_s_1_2_2(or_201_cse, mux_tmp_153, fsm_output[5]);
  assign mux_174_nl = MUX_s_1_2_2(mux_tmp_103, nand_100_cse, fsm_output[6]);
  assign mux_175_nl = MUX_s_1_2_2(or_765_cse, (mux_174_nl), fsm_output[2]);
  assign mux_176_nl = MUX_s_1_2_2((mux_175_nl), or_169_cse, fsm_output[5]);
  assign mux_178_nl = MUX_s_1_2_2((mux_177_nl), (mux_176_nl), fsm_output[1]);
  assign mux_180_nl = MUX_s_1_2_2((mux_179_nl), (mux_178_nl), fsm_output[4]);
  assign nand_12_nl = ~((fsm_output[5]) & (~ mux_tmp_153));
  assign or_198_nl = (fsm_output[5]) | mux_tmp_153;
  assign mux_173_nl = MUX_s_1_2_2((nand_12_nl), (or_198_nl), fsm_output[1]);
  assign or_199_nl = (fsm_output[4]) | (mux_173_nl);
  assign mux_181_nl = MUX_s_1_2_2((mux_180_nl), (or_199_nl), fsm_output[0]);
  assign nor_201_nl = ~((mux_181_nl) | (fsm_output[8]));
  assign or_213_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[6]);
  assign mux_192_nl = MUX_s_1_2_2((or_213_nl), or_176_cse, fsm_output[2]);
  assign or_214_nl = (fsm_output[1]) | (mux_192_nl);
  assign or_212_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[3])
      | (fsm_output[6]);
  assign mux_193_nl = MUX_s_1_2_2((or_214_nl), (or_212_nl), fsm_output[4]);
  assign or_921_nl = (fsm_output[4]) | (~ (fsm_output[1])) | mux_142_cse;
  assign mux_194_nl = MUX_s_1_2_2((mux_193_nl), (or_921_nl), fsm_output[5]);
  assign or_922_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (~ (fsm_output[6]));
  assign mux_186_nl = MUX_s_1_2_2((fsm_output[6]), (~ (fsm_output[6])), fsm_output[3]);
  assign mux_187_nl = MUX_s_1_2_2(or_827_cse, (mux_186_nl), fsm_output[7]);
  assign mux_188_nl = MUX_s_1_2_2(or_176_cse, (mux_187_nl), fsm_output[2]);
  assign mux_189_nl = MUX_s_1_2_2(or_201_cse, (mux_188_nl), fsm_output[1]);
  assign mux_190_nl = MUX_s_1_2_2((or_922_nl), (mux_189_nl), fsm_output[4]);
  assign or_207_nl = (fsm_output[1]) | nand_111_cse;
  assign mux_184_nl = MUX_s_1_2_2(mux_142_cse, or_169_cse, fsm_output[1]);
  assign mux_185_nl = MUX_s_1_2_2((or_207_nl), (mux_184_nl), fsm_output[4]);
  assign mux_191_nl = MUX_s_1_2_2((mux_190_nl), (mux_185_nl), fsm_output[5]);
  assign mux_195_nl = MUX_s_1_2_2((mux_194_nl), (mux_191_nl), fsm_output[0]);
  assign nor_200_nl = ~((mux_195_nl) | (fsm_output[8]));
  assign or_219_nl = (fsm_output[5:4]!=2'b10) | mux_210_cse;
  assign mux_200_nl = MUX_s_1_2_2(or_222_cse, (or_219_nl), fsm_output[1]);
  assign mux_208_nl = MUX_s_1_2_2(mux_207_cse, (mux_200_nl), fsm_output[0]);
  assign nor_199_nl = ~((mux_208_nl) | (fsm_output[8]));
  assign nand_16_nl = ~((fsm_output[5]) & (~ mux_199_cse));
  assign mux_220_nl = MUX_s_1_2_2((nand_16_nl), or_222_cse, fsm_output[1]);
  assign mux_221_nl = MUX_s_1_2_2((mux_220_nl), mux_207_cse, fsm_output[0]);
  assign nor_198_nl = ~((mux_221_nl) | (fsm_output[8]));
  assign nand_132_nl = ~((fsm_output[2]) & (fsm_output[6]) & (~ (fsm_output[0]))
      & (fsm_output[4]));
  assign mux_231_nl = MUX_s_1_2_2(or_tmp_213, (nand_132_nl), fsm_output[7]);
  assign or_248_nl = (fsm_output[3]) | (mux_231_nl);
  assign or_245_nl = (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[0]) | (~
      (fsm_output[4]));
  assign mux_229_nl = MUX_s_1_2_2(or_tmp_219, (or_245_nl), fsm_output[7]);
  assign mux_230_nl = MUX_s_1_2_2((mux_229_nl), mux_tmp_206, fsm_output[3]);
  assign mux_232_nl = MUX_s_1_2_2((or_248_nl), (mux_230_nl), fsm_output[5]);
  assign or_241_nl = (~ (fsm_output[2])) | (~ (fsm_output[6])) | (fsm_output[0])
      | (fsm_output[4]);
  assign mux_226_nl = MUX_s_1_2_2(or_tmp_219, (or_241_nl), fsm_output[7]);
  assign mux_227_nl = MUX_s_1_2_2((mux_226_nl), mux_tmp_206, fsm_output[3]);
  assign or_238_nl = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[0]) | (fsm_output[4]);
  assign mux_222_nl = MUX_s_1_2_2((or_238_nl), or_tmp_213, fsm_output[7]);
  assign nand_127_nl = ~((fsm_output[7]) & (fsm_output[2]) & (fsm_output[6]) & (~
      (fsm_output[0])) & (fsm_output[4]));
  assign mux_223_nl = MUX_s_1_2_2((mux_222_nl), (nand_127_nl), fsm_output[3]);
  assign mux_228_nl = MUX_s_1_2_2((mux_227_nl), (mux_223_nl), fsm_output[5]);
  assign mux_233_nl = MUX_s_1_2_2((mux_232_nl), (mux_228_nl), fsm_output[1]);
  assign nor_197_nl = ~((mux_233_nl) | (fsm_output[8]));
  assign or_261_nl = (~ (fsm_output[2])) | (fsm_output[6]) | nand_100_cse;
  assign mux_246_nl = MUX_s_1_2_2((or_261_nl), mux_245_cse, fsm_output[4]);
  assign or_938_nl = (fsm_output[5]) | (mux_246_nl);
  assign mux_244_nl = MUX_s_1_2_2(mux_tmp_217, or_220_cse, fsm_output[4]);
  assign nand_124_nl = ~((fsm_output[5]) & (~ (mux_244_nl)));
  assign mux_247_nl = MUX_s_1_2_2((or_938_nl), (nand_124_nl), fsm_output[1]);
  assign or_256_nl = (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[7]) | (fsm_output[3]);
  assign mux_241_nl = MUX_s_1_2_2((or_256_nl), nand_62_cse, fsm_output[4]);
  assign mux_240_nl = MUX_s_1_2_2(mux_239_cse, or_765_cse, fsm_output[2]);
  assign nand_18_nl = ~((fsm_output[4]) & (~ (mux_240_nl)));
  assign mux_242_nl = MUX_s_1_2_2((mux_241_nl), (nand_18_nl), fsm_output[5]);
  assign mux_237_nl = MUX_s_1_2_2(nand_62_cse, mux_tmp_217, fsm_output[4]);
  assign or_939_nl = (fsm_output[2]) | mux_234_cse;
  assign mux_235_nl = MUX_s_1_2_2((or_939_nl), nand_111_cse, fsm_output[4]);
  assign mux_238_nl = MUX_s_1_2_2((mux_237_nl), (mux_235_nl), fsm_output[5]);
  assign mux_243_nl = MUX_s_1_2_2((mux_242_nl), (mux_238_nl), fsm_output[1]);
  assign mux_248_nl = MUX_s_1_2_2((mux_247_nl), (mux_243_nl), fsm_output[0]);
  assign nor_196_nl = ~((mux_248_nl) | (fsm_output[8]));
  assign or_283_nl = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[6]);
  assign mux_256_nl = MUX_s_1_2_2((or_283_nl), mux_tmp_232, fsm_output[5]);
  assign or_282_nl = (fsm_output[5]) | (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), (or_282_nl), fsm_output[1]);
  assign or_280_nl = (fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_258_nl = MUX_s_1_2_2((mux_257_nl), (or_280_nl), fsm_output[7]);
  assign nor_138_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[6])));
  assign nor_139_nl = ~((fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[6])));
  assign mux_255_nl = MUX_s_1_2_2((nor_138_nl), (nor_139_nl), fsm_output[5]);
  assign nand_20_nl = ~((fsm_output[7]) & (fsm_output[1]) & (mux_255_nl));
  assign mux_259_nl = MUX_s_1_2_2((mux_258_nl), (nand_20_nl), fsm_output[4]);
  assign or_274_nl = (~ (fsm_output[7])) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[2])
      | (fsm_output[8]) | (~ (fsm_output[6]));
  assign mux_254_nl = MUX_s_1_2_2((or_274_nl), mux_tmp_231, fsm_output[4]);
  assign mux_260_nl = MUX_s_1_2_2((mux_259_nl), (mux_254_nl), fsm_output[3]);
  assign or_271_nl = (fsm_output[5]) | mux_tmp_232;
  assign mux_252_nl = MUX_s_1_2_2((or_271_nl), or_tmp_239, fsm_output[1]);
  assign or_272_nl = (~ (fsm_output[4])) | (fsm_output[7]) | (mux_252_nl);
  assign or_267_nl = (fsm_output[4]) | mux_tmp_231;
  assign mux_253_nl = MUX_s_1_2_2((or_272_nl), (or_267_nl), fsm_output[3]);
  assign mux_261_nl = MUX_s_1_2_2((mux_260_nl), (mux_253_nl), fsm_output[0]);
  assign or_300_nl = (~ (fsm_output[5])) | (~ (fsm_output[2])) | (fsm_output[6])
      | (~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[3]));
  assign nand_21_nl = ~((fsm_output[5]) & (~ mux_tmp_253));
  assign mux_274_nl = MUX_s_1_2_2((or_300_nl), (nand_21_nl), fsm_output[4]);
  assign or_298_nl = (fsm_output[5]) | mux_tmp_253;
  assign mux_273_nl = MUX_s_1_2_2(or_tmp_268, (or_298_nl), fsm_output[4]);
  assign mux_275_nl = MUX_s_1_2_2((mux_274_nl), (mux_273_nl), fsm_output[1]);
  assign or_295_nl = (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[3]);
  assign mux_268_nl = MUX_s_1_2_2((or_295_nl), or_tmp_264, fsm_output[6]);
  assign or_296_nl = (fsm_output[2]) | (mux_268_nl);
  assign or_293_nl = (fsm_output[7]) | (fsm_output[8]) | (fsm_output[3]);
  assign mux_266_nl = MUX_s_1_2_2((or_293_nl), or_tmp_262, fsm_output[6]);
  assign mux_267_nl = MUX_s_1_2_2(or_tmp_270, (mux_266_nl), fsm_output[2]);
  assign mux_269_nl = MUX_s_1_2_2((or_296_nl), (mux_267_nl), fsm_output[5]);
  assign mux_270_nl = MUX_s_1_2_2((mux_269_nl), or_tmp_268, fsm_output[4]);
  assign or_290_nl = (fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[7])
      | (fsm_output[8]) | (fsm_output[3]);
  assign or_289_nl = (~ (fsm_output[2])) | (~ (fsm_output[6])) | (~ (fsm_output[7]))
      | (fsm_output[8]) | (fsm_output[3]);
  assign mux_262_nl = MUX_s_1_2_2(or_tmp_264, or_tmp_262, fsm_output[6]);
  assign or_285_nl = (~ (fsm_output[6])) | (fsm_output[7]) | (fsm_output[8]) | (~
      (fsm_output[3]));
  assign mux_263_nl = MUX_s_1_2_2((mux_262_nl), (or_285_nl), fsm_output[2]);
  assign mux_264_nl = MUX_s_1_2_2((or_289_nl), (mux_263_nl), fsm_output[5]);
  assign mux_265_nl = MUX_s_1_2_2((or_290_nl), (mux_264_nl), fsm_output[4]);
  assign mux_271_nl = MUX_s_1_2_2((mux_270_nl), (mux_265_nl), fsm_output[1]);
  assign mux_276_nl = MUX_s_1_2_2((mux_275_nl), (mux_271_nl), fsm_output[0]);
  assign or_312_nl = (fsm_output[6]) | (~ (fsm_output[7])) | (fsm_output[3]);
  assign mux_287_nl = MUX_s_1_2_2((or_312_nl), or_187_cse, fsm_output[2]);
  assign or_313_nl = (fsm_output[5]) | (mux_287_nl);
  assign nand_23_nl = ~((fsm_output[2]) & (~ mux_239_cse));
  assign mux_286_nl = MUX_s_1_2_2(or_169_cse, (nand_23_nl), fsm_output[5]);
  assign mux_288_nl = MUX_s_1_2_2((or_313_nl), (mux_286_nl), fsm_output[4]);
  assign mux_282_nl = MUX_s_1_2_2(or_187_cse, mux_234_cse, fsm_output[2]);
  assign mux_283_nl = MUX_s_1_2_2(or_169_cse, (mux_282_nl), fsm_output[5]);
  assign mux_284_nl = MUX_s_1_2_2((mux_283_nl), or_tmp_282, fsm_output[4]);
  assign mux_289_nl = MUX_s_1_2_2((mux_288_nl), (mux_284_nl), fsm_output[1]);
  assign or_308_nl = (~ (fsm_output[5])) | (~ (fsm_output[2])) | (fsm_output[6])
      | nand_100_cse;
  assign nand_22_nl = ~((fsm_output[5]) & (~ mux_245_cse));
  assign mux_279_nl = MUX_s_1_2_2((or_308_nl), (nand_22_nl), fsm_output[4]);
  assign or_304_nl = (fsm_output[5]) | mux_245_cse;
  assign mux_278_nl = MUX_s_1_2_2(or_tmp_282, (or_304_nl), fsm_output[4]);
  assign mux_280_nl = MUX_s_1_2_2((mux_279_nl), (mux_278_nl), fsm_output[1]);
  assign mux_290_nl = MUX_s_1_2_2((mux_289_nl), (mux_280_nl), fsm_output[0]);
  assign or_301_nl = (fsm_output[7:0]!=8'b00000010);
  assign mux_291_nl = MUX_s_1_2_2((mux_290_nl), (or_301_nl), fsm_output[8]);
  assign nand_122_nl = ~((fsm_output[4]) & (~ mux_tmp_275));
  assign nand_123_nl = ~((fsm_output[5]) & (fsm_output[1]) & (fsm_output[2]) & (fsm_output[7])
      & (~ (fsm_output[6])));
  assign or_935_nl = (fsm_output[5]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[7])
      | (fsm_output[6]);
  assign mux_296_nl = MUX_s_1_2_2((nand_123_nl), (or_935_nl), fsm_output[4]);
  assign mux_297_nl = MUX_s_1_2_2((nand_122_nl), (mux_296_nl), fsm_output[3]);
  assign or_936_nl = (fsm_output[4]) | mux_tmp_275;
  assign or_937_nl = (~ (fsm_output[4])) | (fsm_output[5]) | (~ (fsm_output[1]))
      | (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign mux_295_nl = MUX_s_1_2_2((or_936_nl), (or_937_nl), fsm_output[3]);
  assign mux_298_nl = MUX_s_1_2_2((mux_297_nl), (mux_295_nl), fsm_output[0]);
  assign nor_195_nl = ~((mux_298_nl) | (fsm_output[8]));
  assign nl_pe_0_0_run_cmp_input_in_rsc_dat = MUX1HOT_v_8_22_2(input_reg_16_15_lpi_2,
      input_reg_16_14_lpi_2, input_reg_16_13_lpi_2, input_reg_16_10_lpi_2, input_reg_16_11_lpi_2,
      input_reg_16_12_lpi_2, ROW_asn_142_itm, (psum_reg_16_2_lpi_2[7:0]), ROW_asn_143_itm,
      ROW_asn_145_itm, ROW_asn_147_itm, ROW_asn_149_itm, ROW_asn_151_itm, ROW_asn_153_itm,
      ROW_asn_155_itm, ROW_asn_157_itm, ROW_asn_159_itm, ROW_asn_161_itm, ROW_asn_163_itm,
      ROW_asn_165_itm, ROW_asn_167_itm, ROW_asn_169_itm, {and_dcpl_12 , and_dcpl_8
      , and_dcpl_42 , and_dcpl_45 , and_dcpl_47 , and_dcpl_51 , (nor_206_nl) , and_dcpl_55
      , (nor_205_nl) , (nor_204_nl) , (nor_203_nl) , (nor_202_nl) , (nor_201_nl)
      , (nor_200_nl) , (nor_199_nl) , (nor_198_nl) , (nor_197_nl) , (nor_196_nl)
      , (~ (mux_261_nl)) , (~ (mux_276_nl)) , (~ (mux_291_nl)) , (nor_195_nl)});
  wire[0:0] and_340_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] and_471_nl;
  wire[0:0] and_343_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] nor_145_nl;
  wire[0:0] nor_146_nl;
  wire[0:0] and_346_nl;
  wire[0:0] mux_108_nl;
  wire [15:0] nl_pe_0_0_run_cmp_psum_in_rsc_dat;
  assign and_471_nl = (fsm_output[7:6]==2'b11);
  assign mux_106_nl = MUX_s_1_2_2(and_dcpl_20, (and_471_nl), fsm_output[2]);
  assign and_340_nl = (mux_106_nl) & (~ (fsm_output[8])) & (~ (fsm_output[4])) &
      and_dcpl_13 & and_463_cse;
  assign nor_145_nl = ~((~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[4]) |
      (fsm_output[7]));
  assign nor_146_nl = ~((fsm_output[2]) | (~((fsm_output[3]) & (fsm_output[4]) &
      (fsm_output[7]))));
  assign mux_107_nl = MUX_s_1_2_2((nor_145_nl), (nor_146_nl), fsm_output[5]);
  assign and_343_nl = (mux_107_nl) & and_dcpl_341 & and_dcpl_1;
  assign mux_108_nl = MUX_s_1_2_2(or_tmp_127, or_tmp_126, fsm_output[5]);
  assign and_346_nl = (~ (mux_108_nl)) & and_dcpl_5 & and_dcpl_14 & and_dcpl_40;
  assign nl_pe_0_0_run_cmp_psum_in_rsc_dat = MUX1HOT_v_16_253_2(psum_reg_15_16_lpi_2,
      psum_reg_15_15_lpi_2, psum_reg_15_14_lpi_2, psum_reg_15_11_lpi_2, psum_reg_15_12_lpi_2,
      psum_reg_15_13_lpi_2, step_output_buf_value_0_sva, psum_reg_1_1_lpi_2, psum_reg_2_1_lpi_2,
      psum_reg_3_1_lpi_2, psum_reg_4_1_lpi_2, psum_reg_5_1_lpi_2, psum_reg_6_1_lpi_2,
      psum_reg_7_1_lpi_2, psum_reg_8_1_lpi_2, psum_reg_9_1_lpi_2, psum_reg_10_1_lpi_2,
      psum_reg_11_1_lpi_2, psum_reg_12_1_lpi_2, psum_reg_13_1_lpi_2, psum_reg_14_1_lpi_2,
      psum_reg_15_1_lpi_2, psum_reg_16_1_lpi_2, psum_reg_1_2_lpi_2, psum_reg_2_2_lpi_2,
      psum_reg_3_2_lpi_2, psum_reg_4_2_lpi_2, psum_reg_5_2_lpi_2, psum_reg_6_2_lpi_2,
      psum_reg_7_2_lpi_2, psum_reg_8_2_lpi_2, psum_reg_9_2_lpi_2, psum_reg_10_2_lpi_2,
      psum_reg_11_2_lpi_2, psum_reg_12_2_lpi_2, psum_reg_13_2_lpi_2, psum_reg_14_2_lpi_2,
      psum_reg_15_2_lpi_2, psum_reg_1_3_lpi_2, psum_reg_2_3_lpi_2, psum_reg_3_3_lpi_2,
      psum_reg_4_3_lpi_2, psum_reg_5_3_lpi_2, psum_reg_6_3_lpi_2, psum_reg_7_3_lpi_2,
      psum_reg_8_3_lpi_2, psum_reg_9_3_lpi_2, psum_reg_10_3_lpi_2, psum_reg_11_3_lpi_2,
      psum_reg_12_3_lpi_2, psum_reg_13_3_lpi_2, psum_reg_14_3_lpi_2, psum_reg_15_3_lpi_2,
      psum_reg_16_10_lpi_2, psum_reg_1_4_lpi_2, psum_reg_2_4_lpi_2, psum_reg_3_4_lpi_2,
      psum_reg_4_4_lpi_2, psum_reg_5_4_lpi_2, psum_reg_6_4_lpi_2, psum_reg_7_4_lpi_2,
      psum_reg_8_4_lpi_2, psum_reg_9_4_lpi_2, psum_reg_10_4_lpi_2, psum_reg_11_4_lpi_2,
      psum_reg_12_4_lpi_2, psum_reg_13_4_lpi_2, psum_reg_14_4_lpi_2, psum_reg_15_4_lpi_2,
      psum_reg_16_4_lpi_2, psum_reg_1_5_lpi_2, psum_reg_2_5_lpi_2, psum_reg_3_5_lpi_2,
      psum_reg_4_5_lpi_2, psum_reg_5_5_lpi_2, psum_reg_6_5_lpi_2, psum_reg_7_5_lpi_2,
      psum_reg_8_5_lpi_2, psum_reg_9_5_lpi_2, psum_reg_10_5_lpi_2, psum_reg_11_5_lpi_2,
      psum_reg_12_5_lpi_2, psum_reg_13_5_lpi_2, psum_reg_14_5_lpi_2, psum_reg_15_5_lpi_2,
      psum_reg_16_5_lpi_2, psum_reg_1_6_lpi_2, psum_reg_2_6_lpi_2, psum_reg_3_6_lpi_2,
      psum_reg_4_6_lpi_2, psum_reg_5_6_lpi_2, psum_reg_6_6_lpi_2, psum_reg_7_6_lpi_2,
      psum_reg_8_6_lpi_2, psum_reg_9_6_lpi_2, psum_reg_10_6_lpi_2, psum_reg_11_6_lpi_2,
      psum_reg_12_6_lpi_2, psum_reg_13_6_lpi_2, psum_reg_14_6_lpi_2, psum_reg_15_6_lpi_2,
      psum_reg_16_6_lpi_2, psum_reg_1_7_lpi_2, psum_reg_2_7_lpi_2, psum_reg_3_7_lpi_2,
      psum_reg_4_7_lpi_2, psum_reg_5_7_lpi_2, psum_reg_6_7_lpi_2, psum_reg_7_7_lpi_2,
      psum_reg_8_7_lpi_2, psum_reg_9_7_lpi_2, psum_reg_10_7_lpi_2, psum_reg_11_7_lpi_2,
      psum_reg_12_7_lpi_2, psum_reg_13_7_lpi_2, psum_reg_14_7_lpi_2, psum_reg_15_7_lpi_2,
      psum_reg_16_7_lpi_2, psum_reg_1_8_lpi_2, psum_reg_2_8_lpi_2, psum_reg_3_8_lpi_2,
      psum_reg_4_8_lpi_2, psum_reg_5_8_lpi_2, psum_reg_6_8_lpi_2, psum_reg_7_8_lpi_2,
      psum_reg_8_8_lpi_2, psum_reg_9_8_lpi_2, psum_reg_10_8_lpi_2, psum_reg_11_8_lpi_2,
      psum_reg_12_8_lpi_2, psum_reg_13_8_lpi_2, psum_reg_14_8_lpi_2, psum_reg_15_8_lpi_2,
      psum_reg_16_8_lpi_2, psum_reg_1_9_lpi_2, psum_reg_2_9_lpi_2, psum_reg_3_9_lpi_2,
      psum_reg_4_9_lpi_2, psum_reg_5_9_lpi_2, psum_reg_6_9_lpi_2, psum_reg_7_9_lpi_2,
      psum_reg_8_9_lpi_2, psum_reg_9_9_lpi_2, psum_reg_10_9_lpi_2, psum_reg_11_9_lpi_2,
      psum_reg_12_9_lpi_2, psum_reg_13_9_lpi_2, psum_reg_14_9_lpi_2, psum_reg_15_9_lpi_2,
      psum_reg_16_9_lpi_2, psum_reg_1_10_lpi_2, psum_reg_2_10_lpi_2, psum_reg_3_10_lpi_2,
      psum_reg_4_10_lpi_2, psum_reg_5_10_lpi_2, psum_reg_6_10_lpi_2, psum_reg_7_10_lpi_2,
      psum_reg_8_10_lpi_2, psum_reg_9_10_lpi_2, psum_reg_10_10_lpi_2, psum_reg_11_10_lpi_2,
      psum_reg_12_10_lpi_2, psum_reg_13_10_lpi_2, psum_reg_14_10_lpi_2, psum_reg_15_10_lpi_2,
      step_accum_fifo_input_15_asn_9_ncse_sva, psum_reg_1_11_lpi_2, psum_reg_2_11_lpi_2,
      psum_reg_3_11_lpi_2, psum_reg_4_11_lpi_2, psum_reg_5_11_lpi_2, psum_reg_6_11_lpi_2,
      psum_reg_7_11_lpi_2, psum_reg_8_11_lpi_2, psum_reg_9_11_lpi_2, psum_reg_10_11_lpi_2,
      psum_reg_11_11_lpi_2, psum_reg_12_11_lpi_2, psum_reg_13_11_lpi_2, psum_reg_14_11_lpi_2,
      psum_reg_1_12_lpi_2, psum_reg_2_12_lpi_2, psum_reg_3_12_lpi_2, psum_reg_4_12_lpi_2,
      psum_reg_5_12_lpi_2, psum_reg_6_12_lpi_2, psum_reg_7_12_lpi_2, psum_reg_8_12_lpi_2,
      psum_reg_9_12_lpi_2, psum_reg_10_12_lpi_2, psum_reg_11_12_lpi_2, psum_reg_12_12_lpi_2,
      psum_reg_13_12_lpi_2, psum_reg_14_12_lpi_2, psum_reg_1_13_lpi_2, psum_reg_2_13_lpi_2,
      psum_reg_3_13_lpi_2, psum_reg_4_13_lpi_2, psum_reg_5_13_lpi_2, psum_reg_6_13_lpi_2,
      psum_reg_7_13_lpi_2, psum_reg_8_13_lpi_2, psum_reg_9_13_lpi_2, psum_reg_10_13_lpi_2,
      psum_reg_11_13_lpi_2, psum_reg_12_13_lpi_2, psum_reg_13_13_lpi_2, psum_reg_14_13_lpi_2,
      step_accum_fifo_input_15_asn_12_ncse_sva, psum_reg_1_14_lpi_2, psum_reg_2_14_lpi_2,
      psum_reg_3_14_lpi_2, psum_reg_4_14_lpi_2, psum_reg_5_14_lpi_2, psum_reg_6_14_lpi_2,
      psum_reg_7_14_lpi_2, psum_reg_8_14_lpi_2, psum_reg_9_14_lpi_2, psum_reg_10_14_lpi_2,
      psum_reg_11_14_lpi_2, psum_reg_12_14_lpi_2, psum_reg_13_14_lpi_2, psum_reg_14_14_lpi_2,
      step_accum_fifo_input_15_asn_13_ncse_sva, psum_reg_1_15_lpi_2, psum_reg_2_15_lpi_2,
      psum_reg_3_15_lpi_2, psum_reg_4_15_lpi_2, psum_reg_5_15_lpi_2, psum_reg_6_15_lpi_2,
      psum_reg_7_15_lpi_2, psum_reg_8_15_lpi_2, psum_reg_9_15_lpi_2, psum_reg_10_15_lpi_2,
      psum_reg_11_15_lpi_2, psum_reg_12_15_lpi_2, psum_reg_13_15_lpi_2, psum_reg_14_15_lpi_2,
      step_accum_fifo_input_15_asn_14_ncse_sva, psum_reg_1_16_lpi_2, psum_reg_2_16_lpi_2,
      psum_reg_3_16_lpi_2, psum_reg_4_16_lpi_2, psum_reg_5_16_lpi_2, psum_reg_6_16_lpi_2,
      psum_reg_7_16_lpi_2, psum_reg_8_16_lpi_2, psum_reg_9_16_lpi_2, psum_reg_10_16_lpi_2,
      psum_reg_11_16_lpi_2, psum_reg_12_16_lpi_2, psum_reg_13_16_lpi_2, psum_reg_14_16_lpi_2,
      {(and_340_nl) , (and_343_nl) , (and_346_nl) , and_dcpl_45 , and_dcpl_47 , and_dcpl_51
      , and_dcpl_53 , and_dcpl_55 , and_dcpl_56 , and_dcpl_57 , and_dcpl_58 , and_dcpl_59
      , and_dcpl_60 , and_dcpl_63 , and_dcpl_64 , and_dcpl_65 , and_dcpl_66 , and_dcpl_67
      , and_dcpl_68 , and_dcpl_69 , and_dcpl_70 , and_dcpl_73 , and_dcpl_74 , and_dcpl_75
      , and_dcpl_76 , and_dcpl_77 , and_dcpl_78 , and_dcpl_79 , and_dcpl_80 , and_dcpl_83
      , and_dcpl_85 , and_dcpl_87 , and_dcpl_89 , and_dcpl_92 , and_dcpl_94 , and_dcpl_96
      , and_dcpl_98 , and_dcpl_99 , and_dcpl_101 , and_dcpl_102 , and_dcpl_103 ,
      and_dcpl_104 , and_dcpl_105 , and_dcpl_106 , and_dcpl_107 , and_dcpl_108 ,
      and_dcpl_109 , and_dcpl_110 , and_dcpl_111 , and_dcpl_112 , and_dcpl_113 ,
      and_dcpl_114 , and_dcpl_115 , and_dcpl_116 , and_dcpl_117 , and_dcpl_118 ,
      and_dcpl_119 , and_dcpl_120 , and_dcpl_121 , and_dcpl_122 , and_dcpl_125 ,
      and_dcpl_126 , and_dcpl_127 , and_dcpl_128 , and_dcpl_129 , and_dcpl_130 ,
      and_dcpl_131 , and_dcpl_132 , and_dcpl_134 , and_dcpl_135 , and_dcpl_136 ,
      and_dcpl_137 , and_dcpl_138 , and_dcpl_139 , and_dcpl_140 , and_dcpl_141 ,
      and_dcpl_143 , and_dcpl_144 , and_dcpl_145 , and_dcpl_146 , and_dcpl_147 ,
      and_dcpl_148 , and_dcpl_149 , and_dcpl_150 , and_dcpl_152 , and_dcpl_153 ,
      and_dcpl_154 , and_dcpl_155 , and_dcpl_156 , and_dcpl_157 , and_dcpl_158 ,
      and_dcpl_159 , and_dcpl_160 , and_dcpl_161 , and_dcpl_162 , and_dcpl_163 ,
      and_dcpl_164 , and_dcpl_165 , and_dcpl_166 , and_dcpl_167 , and_dcpl_168 ,
      and_dcpl_169 , and_dcpl_170 , and_dcpl_171 , and_dcpl_172 , and_dcpl_173 ,
      and_dcpl_174 , and_dcpl_175 , and_dcpl_176 , and_dcpl_177 , and_dcpl_178 ,
      and_dcpl_179 , and_dcpl_180 , and_dcpl_181 , and_dcpl_182 , and_dcpl_183 ,
      and_dcpl_184 , and_dcpl_185 , and_dcpl_186 , and_dcpl_187 , and_dcpl_188 ,
      and_dcpl_189 , and_dcpl_190 , and_dcpl_191 , and_dcpl_195 , and_dcpl_196 ,
      and_dcpl_197 , and_dcpl_198 , and_dcpl_199 , and_dcpl_200 , and_dcpl_201 ,
      and_dcpl_202 , and_dcpl_204 , and_dcpl_205 , and_dcpl_206 , and_dcpl_207 ,
      and_dcpl_208 , and_dcpl_209 , and_dcpl_210 , and_dcpl_211 , and_dcpl_213 ,
      and_dcpl_214 , and_dcpl_215 , and_dcpl_216 , and_dcpl_217 , and_dcpl_218 ,
      and_dcpl_219 , and_dcpl_220 , and_dcpl_222 , and_dcpl_223 , and_dcpl_224 ,
      and_dcpl_225 , and_dcpl_226 , and_dcpl_227 , and_dcpl_228 , and_dcpl_229 ,
      and_dcpl_230 , and_dcpl_231 , and_dcpl_232 , and_dcpl_233 , and_dcpl_234 ,
      and_dcpl_235 , and_dcpl_236 , and_dcpl_237 , and_dcpl_238 , and_dcpl_239 ,
      and_dcpl_240 , and_dcpl_241 , and_dcpl_242 , and_dcpl_243 , and_dcpl_244 ,
      and_dcpl_245 , and_dcpl_246 , and_dcpl_247 , and_dcpl_248 , and_dcpl_249 ,
      and_dcpl_250 , and_dcpl_251 , and_dcpl_252 , and_dcpl_253 , and_dcpl_255 ,
      and_dcpl_256 , and_dcpl_257 , and_dcpl_258 , and_dcpl_259 , and_dcpl_260 ,
      and_dcpl_261 , and_dcpl_264 , and_dcpl_265 , and_dcpl_266 , and_dcpl_267 ,
      and_dcpl_268 , and_dcpl_269 , and_dcpl_270 , and_dcpl_273 , and_dcpl_274 ,
      and_dcpl_275 , and_dcpl_276 , and_dcpl_277 , and_dcpl_278 , and_dcpl_279 ,
      and_dcpl_280 , and_dcpl_282 , and_dcpl_283 , and_dcpl_284 , and_dcpl_285 ,
      and_dcpl_286 , and_dcpl_287 , and_dcpl_288 , and_dcpl_289 , and_dcpl_291 ,
      and_dcpl_292 , and_dcpl_293 , and_dcpl_294 , and_dcpl_295 , and_dcpl_296 ,
      and_dcpl_297 , and_dcpl_298 , and_dcpl_299 , and_dcpl_300 , and_dcpl_301 ,
      and_dcpl_302 , and_dcpl_303 , and_dcpl_304 , and_dcpl_305 , and_dcpl_306 ,
      and_dcpl_307 , and_dcpl_308 , and_dcpl_309 , and_dcpl_310 , and_dcpl_311 ,
      and_dcpl_312 , and_dcpl_313 , and_dcpl_314 , and_dcpl_315 , and_dcpl_316 ,
      and_dcpl_317 , and_dcpl_318 , and_dcpl_319 , and_dcpl_320 , and_dcpl_321 ,
      and_dcpl_322 , and_dcpl_323 , and_dcpl_324 , and_dcpl_325 , and_dcpl_326 ,
      and_dcpl_327 , and_dcpl_328 , and_dcpl_329 , and_dcpl_330 , and_dcpl_334 ,
      and_dcpl_335 , and_dcpl_336});
  wire[0:0] and_39_nl;
  wire [7:0] nl_pe_0_0_run_cmp_weight_rsc_dat;
  assign and_39_nl = (~(operator_16_false_slc_operator_16_false_acc_12_svs & (step_step_sva[3:0]==4'b1111)))
      & and_dcpl_5 & and_dcpl_14 & and_dcpl_29 & and_dcpl_35;
  assign nl_pe_0_0_run_cmp_weight_rsc_dat = MUX1HOT_v_8_257_2((weight_rsci_idat_mxwt[127:120]),
      weight_reg_15_15_lpi_2, weight_reg_15_14_lpi_2, weight_reg_15_13_lpi_2, weight_reg_15_10_lpi_2,
      weight_reg_15_11_lpi_2, weight_reg_15_12_lpi_2, weight_reg_0_0_lpi_2, weight_reg_1_0_lpi_2,
      weight_reg_2_0_lpi_2, weight_reg_3_0_lpi_2, weight_reg_4_0_lpi_2, weight_reg_5_0_lpi_2,
      weight_reg_6_0_lpi_2, weight_reg_7_0_lpi_2, weight_reg_8_0_lpi_2, weight_reg_9_0_lpi_2,
      weight_reg_10_0_lpi_2, weight_reg_11_0_lpi_2, weight_reg_12_0_lpi_2, weight_reg_13_0_lpi_2,
      weight_reg_14_0_lpi_2, weight_reg_15_0_lpi_2, weight_reg_0_1_lpi_2, weight_reg_1_1_lpi_2,
      weight_reg_2_1_lpi_2, weight_reg_3_1_lpi_2, weight_reg_4_1_lpi_2, weight_reg_5_1_lpi_2,
      weight_reg_6_1_lpi_2, weight_reg_7_1_lpi_2, weight_reg_8_1_lpi_2, weight_reg_9_1_lpi_2,
      weight_reg_10_1_lpi_2, weight_reg_11_1_lpi_2, weight_reg_12_1_lpi_2, weight_reg_13_1_lpi_2,
      weight_reg_14_1_lpi_2, weight_reg_15_1_lpi_2, weight_reg_0_2_lpi_2, weight_reg_1_2_lpi_2,
      weight_reg_2_2_lpi_2, weight_reg_3_2_lpi_2, weight_reg_4_2_lpi_2, weight_reg_5_2_lpi_2,
      weight_reg_6_2_lpi_2, weight_reg_7_2_lpi_2, weight_reg_8_2_lpi_2, weight_reg_9_2_lpi_2,
      weight_reg_10_2_lpi_2, weight_reg_11_2_lpi_2, weight_reg_12_2_lpi_2, weight_reg_13_2_lpi_2,
      weight_reg_14_2_lpi_2, weight_reg_15_2_lpi_2, weight_reg_0_3_lpi_2, weight_reg_1_3_lpi_2,
      weight_reg_2_3_lpi_2, weight_reg_3_3_lpi_2, weight_reg_4_3_lpi_2, weight_reg_5_3_lpi_2,
      weight_reg_6_3_lpi_2, weight_reg_7_3_lpi_2, weight_reg_8_3_lpi_2, weight_reg_9_3_lpi_2,
      weight_reg_10_3_lpi_2, weight_reg_11_3_lpi_2, weight_reg_12_3_lpi_2, weight_reg_13_3_lpi_2,
      weight_reg_14_3_lpi_2, weight_reg_15_3_lpi_2, weight_reg_0_4_lpi_2, weight_reg_1_4_lpi_2,
      weight_reg_2_4_lpi_2, weight_reg_3_4_lpi_2, weight_reg_4_4_lpi_2, weight_reg_5_4_lpi_2,
      weight_reg_6_4_lpi_2, weight_reg_7_4_lpi_2, weight_reg_8_4_lpi_2, weight_reg_9_4_lpi_2,
      weight_reg_10_4_lpi_2, weight_reg_11_4_lpi_2, weight_reg_12_4_lpi_2, weight_reg_13_4_lpi_2,
      weight_reg_14_4_lpi_2, weight_reg_15_4_lpi_2, weight_reg_0_5_lpi_2, weight_reg_1_5_lpi_2,
      weight_reg_2_5_lpi_2, weight_reg_3_5_lpi_2, weight_reg_4_5_lpi_2, weight_reg_5_5_lpi_2,
      weight_reg_6_5_lpi_2, weight_reg_7_5_lpi_2, weight_reg_8_5_lpi_2, weight_reg_9_5_lpi_2,
      weight_reg_10_5_lpi_2, weight_reg_11_5_lpi_2, weight_reg_12_5_lpi_2, weight_reg_13_5_lpi_2,
      weight_reg_14_5_lpi_2, weight_reg_15_5_lpi_2, weight_reg_0_6_lpi_2, weight_reg_1_6_lpi_2,
      weight_reg_2_6_lpi_2, weight_reg_3_6_lpi_2, weight_reg_4_6_lpi_2, weight_reg_5_6_lpi_2,
      weight_reg_6_6_lpi_2, weight_reg_7_6_lpi_2, weight_reg_8_6_lpi_2, weight_reg_9_6_lpi_2,
      weight_reg_10_6_lpi_2, weight_reg_11_6_lpi_2, weight_reg_12_6_lpi_2, weight_reg_13_6_lpi_2,
      weight_reg_14_6_lpi_2, weight_reg_15_6_lpi_2, weight_reg_0_7_lpi_2, weight_reg_1_7_lpi_2,
      weight_reg_2_7_lpi_2, weight_reg_3_7_lpi_2, weight_reg_4_7_lpi_2, weight_reg_5_7_lpi_2,
      weight_reg_6_7_lpi_2, weight_reg_7_7_lpi_2, weight_reg_8_7_lpi_2, weight_reg_9_7_lpi_2,
      weight_reg_10_7_lpi_2, weight_reg_11_7_lpi_2, weight_reg_12_7_lpi_2, weight_reg_13_7_lpi_2,
      weight_reg_14_7_lpi_2, weight_reg_15_7_lpi_2, weight_reg_0_8_lpi_2, weight_reg_1_8_lpi_2,
      weight_reg_2_8_lpi_2, weight_reg_3_8_lpi_2, weight_reg_4_8_lpi_2, weight_reg_5_8_lpi_2,
      weight_reg_6_8_lpi_2, weight_reg_7_8_lpi_2, weight_reg_8_8_lpi_2, weight_reg_9_8_lpi_2,
      weight_reg_10_8_lpi_2, weight_reg_11_8_lpi_2, weight_reg_12_8_lpi_2, weight_reg_13_8_lpi_2,
      weight_reg_14_8_lpi_2, weight_reg_15_8_lpi_2, weight_reg_0_9_lpi_2, weight_reg_1_9_lpi_2,
      weight_reg_2_9_lpi_2, weight_reg_3_9_lpi_2, weight_reg_4_9_lpi_2, weight_reg_5_9_lpi_2,
      weight_reg_6_9_lpi_2, weight_reg_7_9_lpi_2, weight_reg_8_9_lpi_2, weight_reg_9_9_lpi_2,
      weight_reg_10_9_lpi_2, weight_reg_11_9_lpi_2, weight_reg_12_9_lpi_2, weight_reg_13_9_lpi_2,
      weight_reg_14_9_lpi_2, weight_reg_15_9_lpi_2, weight_reg_0_10_lpi_2, weight_reg_1_10_lpi_2,
      weight_reg_2_10_lpi_2, weight_reg_3_10_lpi_2, weight_reg_4_10_lpi_2, weight_reg_5_10_lpi_2,
      weight_reg_6_10_lpi_2, weight_reg_7_10_lpi_2, weight_reg_8_10_lpi_2, weight_reg_9_10_lpi_2,
      weight_reg_10_10_lpi_2, weight_reg_11_10_lpi_2, weight_reg_12_10_lpi_2, weight_reg_13_10_lpi_2,
      weight_reg_14_10_lpi_2, weight_reg_0_11_lpi_2, weight_reg_1_11_lpi_2, weight_reg_2_11_lpi_2,
      weight_reg_3_11_lpi_2, weight_reg_4_11_lpi_2, weight_reg_5_11_lpi_2, weight_reg_6_11_lpi_2,
      weight_reg_7_11_lpi_2, weight_reg_8_11_lpi_2, weight_reg_9_11_lpi_2, weight_reg_10_11_lpi_2,
      weight_reg_11_11_lpi_2, weight_reg_12_11_lpi_2, weight_reg_13_11_lpi_2, weight_reg_14_11_lpi_2,
      weight_reg_0_12_lpi_2, weight_reg_1_12_lpi_2, weight_reg_2_12_lpi_2, weight_reg_3_12_lpi_2,
      weight_reg_4_12_lpi_2, weight_reg_5_12_lpi_2, weight_reg_6_12_lpi_2, weight_reg_7_12_lpi_2,
      weight_reg_8_12_lpi_2, weight_reg_9_12_lpi_2, weight_reg_10_12_lpi_2, weight_reg_11_12_lpi_2,
      weight_reg_12_12_lpi_2, weight_reg_13_12_lpi_2, weight_reg_14_12_lpi_2, weight_reg_0_13_lpi_2,
      weight_reg_1_13_lpi_2, weight_reg_2_13_lpi_2, weight_reg_3_13_lpi_2, weight_reg_4_13_lpi_2,
      weight_reg_5_13_lpi_2, weight_reg_6_13_lpi_2, weight_reg_7_13_lpi_2, weight_reg_8_13_lpi_2,
      weight_reg_9_13_lpi_2, weight_reg_10_13_lpi_2, weight_reg_11_13_lpi_2, weight_reg_12_13_lpi_2,
      weight_reg_13_13_lpi_2, weight_reg_14_13_lpi_2, weight_reg_0_14_lpi_2, weight_reg_1_14_lpi_2,
      weight_reg_2_14_lpi_2, weight_reg_3_14_lpi_2, weight_reg_4_14_lpi_2, weight_reg_5_14_lpi_2,
      weight_reg_6_14_lpi_2, weight_reg_7_14_lpi_2, weight_reg_8_14_lpi_2, weight_reg_9_14_lpi_2,
      weight_reg_10_14_lpi_2, weight_reg_11_14_lpi_2, weight_reg_12_14_lpi_2, weight_reg_13_14_lpi_2,
      weight_reg_14_14_lpi_2, weight_reg_0_15_lpi_2, weight_reg_1_15_lpi_2, weight_reg_2_15_lpi_2,
      weight_reg_3_15_lpi_2, weight_reg_4_15_lpi_2, weight_reg_5_15_lpi_2, weight_reg_6_15_lpi_2,
      weight_reg_7_15_lpi_2, weight_reg_8_15_lpi_2, weight_reg_9_15_lpi_2, weight_reg_10_15_lpi_2,
      weight_reg_11_15_lpi_2, weight_reg_12_15_lpi_2, weight_reg_13_15_lpi_2, weight_reg_14_15_lpi_2,
      {and_dcpl_33 , (and_39_nl) , and_dcpl_8 , and_dcpl_42 , and_dcpl_45 , and_dcpl_47
      , and_dcpl_51 , and_dcpl_53 , and_dcpl_55 , and_dcpl_56 , and_dcpl_57 , and_dcpl_58
      , and_dcpl_59 , and_dcpl_60 , and_dcpl_63 , and_dcpl_64 , and_dcpl_65 , and_dcpl_66
      , and_dcpl_67 , and_dcpl_68 , and_dcpl_69 , and_dcpl_70 , and_dcpl_73 , and_dcpl_74
      , and_dcpl_75 , and_dcpl_76 , and_dcpl_77 , and_dcpl_78 , and_dcpl_79 , and_dcpl_80
      , and_dcpl_83 , and_dcpl_85 , and_dcpl_87 , and_dcpl_89 , and_dcpl_92 , and_dcpl_94
      , and_dcpl_96 , and_dcpl_98 , and_dcpl_99 , and_dcpl_100 , and_dcpl_101 , and_dcpl_102
      , and_dcpl_103 , and_dcpl_104 , and_dcpl_105 , and_dcpl_106 , and_dcpl_107
      , and_dcpl_108 , and_dcpl_109 , and_dcpl_110 , and_dcpl_111 , and_dcpl_112
      , and_dcpl_113 , and_dcpl_114 , and_dcpl_115 , and_dcpl_116 , and_dcpl_117
      , and_dcpl_118 , and_dcpl_119 , and_dcpl_120 , and_dcpl_121 , and_dcpl_122
      , and_dcpl_125 , and_dcpl_126 , and_dcpl_127 , and_dcpl_128 , and_dcpl_129
      , and_dcpl_130 , and_dcpl_131 , and_dcpl_132 , and_dcpl_134 , and_dcpl_135
      , and_dcpl_136 , and_dcpl_137 , and_dcpl_138 , and_dcpl_139 , and_dcpl_140
      , and_dcpl_141 , and_dcpl_143 , and_dcpl_144 , and_dcpl_145 , and_dcpl_146
      , and_dcpl_147 , and_dcpl_148 , and_dcpl_149 , and_dcpl_150 , and_dcpl_152
      , and_dcpl_153 , and_dcpl_154 , and_dcpl_155 , and_dcpl_156 , and_dcpl_157
      , and_dcpl_158 , and_dcpl_159 , and_dcpl_160 , and_dcpl_161 , and_dcpl_162
      , and_dcpl_163 , and_dcpl_164 , and_dcpl_165 , and_dcpl_166 , and_dcpl_167
      , and_dcpl_168 , and_dcpl_169 , and_dcpl_170 , and_dcpl_171 , and_dcpl_172
      , and_dcpl_173 , and_dcpl_174 , and_dcpl_175 , and_dcpl_176 , and_dcpl_177
      , and_dcpl_178 , and_dcpl_179 , and_dcpl_180 , and_dcpl_181 , and_dcpl_182
      , and_dcpl_183 , and_dcpl_184 , and_dcpl_185 , and_dcpl_186 , and_dcpl_187
      , and_dcpl_188 , and_dcpl_189 , and_dcpl_190 , and_dcpl_191 , and_dcpl_195
      , and_dcpl_196 , and_dcpl_197 , and_dcpl_198 , and_dcpl_199 , and_dcpl_200
      , and_dcpl_201 , and_dcpl_202 , and_dcpl_204 , and_dcpl_205 , and_dcpl_206
      , and_dcpl_207 , and_dcpl_208 , and_dcpl_209 , and_dcpl_210 , and_dcpl_211
      , and_dcpl_213 , and_dcpl_214 , and_dcpl_215 , and_dcpl_216 , and_dcpl_217
      , and_dcpl_218 , and_dcpl_219 , and_dcpl_220 , and_dcpl_222 , and_dcpl_223
      , and_dcpl_224 , and_dcpl_225 , and_dcpl_226 , and_dcpl_227 , and_dcpl_228
      , and_dcpl_229 , and_dcpl_230 , and_dcpl_231 , and_dcpl_232 , and_dcpl_233
      , and_dcpl_234 , and_dcpl_235 , and_dcpl_236 , and_dcpl_237 , and_dcpl_238
      , and_dcpl_239 , and_dcpl_240 , and_dcpl_241 , and_dcpl_242 , and_dcpl_243
      , and_dcpl_244 , and_dcpl_245 , and_dcpl_246 , and_dcpl_247 , and_dcpl_248
      , and_dcpl_249 , and_dcpl_250 , and_dcpl_251 , and_dcpl_252 , and_dcpl_253
      , and_dcpl_254 , and_dcpl_255 , and_dcpl_256 , and_dcpl_257 , and_dcpl_258
      , and_dcpl_259 , and_dcpl_260 , and_dcpl_261 , and_dcpl_264 , and_dcpl_265
      , and_dcpl_266 , and_dcpl_267 , and_dcpl_268 , and_dcpl_269 , and_dcpl_270
      , and_dcpl_271 , and_dcpl_273 , and_dcpl_274 , and_dcpl_275 , and_dcpl_276
      , and_dcpl_277 , and_dcpl_278 , and_dcpl_279 , and_dcpl_280 , and_dcpl_282
      , and_dcpl_283 , and_dcpl_284 , and_dcpl_285 , and_dcpl_286 , and_dcpl_287
      , and_dcpl_288 , and_dcpl_289 , and_dcpl_291 , and_dcpl_292 , and_dcpl_293
      , and_dcpl_294 , and_dcpl_295 , and_dcpl_296 , and_dcpl_297 , and_dcpl_298
      , and_dcpl_299 , and_dcpl_300 , and_dcpl_301 , and_dcpl_302 , and_dcpl_303
      , and_dcpl_304 , and_dcpl_305 , and_dcpl_306 , and_dcpl_307 , and_dcpl_308
      , and_dcpl_309 , and_dcpl_310 , and_dcpl_311 , and_dcpl_312 , and_dcpl_313
      , and_dcpl_314 , and_dcpl_315 , and_dcpl_316 , and_dcpl_317 , and_dcpl_318
      , and_dcpl_319 , and_dcpl_320 , and_dcpl_321 , and_dcpl_322 , and_dcpl_323
      , and_dcpl_324 , and_dcpl_325 , and_dcpl_326 , and_dcpl_327 , and_dcpl_328
      , and_dcpl_329 , and_dcpl_330 , and_dcpl_334 , and_dcpl_335 , and_dcpl_336});
  wire [0:0] nl_pe_0_0_run_cmp_ccs_ccore_start_rsc_dat;
  assign nl_pe_0_0_run_cmp_ccs_ccore_start_rsc_dat = (or_94_cse | or_52_cse | or_dcpl_14
      | and_463_cse) ^ (fsm_output[8]);
  wire[15:0] step_if_2_step_if_2_and_nl;
  wire[0:0] step_if_2_aelse_1_not_31_nl;
  wire [15:0] nl_accum_fifo_0_run_cmp_input_rsc_dat;
  assign step_if_2_aelse_1_not_31_nl = ~ operator_16_false_slc_operator_16_false_acc_12_svs;
  assign step_if_2_step_if_2_and_nl = MUX_v_16_2_2(16'b0000000000000000, accumulation_buffer_rsc_0_0_i_dout_d_mxwt,
      (step_if_2_aelse_1_not_31_nl));
  assign nl_accum_fifo_0_run_cmp_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_16_lpi_2,
      (step_if_2_step_if_2_and_nl), and_dcpl_8);
  wire[0:0] mux_101_nl;
  wire[0:0] mux_100_nl;
  wire [0:0] nl_accum_fifo_0_run_cmp_ccs_ccore_start_rsc_dat;
  assign mux_100_nl = MUX_s_1_2_2(or_tmp_121, or_47_cse, fsm_output[1]);
  assign mux_101_nl = MUX_s_1_2_2(or_tmp_122, (mux_100_nl), fsm_output[0]);
  assign nl_accum_fifo_0_run_cmp_ccs_ccore_start_rsc_dat = (~ (mux_101_nl)) & (~
      (fsm_output[7])) & and_dcpl_15;
  wire [7:0] nl_input_fifo_0_run_cmp_input_rsc_dat;
  assign nl_input_fifo_0_run_cmp_input_rsc_dat = step_in_col_value_lpi_2_dfm_mx0[7:0];
  wire [255:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat
      = {output_rsci_idat_255_240 , output_rsci_idat_239_224 , output_rsci_idat_223_208
      , output_rsci_idat_207_192 , output_rsci_idat_191_176 , output_rsci_idat_175_160
      , output_rsci_idat_159_144 , output_rsci_idat_143_128 , output_rsci_idat_127_112
      , output_rsci_idat_111_96 , output_rsci_idat_95_80 , output_rsci_idat_79_64
      , output_rsci_idat_63_48 , output_rsci_idat_47_32 , output_rsci_idat_31_16
      , output_rsci_idat_15_0};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [11:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_addr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_addr_d_run
      = {6'b0, operator_16_false_mux_rmff};
  wire [0:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp_inst_ensig_cgo_iro_45;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp_inst_ensig_cgo_iro_45
      = ~ mux_302_itm;
  wire [0:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_inst_step_C_0_tr0;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_inst_step_C_0_tr0
      = ~ operator_32_false_acc_itm_31_1;
  Fifo_ODTYPE_16  accum_fifo_15_rsci (
      .input_rsc_dat(nl_accum_fifo_15_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_15_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_16  output_fifo_0_rsci (
      .input_rsc_dat(nl_output_fifo_0_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_0_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_15  accum_fifo_14_rsci (
      .input_rsc_dat(nl_accum_fifo_14_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_15  output_fifo_1_rsci (
      .input_rsc_dat(nl_output_fifo_1_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_14  accum_fifo_13_rsci (
      .input_rsc_dat(nl_accum_fifo_13_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_14  output_fifo_2_rsci (
      .input_rsc_dat(nl_output_fifo_2_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_13  accum_fifo_12_rsci (
      .input_rsc_dat(nl_accum_fifo_12_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_13  output_fifo_3_rsci (
      .input_rsc_dat(nl_output_fifo_3_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_12  accum_fifo_11_rsci (
      .input_rsc_dat(nl_accum_fifo_11_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_12  output_fifo_4_rsci (
      .input_rsc_dat(nl_output_fifo_4_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_11  accum_fifo_10_rsci (
      .input_rsc_dat(nl_accum_fifo_10_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_11  output_fifo_5_rsci (
      .input_rsc_dat(nl_output_fifo_5_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_10  accum_fifo_9_rsci (
      .input_rsc_dat(nl_accum_fifo_9_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_10  output_fifo_6_rsci (
      .input_rsc_dat(nl_output_fifo_6_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_9  accum_fifo_8_rsci (
      .input_rsc_dat(nl_accum_fifo_8_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_9  output_fifo_7_rsci (
      .input_rsc_dat(nl_output_fifo_7_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_8  accum_fifo_7_rsci (
      .input_rsc_dat(nl_accum_fifo_7_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_8  output_fifo_8_rsci (
      .input_rsc_dat(nl_output_fifo_8_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_7  accum_fifo_6_rsci (
      .input_rsc_dat(nl_accum_fifo_6_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_7  output_fifo_9_rsci (
      .input_rsc_dat(nl_output_fifo_9_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_6  accum_fifo_5_rsci (
      .input_rsc_dat(nl_accum_fifo_5_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_6  output_fifo_10_rsci (
      .input_rsc_dat(nl_output_fifo_10_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_5  accum_fifo_4_rsci (
      .input_rsc_dat(nl_accum_fifo_4_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_5  output_fifo_11_rsci (
      .input_rsc_dat(nl_output_fifo_11_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_4  accum_fifo_3_rsci (
      .input_rsc_dat(nl_accum_fifo_3_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_4  output_fifo_12_rsci (
      .input_rsc_dat(nl_output_fifo_12_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_3  accum_fifo_2_rsci (
      .input_rsc_dat(nl_accum_fifo_2_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_3  output_fifo_13_rsci (
      .input_rsc_dat(nl_output_fifo_13_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_ODTYPE_2  accum_fifo_1_rsci (
      .input_rsc_dat(nl_accum_fifo_1_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_8)
    );
  Fifo_ODTYPE_2  output_fifo_14_rsci (
      .input_rsc_dat(nl_output_fifo_14_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_362)
    );
  Fifo_IDTYPE_16  input_fifo_15_rsci (
      .input_rsc_dat(nl_input_fifo_15_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_15_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_15  input_fifo_14_rsci (
      .input_rsc_dat(nl_input_fifo_14_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_14  input_fifo_13_rsci (
      .input_rsc_dat(nl_input_fifo_13_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_13  input_fifo_12_rsci (
      .input_rsc_dat(nl_input_fifo_12_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_12  input_fifo_11_rsci (
      .input_rsc_dat(nl_input_fifo_11_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_11  input_fifo_10_rsci (
      .input_rsc_dat(nl_input_fifo_10_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_10  input_fifo_9_rsci (
      .input_rsc_dat(nl_input_fifo_9_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_9  input_fifo_8_rsci (
      .input_rsc_dat(nl_input_fifo_8_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_8  input_fifo_7_rsci (
      .input_rsc_dat(nl_input_fifo_7_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_7  input_fifo_6_rsci (
      .input_rsc_dat(nl_input_fifo_6_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_6  input_fifo_5_rsci (
      .input_rsc_dat(nl_input_fifo_5_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_5  input_fifo_4_rsci (
      .input_rsc_dat(nl_input_fifo_4_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_4  input_fifo_3_rsci (
      .input_rsc_dat(nl_input_fifo_3_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_3  input_fifo_2_rsci (
      .input_rsc_dat(nl_input_fifo_2_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  Fifo_IDTYPE_2  input_fifo_1_rsci (
      .input_rsc_dat(nl_input_fifo_1_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(pe_0_0_run_cmp_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(nl_pe_0_0_run_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  Fifo_ODTYPE_1  accum_fifo_0_run_cmp (
      .input_rsc_dat(nl_accum_fifo_0_run_cmp_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_0_run_cmp_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_0_run_cmp_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(nl_accum_fifo_0_run_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  Fifo_IDTYPE_1  input_fifo_0_run_cmp (
      .input_rsc_dat(nl_input_fifo_0_run_cmp_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_0_run_cmp_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_12)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .run_wen(run_wen),
      .input_rsci_oswt(reg_input_rsci_irdy_run_psct_cse),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weight_rsc_dat(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .run_wen(run_wen),
      .weight_rsci_oswt(reg_weight_rsci_irdy_run_psct_cse),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_idat_mxwt(weight_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .run_wen(run_wen),
      .output_rsci_oswt(reg_output_rsci_ivld_run_psct_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_idat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat[255:0])
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_loopIndicesIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(reg_loopIndicesIn_rsci_irdy_run_psct_cse),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_0_i_web_d(accumulation_buffer_rsc_0_0_i_web_d_reg),
      .accumulation_buffer_rsc_0_0_i_addr_d(accumulation_buffer_rsc_0_0_i_addr_d_reg),
      .accumulation_buffer_rsc_0_0_i_dout_d(accumulation_buffer_rsc_0_0_i_dout_d),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_0_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_0_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_0_i_dout_d_mxwt(accumulation_buffer_rsc_0_0_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_0_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_0_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_1_i_web_d(accumulation_buffer_rsc_0_1_i_web_d_reg),
      .accumulation_buffer_rsc_0_1_i_addr_d(accumulation_buffer_rsc_0_1_i_addr_d_reg),
      .accumulation_buffer_rsc_0_1_i_dout_d(accumulation_buffer_rsc_0_1_i_dout_d),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_1_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_1_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_1_i_dout_d_mxwt(accumulation_buffer_rsc_0_1_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_1_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_1_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_2_i_web_d(accumulation_buffer_rsc_0_2_i_web_d_reg),
      .accumulation_buffer_rsc_0_2_i_addr_d(accumulation_buffer_rsc_0_2_i_addr_d_reg),
      .accumulation_buffer_rsc_0_2_i_dout_d(accumulation_buffer_rsc_0_2_i_dout_d),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_2_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_2_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_2_i_dout_d_mxwt(accumulation_buffer_rsc_0_2_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_2_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_2_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_3_i_web_d(accumulation_buffer_rsc_0_3_i_web_d_reg),
      .accumulation_buffer_rsc_0_3_i_addr_d(accumulation_buffer_rsc_0_3_i_addr_d_reg),
      .accumulation_buffer_rsc_0_3_i_dout_d(accumulation_buffer_rsc_0_3_i_dout_d),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_3_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_3_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_3_i_dout_d_mxwt(accumulation_buffer_rsc_0_3_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_3_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_3_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_4_i_web_d(accumulation_buffer_rsc_0_4_i_web_d_reg),
      .accumulation_buffer_rsc_0_4_i_addr_d(accumulation_buffer_rsc_0_4_i_addr_d_reg),
      .accumulation_buffer_rsc_0_4_i_dout_d(accumulation_buffer_rsc_0_4_i_dout_d),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_4_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_4_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_4_i_dout_d_mxwt(accumulation_buffer_rsc_0_4_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_4_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_4_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_5_i_web_d(accumulation_buffer_rsc_0_5_i_web_d_reg),
      .accumulation_buffer_rsc_0_5_i_addr_d(accumulation_buffer_rsc_0_5_i_addr_d_reg),
      .accumulation_buffer_rsc_0_5_i_dout_d(accumulation_buffer_rsc_0_5_i_dout_d),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_5_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_5_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_5_i_dout_d_mxwt(accumulation_buffer_rsc_0_5_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_5_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_5_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_6_i_web_d(accumulation_buffer_rsc_0_6_i_web_d_reg),
      .accumulation_buffer_rsc_0_6_i_addr_d(accumulation_buffer_rsc_0_6_i_addr_d_reg),
      .accumulation_buffer_rsc_0_6_i_dout_d(accumulation_buffer_rsc_0_6_i_dout_d),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_6_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_6_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_6_i_dout_d_mxwt(accumulation_buffer_rsc_0_6_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_6_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_6_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_7_i_web_d(accumulation_buffer_rsc_0_7_i_web_d_reg),
      .accumulation_buffer_rsc_0_7_i_addr_d(accumulation_buffer_rsc_0_7_i_addr_d_reg),
      .accumulation_buffer_rsc_0_7_i_dout_d(accumulation_buffer_rsc_0_7_i_dout_d),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_7_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_7_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_7_i_dout_d_mxwt(accumulation_buffer_rsc_0_7_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_7_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_7_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_8_i_web_d(accumulation_buffer_rsc_0_8_i_web_d_reg),
      .accumulation_buffer_rsc_0_8_i_addr_d(accumulation_buffer_rsc_0_8_i_addr_d_reg),
      .accumulation_buffer_rsc_0_8_i_dout_d(accumulation_buffer_rsc_0_8_i_dout_d),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_8_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_8_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_8_i_dout_d_mxwt(accumulation_buffer_rsc_0_8_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_8_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_8_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_9_i_web_d(accumulation_buffer_rsc_0_9_i_web_d_reg),
      .accumulation_buffer_rsc_0_9_i_addr_d(accumulation_buffer_rsc_0_9_i_addr_d_reg),
      .accumulation_buffer_rsc_0_9_i_dout_d(accumulation_buffer_rsc_0_9_i_dout_d),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_9_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_9_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_9_i_dout_d_mxwt(accumulation_buffer_rsc_0_9_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_9_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_9_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_10_i_web_d(accumulation_buffer_rsc_0_10_i_web_d_reg),
      .accumulation_buffer_rsc_0_10_i_addr_d(accumulation_buffer_rsc_0_10_i_addr_d_reg),
      .accumulation_buffer_rsc_0_10_i_dout_d(accumulation_buffer_rsc_0_10_i_dout_d),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_10_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_10_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_10_i_dout_d_mxwt(accumulation_buffer_rsc_0_10_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_10_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_10_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_11_i_web_d(accumulation_buffer_rsc_0_11_i_web_d_reg),
      .accumulation_buffer_rsc_0_11_i_addr_d(accumulation_buffer_rsc_0_11_i_addr_d_reg),
      .accumulation_buffer_rsc_0_11_i_dout_d(accumulation_buffer_rsc_0_11_i_dout_d),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_11_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_11_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_11_i_dout_d_mxwt(accumulation_buffer_rsc_0_11_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_11_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_11_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_12_i_web_d(accumulation_buffer_rsc_0_12_i_web_d_reg),
      .accumulation_buffer_rsc_0_12_i_addr_d(accumulation_buffer_rsc_0_12_i_addr_d_reg),
      .accumulation_buffer_rsc_0_12_i_dout_d(accumulation_buffer_rsc_0_12_i_dout_d),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_12_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_12_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_12_i_dout_d_mxwt(accumulation_buffer_rsc_0_12_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_12_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_12_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_13_i_web_d(accumulation_buffer_rsc_0_13_i_web_d_reg),
      .accumulation_buffer_rsc_0_13_i_addr_d(accumulation_buffer_rsc_0_13_i_addr_d_reg),
      .accumulation_buffer_rsc_0_13_i_dout_d(accumulation_buffer_rsc_0_13_i_dout_d),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_13_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_13_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_13_i_dout_d_mxwt(accumulation_buffer_rsc_0_13_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_13_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_13_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_14_i_web_d(accumulation_buffer_rsc_0_14_i_web_d_reg),
      .accumulation_buffer_rsc_0_14_i_addr_d(accumulation_buffer_rsc_0_14_i_addr_d_reg),
      .accumulation_buffer_rsc_0_14_i_dout_d(accumulation_buffer_rsc_0_14_i_dout_d),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_14_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_14_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_14_i_dout_d_mxwt(accumulation_buffer_rsc_0_14_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_14_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_14_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_15_i_web_d(accumulation_buffer_rsc_0_15_i_web_d_reg),
      .accumulation_buffer_rsc_0_15_i_addr_d(accumulation_buffer_rsc_0_15_i_addr_d_reg),
      .accumulation_buffer_rsc_0_15_i_dout_d(accumulation_buffer_rsc_0_15_i_dout_d),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_15_i_oswt(reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse),
      .accumulation_buffer_rsc_0_15_i_addr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_addr_d_run[11:0]),
      .accumulation_buffer_rsc_0_15_i_dout_d_mxwt(accumulation_buffer_rsc_0_15_i_dout_d_mxwt),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct(and_377_rmff),
      .accumulation_buffer_rsc_0_15_i_web_d_run_psct_pff(and_372_rmff),
      .accumulation_buffer_rsc_0_15_i_oswt_pff(and_380_rmff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp_inst
      (
      .ensig_cgo_iro(and_368_rmff),
      .ensig_cgo_iro_1(and_364_rmff),
      .ensig_cgo_iro_30(and_17_rmff),
      .ensig_cgo_iro_45(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp_inst_ensig_cgo_iro_45[0:0]),
      .ensig_cgo_iro_46(and_23_rmff),
      .run_wen(run_wen),
      .ensig_cgo(reg_ensig_cgo_28_cse),
      .accum_fifo_15_rsci_ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ensig_cgo_1(reg_ensig_cgo_29_cse),
      .output_fifo_0_rsci_ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ensig_cgo_30(reg_ensig_cgo_47_cse),
      .input_fifo_15_rsci_ccs_ccore_en(input_fifo_15_rsci_ccs_ccore_en),
      .ensig_cgo_45(reg_ensig_cgo_45_cse),
      .pe_0_0_run_cmp_ccs_ccore_en(pe_0_0_run_cmp_ccs_ccore_en),
      .ensig_cgo_46(reg_ensig_cgo_46_cse),
      .accum_fifo_0_run_cmp_ccs_ccore_en(accum_fifo_0_run_cmp_ccs_ccore_en)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .step_C_0_tr0(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_inst_step_C_0_tr0[0:0])
    );
  assign operator_16_false_mux_rmff = MUX_v_6_2_2((step_step_sva[5:0]), (ROW_asn_142_itm[5:0]),
      and_dcpl_8);
  assign output_and_cse = run_wen & (~(or_dcpl_10 | (fsm_output[6:2]!=5'b00000) |
      or_dcpl_4 | operator_16_false_slc_operator_16_false_acc_16_itm | (~(step_if_3_step_if_3_if_step_if_3_if_nor_tmp
      & step_if_3_aif_step_if_3_aelse_step_if_3_aelse_nor_tmp & step_if_3_aif_1_step_if_3_aelse_1_step_if_3_aelse_1_nor_tmp))));
  assign and_17_rmff = (~ mux_tmp_80) & and_dcpl_5 & and_dcpl_15;
  assign or_137_nl = (~ (fsm_output[2])) | (fsm_output[8]);
  assign mux_103_nl = MUX_s_1_2_2((or_137_nl), or_tmp_121, fsm_output[1]);
  assign mux_104_nl = MUX_s_1_2_2(or_tmp_122, (mux_103_nl), operator_32_false_acc_itm_31_1);
  assign mux_102_nl = MUX_s_1_2_2((fsm_output[8]), or_47_cse, fsm_output[1]);
  assign mux_105_nl = MUX_s_1_2_2((mux_104_nl), (mux_102_nl), fsm_output[0]);
  assign and_23_rmff = (~ (mux_105_nl)) & and_dcpl_20 & (~ (fsm_output[4])) & and_dcpl_13;
  assign nand_111_cse = ~((fsm_output[2]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[3]));
  assign or_169_cse = (fsm_output[2]) | (~((fsm_output[6]) & (fsm_output[7]) & (fsm_output[3])));
  assign mux_130_cse = MUX_s_1_2_2(nand_111_cse, or_169_cse, fsm_output[5]);
  assign or_170_cse = (fsm_output[1]) | mux_130_cse;
  assign or_186_cse = (fsm_output[5]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~
      (fsm_output[6])) | (fsm_output[3]);
  assign or_201_cse = (fsm_output[2]) | (~ (fsm_output[6])) | (~ (fsm_output[7]))
      | (fsm_output[3]);
  assign nand_94_cse = ~((fsm_output[6]) & (fsm_output[7]) & (fsm_output[2]));
  assign or_187_cse = (fsm_output[7]) | (~ (fsm_output[6])) | (fsm_output[3]);
  assign or_220_cse = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[2]);
  assign or_228_cse = (fsm_output[6]) | (~((fsm_output[7]) & (fsm_output[2])));
  assign nand_100_cse = ~((fsm_output[7]) & (fsm_output[3]));
  assign mux_111_cse = MUX_s_1_2_2(or_tmp_129, or_tmp_133, fsm_output[6]);
  assign mux_109_cse = MUX_s_1_2_2(or_tmp_130, or_tmp_129, fsm_output[6]);
  assign mux_239_cse = MUX_s_1_2_2(nand_100_cse, or_tmp_225, fsm_output[6]);
  assign or_250_nl = (fsm_output[7]) | (fsm_output[3]);
  assign mux_234_cse = MUX_s_1_2_2((or_250_nl), or_tmp_225, fsm_output[6]);
  assign or_258_nl = (fsm_output[6]) | (fsm_output[7]) | (fsm_output[3]);
  assign mux_245_cse = MUX_s_1_2_2(or_187_cse, (or_258_nl), fsm_output[2]);
  assign or_176_cse = (fsm_output[7]) | (~((fsm_output[6]) & (fsm_output[3])));
  assign mux_142_cse = MUX_s_1_2_2(or_176_cse, mux_tmp_118, fsm_output[2]);
  assign or_177_cse = (fsm_output[5]) | mux_142_cse;
  assign mux_159_nl = MUX_s_1_2_2(mux_tmp_118, or_187_cse, fsm_output[2]);
  assign nand_10_cse = ~((fsm_output[5]) & (~ (mux_159_nl)));
  assign mux_210_cse = MUX_s_1_2_2(or_228_cse, mux_109_cse, fsm_output[3]);
  assign mux_143_nl = MUX_s_1_2_2(or_177_cse, nand_10_cse, fsm_output[1]);
  assign or_178_cse = (fsm_output[4]) | (mux_143_nl);
  assign mux_155_nl = MUX_s_1_2_2(or_186_cse, mux_130_cse, fsm_output[1]);
  assign mux_149_nl = MUX_s_1_2_2((fsm_output[3]), (~ (fsm_output[3])), fsm_output[6]);
  assign mux_150_nl = MUX_s_1_2_2(or_827_cse, (mux_149_nl), fsm_output[7]);
  assign mux_151_nl = MUX_s_1_2_2(or_176_cse, (mux_150_nl), fsm_output[2]);
  assign mux_152_nl = MUX_s_1_2_2((mux_151_nl), or_169_cse, fsm_output[5]);
  assign mux_153_nl = MUX_s_1_2_2((mux_152_nl), nand_10_cse, fsm_output[1]);
  assign mux_156_cse = MUX_s_1_2_2((mux_155_nl), (mux_153_nl), fsm_output[4]);
  assign or_225_nl = (fsm_output[3]) | nand_94_cse;
  assign mux_205_nl = MUX_s_1_2_2((or_225_nl), nand_tmp_14, fsm_output[4]);
  assign nor_143_nl = ~((fsm_output[3]) | mux_111_cse);
  assign mux_204_nl = MUX_s_1_2_2((nor_143_nl), nor_tmp_41, fsm_output[4]);
  assign mux_206_nl = MUX_s_1_2_2((mux_205_nl), (~ (mux_204_nl)), fsm_output[5]);
  assign or_223_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[6]))
      | (~ (fsm_output[7])) | (fsm_output[2]);
  assign mux_201_nl = MUX_s_1_2_2((~ nor_tmp_41), mux_210_cse, fsm_output[4]);
  assign mux_202_nl = MUX_s_1_2_2((or_223_nl), (mux_201_nl), fsm_output[5]);
  assign mux_207_cse = MUX_s_1_2_2((mux_206_nl), (mux_202_nl), fsm_output[1]);
  assign mux_199_cse = MUX_s_1_2_2(nand_tmp_14, or_220_cse, fsm_output[4]);
  assign or_222_cse = (fsm_output[5]) | mux_199_cse;
  assign mux_302_itm = MUX_s_1_2_2(mux_tmp_282, mux_tmp_280, and_463_cse);
  assign and_364_rmff = and_dcpl_7 & and_dcpl_360 & (operator_32_false_acc_itm_31_1
      | (fsm_output[0]));
  assign and_368_rmff = and_dcpl_31 & (~ (fsm_output[3])) & (fsm_output[2]) & (~
      (fsm_output[5])) & (~ (fsm_output[1]));
  assign and_372_rmff = and_dcpl_7 & and_dcpl_2 & (fsm_output[1:0]==2'b00) & (~ operator_16_false_slc_operator_16_false_acc_16_itm);
  assign and_377_rmff = and_dcpl_376 & and_dcpl_35 & step_if_1_acc_cse_32 & (~ step_if_2_if_step_if_2_if_and_tmp);
  assign or_329_nl = (fsm_output[2:0]!=3'b100);
  assign mux_303_nl = MUX_s_1_2_2((or_329_nl), mux_tmp_80, step_if_1_acc_cse_32);
  assign nand_84_nl = ~(step_if_1_acc_cse_32 & (fsm_output[2:0]==3'b011));
  assign mux_304_nl = MUX_s_1_2_2((mux_303_nl), (nand_84_nl), operator_16_false_slc_operator_16_false_acc_16_itm);
  assign or_326_nl = operator_16_false_slc_operator_16_false_acc_16_itm | (fsm_output[2:0]!=3'b100);
  assign mux_305_nl = MUX_s_1_2_2((mux_304_nl), (or_326_nl), step_if_2_if_step_if_2_if_and_tmp);
  assign and_380_rmff = (~ (mux_305_nl)) & and_dcpl_6 & and_dcpl_4 & (~ (fsm_output[5]));
  assign or_338_cse = (fsm_output[7:3]!=5'b00000);
  assign nor_133_cse = ~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[8]));
  assign nor_150_cse = ~((fsm_output[7:2]!=6'b000000));
  assign mux_306_cse = MUX_s_1_2_2(nor_133_cse, (fsm_output[8]), or_338_cse);
  assign input_reg_and_1_cse = run_wen & (~(or_dcpl_66 | or_dcpl_57));
  assign input_reg_and_2_cse = run_wen & (~(or_dcpl_66 | or_dcpl_59));
  assign input_reg_and_3_cse = run_wen & (~(or_dcpl_66 | or_dcpl_61));
  assign input_reg_and_4_cse = run_wen & (~(or_dcpl_66 | or_dcpl_63));
  assign input_reg_and_5_cse = run_wen & (~(or_dcpl_76 | or_dcpl_44));
  assign input_reg_and_6_cse = run_wen & (~(or_dcpl_76 | or_dcpl_50));
  assign input_reg_and_7_cse = run_wen & (~(or_dcpl_76 | or_dcpl_52));
  assign input_reg_and_8_cse = run_wen & (~(or_dcpl_76 | or_dcpl_54));
  assign input_reg_and_9_cse = run_wen & (~(or_dcpl_76 | or_dcpl_57));
  assign input_reg_and_10_cse = run_wen & (~(or_dcpl_76 | or_dcpl_59));
  assign input_reg_and_11_cse = run_wen & (~(or_dcpl_76 | or_dcpl_61));
  assign input_reg_and_12_cse = run_wen & (~(or_dcpl_76 | or_dcpl_63));
  assign input_reg_and_13_cse = run_wen & (~(or_dcpl_85 | or_dcpl_44));
  assign input_reg_and_14_cse = run_wen & (~(or_dcpl_85 | or_dcpl_50));
  assign input_reg_and_16_cse = run_wen & (~(or_dcpl_85 | or_dcpl_54));
  assign input_reg_and_17_cse = run_wen & (~(or_dcpl_85 | or_dcpl_57));
  assign input_reg_and_18_cse = run_wen & (~(or_dcpl_85 | or_dcpl_59));
  assign input_reg_and_19_cse = run_wen & (~(or_dcpl_85 | or_dcpl_61));
  assign input_reg_and_20_cse = run_wen & (~(or_dcpl_85 | or_dcpl_63));
  assign input_reg_and_21_cse = run_wen & (~(or_dcpl_48 | or_dcpl_95));
  assign input_reg_and_22_cse = run_wen & (~(or_dcpl_48 | or_dcpl_97));
  assign input_reg_and_23_cse = run_wen & (~(or_dcpl_48 | or_dcpl_99));
  assign input_reg_and_24_cse = run_wen & (~(or_dcpl_48 | or_dcpl_101));
  assign input_reg_and_25_cse = run_wen & (~(or_dcpl_48 | or_dcpl_103));
  assign input_reg_and_26_cse = run_wen & (~(or_dcpl_48 | or_dcpl_32));
  assign input_reg_and_27_cse = run_wen & (~(or_dcpl_48 | or_dcpl_38));
  assign input_reg_and_28_cse = run_wen & (~(or_dcpl_48 | or_dcpl_41));
  assign input_reg_and_29_cse = run_wen & (~(or_dcpl_66 | or_dcpl_95));
  assign input_reg_and_30_cse = run_wen & (~(or_dcpl_66 | or_dcpl_97));
  assign input_reg_and_31_cse = run_wen & (~(or_dcpl_66 | or_dcpl_99));
  assign input_reg_and_32_cse = run_wen & (~(or_dcpl_66 | or_dcpl_101));
  assign input_reg_and_33_cse = run_wen & (~(or_dcpl_66 | or_dcpl_103));
  assign input_reg_and_34_cse = run_wen & (~(or_dcpl_66 | or_dcpl_32));
  assign input_reg_and_35_cse = run_wen & (~(or_dcpl_66 | or_dcpl_38));
  assign input_reg_and_36_cse = run_wen & (~(or_dcpl_66 | or_dcpl_41));
  assign input_reg_and_37_cse = run_wen & (~(or_dcpl_76 | or_dcpl_95));
  assign input_reg_and_38_cse = run_wen & (~(or_dcpl_76 | or_dcpl_97));
  assign input_reg_and_39_cse = run_wen & (~(or_dcpl_76 | or_dcpl_99));
  assign input_reg_and_40_cse = run_wen & (~(or_dcpl_76 | or_dcpl_101));
  assign input_reg_and_41_cse = run_wen & (~(or_dcpl_76 | or_dcpl_103));
  assign input_reg_and_42_cse = run_wen & (~(or_dcpl_76 | or_dcpl_32));
  assign input_reg_and_43_cse = run_wen & (~(or_dcpl_76 | or_dcpl_38));
  assign input_reg_and_44_cse = run_wen & (~(or_dcpl_76 | or_dcpl_41));
  assign input_reg_and_45_cse = run_wen & (~(or_dcpl_85 | or_dcpl_95));
  assign input_reg_and_46_cse = run_wen & (~(or_dcpl_85 | or_dcpl_97));
  assign input_reg_and_47_cse = run_wen & (~(or_dcpl_85 | or_dcpl_99));
  assign input_reg_and_48_cse = run_wen & (~(or_dcpl_85 | or_dcpl_101));
  assign input_reg_and_49_cse = run_wen & (~(or_dcpl_85 | or_dcpl_103));
  assign input_reg_and_50_cse = run_wen & (~(or_dcpl_85 | or_dcpl_32));
  assign input_reg_and_51_cse = run_wen & (~(or_dcpl_85 | or_dcpl_38));
  assign input_reg_and_52_cse = run_wen & (~(or_dcpl_85 | or_dcpl_41));
  assign input_reg_and_53_cse = run_wen & (~(or_dcpl_133 | or_dcpl_44));
  assign input_reg_and_54_cse = run_wen & (~(or_dcpl_133 | or_dcpl_50));
  assign input_reg_and_55_cse = run_wen & (~(or_dcpl_133 | or_dcpl_52));
  assign input_reg_and_56_cse = run_wen & (~(or_dcpl_133 | or_dcpl_54));
  assign input_reg_and_57_cse = run_wen & (~(or_dcpl_133 | or_dcpl_57));
  assign input_reg_and_58_cse = run_wen & (~(or_dcpl_133 | or_dcpl_59));
  assign input_reg_and_59_cse = run_wen & (~(or_dcpl_133 | or_dcpl_61));
  assign input_reg_and_60_cse = run_wen & (~(or_dcpl_133 | or_dcpl_63));
  assign input_reg_and_61_cse = run_wen & (~(or_dcpl_142 | or_dcpl_44));
  assign input_reg_and_62_cse = run_wen & (~(or_dcpl_142 | or_dcpl_50));
  assign input_reg_and_63_cse = run_wen & (~(or_dcpl_142 | or_dcpl_52));
  assign input_reg_and_64_cse = run_wen & (~(or_dcpl_142 | or_dcpl_54));
  assign input_reg_and_65_cse = run_wen & (~(or_dcpl_142 | or_dcpl_57));
  assign input_reg_and_66_cse = run_wen & (~(or_dcpl_142 | or_dcpl_59));
  assign input_reg_and_67_cse = run_wen & (~(or_dcpl_142 | or_dcpl_61));
  assign input_reg_and_68_cse = run_wen & (~(or_dcpl_142 | or_dcpl_63));
  assign input_reg_and_69_cse = run_wen & (~(or_dcpl_151 | or_dcpl_44));
  assign input_reg_and_70_cse = run_wen & (~(or_dcpl_151 | or_dcpl_50));
  assign input_reg_and_71_cse = run_wen & (~(or_dcpl_151 | or_dcpl_52));
  assign input_reg_and_72_cse = run_wen & (~(or_dcpl_151 | or_dcpl_54));
  assign input_reg_and_73_cse = run_wen & (~(or_dcpl_151 | or_dcpl_57));
  assign input_reg_and_74_cse = run_wen & (~(or_dcpl_151 | or_dcpl_59));
  assign input_reg_and_75_cse = run_wen & (~(or_dcpl_151 | or_dcpl_63));
  assign input_reg_and_76_cse = run_wen & (~(or_dcpl_159 | or_dcpl_44));
  assign input_reg_and_77_cse = run_wen & (~(or_dcpl_159 | or_dcpl_50));
  assign input_reg_and_78_cse = run_wen & (~(or_dcpl_159 | or_dcpl_52));
  assign input_reg_and_79_cse = run_wen & (~(or_dcpl_159 | or_dcpl_54));
  assign input_reg_and_80_cse = run_wen & (~(or_dcpl_159 | or_dcpl_57));
  assign input_reg_and_81_cse = run_wen & (~(or_dcpl_159 | or_dcpl_59));
  assign input_reg_and_82_cse = run_wen & (~(or_dcpl_159 | or_dcpl_61));
  assign input_reg_and_83_cse = run_wen & (~(or_dcpl_159 | or_dcpl_63));
  assign input_reg_and_84_cse = run_wen & (~(or_dcpl_133 | or_dcpl_95));
  assign input_reg_and_85_cse = run_wen & (~(or_dcpl_133 | or_dcpl_97));
  assign input_reg_and_86_cse = run_wen & (~(or_dcpl_133 | or_dcpl_99));
  assign input_reg_and_87_cse = run_wen & (~(or_dcpl_133 | or_dcpl_101));
  assign input_reg_and_88_cse = run_wen & (~(or_dcpl_133 | or_dcpl_103));
  assign input_reg_and_89_cse = run_wen & (~(or_dcpl_133 | or_dcpl_32));
  assign input_reg_and_91_cse = run_wen & (~(or_dcpl_133 | or_dcpl_41));
  assign input_reg_and_92_cse = run_wen & (~(or_dcpl_142 | or_dcpl_95));
  assign input_reg_and_93_cse = run_wen & (~(or_dcpl_142 | or_dcpl_97));
  assign input_reg_and_94_cse = run_wen & (~(or_dcpl_142 | or_dcpl_99));
  assign input_reg_and_95_cse = run_wen & (~(or_dcpl_142 | or_dcpl_101));
  assign input_reg_and_96_cse = run_wen & (~(or_dcpl_142 | or_dcpl_103));
  assign input_reg_and_97_cse = run_wen & (~(or_dcpl_142 | or_dcpl_32));
  assign input_reg_and_98_cse = run_wen & (~(or_dcpl_142 | or_dcpl_38));
  assign input_reg_and_99_cse = run_wen & (~(or_dcpl_142 | or_dcpl_41));
  assign input_reg_and_100_cse = run_wen & (~(or_dcpl_151 | or_dcpl_95));
  assign input_reg_and_101_cse = run_wen & (~(or_dcpl_151 | or_dcpl_97));
  assign input_reg_and_102_cse = run_wen & (~(or_dcpl_151 | or_dcpl_99));
  assign input_reg_and_103_cse = run_wen & (~(or_dcpl_151 | or_dcpl_101));
  assign input_reg_and_104_cse = run_wen & (~(or_dcpl_151 | or_dcpl_103));
  assign input_reg_and_105_cse = run_wen & (~(or_dcpl_151 | or_dcpl_32));
  assign input_reg_and_107_cse = run_wen & (~(or_dcpl_151 | or_dcpl_41));
  assign input_reg_and_108_cse = run_wen & (~(or_dcpl_159 | or_dcpl_95));
  assign input_reg_and_109_cse = run_wen & (~(or_dcpl_159 | or_dcpl_97));
  assign input_reg_and_110_cse = run_wen & (~(or_dcpl_159 | or_dcpl_99));
  assign input_reg_and_111_cse = run_wen & (~(or_dcpl_159 | or_dcpl_101));
  assign input_reg_and_112_cse = run_wen & (~(or_dcpl_159 | or_dcpl_103));
  assign input_reg_and_113_cse = run_wen & (~(or_dcpl_159 | or_dcpl_32));
  assign input_reg_and_114_cse = run_wen & (~(or_dcpl_159 | or_dcpl_38));
  assign input_reg_and_115_cse = run_wen & (~(or_dcpl_159 | or_dcpl_41));
  assign input_reg_and_116_cse = run_wen & (~(or_dcpl_201 | or_dcpl_44));
  assign input_reg_and_117_cse = run_wen & (~(or_dcpl_201 | or_dcpl_50));
  assign input_reg_and_118_cse = run_wen & (~(or_dcpl_201 | or_dcpl_52));
  assign input_reg_and_119_cse = run_wen & (~(or_dcpl_201 | or_dcpl_54));
  assign input_reg_and_120_cse = run_wen & (~(or_dcpl_201 | or_dcpl_57));
  assign input_reg_and_121_cse = run_wen & (~(or_dcpl_201 | or_dcpl_59));
  assign input_reg_and_123_cse = run_wen & (~(or_dcpl_201 | or_dcpl_63));
  assign input_reg_and_124_cse = run_wen & (~(or_dcpl_210 | or_dcpl_44));
  assign input_reg_and_125_cse = run_wen & (~(or_dcpl_210 | or_dcpl_50));
  assign input_reg_and_126_cse = run_wen & (~(or_dcpl_210 | or_dcpl_52));
  assign input_reg_and_127_cse = run_wen & (~(or_dcpl_210 | or_dcpl_54));
  assign input_reg_and_128_cse = run_wen & (~(or_dcpl_210 | or_dcpl_57));
  assign input_reg_and_129_cse = run_wen & (~(or_dcpl_210 | or_dcpl_59));
  assign input_reg_and_130_cse = run_wen & (~(or_dcpl_210 | or_dcpl_61));
  assign input_reg_and_131_cse = run_wen & (~(or_dcpl_210 | or_dcpl_63));
  assign input_reg_and_132_cse = run_wen & (~(or_dcpl_219 | or_dcpl_44));
  assign input_reg_and_133_cse = run_wen & (~(or_dcpl_219 | or_dcpl_50));
  assign input_reg_and_134_cse = run_wen & (~(or_dcpl_219 | or_dcpl_52));
  assign input_reg_and_135_cse = run_wen & (~(or_dcpl_219 | or_dcpl_54));
  assign input_reg_and_136_cse = run_wen & (~(or_dcpl_219 | or_dcpl_57));
  assign input_reg_and_137_cse = run_wen & (~(or_dcpl_219 | or_dcpl_59));
  assign input_reg_and_139_cse = run_wen & (~(or_dcpl_219 | or_dcpl_63));
  assign input_reg_and_140_cse = run_wen & (~(or_dcpl_228 | or_dcpl_44));
  assign input_reg_and_141_cse = run_wen & (~(or_dcpl_228 | or_dcpl_50));
  assign input_reg_and_142_cse = run_wen & (~(or_dcpl_228 | or_dcpl_52));
  assign input_reg_and_143_cse = run_wen & (~(or_dcpl_228 | or_dcpl_54));
  assign input_reg_and_144_cse = run_wen & (~(or_dcpl_228 | or_dcpl_57));
  assign input_reg_and_145_cse = run_wen & (~(or_dcpl_228 | or_dcpl_59));
  assign input_reg_and_146_cse = run_wen & (~(or_dcpl_228 | or_dcpl_61));
  assign input_reg_and_147_cse = run_wen & (~(or_dcpl_228 | or_dcpl_63));
  assign input_reg_and_148_cse = run_wen & (~(or_dcpl_201 | or_dcpl_95));
  assign input_reg_and_149_cse = run_wen & (~(or_dcpl_201 | or_dcpl_97));
  assign input_reg_and_150_cse = run_wen & (~(or_dcpl_201 | or_dcpl_99));
  assign input_reg_and_151_cse = run_wen & (~(or_dcpl_201 | or_dcpl_101));
  assign input_reg_and_152_cse = run_wen & (~(or_dcpl_201 | or_dcpl_103));
  assign input_reg_and_153_cse = run_wen & (~(or_dcpl_201 | or_dcpl_32));
  assign input_reg_and_155_cse = run_wen & (~(or_dcpl_201 | or_dcpl_41));
  assign input_reg_and_156_cse = run_wen & (~(or_dcpl_210 | or_dcpl_95));
  assign input_reg_and_157_cse = run_wen & (~(or_dcpl_210 | or_dcpl_97));
  assign input_reg_and_158_cse = run_wen & (~(or_dcpl_210 | or_dcpl_99));
  assign input_reg_and_159_cse = run_wen & (~(or_dcpl_210 | or_dcpl_101));
  assign input_reg_and_160_cse = run_wen & (~(or_dcpl_210 | or_dcpl_103));
  assign input_reg_and_161_cse = run_wen & (~(or_dcpl_210 | or_dcpl_32));
  assign input_reg_and_162_cse = run_wen & (~(or_dcpl_210 | or_dcpl_38));
  assign input_reg_and_163_cse = run_wen & (~(or_dcpl_210 | or_dcpl_41));
  assign input_reg_and_164_cse = run_wen & (~(or_dcpl_219 | or_dcpl_95));
  assign input_reg_and_165_cse = run_wen & (~(or_dcpl_219 | or_dcpl_97));
  assign input_reg_and_166_cse = run_wen & (~(or_dcpl_219 | or_dcpl_99));
  assign input_reg_and_167_cse = run_wen & (~(or_dcpl_219 | or_dcpl_101));
  assign input_reg_and_168_cse = run_wen & (~(or_dcpl_219 | or_dcpl_103));
  assign input_reg_and_169_cse = run_wen & (~(or_dcpl_219 | or_dcpl_32));
  assign input_reg_and_171_cse = run_wen & (~(or_dcpl_219 | or_dcpl_41));
  assign input_reg_and_172_cse = run_wen & (~(or_dcpl_228 | or_dcpl_95));
  assign input_reg_and_173_cse = run_wen & (~(or_dcpl_228 | or_dcpl_97));
  assign input_reg_and_174_cse = run_wen & (~(or_dcpl_228 | or_dcpl_99));
  assign input_reg_and_175_cse = run_wen & (~(or_dcpl_228 | or_dcpl_101));
  assign input_reg_and_176_cse = run_wen & (~(or_dcpl_228 | or_dcpl_103));
  assign input_reg_and_177_cse = run_wen & (~(or_dcpl_228 | or_dcpl_32));
  assign input_reg_and_178_cse = run_wen & (~(or_dcpl_228 | or_dcpl_38));
  assign input_reg_and_179_cse = run_wen & (~(or_dcpl_228 | or_dcpl_41));
  assign input_reg_and_180_cse = run_wen & (~(or_dcpl_269 | or_dcpl_44));
  assign input_reg_and_181_cse = run_wen & (~(or_dcpl_269 | or_dcpl_50));
  assign input_reg_and_182_cse = run_wen & (~(or_dcpl_269 | or_dcpl_52));
  assign input_reg_and_183_cse = run_wen & (~(or_dcpl_269 | or_dcpl_54));
  assign input_reg_and_184_cse = run_wen & (~(or_dcpl_269 | or_dcpl_57));
  assign input_reg_and_185_cse = run_wen & (~(or_dcpl_269 | or_dcpl_59));
  assign input_reg_and_187_cse = run_wen & (~(or_dcpl_269 | or_dcpl_63));
  assign input_reg_and_188_cse = run_wen & (~(or_dcpl_278 | or_dcpl_44));
  assign input_reg_and_189_cse = run_wen & (~(or_dcpl_278 | or_dcpl_50));
  assign input_reg_and_190_cse = run_wen & (~(or_dcpl_278 | or_dcpl_52));
  assign input_reg_and_191_cse = run_wen & (~(or_dcpl_278 | or_dcpl_54));
  assign input_reg_and_192_cse = run_wen & (~(or_dcpl_278 | or_dcpl_57));
  assign input_reg_and_193_cse = run_wen & (~(or_dcpl_278 | or_dcpl_59));
  assign input_reg_and_194_cse = run_wen & (~(or_dcpl_278 | or_dcpl_61));
  assign input_reg_and_195_cse = run_wen & (~(or_dcpl_278 | or_dcpl_63));
  assign input_reg_and_196_cse = run_wen & (~(or_dcpl_287 | or_dcpl_44));
  assign input_reg_and_197_cse = run_wen & (~(or_dcpl_287 | or_dcpl_50));
  assign input_reg_and_198_cse = run_wen & (~(or_dcpl_287 | or_dcpl_52));
  assign input_reg_and_199_cse = run_wen & (~(or_dcpl_287 | or_dcpl_54));
  assign input_reg_and_200_cse = run_wen & (~(or_dcpl_287 | or_dcpl_57));
  assign input_reg_and_201_cse = run_wen & (~(or_dcpl_287 | or_dcpl_59));
  assign input_reg_and_203_cse = run_wen & (~(or_dcpl_287 | or_dcpl_63));
  assign input_reg_and_204_cse = run_wen & (~(or_dcpl_29 | or_dcpl_44));
  assign input_reg_and_205_cse = run_wen & (~(or_dcpl_29 | or_dcpl_50));
  assign input_reg_and_206_cse = run_wen & (~(or_dcpl_29 | or_dcpl_52));
  assign input_reg_and_207_cse = run_wen & (~(or_dcpl_29 | or_dcpl_54));
  assign input_reg_and_208_cse = run_wen & (~(or_dcpl_29 | or_dcpl_57));
  assign input_reg_and_209_cse = run_wen & (~(or_dcpl_29 | or_dcpl_59));
  assign input_reg_and_210_cse = run_wen & (~(or_dcpl_29 | or_dcpl_61));
  assign input_reg_and_211_cse = run_wen & (~(or_dcpl_29 | or_dcpl_63));
  assign input_reg_and_212_cse = run_wen & (~(or_dcpl_269 | or_dcpl_95));
  assign input_reg_and_213_cse = run_wen & (~(or_dcpl_269 | or_dcpl_97));
  assign input_reg_and_214_cse = run_wen & (~(or_dcpl_269 | or_dcpl_99));
  assign input_reg_and_215_cse = run_wen & (~(or_dcpl_269 | or_dcpl_101));
  assign input_reg_and_216_cse = run_wen & (~(or_dcpl_269 | or_dcpl_103));
  assign input_reg_and_217_cse = run_wen & (~(or_dcpl_269 | or_dcpl_32));
  assign input_reg_and_219_cse = run_wen & (~(or_dcpl_269 | or_dcpl_41));
  assign input_reg_and_220_cse = run_wen & (~(or_dcpl_278 | or_dcpl_95));
  assign input_reg_and_221_cse = run_wen & (~(or_dcpl_278 | or_dcpl_97));
  assign input_reg_and_222_cse = run_wen & (~(or_dcpl_278 | or_dcpl_99));
  assign input_reg_and_223_cse = run_wen & (~(or_dcpl_278 | or_dcpl_101));
  assign input_reg_and_224_cse = run_wen & (~(or_dcpl_278 | or_dcpl_103));
  assign input_reg_and_225_cse = run_wen & (~(or_dcpl_278 | or_dcpl_32));
  assign input_reg_and_226_cse = run_wen & (~(or_dcpl_278 | or_dcpl_38));
  assign input_reg_and_227_cse = run_wen & (~(or_dcpl_278 | or_dcpl_41));
  assign input_reg_and_228_cse = run_wen & (~(or_dcpl_287 | or_dcpl_95));
  assign input_reg_and_229_cse = run_wen & (~(or_dcpl_287 | or_dcpl_97));
  assign input_reg_and_230_cse = run_wen & (~(or_dcpl_287 | or_dcpl_99));
  assign input_reg_and_231_cse = run_wen & (~(or_dcpl_287 | or_dcpl_101));
  assign input_reg_and_232_cse = run_wen & (~(or_dcpl_287 | or_dcpl_103));
  assign input_reg_and_233_cse = run_wen & (~(or_dcpl_287 | or_dcpl_32));
  assign or_645_cse = (fsm_output[7:4]!=4'b0000);
  assign input_reg_and_239_cse = run_wen & (~(or_dcpl_29 | or_dcpl_99));
  assign and_443_m1c = and_dcpl_7 & and_dcpl_54;
  assign or_47_cse = (~ (fsm_output[8])) | (fsm_output[2]);
  assign or_52_cse = (fsm_output[4:3]!=2'b00);
  assign and_cse = (fsm_output[4:3]==2'b11);
  assign nor_174_cse = ~((~((fsm_output[2:1]!=2'b00))) | (fsm_output[8]));
  assign or_674_nl = (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_322_cse = MUX_s_1_2_2(nor_133_cse, (or_674_nl), fsm_output[2]);
  assign or_58_cse = (fsm_output[4]) | (fsm_output[7]);
  assign or_55_cse = (fsm_output[6:5]!=2'b00);
  assign or_94_cse = (fsm_output[7:6]!=2'b00);
  assign operator_16_false_and_1_cse = run_wen & (~(or_dcpl_29 | or_dcpl_32)) & operator_32_false_acc_itm_31_1;
  assign or_743_cse = (fsm_output[6]) | mux_tmp_103;
  assign mux_377_cse = MUX_s_1_2_2(or_743_cse, or_187_cse, fsm_output[2]);
  assign or_765_cse = (~ (fsm_output[6])) | (fsm_output[7]) | (~ (fsm_output[3]));
  assign mux_434_cse = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[6]);
  assign or_827_cse = (fsm_output[6]) | (~ (fsm_output[3]));
  assign nand_62_cse = ~((fsm_output[7]) & (fsm_output[2]) & (fsm_output[6]) & (~
      (fsm_output[3])));
  assign and_463_cse = (fsm_output[1:0]==2'b11);
  assign nl_step_if_1_acc_nl = ({17'b10000000000000000 , step_step_sva}) + conv_u2u_32_33(~
      step_mul_itm) + 33'b000000000000000000000000000000001;
  assign step_if_1_acc_nl = nl_step_if_1_acc_nl[32:0];
  assign step_if_1_acc_itm_32_1 = readslicef_33_1_32((step_if_1_acc_nl));
  assign nl_operator_16_false_acc_nl_1 = conv_u2u_12_13(step_step_sva[15:4]) + 13'b1111111111111;
  assign operator_16_false_acc_nl_1 = nl_operator_16_false_acc_nl_1[12:0];
  assign operator_16_false_acc_itm_12_1 = readslicef_13_1_12((operator_16_false_acc_nl_1));
  assign step_if_2_if_step_if_2_if_and_tmp = (loopIndicesIn_crt_sva==48'b000000000000000000000000000000000000000000000000);
  assign step_mul_itm = conv_u2u_32_32((paramsIn_crt_sva_127_32[31:16]) * (paramsIn_crt_sva_127_32[15:0]));
  assign step_in_col_value_lpi_2_dfm_mx0 = MUX_v_128_2_2(step_in_col_value_lpi_2,
      input_rsci_idat_mxwt, step_if_1_acc_cse_32);
  assign nl_operator_16_false_3_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_sva_127_32[95:80])
      + 17'b11111111111111111;
  assign operator_16_false_3_acc_psp_sva_1 = nl_operator_16_false_3_acc_psp_sva_1[16:0];
  assign nl_operator_16_false_2_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_sva_127_32[79:64])
      + 17'b11111111111111111;
  assign operator_16_false_2_acc_psp_sva_1 = nl_operator_16_false_2_acc_psp_sva_1[16:0];
  assign nl_operator_16_false_1_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_sva_127_32[63:48])
      + 17'b11111111111111111;
  assign operator_16_false_1_acc_psp_sva_1 = nl_operator_16_false_1_acc_psp_sva_1[16:0];
  assign step_if_3_aif_1_step_if_3_aelse_1_step_if_3_aelse_1_nor_tmp = ~(((loopIndicesIn_crt_sva[47:32])
      != (operator_16_false_3_acc_psp_sva_1[15:0])) | (operator_16_false_3_acc_psp_sva_1[16]));
  assign step_if_3_aif_step_if_3_aelse_step_if_3_aelse_nor_tmp = ~(((loopIndicesIn_crt_sva[31:16])
      != (operator_16_false_2_acc_psp_sva_1[15:0])) | (operator_16_false_2_acc_psp_sva_1[16]));
  assign step_if_3_step_if_3_if_step_if_3_if_nor_tmp = ~(((loopIndicesIn_crt_sva[15:0])
      != (operator_16_false_1_acc_psp_sva_1[15:0])) | (operator_16_false_1_acc_psp_sva_1[16]));
  assign and_dcpl_1 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_2 = (fsm_output[2]) & (~ (fsm_output[5]));
  assign and_dcpl_3 = and_dcpl_2 & and_dcpl_1;
  assign and_dcpl_4 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_5 = ~((fsm_output[8:7]!=2'b00));
  assign and_dcpl_6 = and_dcpl_5 & (~ (fsm_output[6]));
  assign and_dcpl_7 = and_dcpl_6 & and_dcpl_4;
  assign and_dcpl_8 = and_dcpl_7 & and_dcpl_3;
  assign or_dcpl_4 = ~((fsm_output[1:0]==2'b11));
  assign or_dcpl_10 = (fsm_output[8:7]!=2'b00);
  assign and_dcpl_10 = ~((fsm_output[2]) | (fsm_output[5]));
  assign and_dcpl_11 = and_dcpl_10 & and_463_cse;
  assign and_dcpl_12 = and_dcpl_7 & and_dcpl_11;
  assign and_dcpl_13 = ~((fsm_output[3]) | (fsm_output[5]));
  assign and_dcpl_14 = ~((fsm_output[6]) | (fsm_output[4]));
  assign and_dcpl_15 = and_dcpl_14 & and_dcpl_13;
  assign or_133_nl = (fsm_output[2:1]!=2'b10);
  assign or_132_nl = (fsm_output[2:1]!=2'b01);
  assign mux_tmp_80 = MUX_s_1_2_2((or_133_nl), (or_132_nl), fsm_output[0]);
  assign or_tmp_121 = (fsm_output[2]) | (fsm_output[8]);
  assign or_tmp_122 = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[8]);
  assign and_dcpl_20 = ~((fsm_output[7:6]!=2'b00));
  assign or_dcpl_14 = (fsm_output[2]) | (fsm_output[5]);
  assign and_dcpl_24 = (step_step_sva[1:0]==2'b11);
  assign and_dcpl_25 = and_dcpl_24 & (step_step_sva[2]);
  assign and_dcpl_27 = and_463_cse & operator_16_false_slc_operator_16_false_acc_12_svs
      & (step_step_sva[3]);
  assign and_dcpl_29 = ~((fsm_output[3:2]!=2'b00));
  assign and_dcpl_31 = and_dcpl_5 & and_dcpl_14;
  assign and_dcpl_32 = and_dcpl_31 & and_dcpl_29 & (~ (fsm_output[5]));
  assign and_dcpl_33 = and_dcpl_32 & and_dcpl_27 & and_dcpl_25;
  assign and_dcpl_34 = (~ (fsm_output[5])) & (fsm_output[1]);
  assign and_dcpl_35 = and_dcpl_34 & (fsm_output[0]);
  assign and_dcpl_40 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_41 = and_dcpl_2 & and_dcpl_40;
  assign and_dcpl_42 = and_dcpl_7 & and_dcpl_41;
  assign and_dcpl_43 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_44 = and_dcpl_2 & and_dcpl_43;
  assign and_dcpl_45 = and_dcpl_7 & and_dcpl_44;
  assign and_dcpl_46 = and_dcpl_2 & and_463_cse;
  assign and_dcpl_47 = and_dcpl_7 & and_dcpl_46;
  assign and_dcpl_48 = and_dcpl_10 & and_dcpl_1;
  assign and_dcpl_49 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_50 = and_dcpl_6 & and_dcpl_49;
  assign and_dcpl_51 = and_dcpl_50 & and_dcpl_48;
  assign and_dcpl_52 = and_dcpl_10 & and_dcpl_40;
  assign and_dcpl_53 = and_dcpl_50 & and_dcpl_52;
  assign and_dcpl_54 = and_dcpl_10 & and_dcpl_43;
  assign and_dcpl_55 = and_dcpl_50 & and_dcpl_54;
  assign and_dcpl_56 = and_dcpl_50 & and_dcpl_11;
  assign and_dcpl_57 = and_dcpl_50 & and_dcpl_3;
  assign and_dcpl_58 = and_dcpl_50 & and_dcpl_41;
  assign and_dcpl_59 = and_dcpl_50 & and_dcpl_44;
  assign and_dcpl_60 = and_dcpl_50 & and_dcpl_46;
  assign and_dcpl_61 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_62 = and_dcpl_6 & and_dcpl_61;
  assign and_dcpl_63 = and_dcpl_62 & and_dcpl_48;
  assign and_dcpl_64 = and_dcpl_62 & and_dcpl_52;
  assign and_dcpl_65 = and_dcpl_62 & and_dcpl_54;
  assign and_dcpl_66 = and_dcpl_62 & and_dcpl_11;
  assign and_dcpl_67 = and_dcpl_62 & and_dcpl_3;
  assign and_dcpl_68 = and_dcpl_62 & and_dcpl_41;
  assign and_dcpl_69 = and_dcpl_62 & and_dcpl_44;
  assign and_dcpl_70 = and_dcpl_62 & and_dcpl_46;
  assign and_dcpl_72 = and_dcpl_6 & and_cse;
  assign and_dcpl_73 = and_dcpl_72 & and_dcpl_48;
  assign and_dcpl_74 = and_dcpl_72 & and_dcpl_52;
  assign and_dcpl_75 = and_dcpl_72 & and_dcpl_54;
  assign and_dcpl_76 = and_dcpl_72 & and_dcpl_11;
  assign and_dcpl_77 = and_dcpl_72 & and_dcpl_3;
  assign and_dcpl_78 = and_dcpl_72 & and_dcpl_41;
  assign and_dcpl_79 = and_dcpl_72 & and_dcpl_44;
  assign and_dcpl_80 = and_dcpl_72 & and_dcpl_46;
  assign and_dcpl_81 = (~ (fsm_output[2])) & (fsm_output[5]);
  assign and_dcpl_82 = and_dcpl_81 & and_dcpl_1;
  assign and_dcpl_83 = and_dcpl_7 & and_dcpl_82;
  assign and_dcpl_84 = and_dcpl_81 & and_dcpl_40;
  assign and_dcpl_85 = and_dcpl_7 & and_dcpl_84;
  assign and_dcpl_86 = and_dcpl_81 & and_dcpl_43;
  assign and_dcpl_87 = and_dcpl_7 & and_dcpl_86;
  assign and_dcpl_88 = and_dcpl_81 & and_463_cse;
  assign and_dcpl_89 = and_dcpl_7 & and_dcpl_88;
  assign and_dcpl_90 = (fsm_output[2]) & (fsm_output[5]);
  assign and_dcpl_91 = and_dcpl_90 & and_dcpl_1;
  assign and_dcpl_92 = and_dcpl_7 & and_dcpl_91;
  assign and_dcpl_93 = and_dcpl_90 & and_dcpl_40;
  assign and_dcpl_94 = and_dcpl_7 & and_dcpl_93;
  assign and_dcpl_95 = and_dcpl_90 & and_dcpl_43;
  assign and_dcpl_96 = and_dcpl_7 & and_dcpl_95;
  assign and_dcpl_97 = and_dcpl_90 & and_463_cse;
  assign and_dcpl_98 = and_dcpl_7 & and_dcpl_97;
  assign and_dcpl_99 = and_dcpl_50 & and_dcpl_82;
  assign and_dcpl_100 = and_dcpl_50 & and_dcpl_84;
  assign and_dcpl_101 = and_dcpl_50 & and_dcpl_86;
  assign and_dcpl_102 = and_dcpl_50 & and_dcpl_88;
  assign and_dcpl_103 = and_dcpl_50 & and_dcpl_91;
  assign and_dcpl_104 = and_dcpl_50 & and_dcpl_93;
  assign and_dcpl_105 = and_dcpl_50 & and_dcpl_95;
  assign and_dcpl_106 = and_dcpl_50 & and_dcpl_97;
  assign and_dcpl_107 = and_dcpl_62 & and_dcpl_82;
  assign and_dcpl_108 = and_dcpl_62 & and_dcpl_84;
  assign and_dcpl_109 = and_dcpl_62 & and_dcpl_86;
  assign and_dcpl_110 = and_dcpl_62 & and_dcpl_88;
  assign and_dcpl_111 = and_dcpl_62 & and_dcpl_91;
  assign and_dcpl_112 = and_dcpl_62 & and_dcpl_93;
  assign and_dcpl_113 = and_dcpl_62 & and_dcpl_95;
  assign and_dcpl_114 = and_dcpl_62 & and_dcpl_97;
  assign and_dcpl_115 = and_dcpl_72 & and_dcpl_82;
  assign and_dcpl_116 = and_dcpl_72 & and_dcpl_84;
  assign and_dcpl_117 = and_dcpl_72 & and_dcpl_86;
  assign and_dcpl_118 = and_dcpl_72 & and_dcpl_88;
  assign and_dcpl_119 = and_dcpl_72 & and_dcpl_91;
  assign and_dcpl_120 = and_dcpl_72 & and_dcpl_93;
  assign and_dcpl_121 = and_dcpl_72 & and_dcpl_95;
  assign and_dcpl_122 = and_dcpl_72 & and_dcpl_97;
  assign and_dcpl_123 = and_dcpl_5 & (fsm_output[6]);
  assign and_dcpl_124 = and_dcpl_123 & and_dcpl_4;
  assign and_dcpl_125 = and_dcpl_124 & and_dcpl_48;
  assign and_dcpl_126 = and_dcpl_124 & and_dcpl_52;
  assign and_dcpl_127 = and_dcpl_124 & and_dcpl_54;
  assign and_dcpl_128 = and_dcpl_124 & and_dcpl_11;
  assign and_dcpl_129 = and_dcpl_124 & and_dcpl_3;
  assign and_dcpl_130 = and_dcpl_124 & and_dcpl_41;
  assign and_dcpl_131 = and_dcpl_124 & and_dcpl_44;
  assign and_dcpl_132 = and_dcpl_124 & and_dcpl_46;
  assign and_dcpl_133 = and_dcpl_123 & and_dcpl_49;
  assign and_dcpl_134 = and_dcpl_133 & and_dcpl_48;
  assign and_dcpl_135 = and_dcpl_133 & and_dcpl_52;
  assign and_dcpl_136 = and_dcpl_133 & and_dcpl_54;
  assign and_dcpl_137 = and_dcpl_133 & and_dcpl_11;
  assign and_dcpl_138 = and_dcpl_133 & and_dcpl_3;
  assign and_dcpl_139 = and_dcpl_133 & and_dcpl_41;
  assign and_dcpl_140 = and_dcpl_133 & and_dcpl_44;
  assign and_dcpl_141 = and_dcpl_133 & and_dcpl_46;
  assign and_dcpl_142 = and_dcpl_123 & and_dcpl_61;
  assign and_dcpl_143 = and_dcpl_142 & and_dcpl_48;
  assign and_dcpl_144 = and_dcpl_142 & and_dcpl_52;
  assign and_dcpl_145 = and_dcpl_142 & and_dcpl_54;
  assign and_dcpl_146 = and_dcpl_142 & and_dcpl_11;
  assign and_dcpl_147 = and_dcpl_142 & and_dcpl_3;
  assign and_dcpl_148 = and_dcpl_142 & and_dcpl_41;
  assign and_dcpl_149 = and_dcpl_142 & and_dcpl_44;
  assign and_dcpl_150 = and_dcpl_142 & and_dcpl_46;
  assign and_dcpl_151 = and_dcpl_123 & and_cse;
  assign and_dcpl_152 = and_dcpl_151 & and_dcpl_48;
  assign and_dcpl_153 = and_dcpl_151 & and_dcpl_52;
  assign and_dcpl_154 = and_dcpl_151 & and_dcpl_54;
  assign and_dcpl_155 = and_dcpl_151 & and_dcpl_11;
  assign and_dcpl_156 = and_dcpl_151 & and_dcpl_3;
  assign and_dcpl_157 = and_dcpl_151 & and_dcpl_41;
  assign and_dcpl_158 = and_dcpl_151 & and_dcpl_44;
  assign and_dcpl_159 = and_dcpl_151 & and_dcpl_46;
  assign and_dcpl_160 = and_dcpl_124 & and_dcpl_82;
  assign and_dcpl_161 = and_dcpl_124 & and_dcpl_84;
  assign and_dcpl_162 = and_dcpl_124 & and_dcpl_86;
  assign and_dcpl_163 = and_dcpl_124 & and_dcpl_88;
  assign and_dcpl_164 = and_dcpl_124 & and_dcpl_91;
  assign and_dcpl_165 = and_dcpl_124 & and_dcpl_93;
  assign and_dcpl_166 = and_dcpl_124 & and_dcpl_95;
  assign and_dcpl_167 = and_dcpl_124 & and_dcpl_97;
  assign and_dcpl_168 = and_dcpl_133 & and_dcpl_82;
  assign and_dcpl_169 = and_dcpl_133 & and_dcpl_84;
  assign and_dcpl_170 = and_dcpl_133 & and_dcpl_86;
  assign and_dcpl_171 = and_dcpl_133 & and_dcpl_88;
  assign and_dcpl_172 = and_dcpl_133 & and_dcpl_91;
  assign and_dcpl_173 = and_dcpl_133 & and_dcpl_93;
  assign and_dcpl_174 = and_dcpl_133 & and_dcpl_95;
  assign and_dcpl_175 = and_dcpl_133 & and_dcpl_97;
  assign and_dcpl_176 = and_dcpl_142 & and_dcpl_82;
  assign and_dcpl_177 = and_dcpl_142 & and_dcpl_84;
  assign and_dcpl_178 = and_dcpl_142 & and_dcpl_86;
  assign and_dcpl_179 = and_dcpl_142 & and_dcpl_88;
  assign and_dcpl_180 = and_dcpl_142 & and_dcpl_91;
  assign and_dcpl_181 = and_dcpl_142 & and_dcpl_93;
  assign and_dcpl_182 = and_dcpl_142 & and_dcpl_95;
  assign and_dcpl_183 = and_dcpl_142 & and_dcpl_97;
  assign and_dcpl_184 = and_dcpl_151 & and_dcpl_82;
  assign and_dcpl_185 = and_dcpl_151 & and_dcpl_84;
  assign and_dcpl_186 = and_dcpl_151 & and_dcpl_86;
  assign and_dcpl_187 = and_dcpl_151 & and_dcpl_88;
  assign and_dcpl_188 = and_dcpl_151 & and_dcpl_91;
  assign and_dcpl_189 = and_dcpl_151 & and_dcpl_93;
  assign and_dcpl_190 = and_dcpl_151 & and_dcpl_95;
  assign and_dcpl_191 = and_dcpl_151 & and_dcpl_97;
  assign and_dcpl_192 = (fsm_output[8:7]==2'b01);
  assign and_dcpl_193 = and_dcpl_192 & (~ (fsm_output[6]));
  assign and_dcpl_194 = and_dcpl_193 & and_dcpl_4;
  assign and_dcpl_195 = and_dcpl_194 & and_dcpl_48;
  assign and_dcpl_196 = and_dcpl_194 & and_dcpl_52;
  assign and_dcpl_197 = and_dcpl_194 & and_dcpl_54;
  assign and_dcpl_198 = and_dcpl_194 & and_dcpl_11;
  assign and_dcpl_199 = and_dcpl_194 & and_dcpl_3;
  assign and_dcpl_200 = and_dcpl_194 & and_dcpl_41;
  assign and_dcpl_201 = and_dcpl_194 & and_dcpl_44;
  assign and_dcpl_202 = and_dcpl_194 & and_dcpl_46;
  assign and_dcpl_203 = and_dcpl_193 & and_dcpl_49;
  assign and_dcpl_204 = and_dcpl_203 & and_dcpl_48;
  assign and_dcpl_205 = and_dcpl_203 & and_dcpl_52;
  assign and_dcpl_206 = and_dcpl_203 & and_dcpl_54;
  assign and_dcpl_207 = and_dcpl_203 & and_dcpl_11;
  assign and_dcpl_208 = and_dcpl_203 & and_dcpl_3;
  assign and_dcpl_209 = and_dcpl_203 & and_dcpl_41;
  assign and_dcpl_210 = and_dcpl_203 & and_dcpl_44;
  assign and_dcpl_211 = and_dcpl_203 & and_dcpl_46;
  assign and_dcpl_212 = and_dcpl_193 & and_dcpl_61;
  assign and_dcpl_213 = and_dcpl_212 & and_dcpl_48;
  assign and_dcpl_214 = and_dcpl_212 & and_dcpl_52;
  assign and_dcpl_215 = and_dcpl_212 & and_dcpl_54;
  assign and_dcpl_216 = and_dcpl_212 & and_dcpl_11;
  assign and_dcpl_217 = and_dcpl_212 & and_dcpl_3;
  assign and_dcpl_218 = and_dcpl_212 & and_dcpl_41;
  assign and_dcpl_219 = and_dcpl_212 & and_dcpl_44;
  assign and_dcpl_220 = and_dcpl_212 & and_dcpl_46;
  assign and_dcpl_221 = and_dcpl_193 & and_cse;
  assign and_dcpl_222 = and_dcpl_221 & and_dcpl_48;
  assign and_dcpl_223 = and_dcpl_221 & and_dcpl_52;
  assign and_dcpl_224 = and_dcpl_221 & and_dcpl_54;
  assign and_dcpl_225 = and_dcpl_221 & and_dcpl_11;
  assign and_dcpl_226 = and_dcpl_221 & and_dcpl_3;
  assign and_dcpl_227 = and_dcpl_221 & and_dcpl_41;
  assign and_dcpl_228 = and_dcpl_221 & and_dcpl_44;
  assign and_dcpl_229 = and_dcpl_221 & and_dcpl_46;
  assign and_dcpl_230 = and_dcpl_194 & and_dcpl_82;
  assign and_dcpl_231 = and_dcpl_194 & and_dcpl_84;
  assign and_dcpl_232 = and_dcpl_194 & and_dcpl_86;
  assign and_dcpl_233 = and_dcpl_194 & and_dcpl_88;
  assign and_dcpl_234 = and_dcpl_194 & and_dcpl_91;
  assign and_dcpl_235 = and_dcpl_194 & and_dcpl_93;
  assign and_dcpl_236 = and_dcpl_194 & and_dcpl_95;
  assign and_dcpl_237 = and_dcpl_194 & and_dcpl_97;
  assign and_dcpl_238 = and_dcpl_203 & and_dcpl_82;
  assign and_dcpl_239 = and_dcpl_203 & and_dcpl_84;
  assign and_dcpl_240 = and_dcpl_203 & and_dcpl_86;
  assign and_dcpl_241 = and_dcpl_203 & and_dcpl_88;
  assign and_dcpl_242 = and_dcpl_203 & and_dcpl_91;
  assign and_dcpl_243 = and_dcpl_203 & and_dcpl_93;
  assign and_dcpl_244 = and_dcpl_203 & and_dcpl_95;
  assign and_dcpl_245 = and_dcpl_203 & and_dcpl_97;
  assign and_dcpl_246 = and_dcpl_212 & and_dcpl_82;
  assign and_dcpl_247 = and_dcpl_212 & and_dcpl_84;
  assign and_dcpl_248 = and_dcpl_212 & and_dcpl_86;
  assign and_dcpl_249 = and_dcpl_212 & and_dcpl_88;
  assign and_dcpl_250 = and_dcpl_212 & and_dcpl_91;
  assign and_dcpl_251 = and_dcpl_212 & and_dcpl_93;
  assign and_dcpl_252 = and_dcpl_212 & and_dcpl_95;
  assign and_dcpl_253 = and_dcpl_212 & and_dcpl_97;
  assign and_dcpl_254 = and_dcpl_221 & and_dcpl_82;
  assign and_dcpl_255 = and_dcpl_221 & and_dcpl_84;
  assign and_dcpl_256 = and_dcpl_221 & and_dcpl_86;
  assign and_dcpl_257 = and_dcpl_221 & and_dcpl_88;
  assign and_dcpl_258 = and_dcpl_221 & and_dcpl_91;
  assign and_dcpl_259 = and_dcpl_221 & and_dcpl_93;
  assign and_dcpl_260 = and_dcpl_221 & and_dcpl_95;
  assign and_dcpl_261 = and_dcpl_221 & and_dcpl_97;
  assign and_dcpl_262 = and_dcpl_192 & (fsm_output[6]);
  assign and_dcpl_263 = and_dcpl_262 & and_dcpl_4;
  assign and_dcpl_264 = and_dcpl_263 & and_dcpl_48;
  assign and_dcpl_265 = and_dcpl_263 & and_dcpl_52;
  assign and_dcpl_266 = and_dcpl_263 & and_dcpl_54;
  assign and_dcpl_267 = and_dcpl_263 & and_dcpl_11;
  assign and_dcpl_268 = and_dcpl_263 & and_dcpl_3;
  assign and_dcpl_269 = and_dcpl_263 & and_dcpl_41;
  assign and_dcpl_270 = and_dcpl_263 & and_dcpl_44;
  assign and_dcpl_271 = and_dcpl_263 & and_dcpl_46;
  assign and_dcpl_272 = and_dcpl_262 & and_dcpl_49;
  assign and_dcpl_273 = and_dcpl_272 & and_dcpl_48;
  assign and_dcpl_274 = and_dcpl_272 & and_dcpl_52;
  assign and_dcpl_275 = and_dcpl_272 & and_dcpl_54;
  assign and_dcpl_276 = and_dcpl_272 & and_dcpl_11;
  assign and_dcpl_277 = and_dcpl_272 & and_dcpl_3;
  assign and_dcpl_278 = and_dcpl_272 & and_dcpl_41;
  assign and_dcpl_279 = and_dcpl_272 & and_dcpl_44;
  assign and_dcpl_280 = and_dcpl_272 & and_dcpl_46;
  assign and_dcpl_281 = and_dcpl_262 & and_dcpl_61;
  assign and_dcpl_282 = and_dcpl_281 & and_dcpl_48;
  assign and_dcpl_283 = and_dcpl_281 & and_dcpl_52;
  assign and_dcpl_284 = and_dcpl_281 & and_dcpl_54;
  assign and_dcpl_285 = and_dcpl_281 & and_dcpl_11;
  assign and_dcpl_286 = and_dcpl_281 & and_dcpl_3;
  assign and_dcpl_287 = and_dcpl_281 & and_dcpl_41;
  assign and_dcpl_288 = and_dcpl_281 & and_dcpl_44;
  assign and_dcpl_289 = and_dcpl_281 & and_dcpl_46;
  assign and_dcpl_290 = and_dcpl_262 & and_cse;
  assign and_dcpl_291 = and_dcpl_290 & and_dcpl_48;
  assign and_dcpl_292 = and_dcpl_290 & and_dcpl_52;
  assign and_dcpl_293 = and_dcpl_290 & and_dcpl_54;
  assign and_dcpl_294 = and_dcpl_290 & and_dcpl_11;
  assign and_dcpl_295 = and_dcpl_290 & and_dcpl_3;
  assign and_dcpl_296 = and_dcpl_290 & and_dcpl_41;
  assign and_dcpl_297 = and_dcpl_290 & and_dcpl_44;
  assign and_dcpl_298 = and_dcpl_290 & and_dcpl_46;
  assign and_dcpl_299 = and_dcpl_263 & and_dcpl_82;
  assign and_dcpl_300 = and_dcpl_263 & and_dcpl_84;
  assign and_dcpl_301 = and_dcpl_263 & and_dcpl_86;
  assign and_dcpl_302 = and_dcpl_263 & and_dcpl_88;
  assign and_dcpl_303 = and_dcpl_263 & and_dcpl_91;
  assign and_dcpl_304 = and_dcpl_263 & and_dcpl_93;
  assign and_dcpl_305 = and_dcpl_263 & and_dcpl_95;
  assign and_dcpl_306 = and_dcpl_263 & and_dcpl_97;
  assign and_dcpl_307 = and_dcpl_272 & and_dcpl_82;
  assign and_dcpl_308 = and_dcpl_272 & and_dcpl_84;
  assign and_dcpl_309 = and_dcpl_272 & and_dcpl_86;
  assign and_dcpl_310 = and_dcpl_272 & and_dcpl_88;
  assign and_dcpl_311 = and_dcpl_272 & and_dcpl_91;
  assign and_dcpl_312 = and_dcpl_272 & and_dcpl_93;
  assign and_dcpl_313 = and_dcpl_272 & and_dcpl_95;
  assign and_dcpl_314 = and_dcpl_272 & and_dcpl_97;
  assign and_dcpl_315 = and_dcpl_281 & and_dcpl_82;
  assign and_dcpl_316 = and_dcpl_281 & and_dcpl_84;
  assign and_dcpl_317 = and_dcpl_281 & and_dcpl_86;
  assign and_dcpl_318 = and_dcpl_281 & and_dcpl_88;
  assign and_dcpl_319 = and_dcpl_281 & and_dcpl_91;
  assign and_dcpl_320 = and_dcpl_281 & and_dcpl_93;
  assign and_dcpl_321 = and_dcpl_281 & and_dcpl_95;
  assign and_dcpl_322 = and_dcpl_281 & and_dcpl_97;
  assign and_dcpl_323 = and_dcpl_290 & and_dcpl_82;
  assign and_dcpl_324 = and_dcpl_290 & and_dcpl_84;
  assign and_dcpl_325 = and_dcpl_290 & and_dcpl_86;
  assign and_dcpl_326 = and_dcpl_290 & and_dcpl_88;
  assign and_dcpl_327 = and_dcpl_290 & and_dcpl_91;
  assign and_dcpl_328 = and_dcpl_290 & and_dcpl_93;
  assign and_dcpl_329 = and_dcpl_290 & and_dcpl_95;
  assign and_dcpl_330 = and_dcpl_290 & and_dcpl_97;
  assign and_dcpl_333 = (fsm_output[8:6]==3'b100) & and_dcpl_4;
  assign and_dcpl_334 = and_dcpl_333 & and_dcpl_48;
  assign and_dcpl_335 = and_dcpl_333 & and_dcpl_52;
  assign and_dcpl_336 = and_dcpl_333 & and_dcpl_54;
  assign and_dcpl_341 = ~((fsm_output[8]) | (fsm_output[6]));
  assign or_tmp_126 = (fsm_output[3:2]!=2'b10);
  assign or_tmp_127 = (fsm_output[3:2]!=2'b01);
  assign or_tmp_129 = (fsm_output[7]) | (fsm_output[2]);
  assign or_tmp_130 = (fsm_output[7]) | (~ (fsm_output[2]));
  assign mux_tmp_91 = MUX_s_1_2_2(nand_94_cse, or_228_cse, fsm_output[3]);
  assign or_tmp_133 = (~ (fsm_output[7])) | (fsm_output[2]);
  assign mux_tmp_93 = MUX_s_1_2_2(or_tmp_133, or_tmp_130, fsm_output[6]);
  assign mux_tmp_103 = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[7]);
  assign nand_tmp_5 = ~((fsm_output[5]) & (~ mux_377_cse));
  assign nor_tmp_20 = (fsm_output[7]) & (fsm_output[3]);
  assign or_848_nl = (fsm_output[6]) | (fsm_output[3]);
  assign mux_tmp_118 = MUX_s_1_2_2(or_827_cse, (or_848_nl), fsm_output[7]);
  assign mux_tmp_153 = MUX_s_1_2_2(or_765_cse, or_743_cse, fsm_output[2]);
  assign nand_tmp_14 = ~((fsm_output[3]) & (~ mux_tmp_93));
  assign nor_tmp_41 = (fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]) & (fsm_output[2]);
  assign or_tmp_213 = (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[0]) | (fsm_output[4]);
  assign mux_tmp_205 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[0]);
  assign nand_17_nl = ~((fsm_output[2]) & (fsm_output[6]) & (~ mux_tmp_205));
  assign or_240_nl = (fsm_output[2]) | (fsm_output[6]) | mux_tmp_205;
  assign mux_tmp_206 = MUX_s_1_2_2((nand_17_nl), (or_240_nl), fsm_output[7]);
  assign or_tmp_219 = (fsm_output[2]) | (fsm_output[6]) | (~((fsm_output[0]) & (fsm_output[4])));
  assign or_tmp_225 = (~ (fsm_output[7])) | (fsm_output[3]);
  assign or_254_nl = (fsm_output[6]) | nand_100_cse;
  assign mux_tmp_217 = MUX_s_1_2_2((or_254_nl), or_765_cse, fsm_output[2]);
  assign or_tmp_239 = (~ (fsm_output[5])) | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[6]);
  assign nand_121_nl = ~((fsm_output[1]) & (fsm_output[5]) & (fsm_output[2]) & (~
      (fsm_output[8])) & (fsm_output[6]));
  assign or_264_nl = (fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[6]);
  assign mux_249_nl = MUX_s_1_2_2((or_264_nl), or_tmp_239, fsm_output[1]);
  assign mux_tmp_231 = MUX_s_1_2_2((nand_121_nl), (mux_249_nl), fsm_output[7]);
  assign or_270_nl = (fsm_output[8]) | (~ (fsm_output[6]));
  assign or_269_nl = (fsm_output[8]) | (fsm_output[6]);
  assign mux_tmp_232 = MUX_s_1_2_2((or_270_nl), (or_269_nl), fsm_output[2]);
  assign or_tmp_262 = (~ (fsm_output[7])) | (fsm_output[8]) | (fsm_output[3]);
  assign or_tmp_264 = (~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[3]));
  assign or_tmp_268 = (fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[6]) | (~
      (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[3]));
  assign or_tmp_270 = (~ (fsm_output[6])) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[3]);
  assign or_297_nl = (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[3]);
  assign mux_tmp_253 = MUX_s_1_2_2(or_tmp_270, (or_297_nl), fsm_output[2]);
  assign or_tmp_282 = (fsm_output[5]) | (~ (fsm_output[2])) | (fsm_output[6]) | nand_100_cse;
  assign or_tmp_292 = (fsm_output[7:6]!=2'b01);
  assign or_906_nl = (fsm_output[7:6]!=2'b10);
  assign mux_293_nl = MUX_s_1_2_2((or_906_nl), or_tmp_292, fsm_output[2]);
  assign or_318_nl = (fsm_output[1]) | (mux_293_nl);
  assign mux_292_nl = MUX_s_1_2_2(or_tmp_292, or_94_cse, fsm_output[2]);
  assign nand_24_nl = ~((fsm_output[1]) & (~ (mux_292_nl)));
  assign mux_tmp_275 = MUX_s_1_2_2((or_318_nl), (nand_24_nl), fsm_output[5]);
  assign or_322_cse = (fsm_output[6:2]!=5'b00000);
  assign and_472_nl = (fsm_output[8:7]==2'b11);
  assign mux_tmp_280 = MUX_s_1_2_2((and_472_nl), (fsm_output[8]), or_322_cse);
  assign mux_300_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[8]);
  assign mux_tmp_282 = MUX_s_1_2_2((mux_300_nl), (fsm_output[8]), or_322_cse);
  assign and_dcpl_360 = and_dcpl_10 & (fsm_output[1]);
  assign and_dcpl_362 = and_dcpl_7 & and_dcpl_360 & operator_32_false_acc_itm_31_1
      & (~ (fsm_output[0]));
  assign and_dcpl_376 = and_dcpl_6 & and_dcpl_4 & (~ (fsm_output[2]));
  assign or_dcpl_28 = or_dcpl_10 | (fsm_output[6]);
  assign or_dcpl_29 = or_dcpl_28 | or_52_cse;
  assign and_dcpl_388 = and_dcpl_34 & operator_32_false_acc_itm_31_1;
  assign and_dcpl_394 = ~((step_step_sva[1:0]!=2'b00));
  assign and_dcpl_395 = and_dcpl_394 & (~ (step_step_sva[2]));
  assign and_dcpl_397 = and_dcpl_32 & and_dcpl_27 & and_dcpl_395;
  assign and_dcpl_399 = and_463_cse & operator_16_false_slc_operator_16_false_acc_12_svs
      & (~ (step_step_sva[3]));
  assign and_dcpl_401 = and_dcpl_32 & and_dcpl_399 & and_dcpl_395;
  assign and_dcpl_405 = (step_step_sva[1:0]==2'b01);
  assign and_dcpl_406 = and_dcpl_405 & (~ (step_step_sva[2]));
  assign and_dcpl_408 = and_dcpl_32 & and_dcpl_27 & and_dcpl_406;
  assign and_dcpl_410 = and_dcpl_32 & and_dcpl_399 & and_dcpl_406;
  assign and_dcpl_411 = (step_step_sva[1:0]==2'b10);
  assign and_dcpl_412 = and_dcpl_411 & (~ (step_step_sva[2]));
  assign and_dcpl_414 = and_dcpl_32 & and_dcpl_27 & and_dcpl_412;
  assign and_dcpl_416 = and_dcpl_32 & and_dcpl_399 & and_dcpl_412;
  assign and_dcpl_417 = and_dcpl_24 & (~ (step_step_sva[2]));
  assign and_dcpl_419 = and_dcpl_32 & and_dcpl_27 & and_dcpl_417;
  assign and_dcpl_421 = and_dcpl_32 & and_dcpl_399 & and_dcpl_417;
  assign and_dcpl_422 = and_dcpl_394 & (step_step_sva[2]);
  assign and_dcpl_424 = and_dcpl_32 & and_dcpl_27 & and_dcpl_422;
  assign and_dcpl_426 = and_dcpl_32 & and_dcpl_399 & and_dcpl_422;
  assign and_dcpl_427 = and_dcpl_405 & (step_step_sva[2]);
  assign and_dcpl_429 = and_dcpl_32 & and_dcpl_27 & and_dcpl_427;
  assign and_dcpl_431 = and_dcpl_32 & and_dcpl_399 & and_dcpl_427;
  assign and_dcpl_432 = and_dcpl_411 & (step_step_sva[2]);
  assign and_dcpl_434 = and_dcpl_32 & and_dcpl_27 & and_dcpl_432;
  assign and_dcpl_436 = and_dcpl_32 & and_dcpl_399 & and_dcpl_432;
  assign and_dcpl_438 = and_dcpl_32 & and_dcpl_399 & and_dcpl_25;
  assign or_dcpl_31 = (fsm_output[1:0]!=2'b10);
  assign or_dcpl_32 = or_dcpl_14 | or_dcpl_31;
  assign or_dcpl_35 = (fsm_output[8:6]!=3'b100) | or_52_cse;
  assign or_dcpl_37 = (fsm_output[1:0]!=2'b01);
  assign or_dcpl_38 = or_dcpl_14 | or_dcpl_37;
  assign or_dcpl_40 = (fsm_output[1:0]!=2'b00);
  assign or_dcpl_41 = or_dcpl_14 | or_dcpl_40;
  assign or_dcpl_43 = ~((fsm_output[2]) & (fsm_output[5]));
  assign or_dcpl_44 = or_dcpl_43 | or_dcpl_4;
  assign or_dcpl_45 = ~((fsm_output[4:3]==2'b11));
  assign or_dcpl_46 = (fsm_output[8:7]!=2'b01);
  assign or_dcpl_47 = or_dcpl_46 | (~ (fsm_output[6]));
  assign or_dcpl_48 = or_dcpl_47 | or_dcpl_45;
  assign or_dcpl_50 = or_dcpl_43 | or_dcpl_31;
  assign or_dcpl_52 = or_dcpl_43 | or_dcpl_37;
  assign or_dcpl_54 = or_dcpl_43 | or_dcpl_40;
  assign or_dcpl_56 = (fsm_output[2]) | (~ (fsm_output[5]));
  assign or_dcpl_57 = or_dcpl_56 | or_dcpl_4;
  assign or_dcpl_59 = or_dcpl_56 | or_dcpl_31;
  assign or_dcpl_61 = or_dcpl_56 | or_dcpl_37;
  assign or_dcpl_63 = or_dcpl_56 | or_dcpl_40;
  assign or_dcpl_65 = (fsm_output[4:3]!=2'b10);
  assign or_dcpl_66 = or_dcpl_47 | or_dcpl_65;
  assign or_dcpl_75 = (fsm_output[4:3]!=2'b01);
  assign or_dcpl_76 = or_dcpl_47 | or_dcpl_75;
  assign or_dcpl_85 = or_dcpl_47 | or_52_cse;
  assign or_dcpl_94 = (~ (fsm_output[2])) | (fsm_output[5]);
  assign or_dcpl_95 = or_dcpl_94 | or_dcpl_4;
  assign or_dcpl_97 = or_dcpl_94 | or_dcpl_31;
  assign or_dcpl_99 = or_dcpl_94 | or_dcpl_37;
  assign or_dcpl_101 = or_dcpl_94 | or_dcpl_40;
  assign or_dcpl_103 = or_dcpl_14 | or_dcpl_4;
  assign or_dcpl_132 = or_dcpl_46 | (fsm_output[6]);
  assign or_dcpl_133 = or_dcpl_132 | or_dcpl_45;
  assign or_dcpl_142 = or_dcpl_132 | or_dcpl_65;
  assign or_dcpl_151 = or_dcpl_132 | or_dcpl_75;
  assign or_dcpl_159 = or_dcpl_132 | or_52_cse;
  assign or_dcpl_200 = or_dcpl_10 | (~ (fsm_output[6]));
  assign or_dcpl_201 = or_dcpl_200 | or_dcpl_45;
  assign or_dcpl_210 = or_dcpl_200 | or_dcpl_65;
  assign or_dcpl_219 = or_dcpl_200 | or_dcpl_75;
  assign or_dcpl_228 = or_dcpl_200 | or_52_cse;
  assign or_dcpl_269 = or_dcpl_28 | or_dcpl_45;
  assign or_dcpl_278 = or_dcpl_28 | or_dcpl_65;
  assign or_dcpl_287 = or_dcpl_28 | or_dcpl_75;
  assign and_dcpl_445 = and_dcpl_341 & (fsm_output[5:4]==2'b00);
  assign mux_355_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[2]);
  assign mux_tmp_337 = MUX_s_1_2_2((mux_355_nl), or_tmp_127, fsm_output[1]);
  assign mux_tmp_345 = MUX_s_1_2_2(mux_tmp_282, mux_tmp_280, fsm_output[1]);
  assign psum_reg_15_16_lpi_2_mx0c2 = and_dcpl_333 & and_dcpl_11;
  assign ROW_asn_142_itm_mx0c0 = and_dcpl_31 & and_dcpl_29 & and_dcpl_34;
  assign nl_operator_32_false_acc_1_nl = conv_u2u_32_33(~ step_mul_itm) + conv_u2u_16_33(step_step_sva);
  assign operator_32_false_acc_1_nl = nl_operator_32_false_acc_1_nl[32:0];
  assign nl_operator_32_false_acc_nl = (readslicef_33_32_1((operator_32_false_acc_1_nl)))
      + 32'b01111111111111111111111111110001;
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[31:0];
  assign operator_32_false_acc_itm_31_1 = readslicef_32_1_31((operator_32_false_acc_nl));
  assign accumulation_buffer_rsc_0_0_i_web_d = accumulation_buffer_rsc_0_0_i_web_d_reg;
  assign accumulation_buffer_rsc_0_0_i_addr_d = accumulation_buffer_rsc_0_0_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_din_d = step_output_buf_value_0_sva;
  assign accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_1_i_web_d = accumulation_buffer_rsc_0_1_i_web_d_reg;
  assign accumulation_buffer_rsc_0_1_i_addr_d = accumulation_buffer_rsc_0_1_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_din_d = psum_reg_16_8_lpi_2;
  assign accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_2_i_web_d = accumulation_buffer_rsc_0_2_i_web_d_reg;
  assign accumulation_buffer_rsc_0_2_i_addr_d = accumulation_buffer_rsc_0_2_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_din_d = psum_reg_15_16_lpi_2;
  assign accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_3_i_web_d = accumulation_buffer_rsc_0_3_i_web_d_reg;
  assign accumulation_buffer_rsc_0_3_i_addr_d = accumulation_buffer_rsc_0_3_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_din_d = psum_reg_16_15_lpi_2;
  assign accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_4_i_web_d = accumulation_buffer_rsc_0_4_i_web_d_reg;
  assign accumulation_buffer_rsc_0_4_i_addr_d = accumulation_buffer_rsc_0_4_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_din_d = psum_reg_16_16_lpi_2;
  assign accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_5_i_web_d = accumulation_buffer_rsc_0_5_i_web_d_reg;
  assign accumulation_buffer_rsc_0_5_i_addr_d = accumulation_buffer_rsc_0_5_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_din_d = psum_reg_16_2_lpi_2;
  assign accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_6_i_web_d = accumulation_buffer_rsc_0_6_i_web_d_reg;
  assign accumulation_buffer_rsc_0_6_i_addr_d = accumulation_buffer_rsc_0_6_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_din_d = psum_reg_16_3_lpi_2;
  assign accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_7_i_web_d = accumulation_buffer_rsc_0_7_i_web_d_reg;
  assign accumulation_buffer_rsc_0_7_i_addr_d = accumulation_buffer_rsc_0_7_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_din_d = psum_reg_16_4_lpi_2;
  assign accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_8_i_web_d = accumulation_buffer_rsc_0_8_i_web_d_reg;
  assign accumulation_buffer_rsc_0_8_i_addr_d = accumulation_buffer_rsc_0_8_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_din_d = psum_reg_16_5_lpi_2;
  assign accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_9_i_web_d = accumulation_buffer_rsc_0_9_i_web_d_reg;
  assign accumulation_buffer_rsc_0_9_i_addr_d = accumulation_buffer_rsc_0_9_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_din_d = psum_reg_16_6_lpi_2;
  assign accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_10_i_web_d = accumulation_buffer_rsc_0_10_i_web_d_reg;
  assign accumulation_buffer_rsc_0_10_i_addr_d = accumulation_buffer_rsc_0_10_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_din_d = psum_reg_16_7_lpi_2;
  assign accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_11_i_web_d = accumulation_buffer_rsc_0_11_i_web_d_reg;
  assign accumulation_buffer_rsc_0_11_i_addr_d = accumulation_buffer_rsc_0_11_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_din_d = psum_reg_16_1_lpi_2;
  assign accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_12_i_web_d = accumulation_buffer_rsc_0_12_i_web_d_reg;
  assign accumulation_buffer_rsc_0_12_i_addr_d = accumulation_buffer_rsc_0_12_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_din_d = psum_reg_16_10_lpi_2;
  assign accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_13_i_web_d = accumulation_buffer_rsc_0_13_i_web_d_reg;
  assign accumulation_buffer_rsc_0_13_i_addr_d = accumulation_buffer_rsc_0_13_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_din_d = psum_reg_16_11_lpi_2;
  assign accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_14_i_web_d = accumulation_buffer_rsc_0_14_i_web_d_reg;
  assign accumulation_buffer_rsc_0_14_i_addr_d = accumulation_buffer_rsc_0_14_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_din_d = psum_reg_16_12_lpi_2;
  assign accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_15_i_web_d = accumulation_buffer_rsc_0_15_i_web_d_reg;
  assign accumulation_buffer_rsc_0_15_i_addr_d = accumulation_buffer_rsc_0_15_i_addr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_din_d = psum_reg_16_14_lpi_2;
  assign accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d = accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  assign accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d = accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_rsci_idat_15_0 <= 16'b0000000000000000;
      output_rsci_idat_31_16 <= 16'b0000000000000000;
      output_rsci_idat_47_32 <= 16'b0000000000000000;
      output_rsci_idat_63_48 <= 16'b0000000000000000;
      output_rsci_idat_79_64 <= 16'b0000000000000000;
      output_rsci_idat_95_80 <= 16'b0000000000000000;
      output_rsci_idat_111_96 <= 16'b0000000000000000;
      output_rsci_idat_127_112 <= 16'b0000000000000000;
      output_rsci_idat_143_128 <= 16'b0000000000000000;
      output_rsci_idat_159_144 <= 16'b0000000000000000;
      output_rsci_idat_175_160 <= 16'b0000000000000000;
      output_rsci_idat_191_176 <= 16'b0000000000000000;
      output_rsci_idat_207_192 <= 16'b0000000000000000;
      output_rsci_idat_223_208 <= 16'b0000000000000000;
      output_rsci_idat_239_224 <= 16'b0000000000000000;
      output_rsci_idat_255_240 <= 16'b0000000000000000;
    end
    else if ( output_and_cse ) begin
      output_rsci_idat_15_0 <= output_fifo_0_rsci_output_rsc_z;
      output_rsci_idat_31_16 <= output_fifo_1_rsci_output_rsc_z;
      output_rsci_idat_47_32 <= output_fifo_2_rsci_output_rsc_z;
      output_rsci_idat_63_48 <= output_fifo_3_rsci_output_rsc_z;
      output_rsci_idat_79_64 <= output_fifo_4_rsci_output_rsc_z;
      output_rsci_idat_95_80 <= output_fifo_5_rsci_output_rsc_z;
      output_rsci_idat_111_96 <= output_fifo_6_rsci_output_rsc_z;
      output_rsci_idat_127_112 <= output_fifo_7_rsci_output_rsc_z;
      output_rsci_idat_143_128 <= output_fifo_8_rsci_output_rsc_z;
      output_rsci_idat_159_144 <= output_fifo_9_rsci_output_rsc_z;
      output_rsci_idat_175_160 <= output_fifo_10_rsci_output_rsc_z;
      output_rsci_idat_191_176 <= output_fifo_11_rsci_output_rsc_z;
      output_rsci_idat_207_192 <= output_fifo_12_rsci_output_rsc_z;
      output_rsci_idat_223_208 <= output_fifo_13_rsci_output_rsc_z;
      output_rsci_idat_239_224 <= output_fifo_14_rsci_output_rsc_z;
      output_rsci_idat_255_240 <= psum_reg_16_14_lpi_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ensig_cgo_47_cse <= 1'b0;
      reg_ensig_cgo_46_cse <= 1'b0;
      reg_ensig_cgo_45_cse <= 1'b0;
      reg_ensig_cgo_29_cse <= 1'b0;
      reg_ensig_cgo_28_cse <= 1'b0;
      reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse <= 1'b0;
      reg_loopIndicesIn_rsci_irdy_run_psct_cse <= 1'b0;
      reg_output_rsci_ivld_run_psct_cse <= 1'b0;
      reg_weight_rsci_irdy_run_psct_cse <= 1'b0;
      reg_input_rsci_irdy_run_psct_cse <= 1'b0;
      psum_reg_16_16_lpi_2 <= 16'b0000000000000000;
      weight_reg_8_15_lpi_2 <= 8'b00000000;
      weight_reg_8_14_lpi_2 <= 8'b00000000;
      weight_reg_8_13_lpi_2 <= 8'b00000000;
      weight_reg_8_12_lpi_2 <= 8'b00000000;
      weight_reg_8_11_lpi_2 <= 8'b00000000;
      weight_reg_8_10_lpi_2 <= 8'b00000000;
      weight_reg_8_9_lpi_2 <= 8'b00000000;
      weight_reg_8_8_lpi_2 <= 8'b00000000;
      weight_reg_8_7_lpi_2 <= 8'b00000000;
      weight_reg_8_6_lpi_2 <= 8'b00000000;
      weight_reg_8_5_lpi_2 <= 8'b00000000;
      weight_reg_8_4_lpi_2 <= 8'b00000000;
      weight_reg_8_3_lpi_2 <= 8'b00000000;
      weight_reg_8_2_lpi_2 <= 8'b00000000;
      weight_reg_8_1_lpi_2 <= 8'b00000000;
      weight_reg_8_0_lpi_2 <= 8'b00000000;
      weight_reg_0_15_lpi_2 <= 8'b00000000;
      weight_reg_0_14_lpi_2 <= 8'b00000000;
      weight_reg_0_13_lpi_2 <= 8'b00000000;
      weight_reg_0_12_lpi_2 <= 8'b00000000;
      weight_reg_0_11_lpi_2 <= 8'b00000000;
      weight_reg_0_10_lpi_2 <= 8'b00000000;
      weight_reg_0_9_lpi_2 <= 8'b00000000;
      weight_reg_0_8_lpi_2 <= 8'b00000000;
      weight_reg_0_7_lpi_2 <= 8'b00000000;
      weight_reg_0_6_lpi_2 <= 8'b00000000;
      weight_reg_0_5_lpi_2 <= 8'b00000000;
      weight_reg_0_4_lpi_2 <= 8'b00000000;
      weight_reg_0_3_lpi_2 <= 8'b00000000;
      weight_reg_0_2_lpi_2 <= 8'b00000000;
      weight_reg_0_1_lpi_2 <= 8'b00000000;
      weight_reg_0_0_lpi_2 <= 8'b00000000;
      weight_reg_9_15_lpi_2 <= 8'b00000000;
      weight_reg_9_14_lpi_2 <= 8'b00000000;
      weight_reg_9_13_lpi_2 <= 8'b00000000;
      weight_reg_9_12_lpi_2 <= 8'b00000000;
      weight_reg_9_11_lpi_2 <= 8'b00000000;
      weight_reg_9_10_lpi_2 <= 8'b00000000;
      weight_reg_9_9_lpi_2 <= 8'b00000000;
      weight_reg_9_8_lpi_2 <= 8'b00000000;
      weight_reg_9_7_lpi_2 <= 8'b00000000;
      weight_reg_9_6_lpi_2 <= 8'b00000000;
      weight_reg_9_5_lpi_2 <= 8'b00000000;
      weight_reg_9_4_lpi_2 <= 8'b00000000;
      weight_reg_9_3_lpi_2 <= 8'b00000000;
      weight_reg_9_2_lpi_2 <= 8'b00000000;
      weight_reg_9_1_lpi_2 <= 8'b00000000;
      weight_reg_9_0_lpi_2 <= 8'b00000000;
      weight_reg_1_15_lpi_2 <= 8'b00000000;
      weight_reg_1_14_lpi_2 <= 8'b00000000;
      weight_reg_1_13_lpi_2 <= 8'b00000000;
      weight_reg_1_12_lpi_2 <= 8'b00000000;
      weight_reg_1_11_lpi_2 <= 8'b00000000;
      weight_reg_1_10_lpi_2 <= 8'b00000000;
      weight_reg_1_9_lpi_2 <= 8'b00000000;
      weight_reg_1_8_lpi_2 <= 8'b00000000;
      weight_reg_1_7_lpi_2 <= 8'b00000000;
      weight_reg_1_6_lpi_2 <= 8'b00000000;
      weight_reg_1_5_lpi_2 <= 8'b00000000;
      weight_reg_1_4_lpi_2 <= 8'b00000000;
      weight_reg_1_3_lpi_2 <= 8'b00000000;
      weight_reg_1_2_lpi_2 <= 8'b00000000;
      weight_reg_1_1_lpi_2 <= 8'b00000000;
      weight_reg_1_0_lpi_2 <= 8'b00000000;
      weight_reg_10_15_lpi_2 <= 8'b00000000;
      weight_reg_10_14_lpi_2 <= 8'b00000000;
      weight_reg_10_13_lpi_2 <= 8'b00000000;
      weight_reg_10_12_lpi_2 <= 8'b00000000;
      weight_reg_10_11_lpi_2 <= 8'b00000000;
      weight_reg_10_10_lpi_2 <= 8'b00000000;
      weight_reg_10_9_lpi_2 <= 8'b00000000;
      weight_reg_10_8_lpi_2 <= 8'b00000000;
      weight_reg_10_7_lpi_2 <= 8'b00000000;
      weight_reg_10_6_lpi_2 <= 8'b00000000;
      weight_reg_10_5_lpi_2 <= 8'b00000000;
      weight_reg_10_4_lpi_2 <= 8'b00000000;
      weight_reg_10_3_lpi_2 <= 8'b00000000;
      weight_reg_10_2_lpi_2 <= 8'b00000000;
      weight_reg_10_1_lpi_2 <= 8'b00000000;
      weight_reg_10_0_lpi_2 <= 8'b00000000;
      weight_reg_2_15_lpi_2 <= 8'b00000000;
      weight_reg_2_14_lpi_2 <= 8'b00000000;
      weight_reg_2_13_lpi_2 <= 8'b00000000;
      weight_reg_2_12_lpi_2 <= 8'b00000000;
      weight_reg_2_11_lpi_2 <= 8'b00000000;
      weight_reg_2_10_lpi_2 <= 8'b00000000;
      weight_reg_2_9_lpi_2 <= 8'b00000000;
      weight_reg_2_8_lpi_2 <= 8'b00000000;
      weight_reg_2_7_lpi_2 <= 8'b00000000;
      weight_reg_2_6_lpi_2 <= 8'b00000000;
      weight_reg_2_5_lpi_2 <= 8'b00000000;
      weight_reg_2_4_lpi_2 <= 8'b00000000;
      weight_reg_2_3_lpi_2 <= 8'b00000000;
      weight_reg_2_2_lpi_2 <= 8'b00000000;
      weight_reg_2_1_lpi_2 <= 8'b00000000;
      weight_reg_2_0_lpi_2 <= 8'b00000000;
      weight_reg_11_15_lpi_2 <= 8'b00000000;
      weight_reg_11_14_lpi_2 <= 8'b00000000;
      weight_reg_11_13_lpi_2 <= 8'b00000000;
      weight_reg_11_12_lpi_2 <= 8'b00000000;
      weight_reg_11_11_lpi_2 <= 8'b00000000;
      weight_reg_11_10_lpi_2 <= 8'b00000000;
      weight_reg_11_9_lpi_2 <= 8'b00000000;
      weight_reg_11_8_lpi_2 <= 8'b00000000;
      weight_reg_11_7_lpi_2 <= 8'b00000000;
      weight_reg_11_6_lpi_2 <= 8'b00000000;
      weight_reg_11_5_lpi_2 <= 8'b00000000;
      weight_reg_11_4_lpi_2 <= 8'b00000000;
      weight_reg_11_3_lpi_2 <= 8'b00000000;
      weight_reg_11_2_lpi_2 <= 8'b00000000;
      weight_reg_11_1_lpi_2 <= 8'b00000000;
      weight_reg_11_0_lpi_2 <= 8'b00000000;
      weight_reg_3_15_lpi_2 <= 8'b00000000;
      weight_reg_3_14_lpi_2 <= 8'b00000000;
      weight_reg_3_13_lpi_2 <= 8'b00000000;
      weight_reg_3_12_lpi_2 <= 8'b00000000;
      weight_reg_3_11_lpi_2 <= 8'b00000000;
      weight_reg_3_10_lpi_2 <= 8'b00000000;
      weight_reg_3_9_lpi_2 <= 8'b00000000;
      weight_reg_3_8_lpi_2 <= 8'b00000000;
      weight_reg_3_7_lpi_2 <= 8'b00000000;
      weight_reg_3_6_lpi_2 <= 8'b00000000;
      weight_reg_3_5_lpi_2 <= 8'b00000000;
      weight_reg_3_4_lpi_2 <= 8'b00000000;
      weight_reg_3_3_lpi_2 <= 8'b00000000;
      weight_reg_3_2_lpi_2 <= 8'b00000000;
      weight_reg_3_1_lpi_2 <= 8'b00000000;
      weight_reg_3_0_lpi_2 <= 8'b00000000;
      weight_reg_12_15_lpi_2 <= 8'b00000000;
      weight_reg_12_14_lpi_2 <= 8'b00000000;
      weight_reg_12_13_lpi_2 <= 8'b00000000;
      weight_reg_12_12_lpi_2 <= 8'b00000000;
      weight_reg_12_11_lpi_2 <= 8'b00000000;
      weight_reg_12_10_lpi_2 <= 8'b00000000;
      weight_reg_12_9_lpi_2 <= 8'b00000000;
      weight_reg_12_8_lpi_2 <= 8'b00000000;
      weight_reg_12_7_lpi_2 <= 8'b00000000;
      weight_reg_12_6_lpi_2 <= 8'b00000000;
      weight_reg_12_5_lpi_2 <= 8'b00000000;
      weight_reg_12_4_lpi_2 <= 8'b00000000;
      weight_reg_12_3_lpi_2 <= 8'b00000000;
      weight_reg_12_2_lpi_2 <= 8'b00000000;
      weight_reg_12_1_lpi_2 <= 8'b00000000;
      weight_reg_12_0_lpi_2 <= 8'b00000000;
      weight_reg_4_15_lpi_2 <= 8'b00000000;
      weight_reg_4_14_lpi_2 <= 8'b00000000;
      weight_reg_4_13_lpi_2 <= 8'b00000000;
      weight_reg_4_12_lpi_2 <= 8'b00000000;
      weight_reg_4_11_lpi_2 <= 8'b00000000;
      weight_reg_4_10_lpi_2 <= 8'b00000000;
      weight_reg_4_9_lpi_2 <= 8'b00000000;
      weight_reg_4_8_lpi_2 <= 8'b00000000;
      weight_reg_4_7_lpi_2 <= 8'b00000000;
      weight_reg_4_6_lpi_2 <= 8'b00000000;
      weight_reg_4_5_lpi_2 <= 8'b00000000;
      weight_reg_4_4_lpi_2 <= 8'b00000000;
      weight_reg_4_3_lpi_2 <= 8'b00000000;
      weight_reg_4_2_lpi_2 <= 8'b00000000;
      weight_reg_4_1_lpi_2 <= 8'b00000000;
      weight_reg_4_0_lpi_2 <= 8'b00000000;
      weight_reg_13_15_lpi_2 <= 8'b00000000;
      weight_reg_13_14_lpi_2 <= 8'b00000000;
      weight_reg_13_13_lpi_2 <= 8'b00000000;
      weight_reg_13_12_lpi_2 <= 8'b00000000;
      weight_reg_13_11_lpi_2 <= 8'b00000000;
      weight_reg_13_10_lpi_2 <= 8'b00000000;
      weight_reg_13_9_lpi_2 <= 8'b00000000;
      weight_reg_13_8_lpi_2 <= 8'b00000000;
      weight_reg_13_7_lpi_2 <= 8'b00000000;
      weight_reg_13_6_lpi_2 <= 8'b00000000;
      weight_reg_13_5_lpi_2 <= 8'b00000000;
      weight_reg_13_4_lpi_2 <= 8'b00000000;
      weight_reg_13_3_lpi_2 <= 8'b00000000;
      weight_reg_13_2_lpi_2 <= 8'b00000000;
      weight_reg_13_1_lpi_2 <= 8'b00000000;
      weight_reg_13_0_lpi_2 <= 8'b00000000;
      weight_reg_5_15_lpi_2 <= 8'b00000000;
      weight_reg_5_14_lpi_2 <= 8'b00000000;
      weight_reg_5_13_lpi_2 <= 8'b00000000;
      weight_reg_5_12_lpi_2 <= 8'b00000000;
      weight_reg_5_11_lpi_2 <= 8'b00000000;
      weight_reg_5_10_lpi_2 <= 8'b00000000;
      weight_reg_5_9_lpi_2 <= 8'b00000000;
      weight_reg_5_8_lpi_2 <= 8'b00000000;
      weight_reg_5_7_lpi_2 <= 8'b00000000;
      weight_reg_5_6_lpi_2 <= 8'b00000000;
      weight_reg_5_5_lpi_2 <= 8'b00000000;
      weight_reg_5_4_lpi_2 <= 8'b00000000;
      weight_reg_5_3_lpi_2 <= 8'b00000000;
      weight_reg_5_2_lpi_2 <= 8'b00000000;
      weight_reg_5_1_lpi_2 <= 8'b00000000;
      weight_reg_5_0_lpi_2 <= 8'b00000000;
      weight_reg_14_15_lpi_2 <= 8'b00000000;
      weight_reg_14_14_lpi_2 <= 8'b00000000;
      weight_reg_14_13_lpi_2 <= 8'b00000000;
      weight_reg_14_12_lpi_2 <= 8'b00000000;
      weight_reg_14_11_lpi_2 <= 8'b00000000;
      weight_reg_14_10_lpi_2 <= 8'b00000000;
      weight_reg_14_9_lpi_2 <= 8'b00000000;
      weight_reg_14_8_lpi_2 <= 8'b00000000;
      weight_reg_14_7_lpi_2 <= 8'b00000000;
      weight_reg_14_6_lpi_2 <= 8'b00000000;
      weight_reg_14_5_lpi_2 <= 8'b00000000;
      weight_reg_14_4_lpi_2 <= 8'b00000000;
      weight_reg_14_3_lpi_2 <= 8'b00000000;
      weight_reg_14_2_lpi_2 <= 8'b00000000;
      weight_reg_14_1_lpi_2 <= 8'b00000000;
      weight_reg_14_0_lpi_2 <= 8'b00000000;
      weight_reg_6_15_lpi_2 <= 8'b00000000;
      weight_reg_6_14_lpi_2 <= 8'b00000000;
      weight_reg_6_13_lpi_2 <= 8'b00000000;
      weight_reg_6_12_lpi_2 <= 8'b00000000;
      weight_reg_6_11_lpi_2 <= 8'b00000000;
      weight_reg_6_10_lpi_2 <= 8'b00000000;
      weight_reg_6_9_lpi_2 <= 8'b00000000;
      weight_reg_6_8_lpi_2 <= 8'b00000000;
      weight_reg_6_7_lpi_2 <= 8'b00000000;
      weight_reg_6_6_lpi_2 <= 8'b00000000;
      weight_reg_6_5_lpi_2 <= 8'b00000000;
      weight_reg_6_4_lpi_2 <= 8'b00000000;
      weight_reg_6_3_lpi_2 <= 8'b00000000;
      weight_reg_6_2_lpi_2 <= 8'b00000000;
      weight_reg_6_1_lpi_2 <= 8'b00000000;
      weight_reg_6_0_lpi_2 <= 8'b00000000;
      weight_reg_15_15_lpi_2 <= 8'b00000000;
      weight_reg_15_14_lpi_2 <= 8'b00000000;
      weight_reg_15_13_lpi_2 <= 8'b00000000;
      weight_reg_15_12_lpi_2 <= 8'b00000000;
      weight_reg_15_11_lpi_2 <= 8'b00000000;
      weight_reg_15_10_lpi_2 <= 8'b00000000;
      weight_reg_15_9_lpi_2 <= 8'b00000000;
      weight_reg_15_8_lpi_2 <= 8'b00000000;
      weight_reg_15_7_lpi_2 <= 8'b00000000;
      weight_reg_15_6_lpi_2 <= 8'b00000000;
      weight_reg_15_5_lpi_2 <= 8'b00000000;
      weight_reg_15_4_lpi_2 <= 8'b00000000;
      weight_reg_15_3_lpi_2 <= 8'b00000000;
      weight_reg_15_2_lpi_2 <= 8'b00000000;
      weight_reg_15_1_lpi_2 <= 8'b00000000;
      weight_reg_15_0_lpi_2 <= 8'b00000000;
      weight_reg_7_15_lpi_2 <= 8'b00000000;
      weight_reg_7_14_lpi_2 <= 8'b00000000;
      weight_reg_7_13_lpi_2 <= 8'b00000000;
      weight_reg_7_12_lpi_2 <= 8'b00000000;
      weight_reg_7_11_lpi_2 <= 8'b00000000;
      weight_reg_7_10_lpi_2 <= 8'b00000000;
      weight_reg_7_9_lpi_2 <= 8'b00000000;
      weight_reg_7_8_lpi_2 <= 8'b00000000;
      weight_reg_7_7_lpi_2 <= 8'b00000000;
      weight_reg_7_6_lpi_2 <= 8'b00000000;
      weight_reg_7_5_lpi_2 <= 8'b00000000;
      weight_reg_7_4_lpi_2 <= 8'b00000000;
      weight_reg_7_3_lpi_2 <= 8'b00000000;
      weight_reg_7_2_lpi_2 <= 8'b00000000;
      weight_reg_7_1_lpi_2 <= 8'b00000000;
      weight_reg_7_0_lpi_2 <= 8'b00000000;
      step_in_col_value_lpi_2 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      psum_reg_16_15_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_14_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_12_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_11_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_10_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_9_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_8_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_7_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_6_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_5_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_4_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_3_lpi_2 <= 16'b0000000000000000;
      psum_reg_16_2_lpi_2 <= 16'b0000000000000000;
      step_output_buf_value_0_sva <= 16'b0000000000000000;
      step_step_sva <= 16'b0000000000000000;
      paramsIn_crt_sva_127_32 <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      loopIndicesIn_crt_sva <= 48'b000000000000000000000000000000000000000000000000;
      operator_16_false_slc_operator_16_false_acc_12_svs <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_ensig_cgo_47_cse <= and_17_rmff;
      reg_ensig_cgo_46_cse <= and_23_rmff;
      reg_ensig_cgo_45_cse <= ~ mux_302_itm;
      reg_ensig_cgo_29_cse <= and_364_rmff;
      reg_ensig_cgo_28_cse <= and_368_rmff;
      reg_accumulation_buffer_rsc_0_15_i_addr_d_run_psct_cse <= and_380_rmff;
      reg_loopIndicesIn_rsci_irdy_run_psct_cse <= ~(or_dcpl_29 | ((fsm_output[1])
          & operator_32_false_acc_itm_31_1) | (fsm_output[2]) | (fsm_output[5]) |
          (fsm_output[0]));
      reg_output_rsci_ivld_run_psct_cse <= and_dcpl_32 & and_463_cse & (~ operator_16_false_slc_operator_16_false_acc_16_itm)
          & step_if_3_step_if_3_if_step_if_3_if_nor_tmp & step_if_3_aif_step_if_3_aelse_step_if_3_aelse_nor_tmp
          & step_if_3_aif_1_step_if_3_aelse_1_step_if_3_aelse_1_nor_tmp;
      reg_weight_rsci_irdy_run_psct_cse <= and_dcpl_376 & and_dcpl_388 & (~ (fsm_output[0]))
          & operator_16_false_acc_itm_12_1;
      reg_input_rsci_irdy_run_psct_cse <= and_dcpl_376 & and_dcpl_388 & (~ (fsm_output[0]))
          & step_if_1_acc_itm_32_1;
      psum_reg_16_16_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_16_lpi_2, output_fifo_4_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_307_nl)) , and_dcpl_12 , and_dcpl_8});
      weight_reg_8_15_lpi_2 <= MUX_v_8_2_2(weight_reg_8_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_397);
      weight_reg_8_14_lpi_2 <= MUX_v_8_2_2(weight_reg_8_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_397);
      weight_reg_8_13_lpi_2 <= MUX_v_8_2_2(weight_reg_8_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_397);
      weight_reg_8_12_lpi_2 <= MUX_v_8_2_2(weight_reg_8_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_397);
      weight_reg_8_11_lpi_2 <= MUX_v_8_2_2(weight_reg_8_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_397);
      weight_reg_8_10_lpi_2 <= MUX_v_8_2_2(weight_reg_8_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_397);
      weight_reg_8_9_lpi_2 <= MUX_v_8_2_2(weight_reg_8_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_397);
      weight_reg_8_8_lpi_2 <= MUX_v_8_2_2(weight_reg_8_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_397);
      weight_reg_8_7_lpi_2 <= MUX_v_8_2_2(weight_reg_8_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_397);
      weight_reg_8_6_lpi_2 <= MUX_v_8_2_2(weight_reg_8_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_397);
      weight_reg_8_5_lpi_2 <= MUX_v_8_2_2(weight_reg_8_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_397);
      weight_reg_8_4_lpi_2 <= MUX_v_8_2_2(weight_reg_8_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_397);
      weight_reg_8_3_lpi_2 <= MUX_v_8_2_2(weight_reg_8_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_397);
      weight_reg_8_2_lpi_2 <= MUX_v_8_2_2(weight_reg_8_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_397);
      weight_reg_8_1_lpi_2 <= MUX_v_8_2_2(weight_reg_8_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_397);
      weight_reg_8_0_lpi_2 <= MUX_v_8_2_2(weight_reg_8_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_397);
      weight_reg_0_15_lpi_2 <= MUX_v_8_2_2(weight_reg_0_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_401);
      weight_reg_0_14_lpi_2 <= MUX_v_8_2_2(weight_reg_0_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_401);
      weight_reg_0_13_lpi_2 <= MUX_v_8_2_2(weight_reg_0_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_401);
      weight_reg_0_12_lpi_2 <= MUX_v_8_2_2(weight_reg_0_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_401);
      weight_reg_0_11_lpi_2 <= MUX_v_8_2_2(weight_reg_0_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_401);
      weight_reg_0_10_lpi_2 <= MUX_v_8_2_2(weight_reg_0_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_401);
      weight_reg_0_9_lpi_2 <= MUX_v_8_2_2(weight_reg_0_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_401);
      weight_reg_0_8_lpi_2 <= MUX_v_8_2_2(weight_reg_0_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_401);
      weight_reg_0_7_lpi_2 <= MUX_v_8_2_2(weight_reg_0_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_401);
      weight_reg_0_6_lpi_2 <= MUX_v_8_2_2(weight_reg_0_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_401);
      weight_reg_0_5_lpi_2 <= MUX_v_8_2_2(weight_reg_0_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_401);
      weight_reg_0_4_lpi_2 <= MUX_v_8_2_2(weight_reg_0_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_401);
      weight_reg_0_3_lpi_2 <= MUX_v_8_2_2(weight_reg_0_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_401);
      weight_reg_0_2_lpi_2 <= MUX_v_8_2_2(weight_reg_0_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_401);
      weight_reg_0_1_lpi_2 <= MUX_v_8_2_2(weight_reg_0_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_401);
      weight_reg_0_0_lpi_2 <= MUX_v_8_2_2(weight_reg_0_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_401);
      weight_reg_9_15_lpi_2 <= MUX_v_8_2_2(weight_reg_9_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_408);
      weight_reg_9_14_lpi_2 <= MUX_v_8_2_2(weight_reg_9_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_408);
      weight_reg_9_13_lpi_2 <= MUX_v_8_2_2(weight_reg_9_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_408);
      weight_reg_9_12_lpi_2 <= MUX_v_8_2_2(weight_reg_9_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_408);
      weight_reg_9_11_lpi_2 <= MUX_v_8_2_2(weight_reg_9_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_408);
      weight_reg_9_10_lpi_2 <= MUX_v_8_2_2(weight_reg_9_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_408);
      weight_reg_9_9_lpi_2 <= MUX_v_8_2_2(weight_reg_9_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_408);
      weight_reg_9_8_lpi_2 <= MUX_v_8_2_2(weight_reg_9_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_408);
      weight_reg_9_7_lpi_2 <= MUX_v_8_2_2(weight_reg_9_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_408);
      weight_reg_9_6_lpi_2 <= MUX_v_8_2_2(weight_reg_9_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_408);
      weight_reg_9_5_lpi_2 <= MUX_v_8_2_2(weight_reg_9_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_408);
      weight_reg_9_4_lpi_2 <= MUX_v_8_2_2(weight_reg_9_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_408);
      weight_reg_9_3_lpi_2 <= MUX_v_8_2_2(weight_reg_9_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_408);
      weight_reg_9_2_lpi_2 <= MUX_v_8_2_2(weight_reg_9_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_408);
      weight_reg_9_1_lpi_2 <= MUX_v_8_2_2(weight_reg_9_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_408);
      weight_reg_9_0_lpi_2 <= MUX_v_8_2_2(weight_reg_9_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_408);
      weight_reg_1_15_lpi_2 <= MUX_v_8_2_2(weight_reg_1_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_410);
      weight_reg_1_14_lpi_2 <= MUX_v_8_2_2(weight_reg_1_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_410);
      weight_reg_1_13_lpi_2 <= MUX_v_8_2_2(weight_reg_1_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_410);
      weight_reg_1_12_lpi_2 <= MUX_v_8_2_2(weight_reg_1_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_410);
      weight_reg_1_11_lpi_2 <= MUX_v_8_2_2(weight_reg_1_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_410);
      weight_reg_1_10_lpi_2 <= MUX_v_8_2_2(weight_reg_1_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_410);
      weight_reg_1_9_lpi_2 <= MUX_v_8_2_2(weight_reg_1_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_410);
      weight_reg_1_8_lpi_2 <= MUX_v_8_2_2(weight_reg_1_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_410);
      weight_reg_1_7_lpi_2 <= MUX_v_8_2_2(weight_reg_1_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_410);
      weight_reg_1_6_lpi_2 <= MUX_v_8_2_2(weight_reg_1_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_410);
      weight_reg_1_5_lpi_2 <= MUX_v_8_2_2(weight_reg_1_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_410);
      weight_reg_1_4_lpi_2 <= MUX_v_8_2_2(weight_reg_1_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_410);
      weight_reg_1_3_lpi_2 <= MUX_v_8_2_2(weight_reg_1_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_410);
      weight_reg_1_2_lpi_2 <= MUX_v_8_2_2(weight_reg_1_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_410);
      weight_reg_1_1_lpi_2 <= MUX_v_8_2_2(weight_reg_1_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_410);
      weight_reg_1_0_lpi_2 <= MUX_v_8_2_2(weight_reg_1_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_410);
      weight_reg_10_15_lpi_2 <= MUX_v_8_2_2(weight_reg_10_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_414);
      weight_reg_10_14_lpi_2 <= MUX_v_8_2_2(weight_reg_10_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_414);
      weight_reg_10_13_lpi_2 <= MUX_v_8_2_2(weight_reg_10_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_414);
      weight_reg_10_12_lpi_2 <= MUX_v_8_2_2(weight_reg_10_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_414);
      weight_reg_10_11_lpi_2 <= MUX_v_8_2_2(weight_reg_10_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_414);
      weight_reg_10_10_lpi_2 <= MUX_v_8_2_2(weight_reg_10_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_414);
      weight_reg_10_9_lpi_2 <= MUX_v_8_2_2(weight_reg_10_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_414);
      weight_reg_10_8_lpi_2 <= MUX_v_8_2_2(weight_reg_10_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_414);
      weight_reg_10_7_lpi_2 <= MUX_v_8_2_2(weight_reg_10_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_414);
      weight_reg_10_6_lpi_2 <= MUX_v_8_2_2(weight_reg_10_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_414);
      weight_reg_10_5_lpi_2 <= MUX_v_8_2_2(weight_reg_10_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_414);
      weight_reg_10_4_lpi_2 <= MUX_v_8_2_2(weight_reg_10_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_414);
      weight_reg_10_3_lpi_2 <= MUX_v_8_2_2(weight_reg_10_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_414);
      weight_reg_10_2_lpi_2 <= MUX_v_8_2_2(weight_reg_10_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_414);
      weight_reg_10_1_lpi_2 <= MUX_v_8_2_2(weight_reg_10_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_414);
      weight_reg_10_0_lpi_2 <= MUX_v_8_2_2(weight_reg_10_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_414);
      weight_reg_2_15_lpi_2 <= MUX_v_8_2_2(weight_reg_2_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_416);
      weight_reg_2_14_lpi_2 <= MUX_v_8_2_2(weight_reg_2_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_416);
      weight_reg_2_13_lpi_2 <= MUX_v_8_2_2(weight_reg_2_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_416);
      weight_reg_2_12_lpi_2 <= MUX_v_8_2_2(weight_reg_2_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_416);
      weight_reg_2_11_lpi_2 <= MUX_v_8_2_2(weight_reg_2_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_416);
      weight_reg_2_10_lpi_2 <= MUX_v_8_2_2(weight_reg_2_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_416);
      weight_reg_2_9_lpi_2 <= MUX_v_8_2_2(weight_reg_2_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_416);
      weight_reg_2_8_lpi_2 <= MUX_v_8_2_2(weight_reg_2_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_416);
      weight_reg_2_7_lpi_2 <= MUX_v_8_2_2(weight_reg_2_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_416);
      weight_reg_2_6_lpi_2 <= MUX_v_8_2_2(weight_reg_2_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_416);
      weight_reg_2_5_lpi_2 <= MUX_v_8_2_2(weight_reg_2_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_416);
      weight_reg_2_4_lpi_2 <= MUX_v_8_2_2(weight_reg_2_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_416);
      weight_reg_2_3_lpi_2 <= MUX_v_8_2_2(weight_reg_2_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_416);
      weight_reg_2_2_lpi_2 <= MUX_v_8_2_2(weight_reg_2_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_416);
      weight_reg_2_1_lpi_2 <= MUX_v_8_2_2(weight_reg_2_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_416);
      weight_reg_2_0_lpi_2 <= MUX_v_8_2_2(weight_reg_2_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_416);
      weight_reg_11_15_lpi_2 <= MUX_v_8_2_2(weight_reg_11_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_419);
      weight_reg_11_14_lpi_2 <= MUX_v_8_2_2(weight_reg_11_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_419);
      weight_reg_11_13_lpi_2 <= MUX_v_8_2_2(weight_reg_11_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_419);
      weight_reg_11_12_lpi_2 <= MUX_v_8_2_2(weight_reg_11_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_419);
      weight_reg_11_11_lpi_2 <= MUX_v_8_2_2(weight_reg_11_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_419);
      weight_reg_11_10_lpi_2 <= MUX_v_8_2_2(weight_reg_11_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_419);
      weight_reg_11_9_lpi_2 <= MUX_v_8_2_2(weight_reg_11_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_419);
      weight_reg_11_8_lpi_2 <= MUX_v_8_2_2(weight_reg_11_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_419);
      weight_reg_11_7_lpi_2 <= MUX_v_8_2_2(weight_reg_11_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_419);
      weight_reg_11_6_lpi_2 <= MUX_v_8_2_2(weight_reg_11_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_419);
      weight_reg_11_5_lpi_2 <= MUX_v_8_2_2(weight_reg_11_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_419);
      weight_reg_11_4_lpi_2 <= MUX_v_8_2_2(weight_reg_11_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_419);
      weight_reg_11_3_lpi_2 <= MUX_v_8_2_2(weight_reg_11_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_419);
      weight_reg_11_2_lpi_2 <= MUX_v_8_2_2(weight_reg_11_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_419);
      weight_reg_11_1_lpi_2 <= MUX_v_8_2_2(weight_reg_11_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_419);
      weight_reg_11_0_lpi_2 <= MUX_v_8_2_2(weight_reg_11_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_419);
      weight_reg_3_15_lpi_2 <= MUX_v_8_2_2(weight_reg_3_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_421);
      weight_reg_3_14_lpi_2 <= MUX_v_8_2_2(weight_reg_3_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_421);
      weight_reg_3_13_lpi_2 <= MUX_v_8_2_2(weight_reg_3_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_421);
      weight_reg_3_12_lpi_2 <= MUX_v_8_2_2(weight_reg_3_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_421);
      weight_reg_3_11_lpi_2 <= MUX_v_8_2_2(weight_reg_3_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_421);
      weight_reg_3_10_lpi_2 <= MUX_v_8_2_2(weight_reg_3_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_421);
      weight_reg_3_9_lpi_2 <= MUX_v_8_2_2(weight_reg_3_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_421);
      weight_reg_3_8_lpi_2 <= MUX_v_8_2_2(weight_reg_3_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_421);
      weight_reg_3_7_lpi_2 <= MUX_v_8_2_2(weight_reg_3_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_421);
      weight_reg_3_6_lpi_2 <= MUX_v_8_2_2(weight_reg_3_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_421);
      weight_reg_3_5_lpi_2 <= MUX_v_8_2_2(weight_reg_3_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_421);
      weight_reg_3_4_lpi_2 <= MUX_v_8_2_2(weight_reg_3_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_421);
      weight_reg_3_3_lpi_2 <= MUX_v_8_2_2(weight_reg_3_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_421);
      weight_reg_3_2_lpi_2 <= MUX_v_8_2_2(weight_reg_3_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_421);
      weight_reg_3_1_lpi_2 <= MUX_v_8_2_2(weight_reg_3_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_421);
      weight_reg_3_0_lpi_2 <= MUX_v_8_2_2(weight_reg_3_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_421);
      weight_reg_12_15_lpi_2 <= MUX_v_8_2_2(weight_reg_12_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_424);
      weight_reg_12_14_lpi_2 <= MUX_v_8_2_2(weight_reg_12_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_424);
      weight_reg_12_13_lpi_2 <= MUX_v_8_2_2(weight_reg_12_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_424);
      weight_reg_12_12_lpi_2 <= MUX_v_8_2_2(weight_reg_12_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_424);
      weight_reg_12_11_lpi_2 <= MUX_v_8_2_2(weight_reg_12_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_424);
      weight_reg_12_10_lpi_2 <= MUX_v_8_2_2(weight_reg_12_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_424);
      weight_reg_12_9_lpi_2 <= MUX_v_8_2_2(weight_reg_12_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_424);
      weight_reg_12_8_lpi_2 <= MUX_v_8_2_2(weight_reg_12_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_424);
      weight_reg_12_7_lpi_2 <= MUX_v_8_2_2(weight_reg_12_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_424);
      weight_reg_12_6_lpi_2 <= MUX_v_8_2_2(weight_reg_12_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_424);
      weight_reg_12_5_lpi_2 <= MUX_v_8_2_2(weight_reg_12_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_424);
      weight_reg_12_4_lpi_2 <= MUX_v_8_2_2(weight_reg_12_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_424);
      weight_reg_12_3_lpi_2 <= MUX_v_8_2_2(weight_reg_12_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_424);
      weight_reg_12_2_lpi_2 <= MUX_v_8_2_2(weight_reg_12_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_424);
      weight_reg_12_1_lpi_2 <= MUX_v_8_2_2(weight_reg_12_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_424);
      weight_reg_12_0_lpi_2 <= MUX_v_8_2_2(weight_reg_12_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_424);
      weight_reg_4_15_lpi_2 <= MUX_v_8_2_2(weight_reg_4_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_426);
      weight_reg_4_14_lpi_2 <= MUX_v_8_2_2(weight_reg_4_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_426);
      weight_reg_4_13_lpi_2 <= MUX_v_8_2_2(weight_reg_4_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_426);
      weight_reg_4_12_lpi_2 <= MUX_v_8_2_2(weight_reg_4_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_426);
      weight_reg_4_11_lpi_2 <= MUX_v_8_2_2(weight_reg_4_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_426);
      weight_reg_4_10_lpi_2 <= MUX_v_8_2_2(weight_reg_4_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_426);
      weight_reg_4_9_lpi_2 <= MUX_v_8_2_2(weight_reg_4_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_426);
      weight_reg_4_8_lpi_2 <= MUX_v_8_2_2(weight_reg_4_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_426);
      weight_reg_4_7_lpi_2 <= MUX_v_8_2_2(weight_reg_4_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_426);
      weight_reg_4_6_lpi_2 <= MUX_v_8_2_2(weight_reg_4_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_426);
      weight_reg_4_5_lpi_2 <= MUX_v_8_2_2(weight_reg_4_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_426);
      weight_reg_4_4_lpi_2 <= MUX_v_8_2_2(weight_reg_4_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_426);
      weight_reg_4_3_lpi_2 <= MUX_v_8_2_2(weight_reg_4_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_426);
      weight_reg_4_2_lpi_2 <= MUX_v_8_2_2(weight_reg_4_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_426);
      weight_reg_4_1_lpi_2 <= MUX_v_8_2_2(weight_reg_4_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_426);
      weight_reg_4_0_lpi_2 <= MUX_v_8_2_2(weight_reg_4_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_426);
      weight_reg_13_15_lpi_2 <= MUX_v_8_2_2(weight_reg_13_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_429);
      weight_reg_13_14_lpi_2 <= MUX_v_8_2_2(weight_reg_13_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_429);
      weight_reg_13_13_lpi_2 <= MUX_v_8_2_2(weight_reg_13_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_429);
      weight_reg_13_12_lpi_2 <= MUX_v_8_2_2(weight_reg_13_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_429);
      weight_reg_13_11_lpi_2 <= MUX_v_8_2_2(weight_reg_13_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_429);
      weight_reg_13_10_lpi_2 <= MUX_v_8_2_2(weight_reg_13_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_429);
      weight_reg_13_9_lpi_2 <= MUX_v_8_2_2(weight_reg_13_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_429);
      weight_reg_13_8_lpi_2 <= MUX_v_8_2_2(weight_reg_13_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_429);
      weight_reg_13_7_lpi_2 <= MUX_v_8_2_2(weight_reg_13_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_429);
      weight_reg_13_6_lpi_2 <= MUX_v_8_2_2(weight_reg_13_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_429);
      weight_reg_13_5_lpi_2 <= MUX_v_8_2_2(weight_reg_13_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_429);
      weight_reg_13_4_lpi_2 <= MUX_v_8_2_2(weight_reg_13_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_429);
      weight_reg_13_3_lpi_2 <= MUX_v_8_2_2(weight_reg_13_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_429);
      weight_reg_13_2_lpi_2 <= MUX_v_8_2_2(weight_reg_13_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_429);
      weight_reg_13_1_lpi_2 <= MUX_v_8_2_2(weight_reg_13_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_429);
      weight_reg_13_0_lpi_2 <= MUX_v_8_2_2(weight_reg_13_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_429);
      weight_reg_5_15_lpi_2 <= MUX_v_8_2_2(weight_reg_5_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_431);
      weight_reg_5_14_lpi_2 <= MUX_v_8_2_2(weight_reg_5_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_431);
      weight_reg_5_13_lpi_2 <= MUX_v_8_2_2(weight_reg_5_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_431);
      weight_reg_5_12_lpi_2 <= MUX_v_8_2_2(weight_reg_5_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_431);
      weight_reg_5_11_lpi_2 <= MUX_v_8_2_2(weight_reg_5_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_431);
      weight_reg_5_10_lpi_2 <= MUX_v_8_2_2(weight_reg_5_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_431);
      weight_reg_5_9_lpi_2 <= MUX_v_8_2_2(weight_reg_5_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_431);
      weight_reg_5_8_lpi_2 <= MUX_v_8_2_2(weight_reg_5_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_431);
      weight_reg_5_7_lpi_2 <= MUX_v_8_2_2(weight_reg_5_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_431);
      weight_reg_5_6_lpi_2 <= MUX_v_8_2_2(weight_reg_5_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_431);
      weight_reg_5_5_lpi_2 <= MUX_v_8_2_2(weight_reg_5_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_431);
      weight_reg_5_4_lpi_2 <= MUX_v_8_2_2(weight_reg_5_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_431);
      weight_reg_5_3_lpi_2 <= MUX_v_8_2_2(weight_reg_5_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_431);
      weight_reg_5_2_lpi_2 <= MUX_v_8_2_2(weight_reg_5_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_431);
      weight_reg_5_1_lpi_2 <= MUX_v_8_2_2(weight_reg_5_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_431);
      weight_reg_5_0_lpi_2 <= MUX_v_8_2_2(weight_reg_5_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_431);
      weight_reg_14_15_lpi_2 <= MUX_v_8_2_2(weight_reg_14_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_434);
      weight_reg_14_14_lpi_2 <= MUX_v_8_2_2(weight_reg_14_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_434);
      weight_reg_14_13_lpi_2 <= MUX_v_8_2_2(weight_reg_14_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_434);
      weight_reg_14_12_lpi_2 <= MUX_v_8_2_2(weight_reg_14_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_434);
      weight_reg_14_11_lpi_2 <= MUX_v_8_2_2(weight_reg_14_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_434);
      weight_reg_14_10_lpi_2 <= MUX_v_8_2_2(weight_reg_14_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_434);
      weight_reg_14_9_lpi_2 <= MUX_v_8_2_2(weight_reg_14_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_434);
      weight_reg_14_8_lpi_2 <= MUX_v_8_2_2(weight_reg_14_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_434);
      weight_reg_14_7_lpi_2 <= MUX_v_8_2_2(weight_reg_14_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_434);
      weight_reg_14_6_lpi_2 <= MUX_v_8_2_2(weight_reg_14_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_434);
      weight_reg_14_5_lpi_2 <= MUX_v_8_2_2(weight_reg_14_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_434);
      weight_reg_14_4_lpi_2 <= MUX_v_8_2_2(weight_reg_14_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_434);
      weight_reg_14_3_lpi_2 <= MUX_v_8_2_2(weight_reg_14_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_434);
      weight_reg_14_2_lpi_2 <= MUX_v_8_2_2(weight_reg_14_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_434);
      weight_reg_14_1_lpi_2 <= MUX_v_8_2_2(weight_reg_14_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_434);
      weight_reg_14_0_lpi_2 <= MUX_v_8_2_2(weight_reg_14_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_434);
      weight_reg_6_15_lpi_2 <= MUX_v_8_2_2(weight_reg_6_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_436);
      weight_reg_6_14_lpi_2 <= MUX_v_8_2_2(weight_reg_6_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_436);
      weight_reg_6_13_lpi_2 <= MUX_v_8_2_2(weight_reg_6_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_436);
      weight_reg_6_12_lpi_2 <= MUX_v_8_2_2(weight_reg_6_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_436);
      weight_reg_6_11_lpi_2 <= MUX_v_8_2_2(weight_reg_6_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_436);
      weight_reg_6_10_lpi_2 <= MUX_v_8_2_2(weight_reg_6_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_436);
      weight_reg_6_9_lpi_2 <= MUX_v_8_2_2(weight_reg_6_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_436);
      weight_reg_6_8_lpi_2 <= MUX_v_8_2_2(weight_reg_6_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_436);
      weight_reg_6_7_lpi_2 <= MUX_v_8_2_2(weight_reg_6_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_436);
      weight_reg_6_6_lpi_2 <= MUX_v_8_2_2(weight_reg_6_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_436);
      weight_reg_6_5_lpi_2 <= MUX_v_8_2_2(weight_reg_6_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_436);
      weight_reg_6_4_lpi_2 <= MUX_v_8_2_2(weight_reg_6_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_436);
      weight_reg_6_3_lpi_2 <= MUX_v_8_2_2(weight_reg_6_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_436);
      weight_reg_6_2_lpi_2 <= MUX_v_8_2_2(weight_reg_6_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_436);
      weight_reg_6_1_lpi_2 <= MUX_v_8_2_2(weight_reg_6_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_436);
      weight_reg_6_0_lpi_2 <= MUX_v_8_2_2(weight_reg_6_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_436);
      weight_reg_15_15_lpi_2 <= MUX_v_8_2_2(weight_reg_15_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_33);
      weight_reg_15_14_lpi_2 <= MUX_v_8_2_2(weight_reg_15_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_33);
      weight_reg_15_13_lpi_2 <= MUX_v_8_2_2(weight_reg_15_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_33);
      weight_reg_15_12_lpi_2 <= MUX_v_8_2_2(weight_reg_15_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_33);
      weight_reg_15_11_lpi_2 <= MUX_v_8_2_2(weight_reg_15_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_33);
      weight_reg_15_10_lpi_2 <= MUX_v_8_2_2(weight_reg_15_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_33);
      weight_reg_15_9_lpi_2 <= MUX_v_8_2_2(weight_reg_15_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_33);
      weight_reg_15_8_lpi_2 <= MUX_v_8_2_2(weight_reg_15_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_33);
      weight_reg_15_7_lpi_2 <= MUX_v_8_2_2(weight_reg_15_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_33);
      weight_reg_15_6_lpi_2 <= MUX_v_8_2_2(weight_reg_15_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_33);
      weight_reg_15_5_lpi_2 <= MUX_v_8_2_2(weight_reg_15_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_33);
      weight_reg_15_4_lpi_2 <= MUX_v_8_2_2(weight_reg_15_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_33);
      weight_reg_15_3_lpi_2 <= MUX_v_8_2_2(weight_reg_15_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_33);
      weight_reg_15_2_lpi_2 <= MUX_v_8_2_2(weight_reg_15_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_33);
      weight_reg_15_1_lpi_2 <= MUX_v_8_2_2(weight_reg_15_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_33);
      weight_reg_15_0_lpi_2 <= MUX_v_8_2_2(weight_reg_15_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_33);
      weight_reg_7_15_lpi_2 <= MUX_v_8_2_2(weight_reg_7_15_lpi_2, (weight_rsci_idat_mxwt[127:120]),
          and_dcpl_438);
      weight_reg_7_14_lpi_2 <= MUX_v_8_2_2(weight_reg_7_14_lpi_2, (weight_rsci_idat_mxwt[119:112]),
          and_dcpl_438);
      weight_reg_7_13_lpi_2 <= MUX_v_8_2_2(weight_reg_7_13_lpi_2, (weight_rsci_idat_mxwt[111:104]),
          and_dcpl_438);
      weight_reg_7_12_lpi_2 <= MUX_v_8_2_2(weight_reg_7_12_lpi_2, (weight_rsci_idat_mxwt[103:96]),
          and_dcpl_438);
      weight_reg_7_11_lpi_2 <= MUX_v_8_2_2(weight_reg_7_11_lpi_2, (weight_rsci_idat_mxwt[95:88]),
          and_dcpl_438);
      weight_reg_7_10_lpi_2 <= MUX_v_8_2_2(weight_reg_7_10_lpi_2, (weight_rsci_idat_mxwt[87:80]),
          and_dcpl_438);
      weight_reg_7_9_lpi_2 <= MUX_v_8_2_2(weight_reg_7_9_lpi_2, (weight_rsci_idat_mxwt[79:72]),
          and_dcpl_438);
      weight_reg_7_8_lpi_2 <= MUX_v_8_2_2(weight_reg_7_8_lpi_2, (weight_rsci_idat_mxwt[71:64]),
          and_dcpl_438);
      weight_reg_7_7_lpi_2 <= MUX_v_8_2_2(weight_reg_7_7_lpi_2, (weight_rsci_idat_mxwt[63:56]),
          and_dcpl_438);
      weight_reg_7_6_lpi_2 <= MUX_v_8_2_2(weight_reg_7_6_lpi_2, (weight_rsci_idat_mxwt[55:48]),
          and_dcpl_438);
      weight_reg_7_5_lpi_2 <= MUX_v_8_2_2(weight_reg_7_5_lpi_2, (weight_rsci_idat_mxwt[47:40]),
          and_dcpl_438);
      weight_reg_7_4_lpi_2 <= MUX_v_8_2_2(weight_reg_7_4_lpi_2, (weight_rsci_idat_mxwt[39:32]),
          and_dcpl_438);
      weight_reg_7_3_lpi_2 <= MUX_v_8_2_2(weight_reg_7_3_lpi_2, (weight_rsci_idat_mxwt[31:24]),
          and_dcpl_438);
      weight_reg_7_2_lpi_2 <= MUX_v_8_2_2(weight_reg_7_2_lpi_2, (weight_rsci_idat_mxwt[23:16]),
          and_dcpl_438);
      weight_reg_7_1_lpi_2 <= MUX_v_8_2_2(weight_reg_7_1_lpi_2, (weight_rsci_idat_mxwt[15:8]),
          and_dcpl_438);
      weight_reg_7_0_lpi_2 <= MUX_v_8_2_2(weight_reg_7_0_lpi_2, (weight_rsci_idat_mxwt[7:0]),
          and_dcpl_438);
      step_in_col_value_lpi_2 <= MUX_v_128_2_2(step_in_col_value_lpi_2, input_rsci_idat_mxwt,
          and_441_nl);
      psum_reg_16_15_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_15_lpi_2, output_fifo_3_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_312_nl)) , and_dcpl_12 , and_dcpl_42});
      psum_reg_16_14_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_14_lpi_2, accum_fifo_0_run_cmp_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(psum_reg_or_4_nl) , (psum_reg_and_242_nl)
          , and_dcpl_45});
      psum_reg_16_12_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_12_lpi_2, output_fifo_14_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_317_nl)) , and_dcpl_12 , and_dcpl_51});
      psum_reg_16_11_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_11_lpi_2, output_fifo_13_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_318_nl)) , and_dcpl_12 , and_dcpl_47});
      psum_reg_16_10_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_10_lpi_2, output_fifo_12_rsci_output_rsc_z,
          accum_fifo_3_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_325_nl))
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_239});
      psum_reg_16_9_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_9_lpi_2, accum_fifo_9_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_329_nl)) , and_dcpl_42 , and_dcpl_223});
      psum_reg_16_8_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_8_lpi_2, output_fifo_1_rsci_output_rsc_z,
          accum_fifo_8_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_333_nl))
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_205});
      psum_reg_16_7_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_7_lpi_2, output_fifo_10_rsci_output_rsc_z,
          accum_fifo_7_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(mux_336_nl)
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_185});
      psum_reg_16_6_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_6_lpi_2, output_fifo_9_rsci_output_rsc_z,
          accum_fifo_6_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_340_nl))
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_169});
      psum_reg_16_5_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_5_lpi_2, output_fifo_8_rsci_output_rsc_z,
          accum_fifo_5_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_344_nl))
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_153});
      psum_reg_16_4_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_4_lpi_2, output_fifo_7_rsci_output_rsc_z,
          accum_fifo_4_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_348_nl))
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_135});
      psum_reg_16_3_lpi_2 <= MUX1HOT_v_16_3_2(psum_reg_16_3_lpi_2, output_fifo_6_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {(~ (mux_350_nl)) , and_dcpl_12 , and_dcpl_116});
      psum_reg_16_2_lpi_2 <= MUX1HOT_v_16_4_2(psum_reg_16_2_lpi_2, output_fifo_5_rsci_output_rsc_z,
          ({8'b00000000 , (step_input_fifo_input_15_mux_nl)}), pe_0_0_run_cmp_psum_out_rsc_z,
          {(~ (mux_354_nl)) , and_dcpl_12 , (and_447_nl) , and_dcpl_100});
      step_output_buf_value_0_sva <= MUX1HOT_v_16_4_2(step_output_buf_value_0_sva,
          output_fifo_0_rsci_output_rsc_z, accum_fifo_0_run_cmp_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z,
          {(~ (mux_363_nl)) , and_dcpl_12 , and_dcpl_42 , and_dcpl_53});
      step_step_sva <= MUX_v_16_2_2(16'b0000000000000000, (step_step_mux_nl), (step_step_not_nl));
      paramsIn_crt_sva_127_32 <= MUX_v_96_2_2(paramsIn_crt_sva_127_32, paramsIn_rsci_idat_mxwt,
          mux_tmp_345);
      loopIndicesIn_crt_sva <= MUX_v_48_2_2(loopIndicesIn_crt_sva, loopIndicesIn_rsci_idat_mxwt,
          mux_tmp_345);
      operator_16_false_slc_operator_16_false_acc_12_svs <= MUX_s_1_2_2(operator_16_false_acc_itm_12_1,
          step_if_2_if_step_if_2_if_and_tmp, and_dcpl_12);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_14_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_35 | or_dcpl_32)) ) begin
      psum_reg_14_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_13_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_35 | or_dcpl_38)) ) begin
      psum_reg_13_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_12_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_35 | or_dcpl_41)) ) begin
      psum_reg_12_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_11_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_44)) ) begin
      psum_reg_11_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_10_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_50)) ) begin
      psum_reg_10_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_9_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_52)) ) begin
      psum_reg_9_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_8_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_54)) ) begin
      psum_reg_8_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_7_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_57)) ) begin
      psum_reg_7_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_6_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_59)) ) begin
      psum_reg_6_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_5_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_61)) ) begin
      psum_reg_5_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_4_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_48 | or_dcpl_63)) ) begin
      psum_reg_4_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_3_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_66 | or_dcpl_44)) ) begin
      psum_reg_3_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_2_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_66 | or_dcpl_50)) ) begin
      psum_reg_2_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_1_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (~(or_dcpl_66 | or_dcpl_52)) ) begin
      psum_reg_1_16_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_15_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_66 | or_dcpl_54)) ) begin
      input_reg_15_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_15_lpi_2 <= 8'b00000000;
      psum_reg_14_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_1_cse ) begin
      input_reg_14_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_15_lpi_2 <= 8'b00000000;
      psum_reg_13_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_2_cse ) begin
      input_reg_13_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_15_lpi_2 <= 8'b00000000;
      psum_reg_12_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_3_cse ) begin
      input_reg_12_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_15_lpi_2 <= 8'b00000000;
      psum_reg_11_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_4_cse ) begin
      input_reg_11_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_15_lpi_2 <= 8'b00000000;
      psum_reg_10_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_5_cse ) begin
      input_reg_10_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_15_lpi_2 <= 8'b00000000;
      psum_reg_9_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_6_cse ) begin
      input_reg_9_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_15_lpi_2 <= 8'b00000000;
      psum_reg_8_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_7_cse ) begin
      input_reg_8_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_15_lpi_2 <= 8'b00000000;
      psum_reg_7_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_8_cse ) begin
      input_reg_7_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_15_lpi_2 <= 8'b00000000;
      psum_reg_6_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_9_cse ) begin
      input_reg_6_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_15_lpi_2 <= 8'b00000000;
      psum_reg_5_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_10_cse ) begin
      input_reg_5_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_15_lpi_2 <= 8'b00000000;
      psum_reg_4_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_11_cse ) begin
      input_reg_4_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_15_lpi_2 <= 8'b00000000;
      psum_reg_3_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_12_cse ) begin
      input_reg_3_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_15_lpi_2 <= 8'b00000000;
      psum_reg_2_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_13_cse ) begin
      input_reg_2_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_15_lpi_2 <= 8'b00000000;
      psum_reg_1_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_14_cse ) begin
      input_reg_1_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_15_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_14_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_85 | or_dcpl_52)) ) begin
      input_reg_15_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_14_lpi_2 <= 8'b00000000;
      psum_reg_14_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_16_cse ) begin
      input_reg_14_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_14_lpi_2 <= 8'b00000000;
      psum_reg_13_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_17_cse ) begin
      input_reg_13_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_14_lpi_2 <= 8'b00000000;
      psum_reg_12_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_18_cse ) begin
      input_reg_12_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_14_lpi_2 <= 8'b00000000;
      psum_reg_11_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_19_cse ) begin
      input_reg_11_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_14_lpi_2 <= 8'b00000000;
      psum_reg_10_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_20_cse ) begin
      input_reg_10_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_14_lpi_2 <= 8'b00000000;
      psum_reg_9_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_21_cse ) begin
      input_reg_9_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_14_lpi_2 <= 8'b00000000;
      psum_reg_8_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_22_cse ) begin
      input_reg_8_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_14_lpi_2 <= 8'b00000000;
      psum_reg_7_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_23_cse ) begin
      input_reg_7_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_14_lpi_2 <= 8'b00000000;
      psum_reg_6_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_24_cse ) begin
      input_reg_6_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_14_lpi_2 <= 8'b00000000;
      psum_reg_5_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_25_cse ) begin
      input_reg_5_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_14_lpi_2 <= 8'b00000000;
      psum_reg_4_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_26_cse ) begin
      input_reg_4_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_14_lpi_2 <= 8'b00000000;
      psum_reg_3_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_27_cse ) begin
      input_reg_3_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_14_lpi_2 <= 8'b00000000;
      psum_reg_2_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_28_cse ) begin
      input_reg_2_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_14_lpi_2 <= 8'b00000000;
      psum_reg_1_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_29_cse ) begin
      input_reg_1_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_14_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_13_lpi_2 <= 8'b00000000;
      psum_reg_15_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_30_cse ) begin
      input_reg_15_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_13_lpi_2 <= 8'b00000000;
      psum_reg_14_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_31_cse ) begin
      input_reg_14_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_13_lpi_2 <= 8'b00000000;
      psum_reg_13_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_32_cse ) begin
      input_reg_13_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_13_lpi_2 <= 8'b00000000;
      psum_reg_12_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_33_cse ) begin
      input_reg_12_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_13_lpi_2 <= 8'b00000000;
      psum_reg_11_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_34_cse ) begin
      input_reg_11_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_13_lpi_2 <= 8'b00000000;
      psum_reg_10_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_35_cse ) begin
      input_reg_10_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_13_lpi_2 <= 8'b00000000;
      psum_reg_9_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_36_cse ) begin
      input_reg_9_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_13_lpi_2 <= 8'b00000000;
      psum_reg_8_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_37_cse ) begin
      input_reg_8_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_13_lpi_2 <= 8'b00000000;
      psum_reg_7_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_38_cse ) begin
      input_reg_7_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_13_lpi_2 <= 8'b00000000;
      psum_reg_6_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_39_cse ) begin
      input_reg_6_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_13_lpi_2 <= 8'b00000000;
      psum_reg_5_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_40_cse ) begin
      input_reg_5_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_13_lpi_2 <= 8'b00000000;
      psum_reg_4_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_41_cse ) begin
      input_reg_4_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_13_lpi_2 <= 8'b00000000;
      psum_reg_3_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_42_cse ) begin
      input_reg_3_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_13_lpi_2 <= 8'b00000000;
      psum_reg_2_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_43_cse ) begin
      input_reg_2_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_13_lpi_2 <= 8'b00000000;
      psum_reg_1_13_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_44_cse ) begin
      input_reg_1_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_13_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_12_lpi_2 <= 8'b00000000;
      psum_reg_15_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_45_cse ) begin
      input_reg_15_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_12_lpi_2 <= 8'b00000000;
      psum_reg_14_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_46_cse ) begin
      input_reg_14_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_12_lpi_2 <= 8'b00000000;
      psum_reg_13_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_47_cse ) begin
      input_reg_13_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_12_lpi_2 <= 8'b00000000;
      psum_reg_12_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_48_cse ) begin
      input_reg_12_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_12_lpi_2 <= 8'b00000000;
      psum_reg_11_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_49_cse ) begin
      input_reg_11_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_12_lpi_2 <= 8'b00000000;
      psum_reg_10_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_50_cse ) begin
      input_reg_10_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_12_lpi_2 <= 8'b00000000;
      psum_reg_9_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_51_cse ) begin
      input_reg_9_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_12_lpi_2 <= 8'b00000000;
      psum_reg_8_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_52_cse ) begin
      input_reg_8_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_12_lpi_2 <= 8'b00000000;
      psum_reg_7_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_53_cse ) begin
      input_reg_7_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_12_lpi_2 <= 8'b00000000;
      psum_reg_6_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_54_cse ) begin
      input_reg_6_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_12_lpi_2 <= 8'b00000000;
      psum_reg_5_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_55_cse ) begin
      input_reg_5_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_12_lpi_2 <= 8'b00000000;
      psum_reg_4_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_56_cse ) begin
      input_reg_4_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_12_lpi_2 <= 8'b00000000;
      psum_reg_3_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_57_cse ) begin
      input_reg_3_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_12_lpi_2 <= 8'b00000000;
      psum_reg_2_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_58_cse ) begin
      input_reg_2_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_12_lpi_2 <= 8'b00000000;
      psum_reg_1_12_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_59_cse ) begin
      input_reg_1_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_12_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_11_lpi_2 <= 8'b00000000;
      psum_reg_15_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_60_cse ) begin
      input_reg_15_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_11_lpi_2 <= 8'b00000000;
      psum_reg_14_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_61_cse ) begin
      input_reg_14_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_11_lpi_2 <= 8'b00000000;
      psum_reg_13_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_62_cse ) begin
      input_reg_13_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_11_lpi_2 <= 8'b00000000;
      psum_reg_12_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_63_cse ) begin
      input_reg_12_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_11_lpi_2 <= 8'b00000000;
      psum_reg_11_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_64_cse ) begin
      input_reg_11_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_11_lpi_2 <= 8'b00000000;
      psum_reg_10_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_65_cse ) begin
      input_reg_10_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_11_lpi_2 <= 8'b00000000;
      psum_reg_9_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_66_cse ) begin
      input_reg_9_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_11_lpi_2 <= 8'b00000000;
      psum_reg_8_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_67_cse ) begin
      input_reg_8_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_11_lpi_2 <= 8'b00000000;
      psum_reg_7_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_68_cse ) begin
      input_reg_7_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_11_lpi_2 <= 8'b00000000;
      psum_reg_6_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_69_cse ) begin
      input_reg_6_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_11_lpi_2 <= 8'b00000000;
      psum_reg_5_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_70_cse ) begin
      input_reg_5_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_11_lpi_2 <= 8'b00000000;
      psum_reg_4_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_71_cse ) begin
      input_reg_4_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_11_lpi_2 <= 8'b00000000;
      psum_reg_3_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_72_cse ) begin
      input_reg_3_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_11_lpi_2 <= 8'b00000000;
      psum_reg_2_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_73_cse ) begin
      input_reg_2_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_11_lpi_2 <= 8'b00000000;
      psum_reg_1_11_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_74_cse ) begin
      input_reg_1_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_11_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_10_lpi_2 <= 8'b00000000;
      psum_reg_15_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_75_cse ) begin
      input_reg_15_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_10_lpi_2 <= 8'b00000000;
      psum_reg_14_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_76_cse ) begin
      input_reg_14_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_10_lpi_2 <= 8'b00000000;
      psum_reg_13_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_77_cse ) begin
      input_reg_13_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_10_lpi_2 <= 8'b00000000;
      psum_reg_12_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_78_cse ) begin
      input_reg_12_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_10_lpi_2 <= 8'b00000000;
      psum_reg_11_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_79_cse ) begin
      input_reg_11_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_10_lpi_2 <= 8'b00000000;
      psum_reg_10_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_80_cse ) begin
      input_reg_10_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_10_lpi_2 <= 8'b00000000;
      psum_reg_9_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_81_cse ) begin
      input_reg_9_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_10_lpi_2 <= 8'b00000000;
      psum_reg_8_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_82_cse ) begin
      input_reg_8_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_10_lpi_2 <= 8'b00000000;
      psum_reg_7_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_83_cse ) begin
      input_reg_7_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_10_lpi_2 <= 8'b00000000;
      psum_reg_6_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_84_cse ) begin
      input_reg_6_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_10_lpi_2 <= 8'b00000000;
      psum_reg_5_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_85_cse ) begin
      input_reg_5_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_10_lpi_2 <= 8'b00000000;
      psum_reg_4_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_86_cse ) begin
      input_reg_4_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_10_lpi_2 <= 8'b00000000;
      psum_reg_3_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_87_cse ) begin
      input_reg_3_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_10_lpi_2 <= 8'b00000000;
      psum_reg_2_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_88_cse ) begin
      input_reg_2_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_10_lpi_2 <= 8'b00000000;
      psum_reg_1_10_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_89_cse ) begin
      input_reg_1_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_10_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_9_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_133 | or_dcpl_38)) ) begin
      input_reg_16_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_9_lpi_2 <= 8'b00000000;
      psum_reg_15_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_91_cse ) begin
      input_reg_15_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_9_lpi_2 <= 8'b00000000;
      psum_reg_14_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_92_cse ) begin
      input_reg_14_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_9_lpi_2 <= 8'b00000000;
      psum_reg_13_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_93_cse ) begin
      input_reg_13_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_9_lpi_2 <= 8'b00000000;
      psum_reg_12_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_94_cse ) begin
      input_reg_12_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_9_lpi_2 <= 8'b00000000;
      psum_reg_11_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_95_cse ) begin
      input_reg_11_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_9_lpi_2 <= 8'b00000000;
      psum_reg_10_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_96_cse ) begin
      input_reg_10_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_9_lpi_2 <= 8'b00000000;
      psum_reg_9_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_97_cse ) begin
      input_reg_9_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_9_lpi_2 <= 8'b00000000;
      psum_reg_8_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_98_cse ) begin
      input_reg_8_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_9_lpi_2 <= 8'b00000000;
      psum_reg_7_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_99_cse ) begin
      input_reg_7_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_9_lpi_2 <= 8'b00000000;
      psum_reg_6_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_100_cse ) begin
      input_reg_6_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_9_lpi_2 <= 8'b00000000;
      psum_reg_5_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_101_cse ) begin
      input_reg_5_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_9_lpi_2 <= 8'b00000000;
      psum_reg_4_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_102_cse ) begin
      input_reg_4_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_9_lpi_2 <= 8'b00000000;
      psum_reg_3_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_103_cse ) begin
      input_reg_3_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_9_lpi_2 <= 8'b00000000;
      psum_reg_2_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_104_cse ) begin
      input_reg_2_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_9_lpi_2 <= 8'b00000000;
      psum_reg_1_9_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_105_cse ) begin
      input_reg_1_9_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_9_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_8_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_151 | or_dcpl_38)) ) begin
      input_reg_16_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_8_lpi_2 <= 8'b00000000;
      psum_reg_15_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_107_cse ) begin
      input_reg_15_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_8_lpi_2 <= 8'b00000000;
      psum_reg_14_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_108_cse ) begin
      input_reg_14_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_8_lpi_2 <= 8'b00000000;
      psum_reg_13_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_109_cse ) begin
      input_reg_13_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_8_lpi_2 <= 8'b00000000;
      psum_reg_12_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_110_cse ) begin
      input_reg_12_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_8_lpi_2 <= 8'b00000000;
      psum_reg_11_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_111_cse ) begin
      input_reg_11_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_8_lpi_2 <= 8'b00000000;
      psum_reg_10_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_112_cse ) begin
      input_reg_10_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_8_lpi_2 <= 8'b00000000;
      psum_reg_9_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_113_cse ) begin
      input_reg_9_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_8_lpi_2 <= 8'b00000000;
      psum_reg_8_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_114_cse ) begin
      input_reg_8_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_8_lpi_2 <= 8'b00000000;
      psum_reg_7_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_115_cse ) begin
      input_reg_7_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_8_lpi_2 <= 8'b00000000;
      psum_reg_6_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_116_cse ) begin
      input_reg_6_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_8_lpi_2 <= 8'b00000000;
      psum_reg_5_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_117_cse ) begin
      input_reg_5_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_8_lpi_2 <= 8'b00000000;
      psum_reg_4_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_118_cse ) begin
      input_reg_4_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_8_lpi_2 <= 8'b00000000;
      psum_reg_3_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_119_cse ) begin
      input_reg_3_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_8_lpi_2 <= 8'b00000000;
      psum_reg_2_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_120_cse ) begin
      input_reg_2_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_8_lpi_2 <= 8'b00000000;
      psum_reg_1_8_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_121_cse ) begin
      input_reg_1_8_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_8_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_7_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_201 | or_dcpl_61)) ) begin
      input_reg_16_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_7_lpi_2 <= 8'b00000000;
      psum_reg_15_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_123_cse ) begin
      input_reg_15_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_7_lpi_2 <= 8'b00000000;
      psum_reg_14_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_124_cse ) begin
      input_reg_14_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_7_lpi_2 <= 8'b00000000;
      psum_reg_13_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_125_cse ) begin
      input_reg_13_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_7_lpi_2 <= 8'b00000000;
      psum_reg_12_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_126_cse ) begin
      input_reg_12_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_7_lpi_2 <= 8'b00000000;
      psum_reg_11_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_127_cse ) begin
      input_reg_11_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_7_lpi_2 <= 8'b00000000;
      psum_reg_10_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_128_cse ) begin
      input_reg_10_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_7_lpi_2 <= 8'b00000000;
      psum_reg_9_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_129_cse ) begin
      input_reg_9_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_7_lpi_2 <= 8'b00000000;
      psum_reg_8_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_130_cse ) begin
      input_reg_8_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_7_lpi_2 <= 8'b00000000;
      psum_reg_7_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_131_cse ) begin
      input_reg_7_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_7_lpi_2 <= 8'b00000000;
      psum_reg_6_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_132_cse ) begin
      input_reg_6_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_7_lpi_2 <= 8'b00000000;
      psum_reg_5_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_133_cse ) begin
      input_reg_5_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_7_lpi_2 <= 8'b00000000;
      psum_reg_4_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_134_cse ) begin
      input_reg_4_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_7_lpi_2 <= 8'b00000000;
      psum_reg_3_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_135_cse ) begin
      input_reg_3_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_7_lpi_2 <= 8'b00000000;
      psum_reg_2_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_136_cse ) begin
      input_reg_2_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_7_lpi_2 <= 8'b00000000;
      psum_reg_1_7_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_137_cse ) begin
      input_reg_1_7_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_7_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_6_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_219 | or_dcpl_61)) ) begin
      input_reg_16_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_6_lpi_2 <= 8'b00000000;
      psum_reg_15_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_139_cse ) begin
      input_reg_15_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_6_lpi_2 <= 8'b00000000;
      psum_reg_14_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_140_cse ) begin
      input_reg_14_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_6_lpi_2 <= 8'b00000000;
      psum_reg_13_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_141_cse ) begin
      input_reg_13_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_6_lpi_2 <= 8'b00000000;
      psum_reg_12_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_142_cse ) begin
      input_reg_12_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_6_lpi_2 <= 8'b00000000;
      psum_reg_11_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_143_cse ) begin
      input_reg_11_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_6_lpi_2 <= 8'b00000000;
      psum_reg_10_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_144_cse ) begin
      input_reg_10_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_6_lpi_2 <= 8'b00000000;
      psum_reg_9_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_145_cse ) begin
      input_reg_9_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_6_lpi_2 <= 8'b00000000;
      psum_reg_8_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_146_cse ) begin
      input_reg_8_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_6_lpi_2 <= 8'b00000000;
      psum_reg_7_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_147_cse ) begin
      input_reg_7_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_6_lpi_2 <= 8'b00000000;
      psum_reg_6_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_148_cse ) begin
      input_reg_6_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_6_lpi_2 <= 8'b00000000;
      psum_reg_5_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_149_cse ) begin
      input_reg_5_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_6_lpi_2 <= 8'b00000000;
      psum_reg_4_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_150_cse ) begin
      input_reg_4_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_6_lpi_2 <= 8'b00000000;
      psum_reg_3_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_151_cse ) begin
      input_reg_3_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_6_lpi_2 <= 8'b00000000;
      psum_reg_2_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_152_cse ) begin
      input_reg_2_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_6_lpi_2 <= 8'b00000000;
      psum_reg_1_6_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_153_cse ) begin
      input_reg_1_6_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_6_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_5_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_201 | or_dcpl_38)) ) begin
      input_reg_16_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_5_lpi_2 <= 8'b00000000;
      psum_reg_15_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_155_cse ) begin
      input_reg_15_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_5_lpi_2 <= 8'b00000000;
      psum_reg_14_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_156_cse ) begin
      input_reg_14_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_5_lpi_2 <= 8'b00000000;
      psum_reg_13_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_157_cse ) begin
      input_reg_13_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_5_lpi_2 <= 8'b00000000;
      psum_reg_12_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_158_cse ) begin
      input_reg_12_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_5_lpi_2 <= 8'b00000000;
      psum_reg_11_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_159_cse ) begin
      input_reg_11_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_5_lpi_2 <= 8'b00000000;
      psum_reg_10_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_160_cse ) begin
      input_reg_10_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_5_lpi_2 <= 8'b00000000;
      psum_reg_9_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_161_cse ) begin
      input_reg_9_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_5_lpi_2 <= 8'b00000000;
      psum_reg_8_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_162_cse ) begin
      input_reg_8_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_5_lpi_2 <= 8'b00000000;
      psum_reg_7_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_163_cse ) begin
      input_reg_7_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_5_lpi_2 <= 8'b00000000;
      psum_reg_6_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_164_cse ) begin
      input_reg_6_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_5_lpi_2 <= 8'b00000000;
      psum_reg_5_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_165_cse ) begin
      input_reg_5_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_5_lpi_2 <= 8'b00000000;
      psum_reg_4_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_166_cse ) begin
      input_reg_4_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_5_lpi_2 <= 8'b00000000;
      psum_reg_3_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_167_cse ) begin
      input_reg_3_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_5_lpi_2 <= 8'b00000000;
      psum_reg_2_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_168_cse ) begin
      input_reg_2_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_5_lpi_2 <= 8'b00000000;
      psum_reg_1_5_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_169_cse ) begin
      input_reg_1_5_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_5_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_4_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_219 | or_dcpl_38)) ) begin
      input_reg_16_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_4_lpi_2 <= 8'b00000000;
      psum_reg_15_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_171_cse ) begin
      input_reg_15_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_4_lpi_2 <= 8'b00000000;
      psum_reg_14_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_172_cse ) begin
      input_reg_14_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_4_lpi_2 <= 8'b00000000;
      psum_reg_13_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_173_cse ) begin
      input_reg_13_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_4_lpi_2 <= 8'b00000000;
      psum_reg_12_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_174_cse ) begin
      input_reg_12_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_4_lpi_2 <= 8'b00000000;
      psum_reg_11_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_175_cse ) begin
      input_reg_11_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_4_lpi_2 <= 8'b00000000;
      psum_reg_10_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_176_cse ) begin
      input_reg_10_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_4_lpi_2 <= 8'b00000000;
      psum_reg_9_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_177_cse ) begin
      input_reg_9_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_4_lpi_2 <= 8'b00000000;
      psum_reg_8_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_178_cse ) begin
      input_reg_8_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_4_lpi_2 <= 8'b00000000;
      psum_reg_7_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_179_cse ) begin
      input_reg_7_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_4_lpi_2 <= 8'b00000000;
      psum_reg_6_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_180_cse ) begin
      input_reg_6_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_4_lpi_2 <= 8'b00000000;
      psum_reg_5_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_181_cse ) begin
      input_reg_5_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_4_lpi_2 <= 8'b00000000;
      psum_reg_4_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_182_cse ) begin
      input_reg_4_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_4_lpi_2 <= 8'b00000000;
      psum_reg_3_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_183_cse ) begin
      input_reg_3_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_4_lpi_2 <= 8'b00000000;
      psum_reg_2_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_184_cse ) begin
      input_reg_2_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_4_lpi_2 <= 8'b00000000;
      psum_reg_1_4_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_185_cse ) begin
      input_reg_1_4_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_4_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_3_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_269 | or_dcpl_61)) ) begin
      input_reg_16_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_3_lpi_2 <= 8'b00000000;
      psum_reg_15_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_187_cse ) begin
      input_reg_15_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_3_lpi_2 <= 8'b00000000;
      psum_reg_14_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_188_cse ) begin
      input_reg_14_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_3_lpi_2 <= 8'b00000000;
      psum_reg_13_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_189_cse ) begin
      input_reg_13_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_3_lpi_2 <= 8'b00000000;
      psum_reg_12_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_190_cse ) begin
      input_reg_12_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_3_lpi_2 <= 8'b00000000;
      psum_reg_11_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_191_cse ) begin
      input_reg_11_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_3_lpi_2 <= 8'b00000000;
      psum_reg_10_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_192_cse ) begin
      input_reg_10_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_3_lpi_2 <= 8'b00000000;
      psum_reg_9_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_193_cse ) begin
      input_reg_9_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_3_lpi_2 <= 8'b00000000;
      psum_reg_8_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_194_cse ) begin
      input_reg_8_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_3_lpi_2 <= 8'b00000000;
      psum_reg_7_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_195_cse ) begin
      input_reg_7_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_3_lpi_2 <= 8'b00000000;
      psum_reg_6_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_196_cse ) begin
      input_reg_6_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_3_lpi_2 <= 8'b00000000;
      psum_reg_5_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_197_cse ) begin
      input_reg_5_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_3_lpi_2 <= 8'b00000000;
      psum_reg_4_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_198_cse ) begin
      input_reg_4_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_3_lpi_2 <= 8'b00000000;
      psum_reg_3_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_199_cse ) begin
      input_reg_3_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_3_lpi_2 <= 8'b00000000;
      psum_reg_2_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_200_cse ) begin
      input_reg_2_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_3_lpi_2 <= 8'b00000000;
      psum_reg_1_3_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_201_cse ) begin
      input_reg_1_3_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_3_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_2_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_287 | or_dcpl_61)) ) begin
      input_reg_16_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_2_lpi_2 <= 8'b00000000;
      psum_reg_15_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_203_cse ) begin
      input_reg_15_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_2_lpi_2 <= 8'b00000000;
      psum_reg_14_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_204_cse ) begin
      input_reg_14_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_2_lpi_2 <= 8'b00000000;
      psum_reg_13_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_205_cse ) begin
      input_reg_13_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_2_lpi_2 <= 8'b00000000;
      psum_reg_12_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_206_cse ) begin
      input_reg_12_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_2_lpi_2 <= 8'b00000000;
      psum_reg_11_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_207_cse ) begin
      input_reg_11_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_2_lpi_2 <= 8'b00000000;
      psum_reg_10_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_208_cse ) begin
      input_reg_10_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_2_lpi_2 <= 8'b00000000;
      psum_reg_9_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_209_cse ) begin
      input_reg_9_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_2_lpi_2 <= 8'b00000000;
      psum_reg_8_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_210_cse ) begin
      input_reg_8_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_2_lpi_2 <= 8'b00000000;
      psum_reg_7_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_211_cse ) begin
      input_reg_7_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_2_lpi_2 <= 8'b00000000;
      psum_reg_6_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_212_cse ) begin
      input_reg_6_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_2_lpi_2 <= 8'b00000000;
      psum_reg_5_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_213_cse ) begin
      input_reg_5_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_2_lpi_2 <= 8'b00000000;
      psum_reg_4_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_214_cse ) begin
      input_reg_4_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_2_lpi_2 <= 8'b00000000;
      psum_reg_3_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_215_cse ) begin
      input_reg_3_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_2_lpi_2 <= 8'b00000000;
      psum_reg_2_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_216_cse ) begin
      input_reg_2_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_2_lpi_2 <= 8'b00000000;
      psum_reg_1_2_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_217_cse ) begin
      input_reg_1_2_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_2_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_1_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_269 | or_dcpl_38)) ) begin
      input_reg_16_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_15_1_lpi_2 <= 8'b00000000;
      psum_reg_15_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_219_cse ) begin
      input_reg_15_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_15_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_14_1_lpi_2 <= 8'b00000000;
      psum_reg_14_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_220_cse ) begin
      input_reg_14_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_14_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_13_1_lpi_2 <= 8'b00000000;
      psum_reg_13_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_221_cse ) begin
      input_reg_13_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_13_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_12_1_lpi_2 <= 8'b00000000;
      psum_reg_12_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_222_cse ) begin
      input_reg_12_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_12_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_11_1_lpi_2 <= 8'b00000000;
      psum_reg_11_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_223_cse ) begin
      input_reg_11_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_11_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_10_1_lpi_2 <= 8'b00000000;
      psum_reg_10_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_224_cse ) begin
      input_reg_10_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_10_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_9_1_lpi_2 <= 8'b00000000;
      psum_reg_9_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_225_cse ) begin
      input_reg_9_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_9_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_8_1_lpi_2 <= 8'b00000000;
      psum_reg_8_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_226_cse ) begin
      input_reg_8_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_8_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_7_1_lpi_2 <= 8'b00000000;
      psum_reg_7_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_227_cse ) begin
      input_reg_7_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_7_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_6_1_lpi_2 <= 8'b00000000;
      psum_reg_6_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_228_cse ) begin
      input_reg_6_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_6_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_5_1_lpi_2 <= 8'b00000000;
      psum_reg_5_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_229_cse ) begin
      input_reg_5_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_5_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_4_1_lpi_2 <= 8'b00000000;
      psum_reg_4_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_230_cse ) begin
      input_reg_4_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_4_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_3_1_lpi_2 <= 8'b00000000;
      psum_reg_3_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_231_cse ) begin
      input_reg_3_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_3_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_2_1_lpi_2 <= 8'b00000000;
      psum_reg_2_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_232_cse ) begin
      input_reg_2_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_2_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_1_1_lpi_2 <= 8'b00000000;
      psum_reg_1_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( input_reg_and_233_cse ) begin
      input_reg_1_1_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      psum_reg_1_1_lpi_2 <= pe_0_0_run_cmp_psum_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_12_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_287 | or_dcpl_41)) ) begin
      input_reg_16_12_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_11_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_29 | or_dcpl_95)) ) begin
      input_reg_16_11_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_10_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_151 | or_dcpl_61)) ) begin
      input_reg_16_10_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_15_14_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (and_dcpl_42 | and_dcpl_304) ) begin
      psum_reg_15_14_lpi_2 <= MUX_v_16_2_2(accum_fifo_2_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z,
          and_dcpl_304);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_13_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_287 | or_dcpl_38)) ) begin
      input_reg_16_13_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_15_15_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (and_dcpl_42 | and_dcpl_319) ) begin
      psum_reg_15_15_lpi_2 <= MUX_v_16_2_2(accum_fifo_11_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z,
          and_dcpl_319);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_14_lpi_2 <= 8'b00000000;
    end
    else if ( run_wen & (~(or_dcpl_29 | or_dcpl_97)) ) begin
      input_reg_16_14_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_15_16_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (and_dcpl_12 | and_dcpl_42 | psum_reg_15_16_lpi_2_mx0c2)
        ) begin
      psum_reg_15_16_lpi_2 <= MUX1HOT_v_16_3_2(output_fifo_2_rsci_output_rsc_z, accum_fifo_12_rsci_output_rsc_z,
          pe_0_0_run_cmp_psum_out_rsc_z, {and_dcpl_12 , and_dcpl_42 , psum_reg_15_16_lpi_2_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_reg_16_15_lpi_2 <= 8'b00000000;
      step_accum_fifo_input_15_asn_14_ncse_sva <= 16'b0000000000000000;
      step_accum_fifo_input_15_asn_13_ncse_sva <= 16'b0000000000000000;
      step_accum_fifo_input_15_asn_12_ncse_sva <= 16'b0000000000000000;
      step_accum_fifo_input_15_asn_9_ncse_sva <= 16'b0000000000000000;
    end
    else if ( input_reg_and_239_cse ) begin
      input_reg_16_15_lpi_2 <= pe_0_0_run_cmp_input_out_rsc_z;
      step_accum_fifo_input_15_asn_14_ncse_sva <= accum_fifo_15_rsci_output_rsc_z;
      step_accum_fifo_input_15_asn_13_ncse_sva <= accum_fifo_14_rsci_output_rsc_z;
      step_accum_fifo_input_15_asn_12_ncse_sva <= accum_fifo_13_rsci_output_rsc_z;
      step_accum_fifo_input_15_asn_9_ncse_sva <= accum_fifo_10_rsci_output_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_16_1_lpi_2 <= 16'b0000000000000000;
    end
    else if ( run_wen & (and_dcpl_362 | and_dcpl_12 | and_dcpl_42 | and_dcpl_74)
        ) begin
      psum_reg_16_1_lpi_2 <= MUX1HOT_v_16_4_2((step_acc_3_nl), output_fifo_11_rsci_output_rsc_z,
          accum_fifo_1_rsci_output_rsc_z, pe_0_0_run_cmp_psum_out_rsc_z, {and_dcpl_362
          , and_dcpl_12 , and_dcpl_42 , and_dcpl_74});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_slc_operator_16_false_acc_16_itm <= 1'b0;
      step_if_1_acc_cse_32 <= 1'b0;
    end
    else if ( operator_16_false_and_1_cse ) begin
      operator_16_false_slc_operator_16_false_acc_16_itm <= readslicef_17_1_16((operator_16_false_acc_nl));
      step_if_1_acc_cse_32 <= step_if_1_acc_itm_32_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_142_itm <= 8'b00000000;
    end
    else if ( run_wen & (ROW_asn_142_itm_mx0c0 | and_dcpl_8 | and_dcpl_55 | and_dcpl_74
        | and_dcpl_99 | and_dcpl_114 | and_dcpl_131 | and_dcpl_148 | and_dcpl_164
        | and_dcpl_179 | and_dcpl_197 | and_dcpl_214 | and_dcpl_230 | and_dcpl_245
        | and_dcpl_259 | and_dcpl_276 | and_dcpl_292 | and_dcpl_306) ) begin
      ROW_asn_142_itm <= MUX1HOT_v_8_18_2(({2'b00 , (operator_16_false_mux_1_nl)}),
          input_fifo_0_run_cmp_output_rsc_z, input_reg_1_1_lpi_2, input_reg_16_1_lpi_2,
          input_reg_15_2_lpi_2, input_reg_14_3_lpi_2, input_reg_13_4_lpi_2, input_reg_12_5_lpi_2,
          input_reg_11_6_lpi_2, input_reg_10_7_lpi_2, input_reg_9_8_lpi_2, input_reg_8_9_lpi_2,
          input_reg_7_10_lpi_2, input_reg_6_11_lpi_2, input_reg_5_12_lpi_2, input_reg_4_13_lpi_2,
          input_reg_3_14_lpi_2, input_reg_2_15_lpi_2, {ROW_asn_142_itm_mx0c0 , and_dcpl_8
          , and_dcpl_55 , and_dcpl_74 , and_dcpl_99 , and_dcpl_114 , and_dcpl_131
          , and_dcpl_148 , and_dcpl_164 , and_dcpl_179 , and_dcpl_197 , and_dcpl_214
          , and_dcpl_230 , and_dcpl_245 , and_dcpl_259 , and_dcpl_276 , and_dcpl_292
          , and_dcpl_306});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_143_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_56 | and_dcpl_75 | and_dcpl_100 |
        and_dcpl_115 | and_dcpl_132 | and_dcpl_149 | and_dcpl_165 | and_dcpl_180
        | and_dcpl_198 | and_dcpl_215 | and_dcpl_231 | and_dcpl_246 | and_dcpl_260
        | and_dcpl_277 | and_dcpl_293 | and_dcpl_307) ) begin
      ROW_asn_143_itm <= MUX1HOT_v_8_17_2(input_fifo_2_rsci_output_rsc_z, input_reg_2_1_lpi_2,
          input_reg_1_2_lpi_2, input_reg_16_2_lpi_2, input_reg_15_3_lpi_2, input_reg_14_4_lpi_2,
          input_reg_13_5_lpi_2, input_reg_12_6_lpi_2, input_reg_11_7_lpi_2, input_reg_10_8_lpi_2,
          input_reg_9_9_lpi_2, input_reg_8_10_lpi_2, input_reg_7_11_lpi_2, input_reg_6_12_lpi_2,
          input_reg_5_13_lpi_2, input_reg_4_14_lpi_2, input_reg_3_15_lpi_2, {and_dcpl_8
          , and_dcpl_56 , and_dcpl_75 , and_dcpl_100 , and_dcpl_115 , and_dcpl_132
          , and_dcpl_149 , and_dcpl_165 , and_dcpl_180 , and_dcpl_198 , and_dcpl_215
          , and_dcpl_231 , and_dcpl_246 , and_dcpl_260 , and_dcpl_277 , and_dcpl_293
          , and_dcpl_307});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_145_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_57 | and_dcpl_76 | and_dcpl_101 |
        and_dcpl_116 | and_dcpl_134 | and_dcpl_150 | and_dcpl_166 | and_dcpl_181
        | and_dcpl_199 | and_dcpl_216 | and_dcpl_232 | and_dcpl_247 | and_dcpl_261
        | and_dcpl_278 | and_dcpl_294 | and_dcpl_308) ) begin
      ROW_asn_145_itm <= MUX1HOT_v_8_17_2(input_fifo_3_rsci_output_rsc_z, input_reg_3_1_lpi_2,
          input_reg_2_2_lpi_2, input_reg_1_3_lpi_2, input_reg_16_3_lpi_2, input_reg_15_4_lpi_2,
          input_reg_14_5_lpi_2, input_reg_13_6_lpi_2, input_reg_12_7_lpi_2, input_reg_11_8_lpi_2,
          input_reg_10_9_lpi_2, input_reg_9_10_lpi_2, input_reg_8_11_lpi_2, input_reg_7_12_lpi_2,
          input_reg_6_13_lpi_2, input_reg_5_14_lpi_2, input_reg_4_15_lpi_2, {and_dcpl_8
          , and_dcpl_57 , and_dcpl_76 , and_dcpl_101 , and_dcpl_116 , and_dcpl_134
          , and_dcpl_150 , and_dcpl_166 , and_dcpl_181 , and_dcpl_199 , and_dcpl_216
          , and_dcpl_232 , and_dcpl_247 , and_dcpl_261 , and_dcpl_278 , and_dcpl_294
          , and_dcpl_308});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_147_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_58 | and_dcpl_77 | and_dcpl_102 |
        and_dcpl_117 | and_dcpl_135 | and_dcpl_152 | and_dcpl_167 | and_dcpl_182
        | and_dcpl_200 | and_dcpl_217 | and_dcpl_233 | and_dcpl_248 | and_dcpl_264
        | and_dcpl_279 | and_dcpl_295 | and_dcpl_309) ) begin
      ROW_asn_147_itm <= MUX1HOT_v_8_17_2(input_fifo_4_rsci_output_rsc_z, input_reg_4_1_lpi_2,
          input_reg_3_2_lpi_2, input_reg_2_3_lpi_2, input_reg_1_4_lpi_2, input_reg_16_4_lpi_2,
          input_reg_15_5_lpi_2, input_reg_14_6_lpi_2, input_reg_13_7_lpi_2, input_reg_12_8_lpi_2,
          input_reg_11_9_lpi_2, input_reg_10_10_lpi_2, input_reg_9_11_lpi_2, input_reg_8_12_lpi_2,
          input_reg_7_13_lpi_2, input_reg_6_14_lpi_2, input_reg_5_15_lpi_2, {and_dcpl_8
          , and_dcpl_58 , and_dcpl_77 , and_dcpl_102 , and_dcpl_117 , and_dcpl_135
          , and_dcpl_152 , and_dcpl_167 , and_dcpl_182 , and_dcpl_200 , and_dcpl_217
          , and_dcpl_233 , and_dcpl_248 , and_dcpl_264 , and_dcpl_279 , and_dcpl_295
          , and_dcpl_309});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_149_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_59 | and_dcpl_78 | and_dcpl_103 |
        and_dcpl_118 | and_dcpl_136 | and_dcpl_153 | and_dcpl_168 | and_dcpl_183
        | and_dcpl_201 | and_dcpl_218 | and_dcpl_234 | and_dcpl_249 | and_dcpl_265
        | and_dcpl_280 | and_dcpl_296 | and_dcpl_310) ) begin
      ROW_asn_149_itm <= MUX1HOT_v_8_17_2(input_fifo_5_rsci_output_rsc_z, input_reg_5_1_lpi_2,
          input_reg_4_2_lpi_2, input_reg_3_3_lpi_2, input_reg_2_4_lpi_2, input_reg_1_5_lpi_2,
          input_reg_16_5_lpi_2, input_reg_15_6_lpi_2, input_reg_14_7_lpi_2, input_reg_13_8_lpi_2,
          input_reg_12_9_lpi_2, input_reg_11_10_lpi_2, input_reg_10_11_lpi_2, input_reg_9_12_lpi_2,
          input_reg_8_13_lpi_2, input_reg_7_14_lpi_2, input_reg_6_15_lpi_2, {and_dcpl_8
          , and_dcpl_59 , and_dcpl_78 , and_dcpl_103 , and_dcpl_118 , and_dcpl_136
          , and_dcpl_153 , and_dcpl_168 , and_dcpl_183 , and_dcpl_201 , and_dcpl_218
          , and_dcpl_234 , and_dcpl_249 , and_dcpl_265 , and_dcpl_280 , and_dcpl_296
          , and_dcpl_310});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_151_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_60 | and_dcpl_79 | and_dcpl_104 |
        and_dcpl_119 | and_dcpl_137 | and_dcpl_154 | and_dcpl_169 | and_dcpl_184
        | and_dcpl_202 | and_dcpl_219 | and_dcpl_235 | and_dcpl_250 | and_dcpl_266
        | and_dcpl_282 | and_dcpl_297 | and_dcpl_311) ) begin
      ROW_asn_151_itm <= MUX1HOT_v_8_17_2(input_fifo_6_rsci_output_rsc_z, input_reg_6_1_lpi_2,
          input_reg_5_2_lpi_2, input_reg_4_3_lpi_2, input_reg_3_4_lpi_2, input_reg_2_5_lpi_2,
          input_reg_1_6_lpi_2, input_reg_16_6_lpi_2, input_reg_15_7_lpi_2, input_reg_14_8_lpi_2,
          input_reg_13_9_lpi_2, input_reg_12_10_lpi_2, input_reg_11_11_lpi_2, input_reg_10_12_lpi_2,
          input_reg_9_13_lpi_2, input_reg_8_14_lpi_2, input_reg_7_15_lpi_2, {and_dcpl_8
          , and_dcpl_60 , and_dcpl_79 , and_dcpl_104 , and_dcpl_119 , and_dcpl_137
          , and_dcpl_154 , and_dcpl_169 , and_dcpl_184 , and_dcpl_202 , and_dcpl_219
          , and_dcpl_235 , and_dcpl_250 , and_dcpl_266 , and_dcpl_282 , and_dcpl_297
          , and_dcpl_311});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_153_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_63 | and_dcpl_80 | and_dcpl_105 |
        and_dcpl_120 | and_dcpl_138 | and_dcpl_155 | and_dcpl_170 | and_dcpl_185
        | and_dcpl_204 | and_dcpl_220 | and_dcpl_236 | and_dcpl_251 | and_dcpl_267
        | and_dcpl_283 | and_dcpl_298 | and_dcpl_312) ) begin
      ROW_asn_153_itm <= MUX1HOT_v_8_17_2(input_fifo_7_rsci_output_rsc_z, input_reg_7_1_lpi_2,
          input_reg_6_2_lpi_2, input_reg_5_3_lpi_2, input_reg_4_4_lpi_2, input_reg_3_5_lpi_2,
          input_reg_2_6_lpi_2, input_reg_1_7_lpi_2, input_reg_16_7_lpi_2, input_reg_15_8_lpi_2,
          input_reg_14_9_lpi_2, input_reg_13_10_lpi_2, input_reg_12_11_lpi_2, input_reg_11_12_lpi_2,
          input_reg_10_13_lpi_2, input_reg_9_14_lpi_2, input_reg_8_15_lpi_2, {and_dcpl_8
          , and_dcpl_63 , and_dcpl_80 , and_dcpl_105 , and_dcpl_120 , and_dcpl_138
          , and_dcpl_155 , and_dcpl_170 , and_dcpl_185 , and_dcpl_204 , and_dcpl_220
          , and_dcpl_236 , and_dcpl_251 , and_dcpl_267 , and_dcpl_283 , and_dcpl_298
          , and_dcpl_312});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_155_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_64 | and_dcpl_83 | and_dcpl_106 |
        and_dcpl_121 | and_dcpl_139 | and_dcpl_156 | and_dcpl_171 | and_dcpl_186
        | and_dcpl_205 | and_dcpl_222 | and_dcpl_237 | and_dcpl_252 | and_dcpl_268
        | and_dcpl_284 | and_dcpl_299 | and_dcpl_313) ) begin
      ROW_asn_155_itm <= MUX1HOT_v_8_17_2(input_fifo_8_rsci_output_rsc_z, input_reg_8_1_lpi_2,
          input_reg_7_2_lpi_2, input_reg_6_3_lpi_2, input_reg_5_4_lpi_2, input_reg_4_5_lpi_2,
          input_reg_3_6_lpi_2, input_reg_2_7_lpi_2, input_reg_1_8_lpi_2, input_reg_16_8_lpi_2,
          input_reg_15_9_lpi_2, input_reg_14_10_lpi_2, input_reg_13_11_lpi_2, input_reg_12_12_lpi_2,
          input_reg_11_13_lpi_2, input_reg_10_14_lpi_2, input_reg_9_15_lpi_2, {and_dcpl_8
          , and_dcpl_64 , and_dcpl_83 , and_dcpl_106 , and_dcpl_121 , and_dcpl_139
          , and_dcpl_156 , and_dcpl_171 , and_dcpl_186 , and_dcpl_205 , and_dcpl_222
          , and_dcpl_237 , and_dcpl_252 , and_dcpl_268 , and_dcpl_284 , and_dcpl_299
          , and_dcpl_313});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_157_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_65 | and_dcpl_85 | and_dcpl_107 |
        and_dcpl_122 | and_dcpl_140 | and_dcpl_157 | and_dcpl_172 | and_dcpl_187
        | and_dcpl_206 | and_dcpl_223 | and_dcpl_238 | and_dcpl_253 | and_dcpl_269
        | and_dcpl_285 | and_dcpl_300 | and_dcpl_314) ) begin
      ROW_asn_157_itm <= MUX1HOT_v_8_17_2(input_fifo_9_rsci_output_rsc_z, input_reg_9_1_lpi_2,
          input_reg_8_2_lpi_2, input_reg_7_3_lpi_2, input_reg_6_4_lpi_2, input_reg_5_5_lpi_2,
          input_reg_4_6_lpi_2, input_reg_3_7_lpi_2, input_reg_2_8_lpi_2, input_reg_1_9_lpi_2,
          input_reg_16_9_lpi_2, input_reg_15_10_lpi_2, input_reg_14_11_lpi_2, input_reg_13_12_lpi_2,
          input_reg_12_13_lpi_2, input_reg_11_14_lpi_2, input_reg_10_15_lpi_2, {and_dcpl_8
          , and_dcpl_65 , and_dcpl_85 , and_dcpl_107 , and_dcpl_122 , and_dcpl_140
          , and_dcpl_157 , and_dcpl_172 , and_dcpl_187 , and_dcpl_206 , and_dcpl_223
          , and_dcpl_238 , and_dcpl_253 , and_dcpl_269 , and_dcpl_285 , and_dcpl_300
          , and_dcpl_314});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_159_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_66 | and_dcpl_87 | and_dcpl_108 |
        and_dcpl_125 | and_dcpl_141 | and_dcpl_158 | and_dcpl_173 | and_dcpl_188
        | and_dcpl_207 | and_dcpl_224 | and_dcpl_240 | and_dcpl_254 | and_dcpl_270
        | and_dcpl_286 | and_dcpl_301 | and_dcpl_315) ) begin
      ROW_asn_159_itm <= MUX1HOT_v_8_17_2(input_fifo_10_rsci_output_rsc_z, input_reg_10_1_lpi_2,
          input_reg_9_2_lpi_2, input_reg_8_3_lpi_2, input_reg_7_4_lpi_2, input_reg_6_5_lpi_2,
          input_reg_5_6_lpi_2, input_reg_4_7_lpi_2, input_reg_3_8_lpi_2, input_reg_2_9_lpi_2,
          input_reg_1_10_lpi_2, input_reg_1_11_lpi_2, input_reg_15_11_lpi_2, input_reg_14_12_lpi_2,
          input_reg_13_13_lpi_2, input_reg_12_14_lpi_2, input_reg_11_15_lpi_2, {and_dcpl_8
          , and_dcpl_66 , and_dcpl_87 , and_dcpl_108 , and_dcpl_125 , and_dcpl_141
          , and_dcpl_158 , and_dcpl_173 , and_dcpl_188 , and_dcpl_207 , and_dcpl_224
          , and_dcpl_240 , and_dcpl_254 , and_dcpl_270 , and_dcpl_286 , and_dcpl_301
          , and_dcpl_315});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_161_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_67 | and_dcpl_89 | and_dcpl_109 |
        and_dcpl_126 | and_dcpl_143 | and_dcpl_159 | and_dcpl_174 | and_dcpl_189
        | and_dcpl_208 | and_dcpl_225 | and_dcpl_241 | and_dcpl_255 | and_dcpl_271
        | and_dcpl_287 | and_dcpl_302 | and_dcpl_316) ) begin
      ROW_asn_161_itm <= MUX1HOT_v_8_17_2(input_fifo_11_rsci_output_rsc_z, input_reg_11_1_lpi_2,
          input_reg_10_2_lpi_2, input_reg_9_3_lpi_2, input_reg_8_4_lpi_2, input_reg_7_5_lpi_2,
          input_reg_6_6_lpi_2, input_reg_5_7_lpi_2, input_reg_4_8_lpi_2, input_reg_3_9_lpi_2,
          input_reg_2_10_lpi_2, input_reg_2_11_lpi_2, input_reg_1_12_lpi_2, input_reg_15_12_lpi_2,
          input_reg_14_13_lpi_2, input_reg_13_14_lpi_2, input_reg_12_15_lpi_2, {and_dcpl_8
          , and_dcpl_67 , and_dcpl_89 , and_dcpl_109 , and_dcpl_126 , and_dcpl_143
          , and_dcpl_159 , and_dcpl_174 , and_dcpl_189 , and_dcpl_208 , and_dcpl_225
          , and_dcpl_241 , and_dcpl_255 , and_dcpl_271 , and_dcpl_287 , and_dcpl_302
          , and_dcpl_316});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_163_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_68 | and_dcpl_92 | and_dcpl_110 |
        and_dcpl_127 | and_dcpl_144 | and_dcpl_160 | and_dcpl_175 | and_dcpl_190
        | and_dcpl_209 | and_dcpl_226 | and_dcpl_242 | and_dcpl_256 | and_dcpl_273
        | and_dcpl_288 | and_dcpl_303 | and_dcpl_317) ) begin
      ROW_asn_163_itm <= MUX1HOT_v_8_17_2(input_fifo_12_rsci_output_rsc_z, input_reg_12_1_lpi_2,
          input_reg_11_2_lpi_2, input_reg_10_3_lpi_2, input_reg_9_4_lpi_2, input_reg_8_5_lpi_2,
          input_reg_7_6_lpi_2, input_reg_6_7_lpi_2, input_reg_5_8_lpi_2, input_reg_4_9_lpi_2,
          input_reg_3_10_lpi_2, input_reg_3_11_lpi_2, input_reg_2_12_lpi_2, input_reg_1_13_lpi_2,
          input_reg_15_13_lpi_2, input_reg_14_14_lpi_2, input_reg_13_15_lpi_2, {and_dcpl_8
          , and_dcpl_68 , and_dcpl_92 , and_dcpl_110 , and_dcpl_127 , and_dcpl_144
          , and_dcpl_160 , and_dcpl_175 , and_dcpl_190 , and_dcpl_209 , and_dcpl_226
          , and_dcpl_242 , and_dcpl_256 , and_dcpl_273 , and_dcpl_288 , and_dcpl_303
          , and_dcpl_317});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_165_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_69 | and_dcpl_94 | and_dcpl_111 |
        and_dcpl_128 | and_dcpl_145 | and_dcpl_161 | and_dcpl_176 | and_dcpl_191
        | and_dcpl_210 | and_dcpl_227 | and_dcpl_243 | and_dcpl_257 | and_dcpl_274
        | and_dcpl_289 | and_dcpl_304 | and_dcpl_318) ) begin
      ROW_asn_165_itm <= MUX1HOT_v_8_17_2(input_fifo_13_rsci_output_rsc_z, input_reg_13_1_lpi_2,
          input_reg_12_2_lpi_2, input_reg_11_3_lpi_2, input_reg_10_4_lpi_2, input_reg_9_5_lpi_2,
          input_reg_8_6_lpi_2, input_reg_7_7_lpi_2, input_reg_6_8_lpi_2, input_reg_5_9_lpi_2,
          input_reg_4_10_lpi_2, input_reg_4_11_lpi_2, input_reg_3_12_lpi_2, input_reg_2_13_lpi_2,
          input_reg_1_14_lpi_2, input_reg_15_14_lpi_2, input_reg_14_15_lpi_2, {and_dcpl_8
          , and_dcpl_69 , and_dcpl_94 , and_dcpl_111 , and_dcpl_128 , and_dcpl_145
          , and_dcpl_161 , and_dcpl_176 , and_dcpl_191 , and_dcpl_210 , and_dcpl_227
          , and_dcpl_243 , and_dcpl_257 , and_dcpl_274 , and_dcpl_289 , and_dcpl_304
          , and_dcpl_318});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_167_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_70 | and_dcpl_96 | and_dcpl_112 |
        and_dcpl_129 | and_dcpl_146 | and_dcpl_162 | and_dcpl_177 | and_dcpl_195
        | and_dcpl_211 | and_dcpl_228 | and_dcpl_244 | and_dcpl_258 | and_dcpl_275
        | and_dcpl_291 | and_dcpl_305 | and_dcpl_319) ) begin
      ROW_asn_167_itm <= MUX1HOT_v_8_17_2(input_fifo_14_rsci_output_rsc_z, input_reg_14_1_lpi_2,
          input_reg_13_2_lpi_2, input_reg_12_3_lpi_2, input_reg_11_4_lpi_2, input_reg_10_5_lpi_2,
          input_reg_9_6_lpi_2, input_reg_8_7_lpi_2, input_reg_7_8_lpi_2, input_reg_6_9_lpi_2,
          input_reg_5_10_lpi_2, input_reg_5_11_lpi_2, input_reg_4_12_lpi_2, input_reg_3_13_lpi_2,
          input_reg_2_14_lpi_2, input_reg_1_15_lpi_2, input_reg_15_15_lpi_2, {and_dcpl_8
          , and_dcpl_70 , and_dcpl_96 , and_dcpl_112 , and_dcpl_129 , and_dcpl_146
          , and_dcpl_162 , and_dcpl_177 , and_dcpl_195 , and_dcpl_211 , and_dcpl_228
          , and_dcpl_244 , and_dcpl_258 , and_dcpl_275 , and_dcpl_291 , and_dcpl_305
          , and_dcpl_319});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROW_asn_169_itm <= 8'b00000000;
    end
    else if ( run_wen & (and_dcpl_8 | and_dcpl_73 | and_dcpl_98 | and_dcpl_113 |
        and_dcpl_130 | and_dcpl_147 | and_dcpl_163 | and_dcpl_178 | and_dcpl_196
        | and_dcpl_213 | and_dcpl_229) ) begin
      ROW_asn_169_itm <= MUX1HOT_v_8_11_2(input_fifo_15_rsci_output_rsc_z, input_reg_15_1_lpi_2,
          input_reg_14_2_lpi_2, input_reg_13_3_lpi_2, input_reg_12_4_lpi_2, input_reg_11_5_lpi_2,
          input_reg_10_6_lpi_2, input_reg_9_7_lpi_2, input_reg_8_8_lpi_2, input_reg_7_9_lpi_2,
          input_reg_6_10_lpi_2, {and_dcpl_8 , and_dcpl_73 , and_dcpl_98 , and_dcpl_113
          , and_dcpl_130 , and_dcpl_147 , and_dcpl_163 , and_dcpl_178 , and_dcpl_196
          , and_dcpl_213 , and_dcpl_229});
    end
  end
  assign or_337_nl = (~((fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[0]) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_307_nl = MUX_s_1_2_2(mux_306_cse, (or_337_nl), fsm_output[2]);
  assign and_441_nl = and_dcpl_7 & and_dcpl_360 & (fsm_output[0]) & step_if_1_acc_cse_32;
  assign or_35_nl = (~((fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_312_nl = MUX_s_1_2_2(mux_306_cse, (or_35_nl), fsm_output[2]);
  assign or_924_nl = (fsm_output[7:2]!=6'b000001);
  assign or_920_nl = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[7]);
  assign mux_313_nl = MUX_s_1_2_2((or_924_nl), (or_920_nl), fsm_output[1]);
  assign mux_314_nl = MUX_s_1_2_2((mux_313_nl), nor_150_cse, fsm_output[8]);
  assign psum_reg_or_4_nl = ((~ operator_32_false_acc_itm_31_1) & and_443_m1c) |
      (mux_314_nl);
  assign psum_reg_and_242_nl = operator_32_false_acc_itm_31_1 & and_443_m1c;
  assign mux_315_nl = MUX_s_1_2_2(nor_133_cse, (fsm_output[8]), or_645_cse);
  assign or_664_nl = (~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[0]) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_316_nl = MUX_s_1_2_2((mux_315_nl), (or_664_nl), fsm_output[3]);
  assign or_662_nl = (~((fsm_output[7:3]!=5'b00000))) | (fsm_output[8]);
  assign mux_317_nl = MUX_s_1_2_2((mux_316_nl), (or_662_nl), fsm_output[2]);
  assign or_669_nl = (fsm_output[2]) | nor_133_cse;
  assign mux_318_nl = MUX_s_1_2_2((or_669_nl), (fsm_output[8]), or_338_cse);
  assign mux_323_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), or_52_cse);
  assign or_51_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[0]) | (fsm_output[8]);
  assign mux_51_nl = MUX_s_1_2_2((fsm_output[8]), (or_51_nl), and_cse);
  assign mux_324_nl = MUX_s_1_2_2((mux_323_nl), (mux_51_nl), fsm_output[5]);
  assign or_676_nl = (fsm_output[6]) | (mux_324_nl);
  assign nand_nl = ~((fsm_output[3]) & nor_174_cse);
  assign mux_49_nl = MUX_s_1_2_2((nand_nl), (fsm_output[8]), fsm_output[4]);
  assign nand_1_nl = ~((fsm_output[5]) & (~ (mux_49_nl)));
  assign mux_50_nl = MUX_s_1_2_2((nand_1_nl), (fsm_output[8]), fsm_output[6]);
  assign mux_325_nl = MUX_s_1_2_2((or_676_nl), (mux_50_nl), fsm_output[7]);
  assign mux_327_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), or_58_cse);
  assign or_57_nl = (~((~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[2])
      | (~ (fsm_output[0])) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_328_nl = MUX_s_1_2_2((mux_327_nl), (or_57_nl), fsm_output[3]);
  assign mux_329_nl = MUX_s_1_2_2((mux_328_nl), (fsm_output[8]), or_55_cse);
  assign mux_331_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), fsm_output[7]);
  assign or_685_nl = (~((~ (fsm_output[7])) | (fsm_output[2]) | (~ (fsm_output[0]))
      | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_332_nl = MUX_s_1_2_2((mux_331_nl), (or_685_nl), fsm_output[3]);
  assign or_67_nl = (fsm_output[6:4]!=3'b000);
  assign mux_333_nl = MUX_s_1_2_2((mux_332_nl), (fsm_output[8]), or_67_nl);
  assign and_461_nl = (fsm_output[6:3]==4'b1111);
  assign nor_117_nl = ~((fsm_output[6:3]!=4'b0000));
  assign mux_334_nl = MUX_s_1_2_2((and_461_nl), (nor_117_nl), fsm_output[1]);
  assign nand_28_nl = ~((fsm_output[0]) & (mux_334_nl));
  assign or_689_nl = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[6]);
  assign mux_335_nl = MUX_s_1_2_2((nand_28_nl), (or_689_nl), fsm_output[2]);
  assign or_918_nl = (fsm_output[7]) | (mux_335_nl);
  assign mux_336_nl = MUX_s_1_2_2((or_918_nl), nor_150_cse, fsm_output[8]);
  assign mux_338_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), or_55_cse);
  assign or_76_nl = (~((~ (fsm_output[5])) | (~ (fsm_output[6])) | (fsm_output[2])
      | (~ (fsm_output[0])) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_339_nl = MUX_s_1_2_2((mux_338_nl), (or_76_nl), fsm_output[3]);
  assign mux_340_nl = MUX_s_1_2_2((mux_339_nl), (fsm_output[8]), or_58_cse);
  assign or_83_nl = (fsm_output[4]) | (fsm_output[6]);
  assign mux_342_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), or_83_nl);
  assign or_82_nl = (~((~ (fsm_output[4])) | (~ (fsm_output[6])) | (fsm_output[2])
      | (~ (fsm_output[0])) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_343_nl = MUX_s_1_2_2((mux_342_nl), (or_82_nl), fsm_output[3]);
  assign or_80_nl = (fsm_output[5]) | (fsm_output[7]);
  assign mux_344_nl = MUX_s_1_2_2((mux_343_nl), (fsm_output[8]), or_80_nl);
  assign mux_346_nl = MUX_s_1_2_2(mux_322_cse, (fsm_output[8]), fsm_output[6]);
  assign or_706_nl = (~((~ (fsm_output[6])) | (fsm_output[2]) | (~ (fsm_output[0]))
      | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_347_nl = MUX_s_1_2_2((mux_346_nl), (or_706_nl), fsm_output[3]);
  assign or_92_nl = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[7]);
  assign mux_348_nl = MUX_s_1_2_2((mux_347_nl), (fsm_output[8]), or_92_nl);
  assign or_714_nl = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[2]) | nor_133_cse;
  assign nand_2_nl = ~((fsm_output[5:4]==2'b11) & nor_174_cse);
  assign mux_349_nl = MUX_s_1_2_2((or_714_nl), (nand_2_nl), fsm_output[3]);
  assign mux_350_nl = MUX_s_1_2_2((mux_349_nl), (fsm_output[8]), or_94_cse);
  assign mux_381_nl = MUX_s_1_2_2(or_tmp_126, or_tmp_127, fsm_output[1]);
  assign mux_382_nl = MUX_s_1_2_2((mux_381_nl), mux_tmp_337, fsm_output[0]);
  assign and_451_nl = (~ (mux_382_nl)) & (~ (fsm_output[7])) & and_dcpl_445;
  assign step_input_fifo_input_15_mux_nl = MUX_v_8_2_2(input_fifo_1_rsci_output_rsc_z,
      (psum_reg_16_2_lpi_2[7:0]), and_451_nl);
  assign or_720_nl = (fsm_output[5]) | nor_133_cse;
  assign or_104_nl = (~ (fsm_output[5])) | (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_351_nl = MUX_s_1_2_2((or_720_nl), (or_104_nl), fsm_output[3]);
  assign or_103_nl = (~ (fsm_output[3])) | (~ (fsm_output[5])) | (fsm_output[8]);
  assign mux_352_nl = MUX_s_1_2_2((mux_351_nl), (or_103_nl), fsm_output[2]);
  assign or_102_nl = (~ (fsm_output[5])) | (fsm_output[8]);
  assign mux_353_nl = MUX_s_1_2_2((mux_352_nl), (or_102_nl), fsm_output[4]);
  assign mux_354_nl = MUX_s_1_2_2((mux_353_nl), (fsm_output[8]), or_94_cse);
  assign and_447_nl = (~ mux_tmp_337) & (~ (fsm_output[7])) & and_dcpl_445;
  assign and_460_nl = or_645_cse & (fsm_output[8]);
  assign nor_168_nl = ~((~ (fsm_output[1])) | (fsm_output[8]));
  assign mux_360_nl = MUX_s_1_2_2((nor_168_nl), (fsm_output[8]), or_645_cse);
  assign mux_361_nl = MUX_s_1_2_2((and_460_nl), (mux_360_nl), fsm_output[0]);
  assign or_729_nl = (~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_362_nl = MUX_s_1_2_2((mux_361_nl), (or_729_nl), fsm_output[2]);
  assign or_727_nl = (~((fsm_output[2]) | (~ (fsm_output[0])) | (fsm_output[4]) |
      (fsm_output[5]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[1]))) | (fsm_output[8]);
  assign mux_363_nl = MUX_s_1_2_2((mux_362_nl), (or_727_nl), fsm_output[3]);
  assign step_step_mux_nl = MUX_v_16_2_2(step_step_sva, psum_reg_16_1_lpi_2, and_dcpl_12);
  assign step_step_not_nl = ~ mux_tmp_345;
  assign nl_step_acc_3_nl = step_step_sva + 16'b0000000000000001;
  assign step_acc_3_nl = nl_step_acc_3_nl[15:0];
  assign nl_operator_16_false_acc_nl = conv_u2s_16_17(step_step_sva) + 17'b11111111111100001;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[16:0];
  assign nl_step_if_3_for_1_operator_16_false_acc_nl = (step_step_sva[5:0]) + 6'b100001;
  assign step_if_3_for_1_operator_16_false_acc_nl = nl_step_if_3_for_1_operator_16_false_acc_nl[5:0];
  assign operator_16_false_mux_1_nl = MUX_v_6_2_2((step_if_3_for_1_operator_16_false_acc_nl),
      (ROW_asn_142_itm[5:0]), and_dcpl_12);

  function automatic [15:0] MUX1HOT_v_16_253_2;
    input [15:0] input_252;
    input [15:0] input_251;
    input [15:0] input_250;
    input [15:0] input_249;
    input [15:0] input_248;
    input [15:0] input_247;
    input [15:0] input_246;
    input [15:0] input_245;
    input [15:0] input_244;
    input [15:0] input_243;
    input [15:0] input_242;
    input [15:0] input_241;
    input [15:0] input_240;
    input [15:0] input_239;
    input [15:0] input_238;
    input [15:0] input_237;
    input [15:0] input_236;
    input [15:0] input_235;
    input [15:0] input_234;
    input [15:0] input_233;
    input [15:0] input_232;
    input [15:0] input_231;
    input [15:0] input_230;
    input [15:0] input_229;
    input [15:0] input_228;
    input [15:0] input_227;
    input [15:0] input_226;
    input [15:0] input_225;
    input [15:0] input_224;
    input [15:0] input_223;
    input [15:0] input_222;
    input [15:0] input_221;
    input [15:0] input_220;
    input [15:0] input_219;
    input [15:0] input_218;
    input [15:0] input_217;
    input [15:0] input_216;
    input [15:0] input_215;
    input [15:0] input_214;
    input [15:0] input_213;
    input [15:0] input_212;
    input [15:0] input_211;
    input [15:0] input_210;
    input [15:0] input_209;
    input [15:0] input_208;
    input [15:0] input_207;
    input [15:0] input_206;
    input [15:0] input_205;
    input [15:0] input_204;
    input [15:0] input_203;
    input [15:0] input_202;
    input [15:0] input_201;
    input [15:0] input_200;
    input [15:0] input_199;
    input [15:0] input_198;
    input [15:0] input_197;
    input [15:0] input_196;
    input [15:0] input_195;
    input [15:0] input_194;
    input [15:0] input_193;
    input [15:0] input_192;
    input [15:0] input_191;
    input [15:0] input_190;
    input [15:0] input_189;
    input [15:0] input_188;
    input [15:0] input_187;
    input [15:0] input_186;
    input [15:0] input_185;
    input [15:0] input_184;
    input [15:0] input_183;
    input [15:0] input_182;
    input [15:0] input_181;
    input [15:0] input_180;
    input [15:0] input_179;
    input [15:0] input_178;
    input [15:0] input_177;
    input [15:0] input_176;
    input [15:0] input_175;
    input [15:0] input_174;
    input [15:0] input_173;
    input [15:0] input_172;
    input [15:0] input_171;
    input [15:0] input_170;
    input [15:0] input_169;
    input [15:0] input_168;
    input [15:0] input_167;
    input [15:0] input_166;
    input [15:0] input_165;
    input [15:0] input_164;
    input [15:0] input_163;
    input [15:0] input_162;
    input [15:0] input_161;
    input [15:0] input_160;
    input [15:0] input_159;
    input [15:0] input_158;
    input [15:0] input_157;
    input [15:0] input_156;
    input [15:0] input_155;
    input [15:0] input_154;
    input [15:0] input_153;
    input [15:0] input_152;
    input [15:0] input_151;
    input [15:0] input_150;
    input [15:0] input_149;
    input [15:0] input_148;
    input [15:0] input_147;
    input [15:0] input_146;
    input [15:0] input_145;
    input [15:0] input_144;
    input [15:0] input_143;
    input [15:0] input_142;
    input [15:0] input_141;
    input [15:0] input_140;
    input [15:0] input_139;
    input [15:0] input_138;
    input [15:0] input_137;
    input [15:0] input_136;
    input [15:0] input_135;
    input [15:0] input_134;
    input [15:0] input_133;
    input [15:0] input_132;
    input [15:0] input_131;
    input [15:0] input_130;
    input [15:0] input_129;
    input [15:0] input_128;
    input [15:0] input_127;
    input [15:0] input_126;
    input [15:0] input_125;
    input [15:0] input_124;
    input [15:0] input_123;
    input [15:0] input_122;
    input [15:0] input_121;
    input [15:0] input_120;
    input [15:0] input_119;
    input [15:0] input_118;
    input [15:0] input_117;
    input [15:0] input_116;
    input [15:0] input_115;
    input [15:0] input_114;
    input [15:0] input_113;
    input [15:0] input_112;
    input [15:0] input_111;
    input [15:0] input_110;
    input [15:0] input_109;
    input [15:0] input_108;
    input [15:0] input_107;
    input [15:0] input_106;
    input [15:0] input_105;
    input [15:0] input_104;
    input [15:0] input_103;
    input [15:0] input_102;
    input [15:0] input_101;
    input [15:0] input_100;
    input [15:0] input_99;
    input [15:0] input_98;
    input [15:0] input_97;
    input [15:0] input_96;
    input [15:0] input_95;
    input [15:0] input_94;
    input [15:0] input_93;
    input [15:0] input_92;
    input [15:0] input_91;
    input [15:0] input_90;
    input [15:0] input_89;
    input [15:0] input_88;
    input [15:0] input_87;
    input [15:0] input_86;
    input [15:0] input_85;
    input [15:0] input_84;
    input [15:0] input_83;
    input [15:0] input_82;
    input [15:0] input_81;
    input [15:0] input_80;
    input [15:0] input_79;
    input [15:0] input_78;
    input [15:0] input_77;
    input [15:0] input_76;
    input [15:0] input_75;
    input [15:0] input_74;
    input [15:0] input_73;
    input [15:0] input_72;
    input [15:0] input_71;
    input [15:0] input_70;
    input [15:0] input_69;
    input [15:0] input_68;
    input [15:0] input_67;
    input [15:0] input_66;
    input [15:0] input_65;
    input [15:0] input_64;
    input [15:0] input_63;
    input [15:0] input_62;
    input [15:0] input_61;
    input [15:0] input_60;
    input [15:0] input_59;
    input [15:0] input_58;
    input [15:0] input_57;
    input [15:0] input_56;
    input [15:0] input_55;
    input [15:0] input_54;
    input [15:0] input_53;
    input [15:0] input_52;
    input [15:0] input_51;
    input [15:0] input_50;
    input [15:0] input_49;
    input [15:0] input_48;
    input [15:0] input_47;
    input [15:0] input_46;
    input [15:0] input_45;
    input [15:0] input_44;
    input [15:0] input_43;
    input [15:0] input_42;
    input [15:0] input_41;
    input [15:0] input_40;
    input [15:0] input_39;
    input [15:0] input_38;
    input [15:0] input_37;
    input [15:0] input_36;
    input [15:0] input_35;
    input [15:0] input_34;
    input [15:0] input_33;
    input [15:0] input_32;
    input [15:0] input_31;
    input [15:0] input_30;
    input [15:0] input_29;
    input [15:0] input_28;
    input [15:0] input_27;
    input [15:0] input_26;
    input [15:0] input_25;
    input [15:0] input_24;
    input [15:0] input_23;
    input [15:0] input_22;
    input [15:0] input_21;
    input [15:0] input_20;
    input [15:0] input_19;
    input [15:0] input_18;
    input [15:0] input_17;
    input [15:0] input_16;
    input [15:0] input_15;
    input [15:0] input_14;
    input [15:0] input_13;
    input [15:0] input_12;
    input [15:0] input_11;
    input [15:0] input_10;
    input [15:0] input_9;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [252:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    result = result | ( input_6 & {16{sel[6]}});
    result = result | ( input_7 & {16{sel[7]}});
    result = result | ( input_8 & {16{sel[8]}});
    result = result | ( input_9 & {16{sel[9]}});
    result = result | ( input_10 & {16{sel[10]}});
    result = result | ( input_11 & {16{sel[11]}});
    result = result | ( input_12 & {16{sel[12]}});
    result = result | ( input_13 & {16{sel[13]}});
    result = result | ( input_14 & {16{sel[14]}});
    result = result | ( input_15 & {16{sel[15]}});
    result = result | ( input_16 & {16{sel[16]}});
    result = result | ( input_17 & {16{sel[17]}});
    result = result | ( input_18 & {16{sel[18]}});
    result = result | ( input_19 & {16{sel[19]}});
    result = result | ( input_20 & {16{sel[20]}});
    result = result | ( input_21 & {16{sel[21]}});
    result = result | ( input_22 & {16{sel[22]}});
    result = result | ( input_23 & {16{sel[23]}});
    result = result | ( input_24 & {16{sel[24]}});
    result = result | ( input_25 & {16{sel[25]}});
    result = result | ( input_26 & {16{sel[26]}});
    result = result | ( input_27 & {16{sel[27]}});
    result = result | ( input_28 & {16{sel[28]}});
    result = result | ( input_29 & {16{sel[29]}});
    result = result | ( input_30 & {16{sel[30]}});
    result = result | ( input_31 & {16{sel[31]}});
    result = result | ( input_32 & {16{sel[32]}});
    result = result | ( input_33 & {16{sel[33]}});
    result = result | ( input_34 & {16{sel[34]}});
    result = result | ( input_35 & {16{sel[35]}});
    result = result | ( input_36 & {16{sel[36]}});
    result = result | ( input_37 & {16{sel[37]}});
    result = result | ( input_38 & {16{sel[38]}});
    result = result | ( input_39 & {16{sel[39]}});
    result = result | ( input_40 & {16{sel[40]}});
    result = result | ( input_41 & {16{sel[41]}});
    result = result | ( input_42 & {16{sel[42]}});
    result = result | ( input_43 & {16{sel[43]}});
    result = result | ( input_44 & {16{sel[44]}});
    result = result | ( input_45 & {16{sel[45]}});
    result = result | ( input_46 & {16{sel[46]}});
    result = result | ( input_47 & {16{sel[47]}});
    result = result | ( input_48 & {16{sel[48]}});
    result = result | ( input_49 & {16{sel[49]}});
    result = result | ( input_50 & {16{sel[50]}});
    result = result | ( input_51 & {16{sel[51]}});
    result = result | ( input_52 & {16{sel[52]}});
    result = result | ( input_53 & {16{sel[53]}});
    result = result | ( input_54 & {16{sel[54]}});
    result = result | ( input_55 & {16{sel[55]}});
    result = result | ( input_56 & {16{sel[56]}});
    result = result | ( input_57 & {16{sel[57]}});
    result = result | ( input_58 & {16{sel[58]}});
    result = result | ( input_59 & {16{sel[59]}});
    result = result | ( input_60 & {16{sel[60]}});
    result = result | ( input_61 & {16{sel[61]}});
    result = result | ( input_62 & {16{sel[62]}});
    result = result | ( input_63 & {16{sel[63]}});
    result = result | ( input_64 & {16{sel[64]}});
    result = result | ( input_65 & {16{sel[65]}});
    result = result | ( input_66 & {16{sel[66]}});
    result = result | ( input_67 & {16{sel[67]}});
    result = result | ( input_68 & {16{sel[68]}});
    result = result | ( input_69 & {16{sel[69]}});
    result = result | ( input_70 & {16{sel[70]}});
    result = result | ( input_71 & {16{sel[71]}});
    result = result | ( input_72 & {16{sel[72]}});
    result = result | ( input_73 & {16{sel[73]}});
    result = result | ( input_74 & {16{sel[74]}});
    result = result | ( input_75 & {16{sel[75]}});
    result = result | ( input_76 & {16{sel[76]}});
    result = result | ( input_77 & {16{sel[77]}});
    result = result | ( input_78 & {16{sel[78]}});
    result = result | ( input_79 & {16{sel[79]}});
    result = result | ( input_80 & {16{sel[80]}});
    result = result | ( input_81 & {16{sel[81]}});
    result = result | ( input_82 & {16{sel[82]}});
    result = result | ( input_83 & {16{sel[83]}});
    result = result | ( input_84 & {16{sel[84]}});
    result = result | ( input_85 & {16{sel[85]}});
    result = result | ( input_86 & {16{sel[86]}});
    result = result | ( input_87 & {16{sel[87]}});
    result = result | ( input_88 & {16{sel[88]}});
    result = result | ( input_89 & {16{sel[89]}});
    result = result | ( input_90 & {16{sel[90]}});
    result = result | ( input_91 & {16{sel[91]}});
    result = result | ( input_92 & {16{sel[92]}});
    result = result | ( input_93 & {16{sel[93]}});
    result = result | ( input_94 & {16{sel[94]}});
    result = result | ( input_95 & {16{sel[95]}});
    result = result | ( input_96 & {16{sel[96]}});
    result = result | ( input_97 & {16{sel[97]}});
    result = result | ( input_98 & {16{sel[98]}});
    result = result | ( input_99 & {16{sel[99]}});
    result = result | ( input_100 & {16{sel[100]}});
    result = result | ( input_101 & {16{sel[101]}});
    result = result | ( input_102 & {16{sel[102]}});
    result = result | ( input_103 & {16{sel[103]}});
    result = result | ( input_104 & {16{sel[104]}});
    result = result | ( input_105 & {16{sel[105]}});
    result = result | ( input_106 & {16{sel[106]}});
    result = result | ( input_107 & {16{sel[107]}});
    result = result | ( input_108 & {16{sel[108]}});
    result = result | ( input_109 & {16{sel[109]}});
    result = result | ( input_110 & {16{sel[110]}});
    result = result | ( input_111 & {16{sel[111]}});
    result = result | ( input_112 & {16{sel[112]}});
    result = result | ( input_113 & {16{sel[113]}});
    result = result | ( input_114 & {16{sel[114]}});
    result = result | ( input_115 & {16{sel[115]}});
    result = result | ( input_116 & {16{sel[116]}});
    result = result | ( input_117 & {16{sel[117]}});
    result = result | ( input_118 & {16{sel[118]}});
    result = result | ( input_119 & {16{sel[119]}});
    result = result | ( input_120 & {16{sel[120]}});
    result = result | ( input_121 & {16{sel[121]}});
    result = result | ( input_122 & {16{sel[122]}});
    result = result | ( input_123 & {16{sel[123]}});
    result = result | ( input_124 & {16{sel[124]}});
    result = result | ( input_125 & {16{sel[125]}});
    result = result | ( input_126 & {16{sel[126]}});
    result = result | ( input_127 & {16{sel[127]}});
    result = result | ( input_128 & {16{sel[128]}});
    result = result | ( input_129 & {16{sel[129]}});
    result = result | ( input_130 & {16{sel[130]}});
    result = result | ( input_131 & {16{sel[131]}});
    result = result | ( input_132 & {16{sel[132]}});
    result = result | ( input_133 & {16{sel[133]}});
    result = result | ( input_134 & {16{sel[134]}});
    result = result | ( input_135 & {16{sel[135]}});
    result = result | ( input_136 & {16{sel[136]}});
    result = result | ( input_137 & {16{sel[137]}});
    result = result | ( input_138 & {16{sel[138]}});
    result = result | ( input_139 & {16{sel[139]}});
    result = result | ( input_140 & {16{sel[140]}});
    result = result | ( input_141 & {16{sel[141]}});
    result = result | ( input_142 & {16{sel[142]}});
    result = result | ( input_143 & {16{sel[143]}});
    result = result | ( input_144 & {16{sel[144]}});
    result = result | ( input_145 & {16{sel[145]}});
    result = result | ( input_146 & {16{sel[146]}});
    result = result | ( input_147 & {16{sel[147]}});
    result = result | ( input_148 & {16{sel[148]}});
    result = result | ( input_149 & {16{sel[149]}});
    result = result | ( input_150 & {16{sel[150]}});
    result = result | ( input_151 & {16{sel[151]}});
    result = result | ( input_152 & {16{sel[152]}});
    result = result | ( input_153 & {16{sel[153]}});
    result = result | ( input_154 & {16{sel[154]}});
    result = result | ( input_155 & {16{sel[155]}});
    result = result | ( input_156 & {16{sel[156]}});
    result = result | ( input_157 & {16{sel[157]}});
    result = result | ( input_158 & {16{sel[158]}});
    result = result | ( input_159 & {16{sel[159]}});
    result = result | ( input_160 & {16{sel[160]}});
    result = result | ( input_161 & {16{sel[161]}});
    result = result | ( input_162 & {16{sel[162]}});
    result = result | ( input_163 & {16{sel[163]}});
    result = result | ( input_164 & {16{sel[164]}});
    result = result | ( input_165 & {16{sel[165]}});
    result = result | ( input_166 & {16{sel[166]}});
    result = result | ( input_167 & {16{sel[167]}});
    result = result | ( input_168 & {16{sel[168]}});
    result = result | ( input_169 & {16{sel[169]}});
    result = result | ( input_170 & {16{sel[170]}});
    result = result | ( input_171 & {16{sel[171]}});
    result = result | ( input_172 & {16{sel[172]}});
    result = result | ( input_173 & {16{sel[173]}});
    result = result | ( input_174 & {16{sel[174]}});
    result = result | ( input_175 & {16{sel[175]}});
    result = result | ( input_176 & {16{sel[176]}});
    result = result | ( input_177 & {16{sel[177]}});
    result = result | ( input_178 & {16{sel[178]}});
    result = result | ( input_179 & {16{sel[179]}});
    result = result | ( input_180 & {16{sel[180]}});
    result = result | ( input_181 & {16{sel[181]}});
    result = result | ( input_182 & {16{sel[182]}});
    result = result | ( input_183 & {16{sel[183]}});
    result = result | ( input_184 & {16{sel[184]}});
    result = result | ( input_185 & {16{sel[185]}});
    result = result | ( input_186 & {16{sel[186]}});
    result = result | ( input_187 & {16{sel[187]}});
    result = result | ( input_188 & {16{sel[188]}});
    result = result | ( input_189 & {16{sel[189]}});
    result = result | ( input_190 & {16{sel[190]}});
    result = result | ( input_191 & {16{sel[191]}});
    result = result | ( input_192 & {16{sel[192]}});
    result = result | ( input_193 & {16{sel[193]}});
    result = result | ( input_194 & {16{sel[194]}});
    result = result | ( input_195 & {16{sel[195]}});
    result = result | ( input_196 & {16{sel[196]}});
    result = result | ( input_197 & {16{sel[197]}});
    result = result | ( input_198 & {16{sel[198]}});
    result = result | ( input_199 & {16{sel[199]}});
    result = result | ( input_200 & {16{sel[200]}});
    result = result | ( input_201 & {16{sel[201]}});
    result = result | ( input_202 & {16{sel[202]}});
    result = result | ( input_203 & {16{sel[203]}});
    result = result | ( input_204 & {16{sel[204]}});
    result = result | ( input_205 & {16{sel[205]}});
    result = result | ( input_206 & {16{sel[206]}});
    result = result | ( input_207 & {16{sel[207]}});
    result = result | ( input_208 & {16{sel[208]}});
    result = result | ( input_209 & {16{sel[209]}});
    result = result | ( input_210 & {16{sel[210]}});
    result = result | ( input_211 & {16{sel[211]}});
    result = result | ( input_212 & {16{sel[212]}});
    result = result | ( input_213 & {16{sel[213]}});
    result = result | ( input_214 & {16{sel[214]}});
    result = result | ( input_215 & {16{sel[215]}});
    result = result | ( input_216 & {16{sel[216]}});
    result = result | ( input_217 & {16{sel[217]}});
    result = result | ( input_218 & {16{sel[218]}});
    result = result | ( input_219 & {16{sel[219]}});
    result = result | ( input_220 & {16{sel[220]}});
    result = result | ( input_221 & {16{sel[221]}});
    result = result | ( input_222 & {16{sel[222]}});
    result = result | ( input_223 & {16{sel[223]}});
    result = result | ( input_224 & {16{sel[224]}});
    result = result | ( input_225 & {16{sel[225]}});
    result = result | ( input_226 & {16{sel[226]}});
    result = result | ( input_227 & {16{sel[227]}});
    result = result | ( input_228 & {16{sel[228]}});
    result = result | ( input_229 & {16{sel[229]}});
    result = result | ( input_230 & {16{sel[230]}});
    result = result | ( input_231 & {16{sel[231]}});
    result = result | ( input_232 & {16{sel[232]}});
    result = result | ( input_233 & {16{sel[233]}});
    result = result | ( input_234 & {16{sel[234]}});
    result = result | ( input_235 & {16{sel[235]}});
    result = result | ( input_236 & {16{sel[236]}});
    result = result | ( input_237 & {16{sel[237]}});
    result = result | ( input_238 & {16{sel[238]}});
    result = result | ( input_239 & {16{sel[239]}});
    result = result | ( input_240 & {16{sel[240]}});
    result = result | ( input_241 & {16{sel[241]}});
    result = result | ( input_242 & {16{sel[242]}});
    result = result | ( input_243 & {16{sel[243]}});
    result = result | ( input_244 & {16{sel[244]}});
    result = result | ( input_245 & {16{sel[245]}});
    result = result | ( input_246 & {16{sel[246]}});
    result = result | ( input_247 & {16{sel[247]}});
    result = result | ( input_248 & {16{sel[248]}});
    result = result | ( input_249 & {16{sel[249]}});
    result = result | ( input_250 & {16{sel[250]}});
    result = result | ( input_251 & {16{sel[251]}});
    result = result | ( input_252 & {16{sel[252]}});
    MUX1HOT_v_16_253_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_11_2;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [10:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    MUX1HOT_v_8_11_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_17_2;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [16:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    MUX1HOT_v_8_17_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_18_2;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [17:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    MUX1HOT_v_8_18_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_22_2;
    input [7:0] input_21;
    input [7:0] input_20;
    input [7:0] input_19;
    input [7:0] input_18;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [21:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    result = result | ( input_18 & {8{sel[18]}});
    result = result | ( input_19 & {8{sel[19]}});
    result = result | ( input_20 & {8{sel[20]}});
    result = result | ( input_21 & {8{sel[21]}});
    MUX1HOT_v_8_22_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_257_2;
    input [7:0] input_256;
    input [7:0] input_255;
    input [7:0] input_254;
    input [7:0] input_253;
    input [7:0] input_252;
    input [7:0] input_251;
    input [7:0] input_250;
    input [7:0] input_249;
    input [7:0] input_248;
    input [7:0] input_247;
    input [7:0] input_246;
    input [7:0] input_245;
    input [7:0] input_244;
    input [7:0] input_243;
    input [7:0] input_242;
    input [7:0] input_241;
    input [7:0] input_240;
    input [7:0] input_239;
    input [7:0] input_238;
    input [7:0] input_237;
    input [7:0] input_236;
    input [7:0] input_235;
    input [7:0] input_234;
    input [7:0] input_233;
    input [7:0] input_232;
    input [7:0] input_231;
    input [7:0] input_230;
    input [7:0] input_229;
    input [7:0] input_228;
    input [7:0] input_227;
    input [7:0] input_226;
    input [7:0] input_225;
    input [7:0] input_224;
    input [7:0] input_223;
    input [7:0] input_222;
    input [7:0] input_221;
    input [7:0] input_220;
    input [7:0] input_219;
    input [7:0] input_218;
    input [7:0] input_217;
    input [7:0] input_216;
    input [7:0] input_215;
    input [7:0] input_214;
    input [7:0] input_213;
    input [7:0] input_212;
    input [7:0] input_211;
    input [7:0] input_210;
    input [7:0] input_209;
    input [7:0] input_208;
    input [7:0] input_207;
    input [7:0] input_206;
    input [7:0] input_205;
    input [7:0] input_204;
    input [7:0] input_203;
    input [7:0] input_202;
    input [7:0] input_201;
    input [7:0] input_200;
    input [7:0] input_199;
    input [7:0] input_198;
    input [7:0] input_197;
    input [7:0] input_196;
    input [7:0] input_195;
    input [7:0] input_194;
    input [7:0] input_193;
    input [7:0] input_192;
    input [7:0] input_191;
    input [7:0] input_190;
    input [7:0] input_189;
    input [7:0] input_188;
    input [7:0] input_187;
    input [7:0] input_186;
    input [7:0] input_185;
    input [7:0] input_184;
    input [7:0] input_183;
    input [7:0] input_182;
    input [7:0] input_181;
    input [7:0] input_180;
    input [7:0] input_179;
    input [7:0] input_178;
    input [7:0] input_177;
    input [7:0] input_176;
    input [7:0] input_175;
    input [7:0] input_174;
    input [7:0] input_173;
    input [7:0] input_172;
    input [7:0] input_171;
    input [7:0] input_170;
    input [7:0] input_169;
    input [7:0] input_168;
    input [7:0] input_167;
    input [7:0] input_166;
    input [7:0] input_165;
    input [7:0] input_164;
    input [7:0] input_163;
    input [7:0] input_162;
    input [7:0] input_161;
    input [7:0] input_160;
    input [7:0] input_159;
    input [7:0] input_158;
    input [7:0] input_157;
    input [7:0] input_156;
    input [7:0] input_155;
    input [7:0] input_154;
    input [7:0] input_153;
    input [7:0] input_152;
    input [7:0] input_151;
    input [7:0] input_150;
    input [7:0] input_149;
    input [7:0] input_148;
    input [7:0] input_147;
    input [7:0] input_146;
    input [7:0] input_145;
    input [7:0] input_144;
    input [7:0] input_143;
    input [7:0] input_142;
    input [7:0] input_141;
    input [7:0] input_140;
    input [7:0] input_139;
    input [7:0] input_138;
    input [7:0] input_137;
    input [7:0] input_136;
    input [7:0] input_135;
    input [7:0] input_134;
    input [7:0] input_133;
    input [7:0] input_132;
    input [7:0] input_131;
    input [7:0] input_130;
    input [7:0] input_129;
    input [7:0] input_128;
    input [7:0] input_127;
    input [7:0] input_126;
    input [7:0] input_125;
    input [7:0] input_124;
    input [7:0] input_123;
    input [7:0] input_122;
    input [7:0] input_121;
    input [7:0] input_120;
    input [7:0] input_119;
    input [7:0] input_118;
    input [7:0] input_117;
    input [7:0] input_116;
    input [7:0] input_115;
    input [7:0] input_114;
    input [7:0] input_113;
    input [7:0] input_112;
    input [7:0] input_111;
    input [7:0] input_110;
    input [7:0] input_109;
    input [7:0] input_108;
    input [7:0] input_107;
    input [7:0] input_106;
    input [7:0] input_105;
    input [7:0] input_104;
    input [7:0] input_103;
    input [7:0] input_102;
    input [7:0] input_101;
    input [7:0] input_100;
    input [7:0] input_99;
    input [7:0] input_98;
    input [7:0] input_97;
    input [7:0] input_96;
    input [7:0] input_95;
    input [7:0] input_94;
    input [7:0] input_93;
    input [7:0] input_92;
    input [7:0] input_91;
    input [7:0] input_90;
    input [7:0] input_89;
    input [7:0] input_88;
    input [7:0] input_87;
    input [7:0] input_86;
    input [7:0] input_85;
    input [7:0] input_84;
    input [7:0] input_83;
    input [7:0] input_82;
    input [7:0] input_81;
    input [7:0] input_80;
    input [7:0] input_79;
    input [7:0] input_78;
    input [7:0] input_77;
    input [7:0] input_76;
    input [7:0] input_75;
    input [7:0] input_74;
    input [7:0] input_73;
    input [7:0] input_72;
    input [7:0] input_71;
    input [7:0] input_70;
    input [7:0] input_69;
    input [7:0] input_68;
    input [7:0] input_67;
    input [7:0] input_66;
    input [7:0] input_65;
    input [7:0] input_64;
    input [7:0] input_63;
    input [7:0] input_62;
    input [7:0] input_61;
    input [7:0] input_60;
    input [7:0] input_59;
    input [7:0] input_58;
    input [7:0] input_57;
    input [7:0] input_56;
    input [7:0] input_55;
    input [7:0] input_54;
    input [7:0] input_53;
    input [7:0] input_52;
    input [7:0] input_51;
    input [7:0] input_50;
    input [7:0] input_49;
    input [7:0] input_48;
    input [7:0] input_47;
    input [7:0] input_46;
    input [7:0] input_45;
    input [7:0] input_44;
    input [7:0] input_43;
    input [7:0] input_42;
    input [7:0] input_41;
    input [7:0] input_40;
    input [7:0] input_39;
    input [7:0] input_38;
    input [7:0] input_37;
    input [7:0] input_36;
    input [7:0] input_35;
    input [7:0] input_34;
    input [7:0] input_33;
    input [7:0] input_32;
    input [7:0] input_31;
    input [7:0] input_30;
    input [7:0] input_29;
    input [7:0] input_28;
    input [7:0] input_27;
    input [7:0] input_26;
    input [7:0] input_25;
    input [7:0] input_24;
    input [7:0] input_23;
    input [7:0] input_22;
    input [7:0] input_21;
    input [7:0] input_20;
    input [7:0] input_19;
    input [7:0] input_18;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [256:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    result = result | ( input_18 & {8{sel[18]}});
    result = result | ( input_19 & {8{sel[19]}});
    result = result | ( input_20 & {8{sel[20]}});
    result = result | ( input_21 & {8{sel[21]}});
    result = result | ( input_22 & {8{sel[22]}});
    result = result | ( input_23 & {8{sel[23]}});
    result = result | ( input_24 & {8{sel[24]}});
    result = result | ( input_25 & {8{sel[25]}});
    result = result | ( input_26 & {8{sel[26]}});
    result = result | ( input_27 & {8{sel[27]}});
    result = result | ( input_28 & {8{sel[28]}});
    result = result | ( input_29 & {8{sel[29]}});
    result = result | ( input_30 & {8{sel[30]}});
    result = result | ( input_31 & {8{sel[31]}});
    result = result | ( input_32 & {8{sel[32]}});
    result = result | ( input_33 & {8{sel[33]}});
    result = result | ( input_34 & {8{sel[34]}});
    result = result | ( input_35 & {8{sel[35]}});
    result = result | ( input_36 & {8{sel[36]}});
    result = result | ( input_37 & {8{sel[37]}});
    result = result | ( input_38 & {8{sel[38]}});
    result = result | ( input_39 & {8{sel[39]}});
    result = result | ( input_40 & {8{sel[40]}});
    result = result | ( input_41 & {8{sel[41]}});
    result = result | ( input_42 & {8{sel[42]}});
    result = result | ( input_43 & {8{sel[43]}});
    result = result | ( input_44 & {8{sel[44]}});
    result = result | ( input_45 & {8{sel[45]}});
    result = result | ( input_46 & {8{sel[46]}});
    result = result | ( input_47 & {8{sel[47]}});
    result = result | ( input_48 & {8{sel[48]}});
    result = result | ( input_49 & {8{sel[49]}});
    result = result | ( input_50 & {8{sel[50]}});
    result = result | ( input_51 & {8{sel[51]}});
    result = result | ( input_52 & {8{sel[52]}});
    result = result | ( input_53 & {8{sel[53]}});
    result = result | ( input_54 & {8{sel[54]}});
    result = result | ( input_55 & {8{sel[55]}});
    result = result | ( input_56 & {8{sel[56]}});
    result = result | ( input_57 & {8{sel[57]}});
    result = result | ( input_58 & {8{sel[58]}});
    result = result | ( input_59 & {8{sel[59]}});
    result = result | ( input_60 & {8{sel[60]}});
    result = result | ( input_61 & {8{sel[61]}});
    result = result | ( input_62 & {8{sel[62]}});
    result = result | ( input_63 & {8{sel[63]}});
    result = result | ( input_64 & {8{sel[64]}});
    result = result | ( input_65 & {8{sel[65]}});
    result = result | ( input_66 & {8{sel[66]}});
    result = result | ( input_67 & {8{sel[67]}});
    result = result | ( input_68 & {8{sel[68]}});
    result = result | ( input_69 & {8{sel[69]}});
    result = result | ( input_70 & {8{sel[70]}});
    result = result | ( input_71 & {8{sel[71]}});
    result = result | ( input_72 & {8{sel[72]}});
    result = result | ( input_73 & {8{sel[73]}});
    result = result | ( input_74 & {8{sel[74]}});
    result = result | ( input_75 & {8{sel[75]}});
    result = result | ( input_76 & {8{sel[76]}});
    result = result | ( input_77 & {8{sel[77]}});
    result = result | ( input_78 & {8{sel[78]}});
    result = result | ( input_79 & {8{sel[79]}});
    result = result | ( input_80 & {8{sel[80]}});
    result = result | ( input_81 & {8{sel[81]}});
    result = result | ( input_82 & {8{sel[82]}});
    result = result | ( input_83 & {8{sel[83]}});
    result = result | ( input_84 & {8{sel[84]}});
    result = result | ( input_85 & {8{sel[85]}});
    result = result | ( input_86 & {8{sel[86]}});
    result = result | ( input_87 & {8{sel[87]}});
    result = result | ( input_88 & {8{sel[88]}});
    result = result | ( input_89 & {8{sel[89]}});
    result = result | ( input_90 & {8{sel[90]}});
    result = result | ( input_91 & {8{sel[91]}});
    result = result | ( input_92 & {8{sel[92]}});
    result = result | ( input_93 & {8{sel[93]}});
    result = result | ( input_94 & {8{sel[94]}});
    result = result | ( input_95 & {8{sel[95]}});
    result = result | ( input_96 & {8{sel[96]}});
    result = result | ( input_97 & {8{sel[97]}});
    result = result | ( input_98 & {8{sel[98]}});
    result = result | ( input_99 & {8{sel[99]}});
    result = result | ( input_100 & {8{sel[100]}});
    result = result | ( input_101 & {8{sel[101]}});
    result = result | ( input_102 & {8{sel[102]}});
    result = result | ( input_103 & {8{sel[103]}});
    result = result | ( input_104 & {8{sel[104]}});
    result = result | ( input_105 & {8{sel[105]}});
    result = result | ( input_106 & {8{sel[106]}});
    result = result | ( input_107 & {8{sel[107]}});
    result = result | ( input_108 & {8{sel[108]}});
    result = result | ( input_109 & {8{sel[109]}});
    result = result | ( input_110 & {8{sel[110]}});
    result = result | ( input_111 & {8{sel[111]}});
    result = result | ( input_112 & {8{sel[112]}});
    result = result | ( input_113 & {8{sel[113]}});
    result = result | ( input_114 & {8{sel[114]}});
    result = result | ( input_115 & {8{sel[115]}});
    result = result | ( input_116 & {8{sel[116]}});
    result = result | ( input_117 & {8{sel[117]}});
    result = result | ( input_118 & {8{sel[118]}});
    result = result | ( input_119 & {8{sel[119]}});
    result = result | ( input_120 & {8{sel[120]}});
    result = result | ( input_121 & {8{sel[121]}});
    result = result | ( input_122 & {8{sel[122]}});
    result = result | ( input_123 & {8{sel[123]}});
    result = result | ( input_124 & {8{sel[124]}});
    result = result | ( input_125 & {8{sel[125]}});
    result = result | ( input_126 & {8{sel[126]}});
    result = result | ( input_127 & {8{sel[127]}});
    result = result | ( input_128 & {8{sel[128]}});
    result = result | ( input_129 & {8{sel[129]}});
    result = result | ( input_130 & {8{sel[130]}});
    result = result | ( input_131 & {8{sel[131]}});
    result = result | ( input_132 & {8{sel[132]}});
    result = result | ( input_133 & {8{sel[133]}});
    result = result | ( input_134 & {8{sel[134]}});
    result = result | ( input_135 & {8{sel[135]}});
    result = result | ( input_136 & {8{sel[136]}});
    result = result | ( input_137 & {8{sel[137]}});
    result = result | ( input_138 & {8{sel[138]}});
    result = result | ( input_139 & {8{sel[139]}});
    result = result | ( input_140 & {8{sel[140]}});
    result = result | ( input_141 & {8{sel[141]}});
    result = result | ( input_142 & {8{sel[142]}});
    result = result | ( input_143 & {8{sel[143]}});
    result = result | ( input_144 & {8{sel[144]}});
    result = result | ( input_145 & {8{sel[145]}});
    result = result | ( input_146 & {8{sel[146]}});
    result = result | ( input_147 & {8{sel[147]}});
    result = result | ( input_148 & {8{sel[148]}});
    result = result | ( input_149 & {8{sel[149]}});
    result = result | ( input_150 & {8{sel[150]}});
    result = result | ( input_151 & {8{sel[151]}});
    result = result | ( input_152 & {8{sel[152]}});
    result = result | ( input_153 & {8{sel[153]}});
    result = result | ( input_154 & {8{sel[154]}});
    result = result | ( input_155 & {8{sel[155]}});
    result = result | ( input_156 & {8{sel[156]}});
    result = result | ( input_157 & {8{sel[157]}});
    result = result | ( input_158 & {8{sel[158]}});
    result = result | ( input_159 & {8{sel[159]}});
    result = result | ( input_160 & {8{sel[160]}});
    result = result | ( input_161 & {8{sel[161]}});
    result = result | ( input_162 & {8{sel[162]}});
    result = result | ( input_163 & {8{sel[163]}});
    result = result | ( input_164 & {8{sel[164]}});
    result = result | ( input_165 & {8{sel[165]}});
    result = result | ( input_166 & {8{sel[166]}});
    result = result | ( input_167 & {8{sel[167]}});
    result = result | ( input_168 & {8{sel[168]}});
    result = result | ( input_169 & {8{sel[169]}});
    result = result | ( input_170 & {8{sel[170]}});
    result = result | ( input_171 & {8{sel[171]}});
    result = result | ( input_172 & {8{sel[172]}});
    result = result | ( input_173 & {8{sel[173]}});
    result = result | ( input_174 & {8{sel[174]}});
    result = result | ( input_175 & {8{sel[175]}});
    result = result | ( input_176 & {8{sel[176]}});
    result = result | ( input_177 & {8{sel[177]}});
    result = result | ( input_178 & {8{sel[178]}});
    result = result | ( input_179 & {8{sel[179]}});
    result = result | ( input_180 & {8{sel[180]}});
    result = result | ( input_181 & {8{sel[181]}});
    result = result | ( input_182 & {8{sel[182]}});
    result = result | ( input_183 & {8{sel[183]}});
    result = result | ( input_184 & {8{sel[184]}});
    result = result | ( input_185 & {8{sel[185]}});
    result = result | ( input_186 & {8{sel[186]}});
    result = result | ( input_187 & {8{sel[187]}});
    result = result | ( input_188 & {8{sel[188]}});
    result = result | ( input_189 & {8{sel[189]}});
    result = result | ( input_190 & {8{sel[190]}});
    result = result | ( input_191 & {8{sel[191]}});
    result = result | ( input_192 & {8{sel[192]}});
    result = result | ( input_193 & {8{sel[193]}});
    result = result | ( input_194 & {8{sel[194]}});
    result = result | ( input_195 & {8{sel[195]}});
    result = result | ( input_196 & {8{sel[196]}});
    result = result | ( input_197 & {8{sel[197]}});
    result = result | ( input_198 & {8{sel[198]}});
    result = result | ( input_199 & {8{sel[199]}});
    result = result | ( input_200 & {8{sel[200]}});
    result = result | ( input_201 & {8{sel[201]}});
    result = result | ( input_202 & {8{sel[202]}});
    result = result | ( input_203 & {8{sel[203]}});
    result = result | ( input_204 & {8{sel[204]}});
    result = result | ( input_205 & {8{sel[205]}});
    result = result | ( input_206 & {8{sel[206]}});
    result = result | ( input_207 & {8{sel[207]}});
    result = result | ( input_208 & {8{sel[208]}});
    result = result | ( input_209 & {8{sel[209]}});
    result = result | ( input_210 & {8{sel[210]}});
    result = result | ( input_211 & {8{sel[211]}});
    result = result | ( input_212 & {8{sel[212]}});
    result = result | ( input_213 & {8{sel[213]}});
    result = result | ( input_214 & {8{sel[214]}});
    result = result | ( input_215 & {8{sel[215]}});
    result = result | ( input_216 & {8{sel[216]}});
    result = result | ( input_217 & {8{sel[217]}});
    result = result | ( input_218 & {8{sel[218]}});
    result = result | ( input_219 & {8{sel[219]}});
    result = result | ( input_220 & {8{sel[220]}});
    result = result | ( input_221 & {8{sel[221]}});
    result = result | ( input_222 & {8{sel[222]}});
    result = result | ( input_223 & {8{sel[223]}});
    result = result | ( input_224 & {8{sel[224]}});
    result = result | ( input_225 & {8{sel[225]}});
    result = result | ( input_226 & {8{sel[226]}});
    result = result | ( input_227 & {8{sel[227]}});
    result = result | ( input_228 & {8{sel[228]}});
    result = result | ( input_229 & {8{sel[229]}});
    result = result | ( input_230 & {8{sel[230]}});
    result = result | ( input_231 & {8{sel[231]}});
    result = result | ( input_232 & {8{sel[232]}});
    result = result | ( input_233 & {8{sel[233]}});
    result = result | ( input_234 & {8{sel[234]}});
    result = result | ( input_235 & {8{sel[235]}});
    result = result | ( input_236 & {8{sel[236]}});
    result = result | ( input_237 & {8{sel[237]}});
    result = result | ( input_238 & {8{sel[238]}});
    result = result | ( input_239 & {8{sel[239]}});
    result = result | ( input_240 & {8{sel[240]}});
    result = result | ( input_241 & {8{sel[241]}});
    result = result | ( input_242 & {8{sel[242]}});
    result = result | ( input_243 & {8{sel[243]}});
    result = result | ( input_244 & {8{sel[244]}});
    result = result | ( input_245 & {8{sel[245]}});
    result = result | ( input_246 & {8{sel[246]}});
    result = result | ( input_247 & {8{sel[247]}});
    result = result | ( input_248 & {8{sel[248]}});
    result = result | ( input_249 & {8{sel[249]}});
    result = result | ( input_250 & {8{sel[250]}});
    result = result | ( input_251 & {8{sel[251]}});
    result = result | ( input_252 & {8{sel[252]}});
    result = result | ( input_253 & {8{sel[253]}});
    result = result | ( input_254 & {8{sel[254]}});
    result = result | ( input_255 & {8{sel[255]}});
    result = result | ( input_256 & {8{sel[256]}});
    MUX1HOT_v_8_257_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [95:0] MUX_v_96_2_2;
    input [95:0] input_0;
    input [95:0] input_1;
    input [0:0] sel;
    reg [95:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_96_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_32_1_31;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_32_1_31 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_16_33 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_33 = {{17{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct (
  clk, arst_n, input_rsc_dat_value, input_rsc_vld, input_rsc_rdy, weight_rsc_dat_value,
      weight_rsc_vld, weight_rsc_rdy, output_rsc_dat_value, output_rsc_vld, output_rsc_rdy,
      paramsIn_rsc_dat_STRIDE, paramsIn_rsc_dat_FY, paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1,
      paramsIn_rsc_dat_OC1, paramsIn_rsc_dat_OX0, paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1,
      paramsIn_rsc_dat_OY1, paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat_fy_idx,
      loopIndicesIn_rsc_dat_fx_idx, loopIndicesIn_rsc_dat_ic1_idx, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat_value;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat_value;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat_value;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] loopIndicesIn_rsc_dat_fy_idx;
  input [15:0] loopIndicesIn_rsc_dat_fx_idx;
  input [15:0] loopIndicesIn_rsc_dat_ic1_idx;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_0_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_0_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_0_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_0_i_dout_d;
  wire accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_1_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_1_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_1_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_1_i_dout_d;
  wire accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_2_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_2_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_2_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_2_i_dout_d;
  wire accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_3_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_3_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_3_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_3_i_dout_d;
  wire accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_4_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_4_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_4_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_4_i_dout_d;
  wire accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_5_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_5_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_5_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_5_i_dout_d;
  wire accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_6_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_6_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_6_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_6_i_dout_d;
  wire accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_7_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_7_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_7_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_7_i_dout_d;
  wire accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_8_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_8_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_8_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_8_i_dout_d;
  wire accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_9_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_9_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_9_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_9_i_dout_d;
  wire accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_10_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_10_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_10_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_10_i_dout_d;
  wire accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_11_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_11_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_11_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_11_i_dout_d;
  wire accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_12_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_12_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_12_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_12_i_dout_d;
  wire accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_13_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_13_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_13_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_13_i_dout_d;
  wire accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_14_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_14_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_14_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_14_i_dout_d;
  wire accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire accumulation_buffer_rsc_0_15_i_web_d;
  wire [11:0] accumulation_buffer_rsc_0_15_i_addr_d;
  wire [15:0] accumulation_buffer_rsc_0_15_i_din_d;
  wire [15:0] accumulation_buffer_rsc_0_15_i_dout_d;
  wire accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d;
  wire accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d;
  wire [15:0] accumulation_buffer_rsc_0_0_dout;
  wire [15:0] accumulation_buffer_rsc_0_0_din;
  wire [11:0] accumulation_buffer_rsc_0_0_addr;
  wire accumulation_buffer_rsc_0_0_web;
  wire accumulation_buffer_rsc_0_0_csb;
  wire [15:0] accumulation_buffer_rsc_0_1_dout;
  wire [15:0] accumulation_buffer_rsc_0_1_din;
  wire [11:0] accumulation_buffer_rsc_0_1_addr;
  wire accumulation_buffer_rsc_0_1_web;
  wire accumulation_buffer_rsc_0_1_csb;
  wire [15:0] accumulation_buffer_rsc_0_2_dout;
  wire [15:0] accumulation_buffer_rsc_0_2_din;
  wire [11:0] accumulation_buffer_rsc_0_2_addr;
  wire accumulation_buffer_rsc_0_2_web;
  wire accumulation_buffer_rsc_0_2_csb;
  wire [15:0] accumulation_buffer_rsc_0_3_dout;
  wire [15:0] accumulation_buffer_rsc_0_3_din;
  wire [11:0] accumulation_buffer_rsc_0_3_addr;
  wire accumulation_buffer_rsc_0_3_web;
  wire accumulation_buffer_rsc_0_3_csb;
  wire [15:0] accumulation_buffer_rsc_0_4_dout;
  wire [15:0] accumulation_buffer_rsc_0_4_din;
  wire [11:0] accumulation_buffer_rsc_0_4_addr;
  wire accumulation_buffer_rsc_0_4_web;
  wire accumulation_buffer_rsc_0_4_csb;
  wire [15:0] accumulation_buffer_rsc_0_5_dout;
  wire [15:0] accumulation_buffer_rsc_0_5_din;
  wire [11:0] accumulation_buffer_rsc_0_5_addr;
  wire accumulation_buffer_rsc_0_5_web;
  wire accumulation_buffer_rsc_0_5_csb;
  wire [15:0] accumulation_buffer_rsc_0_6_dout;
  wire [15:0] accumulation_buffer_rsc_0_6_din;
  wire [11:0] accumulation_buffer_rsc_0_6_addr;
  wire accumulation_buffer_rsc_0_6_web;
  wire accumulation_buffer_rsc_0_6_csb;
  wire [15:0] accumulation_buffer_rsc_0_7_dout;
  wire [15:0] accumulation_buffer_rsc_0_7_din;
  wire [11:0] accumulation_buffer_rsc_0_7_addr;
  wire accumulation_buffer_rsc_0_7_web;
  wire accumulation_buffer_rsc_0_7_csb;
  wire [15:0] accumulation_buffer_rsc_0_8_dout;
  wire [15:0] accumulation_buffer_rsc_0_8_din;
  wire [11:0] accumulation_buffer_rsc_0_8_addr;
  wire accumulation_buffer_rsc_0_8_web;
  wire accumulation_buffer_rsc_0_8_csb;
  wire [15:0] accumulation_buffer_rsc_0_9_dout;
  wire [15:0] accumulation_buffer_rsc_0_9_din;
  wire [11:0] accumulation_buffer_rsc_0_9_addr;
  wire accumulation_buffer_rsc_0_9_web;
  wire accumulation_buffer_rsc_0_9_csb;
  wire [15:0] accumulation_buffer_rsc_0_10_dout;
  wire [15:0] accumulation_buffer_rsc_0_10_din;
  wire [11:0] accumulation_buffer_rsc_0_10_addr;
  wire accumulation_buffer_rsc_0_10_web;
  wire accumulation_buffer_rsc_0_10_csb;
  wire [15:0] accumulation_buffer_rsc_0_11_dout;
  wire [15:0] accumulation_buffer_rsc_0_11_din;
  wire [11:0] accumulation_buffer_rsc_0_11_addr;
  wire accumulation_buffer_rsc_0_11_web;
  wire accumulation_buffer_rsc_0_11_csb;
  wire [15:0] accumulation_buffer_rsc_0_12_dout;
  wire [15:0] accumulation_buffer_rsc_0_12_din;
  wire [11:0] accumulation_buffer_rsc_0_12_addr;
  wire accumulation_buffer_rsc_0_12_web;
  wire accumulation_buffer_rsc_0_12_csb;
  wire [15:0] accumulation_buffer_rsc_0_13_dout;
  wire [15:0] accumulation_buffer_rsc_0_13_din;
  wire [11:0] accumulation_buffer_rsc_0_13_addr;
  wire accumulation_buffer_rsc_0_13_web;
  wire accumulation_buffer_rsc_0_13_csb;
  wire [15:0] accumulation_buffer_rsc_0_14_dout;
  wire [15:0] accumulation_buffer_rsc_0_14_din;
  wire [11:0] accumulation_buffer_rsc_0_14_addr;
  wire accumulation_buffer_rsc_0_14_web;
  wire accumulation_buffer_rsc_0_14_csb;
  wire [15:0] accumulation_buffer_rsc_0_15_dout;
  wire [15:0] accumulation_buffer_rsc_0_15_din;
  wire [11:0] accumulation_buffer_rsc_0_15_addr;
  wire accumulation_buffer_rsc_0_15_web;
  wire accumulation_buffer_rsc_0_15_csb;
  wire [255:0] output_rsc_dat;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat
      = {paramsIn_rsc_dat_STRIDE , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1
      , paramsIn_rsc_dat_OC1 , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1
      , paramsIn_rsc_dat_OY1};
  wire [47:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat
      = {loopIndicesIn_rsc_dat_fy_idx , loopIndicesIn_rsc_dat_fx_idx , loopIndicesIn_rsc_dat_ic1_idx};
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_0_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_0_csb),
      .web(accumulation_buffer_rsc_0_0_web),
      .addr(accumulation_buffer_rsc_0_0_addr),
      .din(accumulation_buffer_rsc_0_0_din),
      .dout(accumulation_buffer_rsc_0_0_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_1_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_1_csb),
      .web(accumulation_buffer_rsc_0_1_web),
      .addr(accumulation_buffer_rsc_0_1_addr),
      .din(accumulation_buffer_rsc_0_1_din),
      .dout(accumulation_buffer_rsc_0_1_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_2_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_2_csb),
      .web(accumulation_buffer_rsc_0_2_web),
      .addr(accumulation_buffer_rsc_0_2_addr),
      .din(accumulation_buffer_rsc_0_2_din),
      .dout(accumulation_buffer_rsc_0_2_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_3_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_3_csb),
      .web(accumulation_buffer_rsc_0_3_web),
      .addr(accumulation_buffer_rsc_0_3_addr),
      .din(accumulation_buffer_rsc_0_3_din),
      .dout(accumulation_buffer_rsc_0_3_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_4_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_4_csb),
      .web(accumulation_buffer_rsc_0_4_web),
      .addr(accumulation_buffer_rsc_0_4_addr),
      .din(accumulation_buffer_rsc_0_4_din),
      .dout(accumulation_buffer_rsc_0_4_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_5_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_5_csb),
      .web(accumulation_buffer_rsc_0_5_web),
      .addr(accumulation_buffer_rsc_0_5_addr),
      .din(accumulation_buffer_rsc_0_5_din),
      .dout(accumulation_buffer_rsc_0_5_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_6_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_6_csb),
      .web(accumulation_buffer_rsc_0_6_web),
      .addr(accumulation_buffer_rsc_0_6_addr),
      .din(accumulation_buffer_rsc_0_6_din),
      .dout(accumulation_buffer_rsc_0_6_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_7_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_7_csb),
      .web(accumulation_buffer_rsc_0_7_web),
      .addr(accumulation_buffer_rsc_0_7_addr),
      .din(accumulation_buffer_rsc_0_7_din),
      .dout(accumulation_buffer_rsc_0_7_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_8_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_8_csb),
      .web(accumulation_buffer_rsc_0_8_web),
      .addr(accumulation_buffer_rsc_0_8_addr),
      .din(accumulation_buffer_rsc_0_8_din),
      .dout(accumulation_buffer_rsc_0_8_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_9_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_9_csb),
      .web(accumulation_buffer_rsc_0_9_web),
      .addr(accumulation_buffer_rsc_0_9_addr),
      .din(accumulation_buffer_rsc_0_9_din),
      .dout(accumulation_buffer_rsc_0_9_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_10_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_10_csb),
      .web(accumulation_buffer_rsc_0_10_web),
      .addr(accumulation_buffer_rsc_0_10_addr),
      .din(accumulation_buffer_rsc_0_10_din),
      .dout(accumulation_buffer_rsc_0_10_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_11_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_11_csb),
      .web(accumulation_buffer_rsc_0_11_web),
      .addr(accumulation_buffer_rsc_0_11_addr),
      .din(accumulation_buffer_rsc_0_11_din),
      .dout(accumulation_buffer_rsc_0_11_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_12_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_12_csb),
      .web(accumulation_buffer_rsc_0_12_web),
      .addr(accumulation_buffer_rsc_0_12_addr),
      .din(accumulation_buffer_rsc_0_12_din),
      .dout(accumulation_buffer_rsc_0_12_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_13_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_13_csb),
      .web(accumulation_buffer_rsc_0_13_web),
      .addr(accumulation_buffer_rsc_0_13_addr),
      .din(accumulation_buffer_rsc_0_13_din),
      .dout(accumulation_buffer_rsc_0_13_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_14_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_14_csb),
      .web(accumulation_buffer_rsc_0_14_web),
      .addr(accumulation_buffer_rsc_0_14_addr),
      .din(accumulation_buffer_rsc_0_14_din),
      .dout(accumulation_buffer_rsc_0_14_dout)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd16),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) accumulation_buffer_rsc_0_15_comp (
      .clk(clk),
      .csb(accumulation_buffer_rsc_0_15_csb),
      .web(accumulation_buffer_rsc_0_15_web),
      .addr(accumulation_buffer_rsc_0_15_addr),
      .din(accumulation_buffer_rsc_0_15_din),
      .dout(accumulation_buffer_rsc_0_15_dout)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_149_16_12_256_16_gen
      accumulation_buffer_rsc_0_0_i (
      .dout(accumulation_buffer_rsc_0_0_dout),
      .din(accumulation_buffer_rsc_0_0_din),
      .addr(accumulation_buffer_rsc_0_0_addr),
      .web(accumulation_buffer_rsc_0_0_web),
      .csb(accumulation_buffer_rsc_0_0_csb),
      .web_d(accumulation_buffer_rsc_0_0_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_0_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_0_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_0_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_150_16_12_256_16_gen
      accumulation_buffer_rsc_0_1_i (
      .dout(accumulation_buffer_rsc_0_1_dout),
      .din(accumulation_buffer_rsc_0_1_din),
      .addr(accumulation_buffer_rsc_0_1_addr),
      .web(accumulation_buffer_rsc_0_1_web),
      .csb(accumulation_buffer_rsc_0_1_csb),
      .web_d(accumulation_buffer_rsc_0_1_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_1_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_1_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_1_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_151_16_12_256_16_gen
      accumulation_buffer_rsc_0_2_i (
      .dout(accumulation_buffer_rsc_0_2_dout),
      .din(accumulation_buffer_rsc_0_2_din),
      .addr(accumulation_buffer_rsc_0_2_addr),
      .web(accumulation_buffer_rsc_0_2_web),
      .csb(accumulation_buffer_rsc_0_2_csb),
      .web_d(accumulation_buffer_rsc_0_2_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_2_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_2_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_2_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_152_16_12_256_16_gen
      accumulation_buffer_rsc_0_3_i (
      .dout(accumulation_buffer_rsc_0_3_dout),
      .din(accumulation_buffer_rsc_0_3_din),
      .addr(accumulation_buffer_rsc_0_3_addr),
      .web(accumulation_buffer_rsc_0_3_web),
      .csb(accumulation_buffer_rsc_0_3_csb),
      .web_d(accumulation_buffer_rsc_0_3_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_3_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_3_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_3_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_153_16_12_256_16_gen
      accumulation_buffer_rsc_0_4_i (
      .dout(accumulation_buffer_rsc_0_4_dout),
      .din(accumulation_buffer_rsc_0_4_din),
      .addr(accumulation_buffer_rsc_0_4_addr),
      .web(accumulation_buffer_rsc_0_4_web),
      .csb(accumulation_buffer_rsc_0_4_csb),
      .web_d(accumulation_buffer_rsc_0_4_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_4_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_4_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_4_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_154_16_12_256_16_gen
      accumulation_buffer_rsc_0_5_i (
      .dout(accumulation_buffer_rsc_0_5_dout),
      .din(accumulation_buffer_rsc_0_5_din),
      .addr(accumulation_buffer_rsc_0_5_addr),
      .web(accumulation_buffer_rsc_0_5_web),
      .csb(accumulation_buffer_rsc_0_5_csb),
      .web_d(accumulation_buffer_rsc_0_5_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_5_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_5_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_5_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_155_16_12_256_16_gen
      accumulation_buffer_rsc_0_6_i (
      .dout(accumulation_buffer_rsc_0_6_dout),
      .din(accumulation_buffer_rsc_0_6_din),
      .addr(accumulation_buffer_rsc_0_6_addr),
      .web(accumulation_buffer_rsc_0_6_web),
      .csb(accumulation_buffer_rsc_0_6_csb),
      .web_d(accumulation_buffer_rsc_0_6_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_6_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_6_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_6_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_156_16_12_256_16_gen
      accumulation_buffer_rsc_0_7_i (
      .dout(accumulation_buffer_rsc_0_7_dout),
      .din(accumulation_buffer_rsc_0_7_din),
      .addr(accumulation_buffer_rsc_0_7_addr),
      .web(accumulation_buffer_rsc_0_7_web),
      .csb(accumulation_buffer_rsc_0_7_csb),
      .web_d(accumulation_buffer_rsc_0_7_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_7_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_7_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_7_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_157_16_12_256_16_gen
      accumulation_buffer_rsc_0_8_i (
      .dout(accumulation_buffer_rsc_0_8_dout),
      .din(accumulation_buffer_rsc_0_8_din),
      .addr(accumulation_buffer_rsc_0_8_addr),
      .web(accumulation_buffer_rsc_0_8_web),
      .csb(accumulation_buffer_rsc_0_8_csb),
      .web_d(accumulation_buffer_rsc_0_8_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_8_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_8_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_8_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_158_16_12_256_16_gen
      accumulation_buffer_rsc_0_9_i (
      .dout(accumulation_buffer_rsc_0_9_dout),
      .din(accumulation_buffer_rsc_0_9_din),
      .addr(accumulation_buffer_rsc_0_9_addr),
      .web(accumulation_buffer_rsc_0_9_web),
      .csb(accumulation_buffer_rsc_0_9_csb),
      .web_d(accumulation_buffer_rsc_0_9_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_9_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_9_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_9_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_159_16_12_256_16_gen
      accumulation_buffer_rsc_0_10_i (
      .dout(accumulation_buffer_rsc_0_10_dout),
      .din(accumulation_buffer_rsc_0_10_din),
      .addr(accumulation_buffer_rsc_0_10_addr),
      .web(accumulation_buffer_rsc_0_10_web),
      .csb(accumulation_buffer_rsc_0_10_csb),
      .web_d(accumulation_buffer_rsc_0_10_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_10_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_10_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_10_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_160_16_12_256_16_gen
      accumulation_buffer_rsc_0_11_i (
      .dout(accumulation_buffer_rsc_0_11_dout),
      .din(accumulation_buffer_rsc_0_11_din),
      .addr(accumulation_buffer_rsc_0_11_addr),
      .web(accumulation_buffer_rsc_0_11_web),
      .csb(accumulation_buffer_rsc_0_11_csb),
      .web_d(accumulation_buffer_rsc_0_11_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_11_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_11_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_11_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_161_16_12_256_16_gen
      accumulation_buffer_rsc_0_12_i (
      .dout(accumulation_buffer_rsc_0_12_dout),
      .din(accumulation_buffer_rsc_0_12_din),
      .addr(accumulation_buffer_rsc_0_12_addr),
      .web(accumulation_buffer_rsc_0_12_web),
      .csb(accumulation_buffer_rsc_0_12_csb),
      .web_d(accumulation_buffer_rsc_0_12_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_12_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_12_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_12_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_162_16_12_256_16_gen
      accumulation_buffer_rsc_0_13_i (
      .dout(accumulation_buffer_rsc_0_13_dout),
      .din(accumulation_buffer_rsc_0_13_din),
      .addr(accumulation_buffer_rsc_0_13_addr),
      .web(accumulation_buffer_rsc_0_13_web),
      .csb(accumulation_buffer_rsc_0_13_csb),
      .web_d(accumulation_buffer_rsc_0_13_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_13_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_13_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_13_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_163_16_12_256_16_gen
      accumulation_buffer_rsc_0_14_i (
      .dout(accumulation_buffer_rsc_0_14_dout),
      .din(accumulation_buffer_rsc_0_14_din),
      .addr(accumulation_buffer_rsc_0_14_addr),
      .web(accumulation_buffer_rsc_0_14_web),
      .csb(accumulation_buffer_rsc_0_14_csb),
      .web_d(accumulation_buffer_rsc_0_14_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_14_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_14_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_14_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_sram_512_128_sram_512_128_rwport_164_16_12_256_16_gen
      accumulation_buffer_rsc_0_15_i (
      .dout(accumulation_buffer_rsc_0_15_dout),
      .din(accumulation_buffer_rsc_0_15_din),
      .addr(accumulation_buffer_rsc_0_15_addr),
      .web(accumulation_buffer_rsc_0_15_web),
      .csb(accumulation_buffer_rsc_0_15_csb),
      .web_d(accumulation_buffer_rsc_0_15_i_web_d),
      .addr_d(accumulation_buffer_rsc_0_15_i_addr_d),
      .din_d(accumulation_buffer_rsc_0_15_i_din_d),
      .dout_d(accumulation_buffer_rsc_0_15_i_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat_value),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .weight_rsc_dat(weight_rsc_dat_value),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .loopIndicesIn_rsc_dat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat[47:0]),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .accumulation_buffer_rsc_0_0_i_web_d(accumulation_buffer_rsc_0_0_i_web_d),
      .accumulation_buffer_rsc_0_0_i_addr_d(accumulation_buffer_rsc_0_0_i_addr_d),
      .accumulation_buffer_rsc_0_0_i_din_d(accumulation_buffer_rsc_0_0_i_din_d),
      .accumulation_buffer_rsc_0_0_i_dout_d(accumulation_buffer_rsc_0_0_i_dout_d),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_0_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_1_i_web_d(accumulation_buffer_rsc_0_1_i_web_d),
      .accumulation_buffer_rsc_0_1_i_addr_d(accumulation_buffer_rsc_0_1_i_addr_d),
      .accumulation_buffer_rsc_0_1_i_din_d(accumulation_buffer_rsc_0_1_i_din_d),
      .accumulation_buffer_rsc_0_1_i_dout_d(accumulation_buffer_rsc_0_1_i_dout_d),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_1_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_2_i_web_d(accumulation_buffer_rsc_0_2_i_web_d),
      .accumulation_buffer_rsc_0_2_i_addr_d(accumulation_buffer_rsc_0_2_i_addr_d),
      .accumulation_buffer_rsc_0_2_i_din_d(accumulation_buffer_rsc_0_2_i_din_d),
      .accumulation_buffer_rsc_0_2_i_dout_d(accumulation_buffer_rsc_0_2_i_dout_d),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_2_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_3_i_web_d(accumulation_buffer_rsc_0_3_i_web_d),
      .accumulation_buffer_rsc_0_3_i_addr_d(accumulation_buffer_rsc_0_3_i_addr_d),
      .accumulation_buffer_rsc_0_3_i_din_d(accumulation_buffer_rsc_0_3_i_din_d),
      .accumulation_buffer_rsc_0_3_i_dout_d(accumulation_buffer_rsc_0_3_i_dout_d),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_3_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_4_i_web_d(accumulation_buffer_rsc_0_4_i_web_d),
      .accumulation_buffer_rsc_0_4_i_addr_d(accumulation_buffer_rsc_0_4_i_addr_d),
      .accumulation_buffer_rsc_0_4_i_din_d(accumulation_buffer_rsc_0_4_i_din_d),
      .accumulation_buffer_rsc_0_4_i_dout_d(accumulation_buffer_rsc_0_4_i_dout_d),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_4_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_5_i_web_d(accumulation_buffer_rsc_0_5_i_web_d),
      .accumulation_buffer_rsc_0_5_i_addr_d(accumulation_buffer_rsc_0_5_i_addr_d),
      .accumulation_buffer_rsc_0_5_i_din_d(accumulation_buffer_rsc_0_5_i_din_d),
      .accumulation_buffer_rsc_0_5_i_dout_d(accumulation_buffer_rsc_0_5_i_dout_d),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_5_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_6_i_web_d(accumulation_buffer_rsc_0_6_i_web_d),
      .accumulation_buffer_rsc_0_6_i_addr_d(accumulation_buffer_rsc_0_6_i_addr_d),
      .accumulation_buffer_rsc_0_6_i_din_d(accumulation_buffer_rsc_0_6_i_din_d),
      .accumulation_buffer_rsc_0_6_i_dout_d(accumulation_buffer_rsc_0_6_i_dout_d),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_6_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_7_i_web_d(accumulation_buffer_rsc_0_7_i_web_d),
      .accumulation_buffer_rsc_0_7_i_addr_d(accumulation_buffer_rsc_0_7_i_addr_d),
      .accumulation_buffer_rsc_0_7_i_din_d(accumulation_buffer_rsc_0_7_i_din_d),
      .accumulation_buffer_rsc_0_7_i_dout_d(accumulation_buffer_rsc_0_7_i_dout_d),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_7_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_8_i_web_d(accumulation_buffer_rsc_0_8_i_web_d),
      .accumulation_buffer_rsc_0_8_i_addr_d(accumulation_buffer_rsc_0_8_i_addr_d),
      .accumulation_buffer_rsc_0_8_i_din_d(accumulation_buffer_rsc_0_8_i_din_d),
      .accumulation_buffer_rsc_0_8_i_dout_d(accumulation_buffer_rsc_0_8_i_dout_d),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_8_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_9_i_web_d(accumulation_buffer_rsc_0_9_i_web_d),
      .accumulation_buffer_rsc_0_9_i_addr_d(accumulation_buffer_rsc_0_9_i_addr_d),
      .accumulation_buffer_rsc_0_9_i_din_d(accumulation_buffer_rsc_0_9_i_din_d),
      .accumulation_buffer_rsc_0_9_i_dout_d(accumulation_buffer_rsc_0_9_i_dout_d),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_9_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_10_i_web_d(accumulation_buffer_rsc_0_10_i_web_d),
      .accumulation_buffer_rsc_0_10_i_addr_d(accumulation_buffer_rsc_0_10_i_addr_d),
      .accumulation_buffer_rsc_0_10_i_din_d(accumulation_buffer_rsc_0_10_i_din_d),
      .accumulation_buffer_rsc_0_10_i_dout_d(accumulation_buffer_rsc_0_10_i_dout_d),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_10_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_11_i_web_d(accumulation_buffer_rsc_0_11_i_web_d),
      .accumulation_buffer_rsc_0_11_i_addr_d(accumulation_buffer_rsc_0_11_i_addr_d),
      .accumulation_buffer_rsc_0_11_i_din_d(accumulation_buffer_rsc_0_11_i_din_d),
      .accumulation_buffer_rsc_0_11_i_dout_d(accumulation_buffer_rsc_0_11_i_dout_d),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_11_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_12_i_web_d(accumulation_buffer_rsc_0_12_i_web_d),
      .accumulation_buffer_rsc_0_12_i_addr_d(accumulation_buffer_rsc_0_12_i_addr_d),
      .accumulation_buffer_rsc_0_12_i_din_d(accumulation_buffer_rsc_0_12_i_din_d),
      .accumulation_buffer_rsc_0_12_i_dout_d(accumulation_buffer_rsc_0_12_i_dout_d),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_12_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_13_i_web_d(accumulation_buffer_rsc_0_13_i_web_d),
      .accumulation_buffer_rsc_0_13_i_addr_d(accumulation_buffer_rsc_0_13_i_addr_d),
      .accumulation_buffer_rsc_0_13_i_din_d(accumulation_buffer_rsc_0_13_i_din_d),
      .accumulation_buffer_rsc_0_13_i_dout_d(accumulation_buffer_rsc_0_13_i_dout_d),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_13_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_14_i_web_d(accumulation_buffer_rsc_0_14_i_web_d),
      .accumulation_buffer_rsc_0_14_i_addr_d(accumulation_buffer_rsc_0_14_i_addr_d),
      .accumulation_buffer_rsc_0_14_i_din_d(accumulation_buffer_rsc_0_14_i_din_d),
      .accumulation_buffer_rsc_0_14_i_dout_d(accumulation_buffer_rsc_0_14_i_dout_d),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_14_i_port_0_rw_ram_ir_internal_WMASK_B_d),
      .accumulation_buffer_rsc_0_15_i_web_d(accumulation_buffer_rsc_0_15_i_web_d),
      .accumulation_buffer_rsc_0_15_i_addr_d(accumulation_buffer_rsc_0_15_i_addr_d),
      .accumulation_buffer_rsc_0_15_i_din_d(accumulation_buffer_rsc_0_15_i_din_d),
      .accumulation_buffer_rsc_0_15_i_dout_d(accumulation_buffer_rsc_0_15_i_dout_d),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_RMASK_B_d),
      .accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_15_i_port_0_rw_ram_ir_internal_WMASK_B_d)
    );
  assign output_rsc_dat_value = output_rsc_dat;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16 (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;


  // Interconnect Declarations
  wire [255:0] output_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE
      = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY
      = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX
      = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1
      = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1
      = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0
      = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0
      = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1
      = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1
      = paramsIn_rsc_dat[15:0];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx
      = loopIndicesIn_rsc_dat[47:32];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx
      = loopIndicesIn_rsc_dat[31:16];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx
      = loopIndicesIn_rsc_dat[15:0];
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat_value(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .weight_rsc_dat_value(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .output_rsc_dat_value(output_rsc_dat_value),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .loopIndicesIn_rsc_dat_fy_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx[15:0]),
      .loopIndicesIn_rsc_dat_fx_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx[15:0]),
      .loopIndicesIn_rsc_dat_ic1_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx[15:0]),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy)
    );
  assign output_rsc_dat = output_rsc_dat_value;
endmodule




//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_in_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_sync_v2 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0
    
    generate 
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data 
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd; 
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
    // synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
    // synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;       // experiment
 
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    // KH assign active = din_vld_int | dout_rdy; // (din_vld & ~din_rdy) | (dout_rdy & ~dout_vld);
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];
             
          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0)) 
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end
        
        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else 
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        if ( peak < count )
          peak = count;
        // synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT 
    generate
    if (ph_clk==1) 
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0) 
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif
   
endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock 
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;
   
    // synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
    // synopsys translate_on

    ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ../WeightDoubleBufferless_384comma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy07
//  Generated date: Sun Feb 23 19:22:11 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    WeightDoublefeSAqem_cns_bctl
// ------------------------------------------------------------------


module WeightDoublefeSAqem_cns_bctl (
  clk, arst_n, paramsIn_rsc_rdy_nweightDoubleBufferWriter, din_rsc_rdy_nweightDoubleBufferWriter,
      dout_rsc_csb_nweightDoubleBufferWriter, dout_rsc_web_nweightDoubleBufferWriter,
      dout_rsc_addr_nweightDoubleBufferWriter, dout_rsc_din_nweightDoubleBufferWriter,
      dout_rsc_dout_nweightDoubleBufferWriter, dout_rsc_req_vz_nweightDoubleBufferWriter,
      paramsIn_rsc_rdy_nweightDoubleBufferReader, din_rsc_csb_nweightDoubleBufferReader,
      din_rsc_web_nweightDoubleBufferReader, din_rsc_addr_nweightDoubleBufferReader,
      din_rsc_din_nweightDoubleBufferReader, din_rsc_dout_nweightDoubleBufferReader,
      din_rsc_req_vz_nweightDoubleBufferReader, dout_rsc_vld_nweightDoubleBufferReader,
      paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud, din_rsc_rdy_nweightDoubleBufferWriter_bud,
      dout_rsc_rls_lz_nweightDoubleBufferWriter_bud, din_rsc_rls_lz_nweightDoubleBufferReader_bud,
      paramsIn_rsc_rdy_nweightDoubleBufferReader_bud, dout_rsc_vld_nweightDoubleBufferReader_bud,
      mem_cns_S0, mem_cns_R0, mem_cns_S1, mem_cns_R1, mem_cns_csb_shi0, mem_cns_csb_shi1,
      mem_cns_web_shi0, mem_cns_web_shi1, mem_cns_addr_shi0, mem_cns_addr_shi1, mem_cns_din_shi0,
      mem_cns_din_shi1, mem_cns_dout_sho0, mem_cns_dout_sho1, mem_cns_S1_pff, mem_cns_S0_pff
);
  input clk;
  input arst_n;
  output paramsIn_rsc_rdy_nweightDoubleBufferWriter;
  output din_rsc_rdy_nweightDoubleBufferWriter;
  input dout_rsc_csb_nweightDoubleBufferWriter;
  input dout_rsc_web_nweightDoubleBufferWriter;
  input [11:0] dout_rsc_addr_nweightDoubleBufferWriter;
  input [127:0] dout_rsc_din_nweightDoubleBufferWriter;
  output [127:0] dout_rsc_dout_nweightDoubleBufferWriter;
  output dout_rsc_req_vz_nweightDoubleBufferWriter;
  output paramsIn_rsc_rdy_nweightDoubleBufferReader;
  input din_rsc_csb_nweightDoubleBufferReader;
  input din_rsc_web_nweightDoubleBufferReader;
  input [11:0] din_rsc_addr_nweightDoubleBufferReader;
  input [127:0] din_rsc_din_nweightDoubleBufferReader;
  output [127:0] din_rsc_dout_nweightDoubleBufferReader;
  output din_rsc_req_vz_nweightDoubleBufferReader;
  output dout_rsc_vld_nweightDoubleBufferReader;
  input paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  input din_rsc_rdy_nweightDoubleBufferWriter_bud;
  input dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  input din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  input paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  input dout_rsc_vld_nweightDoubleBufferReader_bud;
  output mem_cns_S0;
  input mem_cns_R0;
  output mem_cns_S1;
  input mem_cns_R1;
  output mem_cns_csb_shi0;
  output mem_cns_csb_shi1;
  output mem_cns_web_shi0;
  output mem_cns_web_shi1;
  output [11:0] mem_cns_addr_shi0;
  output [11:0] mem_cns_addr_shi1;
  output [127:0] mem_cns_din_shi0;
  output [127:0] mem_cns_din_shi1;
  input [127:0] mem_cns_dout_sho0;
  input [127:0] mem_cns_dout_sho1;
  output mem_cns_S1_pff;
  output mem_cns_S0_pff;


  // Interconnect Declarations
  wire mem_cns_PC0;
  reg mem_cns_ppidx;
  reg [1:0] mem_cns_ppown;
  wire mem_cns_PC1;
  reg mem_cns_ppidx_1;
  reg [1:0] mem_cns_ppown_1;
  wire mem_cns_ppsel_1_pff;
  wire [1:0] mem_acc_1_rmff;
  wire [3:0] nl_mem_acc_1_rmff;
  wire mem_xor_1_rmff;
  wire mem_or_cse_pff;
  wire [1:0] mem_acc_rmff;
  wire [3:0] nl_mem_acc_rmff;
  wire mem_xor_rmff;
  wire mem_cns_ppsel_3_pff;
  wire mem_or_6_cse_pff;

  wire[0:0] mem_mux_11_nl;
  wire[0:0] mem_mux_13_nl;
  wire[0:0] mem_mux_10_nl;
  wire[0:0] mem_mux_12_nl;

  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsc_rdy_nweightDoubleBufferWriter = paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  assign din_rsc_rdy_nweightDoubleBufferWriter = din_rsc_rdy_nweightDoubleBufferWriter_bud;
  assign paramsIn_rsc_rdy_nweightDoubleBufferReader = paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  assign dout_rsc_vld_nweightDoubleBufferReader = dout_rsc_vld_nweightDoubleBufferReader_bud;
  assign dout_rsc_req_vz_nweightDoubleBufferWriter = mem_cns_R0;
  assign din_rsc_req_vz_nweightDoubleBufferReader = mem_cns_R1;
  assign mem_xor_rmff = mem_cns_ppidx ^ mem_cns_PC0;
  assign nl_mem_acc_rmff = mem_cns_ppown + conv_u2u_1_2(mem_cns_PC0) + conv_s2u_1_2(mem_cns_PC1);
  assign mem_acc_rmff = nl_mem_acc_rmff[1:0];
  assign mem_cns_PC0 = mem_cns_S0 & dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  assign mem_xor_1_rmff = mem_cns_ppidx_1 ^ mem_cns_PC1;
  assign nl_mem_acc_1_rmff = mem_cns_ppown_1 + conv_u2u_1_2(mem_cns_PC1) + conv_s2u_1_2(mem_cns_PC0);
  assign mem_acc_1_rmff = nl_mem_acc_1_rmff[1:0];
  assign mem_cns_PC1 = mem_cns_S1 & din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  assign dout_rsc_dout_nweightDoubleBufferWriter = MUX_v_128_2_2(mem_cns_dout_sho0,
      mem_cns_dout_sho1, mem_cns_ppidx);
  assign din_rsc_dout_nweightDoubleBufferReader = MUX_v_128_2_2(mem_cns_dout_sho0,
      mem_cns_dout_sho1, mem_cns_ppidx_1);
  assign mem_mux_11_nl = MUX_s_1_2_2((~ dout_rsc_csb_nweightDoubleBufferWriter),
      (~ din_rsc_csb_nweightDoubleBufferReader), mem_cns_ppsel_1_pff);
  assign mem_cns_csb_shi0 = ~((mem_mux_11_nl) & mem_or_cse_pff);
  assign mem_cns_S1 = (mem_cns_ppown_1!=2'b00);
  assign mem_cns_S1_pff = (mem_acc_1_rmff!=2'b00);
  assign mem_cns_ppsel_1_pff = mem_cns_S1_pff & (~ mem_xor_1_rmff);
  assign mem_cns_S0 = ~((mem_cns_ppown==2'b10));
  assign mem_cns_S0_pff = ~((mem_acc_rmff==2'b10));
  assign mem_or_cse_pff = (mem_cns_S0_pff & (~ mem_xor_rmff)) | mem_cns_ppsel_1_pff;
  assign mem_mux_13_nl = MUX_s_1_2_2((~ dout_rsc_web_nweightDoubleBufferWriter),
      (~ din_rsc_web_nweightDoubleBufferReader), mem_cns_ppsel_1_pff);
  assign mem_cns_web_shi0 = ~((mem_mux_13_nl) & mem_or_cse_pff);
  assign mem_cns_addr_shi0 = MUX_v_12_2_2(dout_rsc_addr_nweightDoubleBufferWriter,
      din_rsc_addr_nweightDoubleBufferReader, mem_cns_ppsel_1_pff);
  assign mem_cns_din_shi0 = MUX_v_128_2_2(dout_rsc_din_nweightDoubleBufferWriter,
      din_rsc_din_nweightDoubleBufferReader, mem_cns_ppsel_1_pff);
  assign mem_mux_10_nl = MUX_s_1_2_2((~ dout_rsc_csb_nweightDoubleBufferWriter),
      (~ din_rsc_csb_nweightDoubleBufferReader), mem_cns_ppsel_3_pff);
  assign mem_cns_csb_shi1 = ~((mem_mux_10_nl) & mem_or_6_cse_pff);
  assign mem_cns_ppsel_3_pff = mem_cns_S1_pff & mem_xor_1_rmff;
  assign mem_or_6_cse_pff = (mem_cns_S0_pff & mem_xor_rmff) | mem_cns_ppsel_3_pff;
  assign mem_mux_12_nl = MUX_s_1_2_2((~ dout_rsc_web_nweightDoubleBufferWriter),
      (~ din_rsc_web_nweightDoubleBufferReader), mem_cns_ppsel_3_pff);
  assign mem_cns_web_shi1 = ~((mem_mux_12_nl) & mem_or_6_cse_pff);
  assign mem_cns_addr_shi1 = MUX_v_12_2_2(dout_rsc_addr_nweightDoubleBufferWriter,
      din_rsc_addr_nweightDoubleBufferReader, mem_cns_ppsel_3_pff);
  assign mem_cns_din_shi1 = MUX_v_128_2_2(dout_rsc_din_nweightDoubleBufferWriter,
      din_rsc_din_nweightDoubleBufferReader, mem_cns_ppsel_3_pff);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mem_cns_ppidx <= 1'b0;
      mem_cns_ppown <= 2'b00;
      mem_cns_ppidx_1 <= 1'b0;
      mem_cns_ppown_1 <= 2'b00;
    end
    else begin
      mem_cns_ppidx <= mem_xor_rmff;
      mem_cns_ppown <= mem_acc_rmff;
      mem_cns_ppidx_1 <= mem_xor_1_rmff;
      mem_cns_ppown_1 <= mem_acc_1_rmff;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier
// ------------------------------------------------------------------


module unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for WeightDoubleBuffer_384_16_16_run_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBuffer_384_16_16_run_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_staller
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_staller (
  run_wen, paramsIn_rsci_wen_comp, weightDoubleBufferWriterParams_cnsi_wen_comp,
      weightDoubleBufferReaderParams_cnsi_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input weightDoubleBufferWriterParams_cnsi_wen_comp;
  input weightDoubleBufferReaderParams_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & weightDoubleBufferWriterParams_cnsi_wen_comp
      & weightDoubleBufferReaderParams_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
    (
  clk, arst_n, weightDoubleBufferReaderParams_cnsi_oswt, weightDoubleBufferReaderParams_cnsi_wen_comp,
      weightDoubleBufferReaderParams_cnsi_biwt, weightDoubleBufferReaderParams_cnsi_bdwt,
      weightDoubleBufferReaderParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  output weightDoubleBufferReaderParams_cnsi_wen_comp;
  input weightDoubleBufferReaderParams_cnsi_biwt;
  input weightDoubleBufferReaderParams_cnsi_bdwt;
  output weightDoubleBufferReaderParams_cnsi_bcwt;
  reg weightDoubleBufferReaderParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferReaderParams_cnsi_wen_comp = (~ weightDoubleBufferReaderParams_cnsi_oswt)
      | weightDoubleBufferReaderParams_cnsi_biwt | weightDoubleBufferReaderParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weightDoubleBufferReaderParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      weightDoubleBufferReaderParams_cnsi_bcwt <= ~((~(weightDoubleBufferReaderParams_cnsi_bcwt
          | weightDoubleBufferReaderParams_cnsi_biwt)) | weightDoubleBufferReaderParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
    (
  run_wen, weightDoubleBufferReaderParams_cnsi_oswt, weightDoubleBufferReaderParams_cnsi_irdy,
      weightDoubleBufferReaderParams_cnsi_biwt, weightDoubleBufferReaderParams_cnsi_bdwt,
      weightDoubleBufferReaderParams_cnsi_bcwt, weightDoubleBufferReaderParams_cnsi_ivld_run_sct
);
  input run_wen;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  input weightDoubleBufferReaderParams_cnsi_irdy;
  output weightDoubleBufferReaderParams_cnsi_biwt;
  output weightDoubleBufferReaderParams_cnsi_bdwt;
  input weightDoubleBufferReaderParams_cnsi_bcwt;
  output weightDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire weightDoubleBufferReaderParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferReaderParams_cnsi_bdwt = weightDoubleBufferReaderParams_cnsi_oswt
      & run_wen;
  assign weightDoubleBufferReaderParams_cnsi_biwt = weightDoubleBufferReaderParams_cnsi_ogwt
      & weightDoubleBufferReaderParams_cnsi_irdy;
  assign weightDoubleBufferReaderParams_cnsi_ogwt = weightDoubleBufferReaderParams_cnsi_oswt
      & (~ weightDoubleBufferReaderParams_cnsi_bcwt);
  assign weightDoubleBufferReaderParams_cnsi_ivld_run_sct = weightDoubleBufferReaderParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
    (
  clk, arst_n, weightDoubleBufferWriterParams_cnsi_oswt, weightDoubleBufferWriterParams_cnsi_wen_comp,
      weightDoubleBufferWriterParams_cnsi_biwt, weightDoubleBufferWriterParams_cnsi_bdwt,
      weightDoubleBufferWriterParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  output weightDoubleBufferWriterParams_cnsi_wen_comp;
  input weightDoubleBufferWriterParams_cnsi_biwt;
  input weightDoubleBufferWriterParams_cnsi_bdwt;
  output weightDoubleBufferWriterParams_cnsi_bcwt;
  reg weightDoubleBufferWriterParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferWriterParams_cnsi_wen_comp = (~ weightDoubleBufferWriterParams_cnsi_oswt)
      | weightDoubleBufferWriterParams_cnsi_biwt | weightDoubleBufferWriterParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weightDoubleBufferWriterParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      weightDoubleBufferWriterParams_cnsi_bcwt <= ~((~(weightDoubleBufferWriterParams_cnsi_bcwt
          | weightDoubleBufferWriterParams_cnsi_biwt)) | weightDoubleBufferWriterParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
    (
  run_wen, weightDoubleBufferWriterParams_cnsi_oswt, weightDoubleBufferWriterParams_cnsi_irdy,
      weightDoubleBufferWriterParams_cnsi_biwt, weightDoubleBufferWriterParams_cnsi_bdwt,
      weightDoubleBufferWriterParams_cnsi_bcwt, weightDoubleBufferWriterParams_cnsi_ivld_run_sct
);
  input run_wen;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  input weightDoubleBufferWriterParams_cnsi_irdy;
  output weightDoubleBufferWriterParams_cnsi_biwt;
  output weightDoubleBufferWriterParams_cnsi_bdwt;
  input weightDoubleBufferWriterParams_cnsi_bcwt;
  output weightDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire weightDoubleBufferWriterParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferWriterParams_cnsi_bdwt = weightDoubleBufferWriterParams_cnsi_oswt
      & run_wen;
  assign weightDoubleBufferWriterParams_cnsi_biwt = weightDoubleBufferWriterParams_cnsi_ogwt
      & weightDoubleBufferWriterParams_cnsi_irdy;
  assign weightDoubleBufferWriterParams_cnsi_ogwt = weightDoubleBufferWriterParams_cnsi_oswt
      & (~ weightDoubleBufferWriterParams_cnsi_bcwt);
  assign weightDoubleBufferWriterParams_cnsi_ivld_run_sct = weightDoubleBufferWriterParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_sram_512_128_sram_512_128_rwport_3_128_12_384_128_gen
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_sram_512_128_sram_512_128_rwport_3_128_12_384_128_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [127:0] dout;
  output [127:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [127:0] din_d;
  output [127:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign dout_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (dout_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_2_tr0, while_while_C_0_tr0, while_while_C_0_tr1,
      while_while_for_for_C_0_tr0, while_while_for_C_1_tr0, while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input main_C_2_tr0;
  input while_while_C_0_tr0;
  input while_while_C_0_tr1;
  input while_while_for_for_C_0_tr0;
  input while_while_for_C_1_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for WeightDoubleBufferWriter_384_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    while_C_0 = 4'd4,
    while_while_C_0 = 4'd5,
    while_while_for_for_C_0 = 4'd6,
    while_while_for_C_0 = 4'd7,
    while_while_for_C_1 = 4'd8,
    while_while_C_1 = 4'd9,
    while_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBufferWriter_384_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 11'b00000001000;
        if ( main_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 11'b00000100000;
        if ( while_while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else if ( while_while_C_0_tr1 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_for_C_0 : begin
        fsm_output = 11'b00001000000;
        if ( while_while_for_for_C_0_tr0 ) begin
          state_var_NS = while_while_for_C_0;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = while_while_for_C_1;
      end
      while_while_for_C_1 : begin
        fsm_output = 11'b00100000000;
        if ( while_while_for_C_1_tr0 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_C_1 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 11'b10000000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_staller
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, din_rsci_wen_comp, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input din_rsci_wen_comp;
  input dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & din_rsci_wen_comp & dout_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
    (
  clk, arst_n, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt, dout_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;
  input dout_rsc_req_obj_biwt;
  input dout_rsc_req_obj_bdwt;
  output dout_rsc_req_obj_bcwt;
  reg dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_wen_comp = (~ dout_rsc_req_obj_oswt) | dout_rsc_req_obj_biwt
      | dout_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_bcwt <= ~((~(dout_rsc_req_obj_bcwt | dout_rsc_req_obj_biwt))
          | dout_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
    (
  run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_vd, dout_rsc_req_obj_biwt, dout_rsc_req_obj_bdwt,
      dout_rsc_req_obj_bcwt
);
  input run_wen;
  input dout_rsc_req_obj_oswt;
  input dout_rsc_req_obj_vd;
  output dout_rsc_req_obj_biwt;
  output dout_rsc_req_obj_bdwt;
  input dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_bdwt = dout_rsc_req_obj_oswt & run_wen;
  assign dout_rsc_req_obj_biwt = dout_rsc_req_obj_oswt & (~ dout_rsc_req_obj_bcwt)
      & dout_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
    (
  run_wten, dout_rsc_rls_obj_iswt0, dout_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input dout_rsc_rls_obj_iswt0;
  output dout_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_rls_obj_ld_run_sct = dout_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl (
  dout_rsci_web_d_run_sct_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_web_d_run_sct_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_web_d_run_sct_pff = dout_rsci_iswt0_pff & (~ run_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp (
  clk, arst_n, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt, din_rsci_biwt,
      din_rsci_bdwt, din_rsci_bcwt, din_rsci_idat
);
  input clk;
  input arst_n;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  output din_rsci_bcwt;
  reg din_rsci_bcwt;
  input [15:0] din_rsci_idat;


  // Interconnect Declarations
  reg [15:0] din_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_idat_mxwt = MUX_v_16_2_2(din_rsci_idat, din_rsci_idat_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_idat_bfwt <= din_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl (
  run_wen, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_bcwt, din_rsci_irdy_run_sct,
      din_rsci_ivld
);
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  input din_rsci_bcwt;
  output din_rsci_irdy_run_sct;
  input din_rsci_ivld;


  // Interconnect Declarations
  wire din_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_ivld;
  assign din_rsci_ogwt = din_rsci_oswt & (~ din_rsci_bcwt);
  assign din_rsci_irdy_run_sct = din_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [73:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [4:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [36:0] reg_paramsIn_rsci_idat_bfwt_ftd_12;
  reg [31:0] reg_paramsIn_rsci_idat_bfwt_ftd_45;
  wire [4:0] paramsIn_rsci_idat_mxwt_opt_116_112;
  wire [36:0] paramsIn_rsci_idat_mxwt_opt_100_64;
  wire [31:0] paramsIn_rsci_idat_mxwt_opt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_116_112 = MUX_v_5_2_2((paramsIn_rsci_idat[116:112]),
      reg_paramsIn_rsci_idat_bfwt_ftd, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_100_64 = MUX_v_37_2_2((paramsIn_rsci_idat[100:64]),
      reg_paramsIn_rsci_idat_bfwt_ftd_12, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_31_0 = MUX_v_32_2_2((paramsIn_rsci_idat[31:0]),
      reg_paramsIn_rsci_idat_bfwt_ftd_45, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {paramsIn_rsci_idat_mxwt_opt_116_112 , paramsIn_rsci_idat_mxwt_opt_100_64
      , paramsIn_rsci_idat_mxwt_opt_31_0};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 5'b00000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_opt_116_112;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= 37'b0000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= paramsIn_rsci_idat_mxwt_opt_100_64;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= paramsIn_rsci_idat_mxwt_opt_31_0;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [36:0] MUX_v_37_2_2;
    input [36:0] input_0;
    input [36:0] input_1;
    input [0:0] sel;
    reg [36:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_37_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_sram_512_128_sram_512_128_rwport_8_128_12_384_128_gen
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_sram_512_128_sram_512_128_rwport_8_128_12_384_128_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [127:0] dout;
  output [127:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [127:0] din_d;
  output [127:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign din_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (din_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_2_tr0, while_while_C_0_tr0, while_while_for_C_0_tr0,
      while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input main_C_2_tr0;
  input while_while_C_0_tr0;
  input while_while_for_C_0_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for WeightDoubleBufferReader_384_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    while_C_0 = 4'd4,
    while_while_C_0 = 4'd5,
    while_while_for_C_0 = 4'd6,
    while_while_C_1 = 4'd7,
    while_C_1 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBufferReader_384_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 9'b000001000;
        if ( main_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 9'b000010000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 9'b000100000;
        if ( while_while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 9'b001000000;
        if ( while_while_for_C_0_tr0 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_C_1 : begin
        fsm_output = 9'b010000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 9'b100000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_staller
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, dout_rsci_wen_comp, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input dout_rsci_wen_comp;
  input din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & dout_rsci_wen_comp & din_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
    (
  clk, arst_n, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt, din_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;
  input din_rsc_req_obj_biwt;
  input din_rsc_req_obj_bdwt;
  output din_rsc_req_obj_bcwt;
  reg din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_wen_comp = (~ din_rsc_req_obj_oswt) | din_rsc_req_obj_biwt
      | din_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_bcwt <= ~((~(din_rsc_req_obj_bcwt | din_rsc_req_obj_biwt))
          | din_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
    (
  run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_vd, din_rsc_req_obj_biwt, din_rsc_req_obj_bdwt,
      din_rsc_req_obj_bcwt
);
  input run_wen;
  input din_rsc_req_obj_oswt;
  input din_rsc_req_obj_vd;
  output din_rsc_req_obj_biwt;
  output din_rsc_req_obj_bdwt;
  input din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_bdwt = din_rsc_req_obj_oswt & run_wen;
  assign din_rsc_req_obj_biwt = din_rsc_req_obj_oswt & (~ din_rsc_req_obj_bcwt) &
      din_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
    (
  run_wten, din_rsc_rls_obj_iswt0, din_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input din_rsc_rls_obj_iswt0;
  output din_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_rls_obj_ld_run_sct = din_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp (
  clk, arst_n, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_bcwt
);
  input clk;
  input arst_n;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;
  output dout_rsci_bcwt;
  reg dout_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl (
  run_wen, dout_rsci_oswt, dout_rsci_irdy, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt,
      dout_rsci_ivld_run_sct
);
  input run_wen;
  input dout_rsci_oswt;
  input dout_rsci_irdy;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  input dout_rsci_bcwt;
  output dout_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dout_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_bdwt = dout_rsci_oswt & run_wen;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_irdy;
  assign dout_rsci_ogwt = dout_rsci_oswt & (~ dout_rsci_bcwt);
  assign dout_rsci_ivld_run_sct = dout_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl (
  run_wen, run_wten, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_addr_d_run_sct_pff,
      din_rsci_oswt_pff
);
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_addr_d_run_sct_pff;
  input din_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = (~ run_wten) & din_rsci_oswt;
  assign din_rsci_addr_d_run_sct_pff = din_rsci_oswt_pff & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp (
  clk, arst_n, din_rsci_addr_d, din_rsci_dout_d, din_rsci_addr_d_run, din_rsci_dout_d_mxwt,
      din_rsci_biwt, din_rsci_bdwt, din_rsci_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  input [11:0] din_rsci_addr_d_run;
  output [127:0] din_rsci_dout_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input din_rsci_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [127:0] din_rsci_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_dout_d_mxwt = MUX_v_128_2_2(din_rsci_dout_d, din_rsci_dout_d_bfwt,
      din_rsci_bcwt);
  assign din_rsci_addr_d = {(~ din_rsci_addr_d_run_sct_pff) , (~ din_rsci_addr_d_run_sct_pff)
      , (~ din_rsci_addr_d_run_sct_pff) , (din_rsci_addr_d_run[8:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_dout_d_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_dout_d_bfwt <= din_rsci_dout_d_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [63:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [31:0] reg_paramsIn_rsci_idat_bfwt_ftd_33;
  wire [63:0] paramsIn_rsci_idat_mxwt_opt_127_64;
  wire [31:0] paramsIn_rsci_idat_mxwt_opt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_127_64 = MUX_v_64_2_2((paramsIn_rsci_idat[127:64]),
      reg_paramsIn_rsci_idat_bfwt_ftd, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_31_0 = MUX_v_32_2_2((paramsIn_rsci_idat[31:0]),
      reg_paramsIn_rsci_idat_bfwt_ftd_33, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {paramsIn_rsci_idat_mxwt_opt_127_64 , paramsIn_rsci_idat_mxwt_opt_31_0};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_opt_127_64;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_33 <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_33 <= paramsIn_rsci_idat_mxwt_opt_31_0;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi (
  clk, arst_n, weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy, run_wen, weightDoubleBufferReaderParams_cnsi_oswt,
      weightDoubleBufferReaderParams_cnsi_wen_comp, weightDoubleBufferReaderParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;
  input run_wen;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  output weightDoubleBufferReaderParams_cnsi_wen_comp;
  input [143:0] weightDoubleBufferReaderParams_cnsi_idat;


  // Interconnect Declarations
  wire weightDoubleBufferReaderParams_cnsi_irdy;
  wire weightDoubleBufferReaderParams_cnsi_biwt;
  wire weightDoubleBufferReaderParams_cnsi_bdwt;
  wire weightDoubleBufferReaderParams_cnsi_bcwt;
  wire weightDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd19),
  .width(32'sd144)) weightDoubleBufferReaderParams_cnsi (
      .irdy(weightDoubleBufferReaderParams_cnsi_irdy),
      .ivld(weightDoubleBufferReaderParams_cnsi_ivld_run_sct),
      .idat(weightDoubleBufferReaderParams_cnsi_idat),
      .rdy(weightDoubleBufferReaderParams_cns_rdy),
      .vld(weightDoubleBufferReaderParams_cns_vld),
      .dat(weightDoubleBufferReaderParams_cns_dat)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weightDoubleBufferReaderParams_cnsi_oswt(weightDoubleBufferReaderParams_cnsi_oswt),
      .weightDoubleBufferReaderParams_cnsi_irdy(weightDoubleBufferReaderParams_cnsi_irdy),
      .weightDoubleBufferReaderParams_cnsi_biwt(weightDoubleBufferReaderParams_cnsi_biwt),
      .weightDoubleBufferReaderParams_cnsi_bdwt(weightDoubleBufferReaderParams_cnsi_bdwt),
      .weightDoubleBufferReaderParams_cnsi_bcwt(weightDoubleBufferReaderParams_cnsi_bcwt),
      .weightDoubleBufferReaderParams_cnsi_ivld_run_sct(weightDoubleBufferReaderParams_cnsi_ivld_run_sct)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferReaderParams_cnsi_oswt(weightDoubleBufferReaderParams_cnsi_oswt),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_biwt(weightDoubleBufferReaderParams_cnsi_biwt),
      .weightDoubleBufferReaderParams_cnsi_bdwt(weightDoubleBufferReaderParams_cnsi_bdwt),
      .weightDoubleBufferReaderParams_cnsi_bcwt(weightDoubleBufferReaderParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi (
  clk, arst_n, weightDoubleBufferWriterParams_cns_dat, weightDoubleBufferWriterParams_cns_vld,
      weightDoubleBufferWriterParams_cns_rdy, run_wen, weightDoubleBufferWriterParams_cnsi_oswt,
      weightDoubleBufferWriterParams_cnsi_wen_comp, weightDoubleBufferWriterParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  input run_wen;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  output weightDoubleBufferWriterParams_cnsi_wen_comp;
  input [143:0] weightDoubleBufferWriterParams_cnsi_idat;


  // Interconnect Declarations
  wire weightDoubleBufferWriterParams_cnsi_irdy;
  wire weightDoubleBufferWriterParams_cnsi_biwt;
  wire weightDoubleBufferWriterParams_cnsi_bdwt;
  wire weightDoubleBufferWriterParams_cnsi_bcwt;
  wire weightDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd18),
  .width(32'sd144)) weightDoubleBufferWriterParams_cnsi (
      .irdy(weightDoubleBufferWriterParams_cnsi_irdy),
      .ivld(weightDoubleBufferWriterParams_cnsi_ivld_run_sct),
      .idat(weightDoubleBufferWriterParams_cnsi_idat),
      .rdy(weightDoubleBufferWriterParams_cns_rdy),
      .vld(weightDoubleBufferWriterParams_cns_vld),
      .dat(weightDoubleBufferWriterParams_cns_dat)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weightDoubleBufferWriterParams_cnsi_oswt(weightDoubleBufferWriterParams_cnsi_oswt),
      .weightDoubleBufferWriterParams_cnsi_irdy(weightDoubleBufferWriterParams_cnsi_irdy),
      .weightDoubleBufferWriterParams_cnsi_biwt(weightDoubleBufferWriterParams_cnsi_biwt),
      .weightDoubleBufferWriterParams_cnsi_bdwt(weightDoubleBufferWriterParams_cnsi_bdwt),
      .weightDoubleBufferWriterParams_cnsi_bcwt(weightDoubleBufferWriterParams_cnsi_bcwt),
      .weightDoubleBufferWriterParams_cnsi_ivld_run_sct(weightDoubleBufferWriterParams_cnsi_ivld_run_sct)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferWriterParams_cnsi_oswt(weightDoubleBufferWriterParams_cnsi_oswt),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_biwt(weightDoubleBufferWriterParams_cnsi_biwt),
      .weightDoubleBufferWriterParams_cnsi_bdwt(weightDoubleBufferWriterParams_cnsi_bdwt),
      .weightDoubleBufferWriterParams_cnsi_bcwt(weightDoubleBufferWriterParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd17),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj (
  clk, arst_n, dout_rsc_req_vz, run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input dout_rsc_req_vz;
  input run_wen;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_rsc_req_obj_vd;
  wire dout_rsc_req_obj_biwt;
  wire dout_rsc_req_obj_bdwt;
  wire dout_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) dout_rsc_req_obj (
      .vd(dout_rsc_req_obj_vd),
      .vz(dout_rsc_req_vz)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
      WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_vd(dout_rsc_req_obj_vd),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj (
  dout_rsc_rls_lz, run_wten, dout_rsc_rls_obj_iswt0
);
  output dout_rsc_rls_lz;
  input run_wten;
  input dout_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) dout_rsc_rls_obj (
      .ld(dout_rsc_rls_obj_ld_run_sct),
      .lz(dout_rsc_rls_lz)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
      WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(dout_rsc_rls_obj_iswt0),
      .dout_rsc_rls_obj_ld_run_sct(dout_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1 (
  dout_rsci_addr_d, dout_rsci_addr_d_run, dout_rsci_web_d_pff, dout_rsci_iswt0_pff,
      run_wten_pff
);
  output [11:0] dout_rsci_addr_d;
  input [11:0] dout_rsci_addr_d_run;
  output dout_rsci_web_d_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;


  // Interconnect Declarations
  wire dout_rsci_web_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl_inst
      (
      .dout_rsci_web_d_run_sct_pff(dout_rsci_web_d_run_sct_iff),
      .dout_rsci_iswt0_pff(dout_rsci_iswt0_pff),
      .run_wten_pff(run_wten_pff)
    );
  assign dout_rsci_web_d_pff = ~ dout_rsci_web_d_run_sct_iff;
  assign dout_rsci_addr_d = {(~ dout_rsci_web_d_run_sct_iff) , (~ dout_rsci_web_d_run_sct_iff)
      , (~ dout_rsci_web_d_run_sct_iff) , (dout_rsci_addr_d_run[8:0])};
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci (
  clk, arst_n, din_rsc_dat, din_rsc_vld, din_rsc_rdy, run_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_bcwt;
  wire din_rsci_irdy_run_sct;
  wire din_rsci_ivld;
  wire [15:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd16)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_irdy_run_sct),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_irdy_run_sct(din_rsci_irdy_run_sct),
      .din_rsci_ivld(din_rsci_ivld)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_idat(din_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [73:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [73:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj (
  clk, arst_n, din_rsc_req_vz, run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input din_rsc_req_vz;
  input run_wen;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_rsc_req_obj_vd;
  wire din_rsc_req_obj_biwt;
  wire din_rsc_req_obj_bdwt;
  wire din_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) din_rsc_req_obj (
      .vd(din_rsc_req_obj_vd),
      .vz(din_rsc_req_vz)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_vd(din_rsc_req_obj_vd),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj (
  din_rsc_rls_lz, run_wten, din_rsc_rls_obj_iswt0
);
  output din_rsc_rls_lz;
  input run_wten;
  input din_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) din_rsc_rls_obj (
      .ld(din_rsc_rls_obj_ld_run_sct),
      .lz(din_rsc_rls_lz)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(din_rsc_rls_obj_iswt0),
      .din_rsc_rls_obj_ld_run_sct(din_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci (
  clk, arst_n, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, run_wen, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_idat
);
  input clk;
  input arst_n;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [127:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_irdy;
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_bcwt;
  wire dout_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd128)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_ivld_run_sct),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_irdy(dout_rsci_irdy),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt),
      .dout_rsci_ivld_run_sct(dout_rsci_ivld_run_sct)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1 (
  clk, arst_n, din_rsci_addr_d, din_rsci_dout_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      run_wen, run_wten, din_rsci_oswt, din_rsci_addr_d_run, din_rsci_dout_d_mxwt,
      din_rsci_oswt_pff
);
  input clk;
  input arst_n;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  input [11:0] din_rsci_addr_d_run;
  output [127:0] din_rsci_dout_d_mxwt;
  input din_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire [11:0] din_rsci_addr_d_reg;
  wire din_rsci_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run;
  assign nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run
      = {3'b000 , (din_rsci_addr_d_run[8:0])};
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_addr_d(din_rsci_addr_d_reg),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_addr_d_run(nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run[11:0]),
      .din_rsci_dout_d_mxwt(din_rsci_dout_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_addr_d_run_sct_pff(din_rsci_addr_d_run_sct_iff)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_addr_d_run_sct_pff(din_rsci_addr_d_run_sct_iff),
      .din_rsci_oswt_pff(din_rsci_oswt_pff)
    );
  assign din_rsci_addr_d = din_rsci_addr_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_addr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [95:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, weightDoubleBufferWriterParams_cns_dat,
      weightDoubleBufferWriterParams_cns_vld, weightDoubleBufferWriterParams_cns_rdy,
      weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire weightDoubleBufferWriterParams_cnsi_wen_comp;
  wire weightDoubleBufferReaderParams_cnsi_wen_comp;
  wire [2:0] fsm_output;
  reg reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse;
  reg [143:0] reg_weightDoubleBufferReaderParams_cnsi_idat_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy),
      .run_wen(run_wen),
      .weightDoubleBufferWriterParams_cnsi_oswt(reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_idat(reg_weightDoubleBufferReaderParams_cnsi_idat_cse)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy),
      .run_wen(run_wen),
      .weightDoubleBufferReaderParams_cnsi_oswt(reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_idat(reg_weightDoubleBufferReaderParams_cnsi_idat_cse)
    );
  WeightDoubleBuffer_384_16_16_run_run_staller WeightDoubleBuffer_384_16_16_run_run_staller_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp)
    );
  WeightDoubleBuffer_384_16_16_run_run_run_fsm WeightDoubleBuffer_384_16_16_run_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_weightDoubleBufferReaderParams_cnsi_idat_cse <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_weightDoubleBufferReaderParams_cnsi_idat_cse <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= fsm_output[1];
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~ (fsm_output[1]);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_req_vz, dout_rsc_rls_lz, dout_rsci_addr_d,
      dout_rsci_din_d, dout_rsci_web_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;
  output [11:0] dout_rsci_addr_d;
  output [127:0] dout_rsci_din_d;
  output dout_rsci_web_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [73:0] paramsIn_rsci_idat_mxwt;
  wire din_rsci_wen_comp;
  wire [15:0] din_rsci_idat_mxwt;
  wire dout_rsc_req_obj_wen_comp;
  wire [10:0] fsm_output;
  wire [3:0] while_while_for_for_acc_1_tmp;
  wire [4:0] nl_while_while_for_for_acc_1_tmp;
  wire and_dcpl_3;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire or_dcpl_19;
  wire and_dcpl_10;
  wire or_dcpl_25;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_34;
  reg exit_while_while_for_sva;
  wire exit_while_sva_mx0;
  reg [2:0] while_while_for_for_oc0_idx_3_0_sva_2_0;
  reg [31:0] reg_paramsIn_crt_sva_116_0_ftd_21;
  reg reg_dout_rsc_req_obj_iswt0_cse;
  reg reg_dout_rsc_rls_obj_ld_run_psct_cse;
  reg reg_din_rsci_irdy_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire dout_rsci_web_d_iff;
  wire [11:0] dout_rsci_addr_d_reg;
  reg [8:0] while_while_for_idx_sva;
  reg [15:0] while_while_for_for_tmp_value_sva;
  reg [7:0] while_while_for_row_value_13_sva;
  reg [7:0] while_while_for_row_value_12_sva;
  reg [7:0] while_while_for_row_value_11_sva;
  reg [7:0] while_while_for_row_value_10_sva;
  reg [7:0] while_while_for_row_value_9_sva;
  reg [7:0] while_while_for_row_value_8_sva;
  reg [7:0] while_while_for_row_value_7_sva;
  reg [7:0] while_while_for_row_value_6_sva;
  reg [7:0] while_while_for_row_value_5_sva;
  reg [7:0] while_while_for_row_value_4_sva;
  reg [7:0] while_while_for_row_value_3_sva;
  reg [7:0] while_while_for_row_value_2_sva;
  reg [7:0] while_while_for_row_value_1_sva;
  reg [7:0] while_while_for_row_value_0_sva;
  reg [4:0] while_current_buffer_size_8_4_sva;
  reg [4:0] block_size_mul_psp_sva;
  wire [9:0] nl_block_size_mul_psp_sva;
  reg [63:0] total_blocks_lpi_3;
  reg [31:0] total_blocks_mul_2_itm;
  reg [47:0] total_blocks_mul_1_itm;
  wire [63:0] total_blocks_sva_1;
  wire [8:0] while_while_for_idx_sva_2;
  wire [9:0] nl_while_while_for_idx_sva_2;
  wire while_while_for_row_value_and_1_cse;
  wire while_while_for_row_value_and_cse;
  wire while_while_for_row_value_and_3_cse;
  wire while_while_for_row_value_and_2_cse;
  wire while_while_for_row_value_and_5_cse;
  wire while_while_for_row_value_and_4_cse;
  wire while_while_for_row_value_and_12_cse;
  wire operator_64_false_1_acc_1_itm_64_1;
  wire while_while_for_acc_2_itm_5_1;
  wire while_while_aelse_acc_itm_5_1;

  wire[63:0] while_while_acc_nl;
  wire[64:0] nl_while_while_acc_nl;
  wire[4:0] while_current_buffer_size_mux_nl;
  wire[4:0] while_while_acc_2_nl;
  wire[5:0] nl_while_while_acc_2_nl;
  wire[0:0] while_current_buffer_size_or_nl;
  wire[5:0] while_while_for_acc_3_nl;
  wire[7:0] nl_while_while_for_acc_3_nl;
  wire[8:0] while_while_for_idx_mux_nl;
  wire[0:0] or_nl;
  wire[0:0] not_60_nl;
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire[64:0] operator_64_false_1_acc_1_nl;
  wire[65:0] nl_operator_64_false_1_acc_1_nl;
  wire[5:0] while_while_for_acc_2_nl;
  wire[6:0] nl_while_while_for_acc_2_nl;
  wire[5:0] while_while_aelse_acc_nl;
  wire[6:0] nl_while_while_aelse_acc_nl;
  wire[5:0] while_while_aelse_acc_1_nl;
  wire[6:0] nl_while_while_aelse_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[4:0] while_while_for_for_1_1_acc_4_nl;
  wire[5:0] nl_while_while_for_for_1_1_acc_4_nl;
  wire [11:0] nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run;
  assign nl_while_while_for_for_1_1_acc_4_nl = while_current_buffer_size_8_4_sva
      + (while_while_for_idx_sva[8:4]);
  assign while_while_for_for_1_1_acc_4_nl = nl_while_while_for_for_1_1_acc_4_nl[4:0];
  assign nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run
      = {3'b000 , (while_while_for_for_1_1_acc_4_nl) , (while_while_for_idx_sva[3:0])};
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff
      = fsm_output[7];
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff
      = ~ run_wen;
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0
      = or_dcpl_19;
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1
      = and_dcpl_3 & (~ while_while_for_acc_2_itm_5_1);
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0
      = while_while_for_for_acc_1_tmp[3];
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci WeightDoubleBufferWriter_384_16_16_run_din_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .run_wen(run_wen),
      .din_rsci_oswt(reg_din_rsci_irdy_run_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1 WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst
      (
      .dout_rsci_addr_d(dout_rsci_addr_d_reg),
      .dout_rsci_addr_d_run(nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run[11:0]),
      .dout_rsci_web_d_pff(dout_rsci_web_d_iff),
      .dout_rsci_iswt0_pff(nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff[0:0]),
      .run_wten_pff(nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff[0:0])
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_inst
      (
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(reg_dout_rsc_rls_obj_ld_run_psct_cse)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(reg_dout_rsc_req_obj_iswt0_cse),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferWriter_384_16_16_run_staller WeightDoubleBufferWriter_384_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferWriter_384_16_16_run_run_fsm WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_2_tr0(exit_while_sva_mx0),
      .while_while_C_0_tr0(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0[0:0]),
      .while_while_C_0_tr1(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1[0:0]),
      .while_while_for_for_C_0_tr0(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0[0:0]),
      .while_while_for_C_1_tr0(exit_while_while_for_sva),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign while_while_for_row_value_and_cse = run_wen & (or_dcpl_7 | or_dcpl_6);
  assign while_while_for_row_value_and_1_cse = run_wen & (or_dcpl_4 | or_dcpl_9);
  assign while_while_for_row_value_and_2_cse = run_wen & (or_dcpl_7 | or_dcpl_9);
  assign while_while_for_row_value_and_3_cse = run_wen & (or_dcpl_4 | or_dcpl_6);
  assign while_while_for_row_value_and_4_cse = run_wen & (or_dcpl_7 | or_dcpl_3);
  assign while_while_for_row_value_and_5_cse = run_wen & (or_dcpl_4 | (while_while_for_for_acc_1_tmp[1:0]!=2'b11));
  assign while_while_for_row_value_and_12_cse = run_wen & (or_dcpl_4 | or_dcpl_3);
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ (readslicef_65_1_64((operator_64_false_acc_1_nl)))),
      (~ operator_64_false_1_acc_1_itm_64_1), fsm_output[10]);
  assign total_blocks_sva_1 = conv_u2u_64_64(total_blocks_mul_1_itm * (reg_paramsIn_crt_sva_116_0_ftd_21[15:0]));
  assign nl_while_while_for_idx_sva_2 = while_while_for_idx_sva + 9'b000000001;
  assign while_while_for_idx_sva_2 = nl_while_while_for_idx_sva_2[8:0];
  assign nl_while_while_for_for_acc_1_tmp = conv_u2s_3_4(while_while_for_for_oc0_idx_3_0_sva_2_0)
      + 4'b0001;
  assign while_while_for_for_acc_1_tmp = nl_while_while_for_for_acc_1_tmp[3:0];
  assign nl_operator_64_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_1_acc_1_nl = nl_operator_64_false_1_acc_1_nl[64:0];
  assign operator_64_false_1_acc_1_itm_64_1 = readslicef_65_1_64((operator_64_false_1_acc_1_nl));
  assign and_dcpl_3 = operator_64_false_1_acc_1_itm_64_1 & (~ while_while_aelse_acc_itm_5_1);
  assign or_dcpl_3 = (while_while_for_for_acc_1_tmp[1:0]!=2'b00);
  assign or_dcpl_4 = (while_while_for_for_acc_1_tmp[3:2]!=2'b00);
  assign or_dcpl_6 = (while_while_for_for_acc_1_tmp[1:0]!=2'b10);
  assign or_dcpl_7 = (while_while_for_for_acc_1_tmp[3:2]!=2'b01);
  assign or_dcpl_9 = (while_while_for_for_acc_1_tmp[1:0]!=2'b01);
  assign or_dcpl_19 = (~ operator_64_false_1_acc_1_itm_64_1) | while_while_aelse_acc_itm_5_1;
  assign and_dcpl_10 = ~((fsm_output[1:0]!=2'b00));
  assign or_dcpl_25 = (while_while_for_for_oc0_idx_3_0_sva_2_0!=3'b110);
  assign or_dcpl_26 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b00);
  assign or_dcpl_27 = or_dcpl_26 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_28 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b10);
  assign or_dcpl_29 = or_dcpl_28 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_30 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b01);
  assign or_dcpl_31 = or_dcpl_30 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign or_dcpl_32 = or_dcpl_28 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign or_dcpl_33 = or_dcpl_30 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_34 = or_dcpl_26 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign nl_while_while_for_acc_2_nl = ({1'b1 , (~ block_size_mul_psp_sva)}) + 6'b000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[5:0];
  assign while_while_for_acc_2_itm_5_1 = readslicef_6_1_5((while_while_for_acc_2_nl));
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_5_6(~ while_current_buffer_size_8_4_sva)
      + conv_u2u_5_6(~ block_size_mul_psp_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[5:0];
  assign nl_while_while_aelse_acc_nl = conv_u2u_5_6(readslicef_6_5_1((while_while_aelse_acc_1_nl)))
      + 6'b101101;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[5:0];
  assign while_while_aelse_acc_itm_5_1 = readslicef_6_1_5((while_while_aelse_acc_nl));
  assign dout_rsci_web_d_pff = dout_rsci_web_d_iff;
  assign dout_rsci_addr_d = dout_rsci_addr_d_reg;
  assign dout_rsci_din_d = {while_while_for_for_tmp_value_sva , while_while_for_row_value_13_sva
      , while_while_for_row_value_12_sva , while_while_for_row_value_11_sva , while_while_for_row_value_10_sva
      , while_while_for_row_value_9_sva , while_while_for_row_value_8_sva , while_while_for_row_value_7_sva
      , while_while_for_row_value_6_sva , while_while_for_row_value_5_sva , while_while_for_row_value_4_sva
      , while_while_for_row_value_3_sva , while_while_for_row_value_2_sva , while_while_for_row_value_1_sva
      , while_while_for_row_value_0_sva};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_din_rsci_irdy_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      total_blocks_mul_2_itm <= 32'b00000000000000000000000000000000;
      total_blocks_mul_1_itm <= 48'b000000000000000000000000000000000000000000000000;
      while_current_buffer_size_8_4_sva <= 5'b00000;
      exit_while_while_for_sva <= 1'b0;
      while_while_for_idx_sva <= 9'b000000000;
      while_while_for_for_oc0_idx_3_0_sva_2_0 <= 3'b000;
    end
    else if ( run_wen ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= ~(exit_while_sva_mx0 | (~((fsm_output[3])
          | (fsm_output[10]))));
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_19 & (fsm_output[5]);
      reg_din_rsci_irdy_run_psct_cse <= (and_dcpl_3 & while_while_for_acc_2_itm_5_1
          & (fsm_output[5])) | ((~ (while_while_for_for_acc_1_tmp[3])) & (fsm_output[6]))
          | ((~ exit_while_while_for_sva) & (fsm_output[8]));
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[3]) | (fsm_output[10])
          | (fsm_output[0]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      total_blocks_mul_2_itm <= conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16]) *
          (paramsIn_rsci_idat_mxwt[15:0]));
      total_blocks_mul_1_itm <= conv_u2u_48_48(total_blocks_mul_2_itm * (reg_paramsIn_crt_sva_116_0_ftd_21[31:16]));
      while_current_buffer_size_8_4_sva <= MUX_v_5_2_2(5'b00000, (while_current_buffer_size_mux_nl),
          (while_current_buffer_size_or_nl));
      exit_while_while_for_sva <= ~ (readslicef_6_1_5((while_while_for_acc_3_nl)));
      while_while_for_idx_sva <= MUX_v_9_2_2(9'b000000000, (while_while_for_idx_mux_nl),
          (not_60_nl));
      while_while_for_for_oc0_idx_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (while_while_for_for_acc_1_tmp[2:0]),
          (fsm_output[6]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_mul_psp_sva <= 5'b00000;
    end
    else if ( run_wen & (~ and_dcpl_10) ) begin
      block_size_mul_psp_sva <= nl_block_size_mul_psp_sva[4:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((fsm_output[2]) | (fsm_output[3]) | (fsm_output[9]) | (~
        and_dcpl_10)) ) begin
      total_blocks_lpi_3 <= MUX_v_64_2_2(total_blocks_sva_1, (while_while_acc_nl),
          fsm_output[9]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_13_sva <= 8'b00000000;
      while_while_for_row_value_12_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_cse ) begin
      while_while_for_row_value_13_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_13_sva, or_dcpl_25);
      while_while_for_row_value_12_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_row_value_12_sva, or_dcpl_25);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_3_sva <= 8'b00000000;
      while_while_for_row_value_2_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_1_cse ) begin
      while_while_for_row_value_3_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_3_sva, or_dcpl_27);
      while_while_for_row_value_2_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_2_sva,
          or_dcpl_27);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_11_sva <= 8'b00000000;
      while_while_for_row_value_10_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_2_cse ) begin
      while_while_for_row_value_11_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_11_sva, or_dcpl_29);
      while_while_for_row_value_10_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_row_value_10_sva, or_dcpl_29);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_5_sva <= 8'b00000000;
      while_while_for_row_value_4_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_3_cse ) begin
      while_while_for_row_value_5_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_5_sva, or_dcpl_31);
      while_while_for_row_value_4_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_4_sva,
          or_dcpl_31);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_9_sva <= 8'b00000000;
      while_while_for_row_value_8_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_4_cse ) begin
      while_while_for_row_value_9_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_9_sva, or_dcpl_32);
      while_while_for_row_value_8_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_8_sva,
          or_dcpl_32);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_7_sva <= 8'b00000000;
      while_while_for_row_value_6_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_5_cse ) begin
      while_while_for_row_value_7_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_7_sva, or_dcpl_33);
      while_while_for_row_value_6_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_6_sva,
          or_dcpl_33);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_1_sva <= 8'b00000000;
      while_while_for_row_value_0_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_12_cse ) begin
      while_while_for_row_value_1_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_1_sva, or_dcpl_34);
      while_while_for_row_value_0_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_0_sva,
          or_dcpl_34);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_tmp_value_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (while_while_for_for_acc_1_tmp[3]) ) begin
      while_while_for_for_tmp_value_sva <= din_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_crt_sva_116_0_ftd_21 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_paramsIn_crt_sva_116_0_ftd_21 <= paramsIn_rsci_idat_mxwt[63:32];
    end
  end
  assign nl_while_while_acc_2_nl = while_current_buffer_size_8_4_sva + block_size_mul_psp_sva;
  assign while_while_acc_2_nl = nl_while_while_acc_2_nl[4:0];
  assign while_current_buffer_size_mux_nl = MUX_v_5_2_2(while_current_buffer_size_8_4_sva,
      (while_while_acc_2_nl), fsm_output[9]);
  assign while_current_buffer_size_or_nl = (fsm_output[9:5]!=5'b00000);
  assign nl_while_while_for_acc_3_nl = ({1'b1 , (while_while_for_idx_sva_2[8:4])})
      + conv_u2u_5_6(~ block_size_mul_psp_sva) + 6'b000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[5:0];
  assign or_nl = (fsm_output[6]) | (fsm_output[8]);
  assign while_while_for_idx_mux_nl = MUX_v_9_2_2(while_while_for_idx_sva_2, while_while_for_idx_sva,
      or_nl);
  assign not_60_nl = ~ (fsm_output[5]);
  assign nl_block_size_mul_psp_sva  = (paramsIn_rsci_idat_mxwt[73:69]) * (paramsIn_rsci_idat_mxwt[68:64]);
  assign nl_while_while_acc_nl = total_blocks_lpi_3 + 64'b1111111111111111111111111111111111111111111111111111111111111111;
  assign while_while_acc_nl = nl_while_while_acc_nl[63:0];

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_6_5_1;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_6_5_1 = tmp[4:0];
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction


  function automatic [63:0] conv_u2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_64 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_req_vz,
      din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, din_rsci_addr_d,
      din_rsci_dout_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [95:0] paramsIn_rsci_idat_mxwt;
  wire [127:0] din_rsci_dout_d_mxwt;
  wire dout_rsci_wen_comp;
  reg [127:0] dout_rsci_idat;
  wire din_rsc_req_obj_wen_comp;
  wire [8:0] fsm_output;
  wire [4:0] while_while_for_for_acc_tmp;
  wire [5:0] nl_while_while_for_for_acc_tmp;
  wire or_dcpl_1;
  wire or_dcpl_4;
  wire or_tmp_13;
  wire or_tmp_22;
  wire exit_while_sva_mx0;
  reg exitL_exit_while_while_for_for_sva;
  reg while_while_for_stage_0;
  reg while_while_for_stage_0_2;
  reg exit_while_while_for_lpi_4_dfm_st_1;
  reg [63:0] reg_paramsIn_crt_sva_127_0_ftd;
  reg reg_din_rsc_req_obj_iswt0_cse;
  reg reg_din_rsc_rls_obj_ld_run_psct_cse;
  reg reg_dout_rsci_ivld_run_psct_cse;
  reg reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire [11:0] din_rsci_addr_d_reg;
  wire and_41_rmff;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  wire [3:0] din_rsci_addr_d_run_3_0_mx1;
  reg [4:0] while_block_count_4_0_sva;
  reg [4:0] block_size_mul_psp_sva;
  reg [31:0] total_blocks_mul_2_itm;
  reg [63:0] total_blocks_lpi_3;
  reg [4:0] while_current_buffer_size_8_4_sva;
  reg [47:0] total_blocks_mul_1_itm;
  reg [3:0] while_while_for_for_r_idx_4_0_lpi_4_3_0;
  wire [63:0] total_blocks_sva_1;
  wire while_while_for_acc_2_itm_32_1;
  wire operator_64_false_1_acc_1_itm_64_1;

  wire[4:0] block_size_mul_nl;
  wire[9:0] nl_block_size_mul_nl;
  wire[31:0] total_blocks_mux1h_2_nl;
  wire[31:0] total_blocks_mul_2_nl;
  wire[31:0] while_while_for_acc_1_nl;
  wire[32:0] nl_while_while_for_acc_1_nl;
  wire[0:0] total_blocks_and_1_nl;
  wire[0:0] total_blocks_and_2_nl;
  wire[0:0] not_nl;
  wire[63:0] while_while_acc_1_nl;
  wire[64:0] nl_while_while_acc_1_nl;
  wire[4:0] while_while_acc_3_nl;
  wire[5:0] nl_while_while_acc_3_nl;
  wire[0:0] while_current_buffer_size_not_1_nl;
  wire[4:0] while_current_buffer_size_mux_1_nl;
  wire[4:0] while_while_acc_nl;
  wire[5:0] nl_while_while_acc_nl;
  wire[0:0] while_block_count_not_nl;
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire[32:0] while_while_for_acc_2_nl;
  wire[34:0] nl_while_while_for_acc_2_nl;
  wire[31:0] while_while_for_mul_nl;
  wire[64:0] operator_64_false_1_acc_1_nl;
  wire[65:0] nl_operator_64_false_1_acc_1_nl;
  wire[5:0] while_while_aelse_acc_nl;
  wire[6:0] nl_while_while_aelse_acc_nl;
  wire[5:0] while_while_aelse_acc_1_nl;
  wire[6:0] nl_while_while_aelse_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[4:0] while_while_for_for_address_acc_nl;
  wire[5:0] nl_while_while_for_for_address_acc_nl;
  wire[4:0] while_while_for_for_address_mul_nl;
  wire[9:0] nl_while_while_for_for_address_mul_nl;
  wire [11:0] nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run;
  assign nl_while_while_for_for_address_mul_nl = while_block_count_4_0_sva * block_size_mul_psp_sva;
  assign while_while_for_for_address_mul_nl = nl_while_while_for_for_address_mul_nl[4:0];
  assign nl_while_while_for_for_address_acc_nl = (while_while_for_for_address_mul_nl)
      + (total_blocks_mul_2_itm[4:0]);
  assign while_while_for_for_address_acc_nl = nl_while_while_for_for_address_acc_nl[4:0];
  assign nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run
      = {3'b000 , (while_while_for_for_address_acc_nl) , din_rsci_addr_d_run_3_0_mx1};
  wire [0:0] nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0;
  assign nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0
      = or_dcpl_4;
  wire [0:0] nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0;
  assign nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0
      = ~(while_while_for_stage_0 | while_while_for_stage_0_2);
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1 WeightDoubleBufferReader_384_16_16_run_din_rsci_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_addr_d(din_rsci_addr_d_reg),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .din_rsci_addr_d_run(nl_WeightDoubleBufferReader_384_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run[11:0]),
      .din_rsci_dout_d_mxwt(din_rsci_dout_d_mxwt),
      .din_rsci_oswt_pff(and_41_rmff)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci WeightDoubleBufferReader_384_16_16_run_dout_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .run_wen(run_wen),
      .dout_rsci_oswt(reg_dout_rsci_ivld_run_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_inst
      (
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(reg_din_rsc_rls_obj_ld_run_psct_cse)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_vz(din_rsc_req_vz),
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(reg_din_rsc_req_obj_iswt0_cse),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferReader_384_16_16_run_staller WeightDoubleBufferReader_384_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferReader_384_16_16_run_run_fsm WeightDoubleBufferReader_384_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_2_tr0(exit_while_sva_mx0),
      .while_while_C_0_tr0(nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0[0:0]),
      .while_while_for_C_0_tr0(nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0[0:0]),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign and_41_rmff = or_dcpl_1 & while_while_for_stage_0 & (fsm_output[6]);
  assign din_rsci_addr_d_run_3_0_mx1 = MUX_v_4_2_2(while_while_for_for_r_idx_4_0_lpi_4_3_0,
      (signext_4_1(~ while_while_for_acc_2_itm_32_1)), exitL_exit_while_while_for_for_sva);
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ (readslicef_65_1_64((operator_64_false_acc_1_nl)))),
      (~ operator_64_false_1_acc_1_itm_64_1), fsm_output[8]);
  assign total_blocks_sva_1 = conv_u2u_64_64(total_blocks_mul_1_itm * (reg_paramsIn_crt_sva_127_0_ftd[15:0]));
  assign while_while_for_mul_nl = conv_u2u_32_32((reg_paramsIn_crt_sva_127_0_ftd[47:32])
      * (reg_paramsIn_crt_sva_127_0_ftd[63:48]));
  assign nl_while_while_for_acc_2_nl = ({1'b1 , total_blocks_mul_2_itm}) + conv_u2u_32_33(~
      (while_while_for_mul_nl)) + 33'b000000000000000000000000000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[32:0];
  assign while_while_for_acc_2_itm_32_1 = readslicef_33_1_32((while_while_for_acc_2_nl));
  assign nl_while_while_for_for_acc_tmp = conv_u2u_4_5(din_rsci_addr_d_run_3_0_mx1)
      + 5'b00001;
  assign while_while_for_for_acc_tmp = nl_while_while_for_for_acc_tmp[4:0];
  assign nl_operator_64_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_1_acc_1_nl = nl_operator_64_false_1_acc_1_nl[64:0];
  assign operator_64_false_1_acc_1_itm_64_1 = readslicef_65_1_64((operator_64_false_1_acc_1_nl));
  assign or_dcpl_1 = (~ exitL_exit_while_while_for_for_sva) | while_while_for_acc_2_itm_32_1;
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_5_6(~ while_current_buffer_size_8_4_sva)
      + conv_u2u_5_6(~ block_size_mul_psp_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[5:0];
  assign nl_while_while_aelse_acc_nl = conv_u2u_5_6(readslicef_6_5_1((while_while_aelse_acc_1_nl)))
      + 6'b101101;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[5:0];
  assign or_dcpl_4 = ~(operator_64_false_1_acc_1_itm_64_1 & (~ (readslicef_6_1_5((while_while_aelse_acc_nl)))));
  assign or_tmp_13 = ~((fsm_output[1:0]!=2'b00));
  assign or_tmp_22 = ~((fsm_output[7:5]!=3'b000));
  assign din_rsci_addr_d = din_rsci_addr_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_din_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_din_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_dout_rsci_ivld_run_psct_cse <= 1'b0;
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      block_size_mul_psp_sva <= 5'b00000;
      total_blocks_mul_2_itm <= 32'b00000000000000000000000000000000;
      total_blocks_mul_1_itm <= 48'b000000000000000000000000000000000000000000000000;
      while_block_count_4_0_sva <= 5'b00000;
      while_while_for_stage_0 <= 1'b0;
      exitL_exit_while_while_for_for_sva <= 1'b0;
      while_while_for_stage_0_2 <= 1'b0;
      reg_paramsIn_crt_sva_127_0_ftd <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_din_rsc_req_obj_iswt0_cse <= ~(exit_while_sva_mx0 | (~((fsm_output[3])
          | (fsm_output[8]))));
      reg_din_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_4 & (fsm_output[5]);
      reg_dout_rsci_ivld_run_psct_cse <= while_while_for_stage_0_2 & (~ exit_while_while_for_lpi_4_dfm_st_1)
          & (fsm_output[6]);
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse <= and_41_rmff;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[3]) | (fsm_output[8])
          | (fsm_output[0]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      block_size_mul_psp_sva <= MUX_v_5_2_2((block_size_mul_nl), block_size_mul_psp_sva,
          or_tmp_13);
      total_blocks_mul_2_itm <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (total_blocks_mux1h_2_nl), (not_nl));
      total_blocks_mul_1_itm <= conv_u2u_48_48(total_blocks_mul_2_itm * (reg_paramsIn_crt_sva_127_0_ftd[31:16]));
      while_block_count_4_0_sva <= MUX_v_5_2_2(5'b00000, (while_current_buffer_size_mux_1_nl),
          (while_block_count_not_nl));
      while_while_for_stage_0 <= ~((~(while_while_for_stage_0 & or_dcpl_1)) & (fsm_output[6]));
      exitL_exit_while_while_for_for_sva <= (while_while_for_for_acc_tmp[4]) | (~
          (fsm_output[6]));
      while_while_for_stage_0_2 <= while_while_for_stage_0 & (fsm_output[6]);
      reg_paramsIn_crt_sva_127_0_ftd <= MUX_v_64_2_2((paramsIn_rsci_idat_mxwt[95:32]),
          reg_paramsIn_crt_sva_127_0_ftd, or_tmp_13);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_idat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ (fsm_output[6])) | (~ while_while_for_stage_0_2) |
        exit_while_while_for_lpi_4_dfm_st_1)) ) begin
      dout_rsci_idat <= din_rsci_dout_d_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[5]) |
        (fsm_output[8]))) ) begin
      total_blocks_lpi_3 <= MUX_v_64_2_2(total_blocks_sva_1, (while_while_acc_1_nl),
          fsm_output[7]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_current_buffer_size_8_4_sva <= 5'b00000;
    end
    else if ( (fsm_output[6:5]==2'b00) & run_wen ) begin
      while_current_buffer_size_8_4_sva <= MUX_v_5_2_2(5'b00000, (while_while_acc_3_nl),
          (while_current_buffer_size_not_1_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_while_while_for_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen & while_while_for_stage_0 ) begin
      exit_while_while_for_lpi_4_dfm_st_1 <= (~ while_while_for_acc_2_itm_32_1) &
          exitL_exit_while_while_for_for_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_r_idx_4_0_lpi_4_3_0 <= 4'b0000;
    end
    else if ( run_wen & or_dcpl_1 & while_while_for_stage_0 & (~ (while_while_for_for_acc_tmp[4]))
        ) begin
      while_while_for_for_r_idx_4_0_lpi_4_3_0 <= while_while_for_for_acc_tmp[3:0];
    end
  end
  assign nl_block_size_mul_nl = (paramsIn_rsci_idat_mxwt[84:80]) * (paramsIn_rsci_idat_mxwt[68:64]);
  assign block_size_mul_nl = nl_block_size_mul_nl[4:0];
  assign total_blocks_mul_2_nl = conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16])
      * (paramsIn_rsci_idat_mxwt[15:0]));
  assign nl_while_while_for_acc_1_nl = total_blocks_mul_2_itm + 32'b00000000000000000000000000000001;
  assign while_while_for_acc_1_nl = nl_while_while_for_acc_1_nl[31:0];
  assign total_blocks_and_1_nl = (~ (while_while_for_for_acc_tmp[4])) & (fsm_output[6]);
  assign total_blocks_and_2_nl = (while_while_for_for_acc_tmp[4]) & (fsm_output[6]);
  assign total_blocks_mux1h_2_nl = MUX1HOT_v_32_3_2((total_blocks_mul_2_nl), total_blocks_mul_2_itm,
      (while_while_for_acc_1_nl), {(fsm_output[1]) , (total_blocks_and_1_nl) , (total_blocks_and_2_nl)});
  assign not_nl = ~ (fsm_output[5]);
  assign nl_while_while_acc_nl = while_block_count_4_0_sva + 5'b00001;
  assign while_while_acc_nl = nl_while_while_acc_nl[4:0];
  assign while_current_buffer_size_mux_1_nl = MUX_v_5_2_2(while_block_count_4_0_sva,
      (while_while_acc_nl), fsm_output[7]);
  assign while_block_count_not_nl = ~ or_tmp_22;
  assign nl_while_while_acc_1_nl = total_blocks_lpi_3 + 64'b1111111111111111111111111111111111111111111111111111111111111111;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[63:0];
  assign nl_while_while_acc_3_nl = while_current_buffer_size_8_4_sva + block_size_mul_psp_sva;
  assign while_while_acc_3_nl = nl_while_while_acc_3_nl[4:0];
  assign while_current_buffer_size_not_1_nl = ~ or_tmp_22;

  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_6_5_1;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_6_5_1 = tmp[4:0];
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction


  function automatic [63:0] conv_u2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_64 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, weightDoubleBufferWriterParams_cns_dat,
      weightDoubleBufferWriterParams_cns_vld, weightDoubleBufferWriterParams_cns_rdy,
      weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;



  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBuffer_384_16_16_run_run WeightDoubleBuffer_384_16_16_run_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_csb, dout_rsc_web, dout_rsc_addr, dout_rsc_din,
      dout_rsc_dout, dout_rsc_req_vz, dout_rsc_rls_lz
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output dout_rsc_csb;
  output dout_rsc_web;
  output [11:0] dout_rsc_addr;
  output [127:0] dout_rsc_din;
  input [127:0] dout_rsc_dout;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;


  // Interconnect Declarations
  wire [11:0] dout_rsci_addr_d;
  wire [127:0] dout_rsci_din_d;
  wire [127:0] dout_rsci_dout_d;
  wire dout_rsci_web_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  assign nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = ~ dout_rsci_web_d_iff;
  WeightDoubleBufferWriter_384_16_16_sram_512_128_sram_512_128_rwport_3_128_12_384_128_gen
      dout_rsci (
      .dout(dout_rsc_dout),
      .din(dout_rsc_din),
      .addr(dout_rsc_addr),
      .web(dout_rsc_web),
      .csb(dout_rsc_csb),
      .web_d(dout_rsci_web_d_iff),
      .addr_d(dout_rsci_addr_d),
      .din_d(dout_rsci_din_d),
      .dout_d(dout_rsci_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d[0:0])
    );
  WeightDoubleBufferWriter_384_16_16_run WeightDoubleBufferWriter_384_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .dout_rsci_addr_d(dout_rsci_addr_d),
      .dout_rsci_din_d(dout_rsci_din_d),
      .dout_rsci_web_d_pff(dout_rsci_web_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_csb,
      din_rsc_web, din_rsc_addr, din_rsc_din, din_rsc_dout, din_rsc_req_vz, din_rsc_rls_lz,
      dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output din_rsc_csb;
  output din_rsc_web;
  output [11:0] din_rsc_addr;
  output [127:0] din_rsc_din;
  input [127:0] din_rsc_dout;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [11:0] din_rsci_addr_d;
  wire [127:0] din_rsci_dout_d;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferReader_384_16_16_sram_512_128_sram_512_128_rwport_8_128_12_384_128_gen
      din_rsci (
      .dout(din_rsc_dout),
      .din(din_rsc_din),
      .addr(din_rsc_addr),
      .web(din_rsc_web),
      .csb(din_rsc_csb),
      .web_d(1'b1),
      .addr_d(din_rsci_addr_d),
      .din_d(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .dout_d(din_rsci_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  WeightDoubleBufferReader_384_16_16_run WeightDoubleBufferReader_384_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_req_vz(din_rsc_req_vz),
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .din_rsci_addr_d(din_rsci_addr_d),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_struct
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_struct (
  clk, arst_n, weights_in_rsc_dat_value, weights_in_rsc_vld, weights_in_rsc_rdy,
      weights_out_rsc_dat_value, weights_out_rsc_vld, weights_out_rsc_rdy, paramsIn_rsc_dat_STRIDE,
      paramsIn_rsc_dat_FY, paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1, paramsIn_rsc_dat_OC1,
      paramsIn_rsc_dat_OX0, paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1, paramsIn_rsc_dat_OY1,
      paramsIn_rsc_vld, paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] weights_in_rsc_dat_value;
  input weights_in_rsc_vld;
  output weights_in_rsc_rdy;
  output [127:0] weights_out_rsc_dat_value;
  output weights_out_rsc_vld;
  input weights_out_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBufferWriter;
  wire paramsIn_rsc_vld_nweightDoubleBufferWriter;
  wire paramsIn_rsc_rdy_nweightDoubleBufferWriter;
  wire din_rsc_rdy_nweightDoubleBufferWriter;
  wire dout_rsc_csb_nweightDoubleBufferWriter;
  wire dout_rsc_web_nweightDoubleBufferWriter;
  wire [11:0] dout_rsc_addr_nweightDoubleBufferWriter;
  wire [127:0] dout_rsc_din_nweightDoubleBufferWriter;
  wire [127:0] dout_rsc_dout_nweightDoubleBufferWriter;
  wire dout_rsc_req_vz_nweightDoubleBufferWriter;
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBufferReader;
  wire paramsIn_rsc_vld_nweightDoubleBufferReader;
  wire paramsIn_rsc_rdy_nweightDoubleBufferReader;
  wire din_rsc_csb_nweightDoubleBufferReader;
  wire din_rsc_web_nweightDoubleBufferReader;
  wire [11:0] din_rsc_addr_nweightDoubleBufferReader;
  wire [127:0] din_rsc_din_nweightDoubleBufferReader;
  wire [127:0] din_rsc_dout_nweightDoubleBufferReader;
  wire din_rsc_req_vz_nweightDoubleBufferReader;
  wire [127:0] dout_rsc_dat_nweightDoubleBufferReader;
  wire dout_rsc_vld_nweightDoubleBufferReader;
  wire [143:0] weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst;
  wire weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst;
  wire [143:0] weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst;
  wire weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst;
  wire paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  wire weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire din_rsc_rdy_nweightDoubleBufferWriter_bud;
  wire dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  wire din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  wire weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire dout_rsc_vld_nweightDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire weightDoubleBufferWriterParams_unc_2;
  wire weightDoubleBufferWriterParams_idle;
  wire mem_cns_R0;
  wire mem_cns_R1;
  wire mem_cns_csb_shi0;
  wire mem_cns_csb_shi1;
  wire mem_cns_web_shi0;
  wire mem_cns_web_shi1;
  wire [11:0] mem_cns_addr_shi0;
  wire [11:0] mem_cns_addr_shi1;
  wire [127:0] mem_cns_din_shi0;
  wire [127:0] mem_cns_din_shi1;
  wire [127:0] mem_cns_dout_sho0;
  wire [127:0] mem_cns_dout_sho1;
  wire weightDoubleBufferReaderParams_unc_2;
  wire weightDoubleBufferReaderParams_idle;
  wire mem_cns_S1_iff;
  wire mem_cns_S0_iff;
  wire mem_cns_S0_dmo;
  wire mem_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat = {paramsIn_rsc_dat_STRIDE
      , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1 , paramsIn_rsc_dat_OC1
      , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1 , paramsIn_rsc_dat_OY1};
  ccs_pipe_v5 #(.rscid(32'sd15),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferWriterParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .din_vld(weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .din(weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBufferWriter),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBufferWriter),
      .dout(paramsIn_rsc_dat_nweightDoubleBufferWriter),
      .sz(weightDoubleBufferWriterParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferWriterParams_idle)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd128),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) mem_cns_comp (
      .clk(clk),
      .csb(mem_cns_csb_shi0),
      .web(mem_cns_web_shi0),
      .addr(mem_cns_addr_shi0),
      .din(mem_cns_din_shi0),
      .dout(mem_cns_dout_sho0)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd128),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) mem_cns_comp_1 (
      .clk(clk),
      .csb(mem_cns_csb_shi1),
      .web(mem_cns_web_shi1),
      .addr(mem_cns_addr_shi1),
      .din(mem_cns_din_shi1),
      .dout(mem_cns_dout_sho1)
    );
  ccs_pipe_v5 #(.rscid(32'sd16),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferReaderParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .din_vld(weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .din(weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBufferReader),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBufferReader),
      .dout(paramsIn_rsc_dat_nweightDoubleBufferReader),
      .sz(weightDoubleBufferReaderParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferReaderParams_idle)
    );
  WeightDoubleBufferWriter_384_16_16 weightDoubleBufferWriter (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBufferWriter),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBufferWriter),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud),
      .din_rsc_dat(weights_in_rsc_dat_value),
      .din_rsc_vld(weights_in_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy_nweightDoubleBufferWriter_bud),
      .dout_rsc_csb(dout_rsc_csb_nweightDoubleBufferWriter),
      .dout_rsc_web(dout_rsc_web_nweightDoubleBufferWriter),
      .dout_rsc_addr(dout_rsc_addr_nweightDoubleBufferWriter),
      .dout_rsc_din(dout_rsc_din_nweightDoubleBufferWriter),
      .dout_rsc_dout(dout_rsc_dout_nweightDoubleBufferWriter),
      .dout_rsc_req_vz(dout_rsc_req_vz_nweightDoubleBufferWriter),
      .dout_rsc_rls_lz(dout_rsc_rls_lz_nweightDoubleBufferWriter_bud)
    );
  WeightDoubleBufferReader_384_16_16 weightDoubleBufferReader (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBufferReader),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBufferReader),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBufferReader_bud),
      .din_rsc_csb(din_rsc_csb_nweightDoubleBufferReader),
      .din_rsc_web(din_rsc_web_nweightDoubleBufferReader),
      .din_rsc_addr(din_rsc_addr_nweightDoubleBufferReader),
      .din_rsc_din(din_rsc_din_nweightDoubleBufferReader),
      .din_rsc_dout(din_rsc_dout_nweightDoubleBufferReader),
      .din_rsc_req_vz(din_rsc_req_vz_nweightDoubleBufferReader),
      .din_rsc_rls_lz(din_rsc_rls_lz_nweightDoubleBufferReader_bud),
      .dout_rsc_dat(dout_rsc_dat_nweightDoubleBufferReader),
      .dout_rsc_vld(dout_rsc_vld_nweightDoubleBufferReader_bud),
      .dout_rsc_rdy(weights_out_rsc_rdy)
    );
  WeightDoubleBuffer_384_16_16_run WeightDoubleBuffer_384_16_16_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst)
    );
  unreg_hier unreg (
      .in_0(mem_cns_S0_iff),
      .out_0(mem_cns_R0)
    );
  unreg_hier unreg_1 (
      .in_0(mem_cns_S1_iff),
      .out_0(mem_cns_R1)
    );
  WeightDoublefeSAqem_cns_bctl WeightDoublefeSAqem_cns_bctl_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_rdy_nweightDoubleBufferWriter(paramsIn_rsc_rdy_nweightDoubleBufferWriter),
      .din_rsc_rdy_nweightDoubleBufferWriter(din_rsc_rdy_nweightDoubleBufferWriter),
      .dout_rsc_csb_nweightDoubleBufferWriter(dout_rsc_csb_nweightDoubleBufferWriter),
      .dout_rsc_web_nweightDoubleBufferWriter(dout_rsc_web_nweightDoubleBufferWriter),
      .dout_rsc_addr_nweightDoubleBufferWriter(dout_rsc_addr_nweightDoubleBufferWriter),
      .dout_rsc_din_nweightDoubleBufferWriter(dout_rsc_din_nweightDoubleBufferWriter),
      .dout_rsc_dout_nweightDoubleBufferWriter(dout_rsc_dout_nweightDoubleBufferWriter),
      .dout_rsc_req_vz_nweightDoubleBufferWriter(dout_rsc_req_vz_nweightDoubleBufferWriter),
      .paramsIn_rsc_rdy_nweightDoubleBufferReader(paramsIn_rsc_rdy_nweightDoubleBufferReader),
      .din_rsc_csb_nweightDoubleBufferReader(din_rsc_csb_nweightDoubleBufferReader),
      .din_rsc_web_nweightDoubleBufferReader(din_rsc_web_nweightDoubleBufferReader),
      .din_rsc_addr_nweightDoubleBufferReader(din_rsc_addr_nweightDoubleBufferReader),
      .din_rsc_din_nweightDoubleBufferReader(din_rsc_din_nweightDoubleBufferReader),
      .din_rsc_dout_nweightDoubleBufferReader(din_rsc_dout_nweightDoubleBufferReader),
      .din_rsc_req_vz_nweightDoubleBufferReader(din_rsc_req_vz_nweightDoubleBufferReader),
      .dout_rsc_vld_nweightDoubleBufferReader(dout_rsc_vld_nweightDoubleBufferReader),
      .paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud(paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud),
      .din_rsc_rdy_nweightDoubleBufferWriter_bud(din_rsc_rdy_nweightDoubleBufferWriter_bud),
      .dout_rsc_rls_lz_nweightDoubleBufferWriter_bud(dout_rsc_rls_lz_nweightDoubleBufferWriter_bud),
      .din_rsc_rls_lz_nweightDoubleBufferReader_bud(din_rsc_rls_lz_nweightDoubleBufferReader_bud),
      .paramsIn_rsc_rdy_nweightDoubleBufferReader_bud(paramsIn_rsc_rdy_nweightDoubleBufferReader_bud),
      .dout_rsc_vld_nweightDoubleBufferReader_bud(dout_rsc_vld_nweightDoubleBufferReader_bud),
      .mem_cns_S0(mem_cns_S0_dmo),
      .mem_cns_R0(mem_cns_R0),
      .mem_cns_S1(mem_cns_S1_dmo),
      .mem_cns_R1(mem_cns_R1),
      .mem_cns_csb_shi0(mem_cns_csb_shi0),
      .mem_cns_csb_shi1(mem_cns_csb_shi1),
      .mem_cns_web_shi0(mem_cns_web_shi0),
      .mem_cns_web_shi1(mem_cns_web_shi1),
      .mem_cns_addr_shi0(mem_cns_addr_shi0),
      .mem_cns_addr_shi1(mem_cns_addr_shi1),
      .mem_cns_din_shi0(mem_cns_din_shi0),
      .mem_cns_din_shi1(mem_cns_din_shi1),
      .mem_cns_dout_sho0(mem_cns_dout_sho0),
      .mem_cns_dout_sho1(mem_cns_dout_sho1),
      .mem_cns_S1_pff(mem_cns_S1_iff),
      .mem_cns_S0_pff(mem_cns_S0_iff)
    );
  assign weights_out_rsc_dat_value = dout_rsc_dat_nweightDoubleBufferReader;
  assign weights_in_rsc_rdy = din_rsc_rdy_nweightDoubleBufferWriter;
  assign weights_out_rsc_vld = dout_rsc_vld_nweightDoubleBufferReader;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16 (
  clk, arst_n, weights_in_rsc_dat, weights_in_rsc_vld, weights_in_rsc_rdy, weights_out_rsc_dat,
      weights_out_rsc_vld, weights_out_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] weights_in_rsc_dat;
  input weights_in_rsc_vld;
  output weights_in_rsc_rdy;
  output [127:0] weights_out_rsc_dat;
  output weights_out_rsc_vld;
  input weights_out_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [127:0] weights_out_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1 = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1 = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0 = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0 = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1 = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1 = paramsIn_rsc_dat[15:0];
  WeightDoubleBuffer_384_16_16_struct WeightDoubleBuffer_384_16_16_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .weights_in_rsc_dat_value(weights_in_rsc_dat),
      .weights_in_rsc_vld(weights_in_rsc_vld),
      .weights_in_rsc_rdy(weights_in_rsc_rdy),
      .weights_out_rsc_dat_value(weights_out_rsc_dat_value),
      .weights_out_rsc_vld(weights_out_rsc_vld),
      .weights_out_rsc_rdy(weights_out_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy)
    );
  assign weights_out_rsc_dat = weights_out_rsc_dat_value;
endmodule




//------> ../InputDoubleBufferless_512comma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy07
//  Generated date: Sun Feb 23 19:20:44 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBDjtfoem_cns_bctl
// ------------------------------------------------------------------


module InputDoubleBDjtfoem_cns_bctl (
  clk, arst_n, paramsIn_rsc_rdy_ninputDoubleBufferWriter, din_rsc_rdy_ninputDoubleBufferWriter,
      dout_rsc_csb_ninputDoubleBufferWriter, dout_rsc_web_ninputDoubleBufferWriter,
      dout_rsc_addr_ninputDoubleBufferWriter, dout_rsc_din_ninputDoubleBufferWriter,
      dout_rsc_dout_ninputDoubleBufferWriter, dout_rsc_req_vz_ninputDoubleBufferWriter,
      paramsIn_rsc_rdy_ninputDoubleBufferReader, din_rsc_csb_ninputDoubleBufferReader,
      din_rsc_web_ninputDoubleBufferReader, din_rsc_addr_ninputDoubleBufferReader,
      din_rsc_din_ninputDoubleBufferReader, din_rsc_dout_ninputDoubleBufferReader,
      din_rsc_req_vz_ninputDoubleBufferReader, dout_rsc_vld_ninputDoubleBufferReader,
      paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud, din_rsc_rdy_ninputDoubleBufferWriter_bud,
      dout_rsc_rls_lz_ninputDoubleBufferWriter_bud, din_rsc_rls_lz_ninputDoubleBufferReader_bud,
      paramsIn_rsc_rdy_ninputDoubleBufferReader_bud, dout_rsc_vld_ninputDoubleBufferReader_bud,
      mem_cns_S0, mem_cns_R0, mem_cns_S1, mem_cns_R1, mem_cns_csb_shi0, mem_cns_csb_shi1,
      mem_cns_web_shi0, mem_cns_web_shi1, mem_cns_addr_shi0, mem_cns_addr_shi1, mem_cns_din_shi0,
      mem_cns_din_shi1, mem_cns_dout_sho0, mem_cns_dout_sho1, mem_cns_S1_pff, mem_cns_S0_pff
);
  input clk;
  input arst_n;
  output paramsIn_rsc_rdy_ninputDoubleBufferWriter;
  output din_rsc_rdy_ninputDoubleBufferWriter;
  input dout_rsc_csb_ninputDoubleBufferWriter;
  input dout_rsc_web_ninputDoubleBufferWriter;
  input [11:0] dout_rsc_addr_ninputDoubleBufferWriter;
  input [127:0] dout_rsc_din_ninputDoubleBufferWriter;
  output [127:0] dout_rsc_dout_ninputDoubleBufferWriter;
  output dout_rsc_req_vz_ninputDoubleBufferWriter;
  output paramsIn_rsc_rdy_ninputDoubleBufferReader;
  input din_rsc_csb_ninputDoubleBufferReader;
  input din_rsc_web_ninputDoubleBufferReader;
  input [11:0] din_rsc_addr_ninputDoubleBufferReader;
  input [127:0] din_rsc_din_ninputDoubleBufferReader;
  output [127:0] din_rsc_dout_ninputDoubleBufferReader;
  output din_rsc_req_vz_ninputDoubleBufferReader;
  output dout_rsc_vld_ninputDoubleBufferReader;
  input paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  input din_rsc_rdy_ninputDoubleBufferWriter_bud;
  input dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  input din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  input paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  input dout_rsc_vld_ninputDoubleBufferReader_bud;
  output mem_cns_S0;
  input mem_cns_R0;
  output mem_cns_S1;
  input mem_cns_R1;
  output mem_cns_csb_shi0;
  output mem_cns_csb_shi1;
  output mem_cns_web_shi0;
  output mem_cns_web_shi1;
  output [11:0] mem_cns_addr_shi0;
  output [11:0] mem_cns_addr_shi1;
  output [127:0] mem_cns_din_shi0;
  output [127:0] mem_cns_din_shi1;
  input [127:0] mem_cns_dout_sho0;
  input [127:0] mem_cns_dout_sho1;
  output mem_cns_S1_pff;
  output mem_cns_S0_pff;


  // Interconnect Declarations
  wire mem_cns_PC0;
  reg mem_cns_ppidx;
  reg [1:0] mem_cns_ppown;
  wire mem_cns_PC1;
  reg mem_cns_ppidx_1;
  reg [1:0] mem_cns_ppown_1;
  wire mem_cns_ppsel_1_pff;
  wire [1:0] mem_acc_1_rmff;
  wire [3:0] nl_mem_acc_1_rmff;
  wire mem_xor_1_rmff;
  wire mem_or_cse_pff;
  wire [1:0] mem_acc_rmff;
  wire [3:0] nl_mem_acc_rmff;
  wire mem_xor_rmff;
  wire mem_cns_ppsel_3_pff;
  wire mem_or_6_cse_pff;

  wire[0:0] mem_mux_11_nl;
  wire[0:0] mem_mux_13_nl;
  wire[0:0] mem_mux_10_nl;
  wire[0:0] mem_mux_12_nl;

  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsc_rdy_ninputDoubleBufferWriter = paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  assign din_rsc_rdy_ninputDoubleBufferWriter = din_rsc_rdy_ninputDoubleBufferWriter_bud;
  assign paramsIn_rsc_rdy_ninputDoubleBufferReader = paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  assign dout_rsc_vld_ninputDoubleBufferReader = dout_rsc_vld_ninputDoubleBufferReader_bud;
  assign dout_rsc_req_vz_ninputDoubleBufferWriter = mem_cns_R0;
  assign din_rsc_req_vz_ninputDoubleBufferReader = mem_cns_R1;
  assign mem_xor_rmff = mem_cns_ppidx ^ mem_cns_PC0;
  assign nl_mem_acc_rmff = mem_cns_ppown + conv_u2u_1_2(mem_cns_PC0) + conv_s2u_1_2(mem_cns_PC1);
  assign mem_acc_rmff = nl_mem_acc_rmff[1:0];
  assign mem_cns_PC0 = mem_cns_S0 & dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  assign mem_xor_1_rmff = mem_cns_ppidx_1 ^ mem_cns_PC1;
  assign nl_mem_acc_1_rmff = mem_cns_ppown_1 + conv_u2u_1_2(mem_cns_PC1) + conv_s2u_1_2(mem_cns_PC0);
  assign mem_acc_1_rmff = nl_mem_acc_1_rmff[1:0];
  assign mem_cns_PC1 = mem_cns_S1 & din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  assign dout_rsc_dout_ninputDoubleBufferWriter = MUX_v_128_2_2(mem_cns_dout_sho0,
      mem_cns_dout_sho1, mem_cns_ppidx);
  assign din_rsc_dout_ninputDoubleBufferReader = MUX_v_128_2_2(mem_cns_dout_sho0,
      mem_cns_dout_sho1, mem_cns_ppidx_1);
  assign mem_mux_11_nl = MUX_s_1_2_2((~ dout_rsc_csb_ninputDoubleBufferWriter), (~
      din_rsc_csb_ninputDoubleBufferReader), mem_cns_ppsel_1_pff);
  assign mem_cns_csb_shi0 = ~((mem_mux_11_nl) & mem_or_cse_pff);
  assign mem_cns_S1 = (mem_cns_ppown_1!=2'b00);
  assign mem_cns_S1_pff = (mem_acc_1_rmff!=2'b00);
  assign mem_cns_ppsel_1_pff = mem_cns_S1_pff & (~ mem_xor_1_rmff);
  assign mem_cns_S0 = ~((mem_cns_ppown==2'b10));
  assign mem_cns_S0_pff = ~((mem_acc_rmff==2'b10));
  assign mem_or_cse_pff = (mem_cns_S0_pff & (~ mem_xor_rmff)) | mem_cns_ppsel_1_pff;
  assign mem_mux_13_nl = MUX_s_1_2_2((~ dout_rsc_web_ninputDoubleBufferWriter), (~
      din_rsc_web_ninputDoubleBufferReader), mem_cns_ppsel_1_pff);
  assign mem_cns_web_shi0 = ~((mem_mux_13_nl) & mem_or_cse_pff);
  assign mem_cns_addr_shi0 = MUX_v_12_2_2(dout_rsc_addr_ninputDoubleBufferWriter,
      din_rsc_addr_ninputDoubleBufferReader, mem_cns_ppsel_1_pff);
  assign mem_cns_din_shi0 = MUX_v_128_2_2(dout_rsc_din_ninputDoubleBufferWriter,
      din_rsc_din_ninputDoubleBufferReader, mem_cns_ppsel_1_pff);
  assign mem_mux_10_nl = MUX_s_1_2_2((~ dout_rsc_csb_ninputDoubleBufferWriter), (~
      din_rsc_csb_ninputDoubleBufferReader), mem_cns_ppsel_3_pff);
  assign mem_cns_csb_shi1 = ~((mem_mux_10_nl) & mem_or_6_cse_pff);
  assign mem_cns_ppsel_3_pff = mem_cns_S1_pff & mem_xor_1_rmff;
  assign mem_or_6_cse_pff = (mem_cns_S0_pff & mem_xor_rmff) | mem_cns_ppsel_3_pff;
  assign mem_mux_12_nl = MUX_s_1_2_2((~ dout_rsc_web_ninputDoubleBufferWriter), (~
      din_rsc_web_ninputDoubleBufferReader), mem_cns_ppsel_3_pff);
  assign mem_cns_web_shi1 = ~((mem_mux_12_nl) & mem_or_6_cse_pff);
  assign mem_cns_addr_shi1 = MUX_v_12_2_2(dout_rsc_addr_ninputDoubleBufferWriter,
      din_rsc_addr_ninputDoubleBufferReader, mem_cns_ppsel_3_pff);
  assign mem_cns_din_shi1 = MUX_v_128_2_2(dout_rsc_din_ninputDoubleBufferWriter,
      din_rsc_din_ninputDoubleBufferReader, mem_cns_ppsel_3_pff);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mem_cns_ppidx <= 1'b0;
      mem_cns_ppown <= 2'b00;
      mem_cns_ppidx_1 <= 1'b0;
      mem_cns_ppown_1 <= 2'b00;
    end
    else begin
      mem_cns_ppidx <= mem_xor_rmff;
      mem_cns_ppown <= mem_acc_rmff;
      mem_cns_ppidx_1 <= mem_xor_1_rmff;
      mem_cns_ppown_1 <= mem_acc_1_rmff;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier
// ------------------------------------------------------------------

/*
module unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule
*/
// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for InputDoubleBuffer_512_16_16_run_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBuffer_512_16_16_run_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_staller
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_staller (
  run_wen, paramsIn_rsci_wen_comp, inputDoubleBufferWriterParams_cnsi_wen_comp, inputDoubleBufferReaderParams_cnsi_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input inputDoubleBufferWriterParams_cnsi_wen_comp;
  input inputDoubleBufferReaderParams_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & inputDoubleBufferWriterParams_cnsi_wen_comp
      & inputDoubleBufferReaderParams_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
    (
  clk, arst_n, inputDoubleBufferReaderParams_cnsi_oswt, inputDoubleBufferReaderParams_cnsi_wen_comp,
      inputDoubleBufferReaderParams_cnsi_biwt, inputDoubleBufferReaderParams_cnsi_bdwt,
      inputDoubleBufferReaderParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  output inputDoubleBufferReaderParams_cnsi_wen_comp;
  input inputDoubleBufferReaderParams_cnsi_biwt;
  input inputDoubleBufferReaderParams_cnsi_bdwt;
  output inputDoubleBufferReaderParams_cnsi_bcwt;
  reg inputDoubleBufferReaderParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferReaderParams_cnsi_wen_comp = (~ inputDoubleBufferReaderParams_cnsi_oswt)
      | inputDoubleBufferReaderParams_cnsi_biwt | inputDoubleBufferReaderParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputDoubleBufferReaderParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      inputDoubleBufferReaderParams_cnsi_bcwt <= ~((~(inputDoubleBufferReaderParams_cnsi_bcwt
          | inputDoubleBufferReaderParams_cnsi_biwt)) | inputDoubleBufferReaderParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
    (
  run_wen, inputDoubleBufferReaderParams_cnsi_oswt, inputDoubleBufferReaderParams_cnsi_irdy,
      inputDoubleBufferReaderParams_cnsi_biwt, inputDoubleBufferReaderParams_cnsi_bdwt,
      inputDoubleBufferReaderParams_cnsi_bcwt, inputDoubleBufferReaderParams_cnsi_ivld_run_sct
);
  input run_wen;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  input inputDoubleBufferReaderParams_cnsi_irdy;
  output inputDoubleBufferReaderParams_cnsi_biwt;
  output inputDoubleBufferReaderParams_cnsi_bdwt;
  input inputDoubleBufferReaderParams_cnsi_bcwt;
  output inputDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire inputDoubleBufferReaderParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferReaderParams_cnsi_bdwt = inputDoubleBufferReaderParams_cnsi_oswt
      & run_wen;
  assign inputDoubleBufferReaderParams_cnsi_biwt = inputDoubleBufferReaderParams_cnsi_ogwt
      & inputDoubleBufferReaderParams_cnsi_irdy;
  assign inputDoubleBufferReaderParams_cnsi_ogwt = inputDoubleBufferReaderParams_cnsi_oswt
      & (~ inputDoubleBufferReaderParams_cnsi_bcwt);
  assign inputDoubleBufferReaderParams_cnsi_ivld_run_sct = inputDoubleBufferReaderParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
    (
  clk, arst_n, inputDoubleBufferWriterParams_cnsi_oswt, inputDoubleBufferWriterParams_cnsi_wen_comp,
      inputDoubleBufferWriterParams_cnsi_biwt, inputDoubleBufferWriterParams_cnsi_bdwt,
      inputDoubleBufferWriterParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  output inputDoubleBufferWriterParams_cnsi_wen_comp;
  input inputDoubleBufferWriterParams_cnsi_biwt;
  input inputDoubleBufferWriterParams_cnsi_bdwt;
  output inputDoubleBufferWriterParams_cnsi_bcwt;
  reg inputDoubleBufferWriterParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferWriterParams_cnsi_wen_comp = (~ inputDoubleBufferWriterParams_cnsi_oswt)
      | inputDoubleBufferWriterParams_cnsi_biwt | inputDoubleBufferWriterParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputDoubleBufferWriterParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      inputDoubleBufferWriterParams_cnsi_bcwt <= ~((~(inputDoubleBufferWriterParams_cnsi_bcwt
          | inputDoubleBufferWriterParams_cnsi_biwt)) | inputDoubleBufferWriterParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
    (
  run_wen, inputDoubleBufferWriterParams_cnsi_oswt, inputDoubleBufferWriterParams_cnsi_irdy,
      inputDoubleBufferWriterParams_cnsi_biwt, inputDoubleBufferWriterParams_cnsi_bdwt,
      inputDoubleBufferWriterParams_cnsi_bcwt, inputDoubleBufferWriterParams_cnsi_ivld_run_sct
);
  input run_wen;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  input inputDoubleBufferWriterParams_cnsi_irdy;
  output inputDoubleBufferWriterParams_cnsi_biwt;
  output inputDoubleBufferWriterParams_cnsi_bdwt;
  input inputDoubleBufferWriterParams_cnsi_bcwt;
  output inputDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire inputDoubleBufferWriterParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferWriterParams_cnsi_bdwt = inputDoubleBufferWriterParams_cnsi_oswt
      & run_wen;
  assign inputDoubleBufferWriterParams_cnsi_biwt = inputDoubleBufferWriterParams_cnsi_ogwt
      & inputDoubleBufferWriterParams_cnsi_irdy;
  assign inputDoubleBufferWriterParams_cnsi_ogwt = inputDoubleBufferWriterParams_cnsi_oswt
      & (~ inputDoubleBufferWriterParams_cnsi_bcwt);
  assign inputDoubleBufferWriterParams_cnsi_ivld_run_sct = inputDoubleBufferWriterParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_sram_512_128_sram_512_128_rwport_3_128_12_512_128_gen
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_sram_512_128_sram_512_128_rwport_3_128_12_512_128_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [127:0] dout;
  output [127:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [127:0] din_d;
  output [127:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire dout_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign dout_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (dout_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_5_tr0, while_while_C_1_tr0, while_while_C_2_tr0,
      while_while_for_for_C_0_tr0, while_while_for_C_1_tr0, while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [15:0] fsm_output;
  reg [15:0] fsm_output;
  input main_C_5_tr0;
  input while_while_C_1_tr0;
  input while_while_C_2_tr0;
  input while_while_for_for_C_0_tr0;
  input while_while_for_C_1_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for InputDoubleBufferWriter_512_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    while_C_0 = 4'd7,
    while_while_C_0 = 4'd8,
    while_while_C_1 = 4'd9,
    while_while_C_2 = 4'd10,
    while_while_for_for_C_0 = 4'd11,
    while_while_for_C_0 = 4'd12,
    while_while_for_C_1 = 4'd13,
    while_while_C_3 = 4'd14,
    while_C_1 = 4'd15;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBufferWriter_512_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 16'b0000000000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 16'b0000000000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 16'b0000000000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 16'b0000000000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 16'b0000000000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 16'b0000000001000000;
        if ( main_C_5_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 16'b0000000010000000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 16'b0000000100000000;
        state_var_NS = while_while_C_1;
      end
      while_while_C_1 : begin
        fsm_output = 16'b0000001000000000;
        if ( while_while_C_1_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_C_2;
        end
      end
      while_while_C_2 : begin
        fsm_output = 16'b0000010000000000;
        if ( while_while_C_2_tr0 ) begin
          state_var_NS = while_while_C_3;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_for_C_0 : begin
        fsm_output = 16'b0000100000000000;
        if ( while_while_for_for_C_0_tr0 ) begin
          state_var_NS = while_while_for_C_0;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 16'b0001000000000000;
        state_var_NS = while_while_for_C_1;
      end
      while_while_for_C_1 : begin
        fsm_output = 16'b0010000000000000;
        if ( while_while_for_C_1_tr0 ) begin
          state_var_NS = while_while_C_3;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_C_3 : begin
        fsm_output = 16'b0100000000000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 16'b1000000000000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 16'b0000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_staller
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, din_rsci_wen_comp, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input din_rsci_wen_comp;
  input dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & din_rsci_wen_comp & dout_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
    (
  clk, arst_n, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt, dout_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;
  input dout_rsc_req_obj_biwt;
  input dout_rsc_req_obj_bdwt;
  output dout_rsc_req_obj_bcwt;
  reg dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_wen_comp = (~ dout_rsc_req_obj_oswt) | dout_rsc_req_obj_biwt
      | dout_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_bcwt <= ~((~(dout_rsc_req_obj_bcwt | dout_rsc_req_obj_biwt))
          | dout_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
    (
  run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_vd, dout_rsc_req_obj_biwt, dout_rsc_req_obj_bdwt,
      dout_rsc_req_obj_bcwt
);
  input run_wen;
  input dout_rsc_req_obj_oswt;
  input dout_rsc_req_obj_vd;
  output dout_rsc_req_obj_biwt;
  output dout_rsc_req_obj_bdwt;
  input dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_bdwt = dout_rsc_req_obj_oswt & run_wen;
  assign dout_rsc_req_obj_biwt = dout_rsc_req_obj_oswt & (~ dout_rsc_req_obj_bcwt)
      & dout_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
    (
  run_wten, dout_rsc_rls_obj_iswt0, dout_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input dout_rsc_rls_obj_iswt0;
  output dout_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_rls_obj_ld_run_sct = dout_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl (
  dout_rsci_web_d_run_sct_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_web_d_run_sct_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_web_d_run_sct_pff = dout_rsci_iswt0_pff & (~ run_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp (
  clk, arst_n, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt, din_rsci_biwt,
      din_rsci_bdwt, din_rsci_bcwt, din_rsci_idat
);
  input clk;
  input arst_n;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  output din_rsci_bcwt;
  reg din_rsci_bcwt;
  input [15:0] din_rsci_idat;


  // Interconnect Declarations
  reg [15:0] din_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_idat_mxwt = MUX_v_16_2_2(din_rsci_idat, din_rsci_idat_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_idat_bfwt <= din_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl (
  run_wen, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_bcwt, din_rsci_irdy_run_sct,
      din_rsci_ivld
);
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  input din_rsci_bcwt;
  output din_rsci_irdy_run_sct;
  input din_rsci_ivld;


  // Interconnect Declarations
  wire din_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_ivld;
  assign din_rsci_ogwt = din_rsci_oswt & (~ din_rsci_bcwt);
  assign din_rsci_irdy_run_sct = din_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [136:0] paramsIn_rsci_idat_bfwt_136_0;
  wire [136:0] paramsIn_rsci_idat_mxwt_opt_136_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_136_0 = MUX_v_137_2_2((paramsIn_rsci_idat[136:0]),
      paramsIn_rsci_idat_bfwt_136_0, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_opt_136_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= paramsIn_rsci_idat_mxwt_opt_136_0;
    end
  end

  function automatic [136:0] MUX_v_137_2_2;
    input [136:0] input_0;
    input [136:0] input_1;
    input [0:0] sel;
    reg [136:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_137_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_sram_512_128_sram_512_128_rwport_8_128_12_512_128_gen
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_sram_512_128_sram_512_128_rwport_8_128_12_512_128_gen
    (
  dout, din, addr, web, csb, web_d, addr_d, din_d, dout_d, port_0_rw_ram_ir_internal_RMASK_B_d,
      port_0_rw_ram_ir_internal_WMASK_B_d
);
  input [127:0] dout;
  output [127:0] din;
  output [11:0] addr;
  output web;
  output csb;
  input web_d;
  input [11:0] addr_d;
  input [127:0] din_d;
  output [127:0] dout_d;
  input port_0_rw_ram_ir_internal_RMASK_B_d;
  input port_0_rw_ram_ir_internal_WMASK_B_d;


  wire din_and_nl;

  // Interconnect Declarations for Component Instantiations 
  assign dout_d = dout;
  assign din = (din_d);
  assign addr = (addr_d);
  assign web = (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign din_and_nl = (~ (port_0_rw_ram_ir_internal_RMASK_B_d)) & (~ (port_0_rw_ram_ir_internal_WMASK_B_d));
  assign csb = (din_and_nl);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_1_tr0, while_while_C_1_tr0, while_while_for_C_0_tr0,
      while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input main_C_1_tr0;
  input while_while_C_1_tr0;
  input while_while_for_C_0_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for InputDoubleBufferReader_512_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    while_C_0 = 4'd3,
    while_while_C_0 = 4'd4,
    while_while_C_1 = 4'd5,
    while_while_for_C_0 = 4'd6,
    while_while_C_2 = 4'd7,
    while_C_1 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBufferReader_512_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        if ( main_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 9'b000001000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 9'b000010000;
        state_var_NS = while_while_C_1;
      end
      while_while_C_1 : begin
        fsm_output = 9'b000100000;
        if ( while_while_C_1_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 9'b001000000;
        if ( while_while_for_C_0_tr0 ) begin
          state_var_NS = while_while_C_2;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_C_2 : begin
        fsm_output = 9'b010000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 9'b100000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_staller
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, dout_rsci_wen_comp, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input dout_rsci_wen_comp;
  input din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & dout_rsci_wen_comp & din_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
    (
  clk, arst_n, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt, din_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;
  input din_rsc_req_obj_biwt;
  input din_rsc_req_obj_bdwt;
  output din_rsc_req_obj_bcwt;
  reg din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_wen_comp = (~ din_rsc_req_obj_oswt) | din_rsc_req_obj_biwt
      | din_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_bcwt <= ~((~(din_rsc_req_obj_bcwt | din_rsc_req_obj_biwt))
          | din_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
    (
  run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_vd, din_rsc_req_obj_biwt, din_rsc_req_obj_bdwt,
      din_rsc_req_obj_bcwt
);
  input run_wen;
  input din_rsc_req_obj_oswt;
  input din_rsc_req_obj_vd;
  output din_rsc_req_obj_biwt;
  output din_rsc_req_obj_bdwt;
  input din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_bdwt = din_rsc_req_obj_oswt & run_wen;
  assign din_rsc_req_obj_biwt = din_rsc_req_obj_oswt & (~ din_rsc_req_obj_bcwt) &
      din_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
    (
  run_wten, din_rsc_rls_obj_iswt0, din_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input din_rsc_rls_obj_iswt0;
  output din_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_rls_obj_ld_run_sct = din_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp (
  clk, arst_n, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_bcwt
);
  input clk;
  input arst_n;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;
  output dout_rsci_bcwt;
  reg dout_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl (
  run_wen, dout_rsci_oswt, dout_rsci_irdy, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt,
      dout_rsci_ivld_run_sct
);
  input run_wen;
  input dout_rsci_oswt;
  input dout_rsci_irdy;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  input dout_rsci_bcwt;
  output dout_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dout_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_bdwt = dout_rsci_oswt & run_wen;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_irdy;
  assign dout_rsci_ogwt = dout_rsci_oswt & (~ dout_rsci_bcwt);
  assign dout_rsci_ivld_run_sct = dout_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl (
  run_wen, run_wten, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_addr_d_run_sct_pff,
      din_rsci_oswt_pff
);
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_addr_d_run_sct_pff;
  input din_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = (~ run_wten) & din_rsci_oswt;
  assign din_rsci_addr_d_run_sct_pff = din_rsci_oswt_pff & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp (
  clk, arst_n, din_rsci_addr_d, din_rsci_dout_d, din_rsci_addr_d_run, din_rsci_dout_d_mxwt,
      din_rsci_biwt, din_rsci_bdwt, din_rsci_addr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  input [11:0] din_rsci_addr_d_run;
  output [127:0] din_rsci_dout_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  input din_rsci_addr_d_run_sct_pff;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [127:0] din_rsci_dout_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_dout_d_mxwt = MUX_v_128_2_2(din_rsci_dout_d, din_rsci_dout_d_bfwt,
      din_rsci_bcwt);
  assign din_rsci_addr_d = {(~ din_rsci_addr_d_run_sct_pff) , (~ din_rsci_addr_d_run_sct_pff)
      , (~ din_rsci_addr_d_run_sct_pff) , (din_rsci_addr_d_run[8:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_dout_d_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_dout_d_bfwt <= din_rsci_dout_d_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [136:0] paramsIn_rsci_idat_bfwt_136_0;
  wire [136:0] paramsIn_rsci_idat_mxwt_opt_136_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_136_0 = MUX_v_137_2_2((paramsIn_rsci_idat[136:0]),
      paramsIn_rsci_idat_bfwt_136_0, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_opt_136_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= paramsIn_rsci_idat_mxwt_opt_136_0;
    end
  end

  function automatic [136:0] MUX_v_137_2_2;
    input [136:0] input_0;
    input [136:0] input_1;
    input [0:0] sel;
    reg [136:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_137_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi (
  clk, arst_n, inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy, run_wen, inputDoubleBufferReaderParams_cnsi_oswt,
      inputDoubleBufferReaderParams_cnsi_wen_comp, inputDoubleBufferReaderParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;
  input run_wen;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  output inputDoubleBufferReaderParams_cnsi_wen_comp;
  input [143:0] inputDoubleBufferReaderParams_cnsi_idat;


  // Interconnect Declarations
  wire inputDoubleBufferReaderParams_cnsi_irdy;
  wire inputDoubleBufferReaderParams_cnsi_biwt;
  wire inputDoubleBufferReaderParams_cnsi_bdwt;
  wire inputDoubleBufferReaderParams_cnsi_bcwt;
  wire inputDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd19),
  .width(32'sd144)) inputDoubleBufferReaderParams_cnsi (
      .irdy(inputDoubleBufferReaderParams_cnsi_irdy),
      .ivld(inputDoubleBufferReaderParams_cnsi_ivld_run_sct),
      .idat(inputDoubleBufferReaderParams_cnsi_idat),
      .rdy(inputDoubleBufferReaderParams_cns_rdy),
      .vld(inputDoubleBufferReaderParams_cns_vld),
      .dat(inputDoubleBufferReaderParams_cns_dat)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputDoubleBufferReaderParams_cnsi_oswt(inputDoubleBufferReaderParams_cnsi_oswt),
      .inputDoubleBufferReaderParams_cnsi_irdy(inputDoubleBufferReaderParams_cnsi_irdy),
      .inputDoubleBufferReaderParams_cnsi_biwt(inputDoubleBufferReaderParams_cnsi_biwt),
      .inputDoubleBufferReaderParams_cnsi_bdwt(inputDoubleBufferReaderParams_cnsi_bdwt),
      .inputDoubleBufferReaderParams_cnsi_bcwt(inputDoubleBufferReaderParams_cnsi_bcwt),
      .inputDoubleBufferReaderParams_cnsi_ivld_run_sct(inputDoubleBufferReaderParams_cnsi_ivld_run_sct)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferReaderParams_cnsi_oswt(inputDoubleBufferReaderParams_cnsi_oswt),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_biwt(inputDoubleBufferReaderParams_cnsi_biwt),
      .inputDoubleBufferReaderParams_cnsi_bdwt(inputDoubleBufferReaderParams_cnsi_bdwt),
      .inputDoubleBufferReaderParams_cnsi_bcwt(inputDoubleBufferReaderParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi (
  clk, arst_n, inputDoubleBufferWriterParams_cns_dat, inputDoubleBufferWriterParams_cns_vld,
      inputDoubleBufferWriterParams_cns_rdy, run_wen, inputDoubleBufferWriterParams_cnsi_oswt,
      inputDoubleBufferWriterParams_cnsi_wen_comp, inputDoubleBufferWriterParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  input run_wen;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  output inputDoubleBufferWriterParams_cnsi_wen_comp;
  input [143:0] inputDoubleBufferWriterParams_cnsi_idat;


  // Interconnect Declarations
  wire inputDoubleBufferWriterParams_cnsi_irdy;
  wire inputDoubleBufferWriterParams_cnsi_biwt;
  wire inputDoubleBufferWriterParams_cnsi_bdwt;
  wire inputDoubleBufferWriterParams_cnsi_bcwt;
  wire inputDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd18),
  .width(32'sd144)) inputDoubleBufferWriterParams_cnsi (
      .irdy(inputDoubleBufferWriterParams_cnsi_irdy),
      .ivld(inputDoubleBufferWriterParams_cnsi_ivld_run_sct),
      .idat(inputDoubleBufferWriterParams_cnsi_idat),
      .rdy(inputDoubleBufferWriterParams_cns_rdy),
      .vld(inputDoubleBufferWriterParams_cns_vld),
      .dat(inputDoubleBufferWriterParams_cns_dat)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputDoubleBufferWriterParams_cnsi_oswt(inputDoubleBufferWriterParams_cnsi_oswt),
      .inputDoubleBufferWriterParams_cnsi_irdy(inputDoubleBufferWriterParams_cnsi_irdy),
      .inputDoubleBufferWriterParams_cnsi_biwt(inputDoubleBufferWriterParams_cnsi_biwt),
      .inputDoubleBufferWriterParams_cnsi_bdwt(inputDoubleBufferWriterParams_cnsi_bdwt),
      .inputDoubleBufferWriterParams_cnsi_bcwt(inputDoubleBufferWriterParams_cnsi_bcwt),
      .inputDoubleBufferWriterParams_cnsi_ivld_run_sct(inputDoubleBufferWriterParams_cnsi_ivld_run_sct)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferWriterParams_cnsi_oswt(inputDoubleBufferWriterParams_cnsi_oswt),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_biwt(inputDoubleBufferWriterParams_cnsi_biwt),
      .inputDoubleBufferWriterParams_cnsi_bdwt(inputDoubleBufferWriterParams_cnsi_bdwt),
      .inputDoubleBufferWriterParams_cnsi_bcwt(inputDoubleBufferWriterParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd17),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj (
  clk, arst_n, dout_rsc_req_vz, run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input dout_rsc_req_vz;
  input run_wen;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_rsc_req_obj_vd;
  wire dout_rsc_req_obj_biwt;
  wire dout_rsc_req_obj_bdwt;
  wire dout_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) dout_rsc_req_obj (
      .vd(dout_rsc_req_obj_vd),
      .vz(dout_rsc_req_vz)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_vd(dout_rsc_req_obj_vd),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj (
  dout_rsc_rls_lz, run_wten, dout_rsc_rls_obj_iswt0
);
  output dout_rsc_rls_lz;
  input run_wten;
  input dout_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) dout_rsc_rls_obj (
      .ld(dout_rsc_rls_obj_ld_run_sct),
      .lz(dout_rsc_rls_lz)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(dout_rsc_rls_obj_iswt0),
      .dout_rsc_rls_obj_ld_run_sct(dout_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsci_1
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsci_1 (
  dout_rsci_addr_d, dout_rsci_addr_d_run, dout_rsci_web_d_pff, dout_rsci_iswt0_pff,
      run_wten_pff
);
  output [11:0] dout_rsci_addr_d;
  input [11:0] dout_rsci_addr_d_run;
  output dout_rsci_web_d_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;


  // Interconnect Declarations
  wire dout_rsci_web_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl_inst
      (
      .dout_rsci_web_d_run_sct_pff(dout_rsci_web_d_run_sct_iff),
      .dout_rsci_iswt0_pff(dout_rsci_iswt0_pff),
      .run_wten_pff(run_wten_pff)
    );
  assign dout_rsci_web_d_pff = ~ dout_rsci_web_d_run_sct_iff;
  assign dout_rsci_addr_d = {(~ dout_rsci_web_d_run_sct_iff) , (~ dout_rsci_web_d_run_sct_iff)
      , (~ dout_rsci_web_d_run_sct_iff) , (dout_rsci_addr_d_run[8:0])};
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci (
  clk, arst_n, din_rsc_dat, din_rsc_vld, din_rsc_rdy, run_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_bcwt;
  wire din_rsci_irdy_run_sct;
  wire din_rsci_ivld;
  wire [15:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd16)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_irdy_run_sct),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_irdy_run_sct(din_rsci_irdy_run_sct),
      .din_rsci_ivld(din_rsci_ivld)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_idat(din_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [136:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj (
  clk, arst_n, din_rsc_req_vz, run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input din_rsc_req_vz;
  input run_wen;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_rsc_req_obj_vd;
  wire din_rsc_req_obj_biwt;
  wire din_rsc_req_obj_bdwt;
  wire din_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) din_rsc_req_obj (
      .vd(din_rsc_req_obj_vd),
      .vz(din_rsc_req_vz)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_vd(din_rsc_req_obj_vd),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj (
  din_rsc_rls_lz, run_wten, din_rsc_rls_obj_iswt0
);
  output din_rsc_rls_lz;
  input run_wten;
  input din_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) din_rsc_rls_obj (
      .ld(din_rsc_rls_obj_ld_run_sct),
      .lz(din_rsc_rls_lz)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(din_rsc_rls_obj_iswt0),
      .din_rsc_rls_obj_ld_run_sct(din_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci (
  clk, arst_n, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, run_wen, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_idat
);
  input clk;
  input arst_n;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [127:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_irdy;
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_bcwt;
  wire dout_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd128)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_ivld_run_sct),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_irdy(dout_rsci_irdy),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt),
      .dout_rsci_ivld_run_sct(dout_rsci_ivld_run_sct)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1 (
  clk, arst_n, din_rsci_addr_d, din_rsci_dout_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d,
      run_wen, run_wten, din_rsci_oswt, din_rsci_addr_d_run, din_rsci_dout_d_mxwt,
      din_rsci_oswt_pff
);
  input clk;
  input arst_n;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  input [11:0] din_rsci_addr_d_run;
  output [127:0] din_rsci_dout_d_mxwt;
  input din_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire [11:0] din_rsci_addr_d_reg;
  wire din_rsci_addr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [11:0] nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run;
  assign nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run
      = {3'b000 , (din_rsci_addr_d_run[8:0])};
  InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_addr_d(din_rsci_addr_d_reg),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_addr_d_run(nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp_inst_din_rsci_addr_d_run[11:0]),
      .din_rsci_dout_d_mxwt(din_rsci_dout_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_addr_d_run_sct_pff(din_rsci_addr_d_run_sct_iff)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_addr_d_run_sct_pff(din_rsci_addr_d_run_sct_iff),
      .din_rsci_oswt_pff(din_rsci_oswt_pff)
    );
  assign din_rsci_addr_d = din_rsci_addr_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_addr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [136:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, inputDoubleBufferWriterParams_cns_dat,
      inputDoubleBufferWriterParams_cns_vld, inputDoubleBufferWriterParams_cns_rdy,
      inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire inputDoubleBufferWriterParams_cnsi_wen_comp;
  wire inputDoubleBufferReaderParams_cnsi_wen_comp;
  wire [2:0] fsm_output;
  reg reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse;
  reg [143:0] reg_inputDoubleBufferReaderParams_cnsi_idat_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy),
      .run_wen(run_wen),
      .inputDoubleBufferWriterParams_cnsi_oswt(reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_idat(reg_inputDoubleBufferReaderParams_cnsi_idat_cse)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld),
      .inputDoubleBufferReaderParams_cns_rdy(inputDoubleBufferReaderParams_cns_rdy),
      .run_wen(run_wen),
      .inputDoubleBufferReaderParams_cnsi_oswt(reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_idat(reg_inputDoubleBufferReaderParams_cnsi_idat_cse)
    );
  InputDoubleBuffer_512_16_16_run_run_staller InputDoubleBuffer_512_16_16_run_run_staller_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp)
    );
  InputDoubleBuffer_512_16_16_run_run_run_fsm InputDoubleBuffer_512_16_16_run_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputDoubleBufferReaderParams_cnsi_idat_cse <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_inputDoubleBufferReaderParams_cnsi_idat_cse <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= fsm_output[1];
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~ (fsm_output[1]);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_req_vz, dout_rsc_rls_lz, dout_rsci_addr_d,
      dout_rsci_din_d, dout_rsci_web_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;
  output [11:0] dout_rsci_addr_d;
  output [127:0] dout_rsci_din_d;
  output dout_rsci_web_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [136:0] paramsIn_rsci_idat_mxwt;
  wire din_rsci_wen_comp;
  wire [15:0] din_rsci_idat_mxwt;
  wire dout_rsc_req_obj_wen_comp;
  wire [15:0] fsm_output;
  wire [3:0] while_while_for_for_acc_1_tmp;
  wire [4:0] nl_while_while_for_for_acc_1_tmp;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_17;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire and_dcpl_11;
  wire or_dcpl_34;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire or_dcpl_38;
  wire or_dcpl_39;
  wire or_dcpl_40;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire or_dcpl_44;
  reg operator_32_false_1_slc_33_svs;
  wire exit_while_sva_mx0;
  reg [2:0] while_while_for_for_ic0_idx_3_0_sva_2_0;
  reg reg_dout_rsc_req_obj_iswt0_cse;
  reg reg_dout_rsc_rls_obj_ld_run_psct_cse;
  reg reg_din_rsci_irdy_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire dout_rsci_web_d_iff;
  wire [11:0] dout_rsci_addr_d_reg;
  reg [15:0] while_while_for_for_tmp_value_sva;
  reg [7:0] while_while_for_column_value_13_sva;
  reg [7:0] while_while_for_column_value_12_sva;
  reg [7:0] while_while_for_column_value_11_sva;
  reg [7:0] while_while_for_column_value_10_sva;
  reg [7:0] while_while_for_column_value_9_sva;
  reg [7:0] while_while_for_column_value_8_sva;
  reg [7:0] while_while_for_column_value_7_sva;
  reg [7:0] while_while_for_column_value_6_sva;
  reg [7:0] while_while_for_column_value_5_sva;
  reg [7:0] while_while_for_column_value_4_sva;
  reg [7:0] while_while_for_column_value_3_sva;
  reg [7:0] while_while_for_column_value_2_sva;
  reg [7:0] while_while_for_column_value_1_sva;
  reg [7:0] while_while_for_column_value_0_sva;
  reg [8:0] block_size_mul_1_itm;
  reg [8:0] operator_16_false_1_acc_itm;
  reg [31:0] total_blocks_lpi_3;
  reg [8:0] block_size_acc_1_itm;
  reg [136:0] paramsIn_crt_sva_136_0;
  wire [8:0] while_while_for_idx_sva_2;
  wire [9:0] nl_while_while_for_idx_sva_2;
  wire [31:0] total_blocks_sva_1;
  wire while_while_for_column_value_and_cse;
  wire while_while_for_column_value_and_2_cse;
  wire while_while_for_column_value_and_1_cse;
  wire while_while_for_column_value_and_4_cse;
  wire while_while_for_column_value_and_3_cse;
  wire while_while_for_column_value_and_6_cse;
  wire while_while_for_column_value_and_5_cse;
  wire operator_32_false_1_acc_1_itm_32_1;
  wire while_while_for_acc_2_itm_9_1;

  wire[8:0] operator_16_false_1_mux1h_4_nl;
  wire[8:0] operator_16_false_1_acc_nl;
  wire[9:0] nl_operator_16_false_1_acc_nl;
  wire[9:0] while_while_aelse_acc_1_nl;
  wire[10:0] nl_while_while_aelse_acc_1_nl;
  wire[0:0] or_59_nl;
  wire[0:0] not_nl;
  wire[8:0] block_size_acc_nl;
  wire[9:0] nl_block_size_acc_nl;
  wire[8:0] block_size_mul_2_nl;
  wire signed [18:0] nl_block_size_mul_2_nl;
  wire[8:0] operator_16_false_acc_nl;
  wire[9:0] nl_operator_16_false_acc_nl;
  wire[8:0] block_size_acc_1_nl;
  wire[9:0] nl_block_size_acc_1_nl;
  wire[8:0] block_size_mul_3_nl;
  wire signed [18:0] nl_block_size_mul_3_nl;
  wire[8:0] block_size_mul_nl;
  wire signed [17:0] nl_block_size_mul_nl;
  wire[8:0] block_size_mux1h_4_nl;
  wire[8:0] block_size_mul_1_nl;
  wire signed [18:0] nl_block_size_mul_1_nl;
  wire[8:0] while_while_acc_1_nl;
  wire[9:0] nl_while_while_acc_1_nl;
  wire[0:0] nor_5_nl;
  wire[0:0] nor_9_nl;
  wire[32:0] operator_32_false_acc_1_nl;
  wire[33:0] nl_operator_32_false_acc_1_nl;
  wire[9:0] while_while_for_acc_3_nl;
  wire[11:0] nl_while_while_for_acc_3_nl;
  wire[31:0] while_while_acc_nl;
  wire[32:0] nl_while_while_acc_nl;
  wire[32:0] operator_32_false_1_acc_1_nl;
  wire[33:0] nl_operator_32_false_1_acc_1_nl;
  wire[9:0] while_while_aelse_acc_nl;
  wire[10:0] nl_while_while_aelse_acc_nl;
  wire[9:0] while_while_for_acc_2_nl;
  wire[10:0] nl_while_while_for_acc_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[8:0] while_while_for_for_1_1_acc_1_nl;
  wire[9:0] nl_while_while_for_for_1_1_acc_1_nl;
  wire [11:0] nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run;
  assign nl_while_while_for_for_1_1_acc_1_nl = block_size_mul_1_itm + operator_16_false_1_acc_itm;
  assign while_while_for_for_1_1_acc_1_nl = nl_while_while_for_for_1_1_acc_1_nl[8:0];
  assign nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run
      = {3'b0, while_while_for_for_1_1_acc_1_nl};
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff;
  assign nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff
      = fsm_output[12];
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff;
  assign nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff =
      ~ run_wen;
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0;
  assign nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0
      = ~ while_while_for_acc_2_itm_9_1;
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0;
  assign nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0
      = while_while_for_for_acc_1_tmp[3];
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci InputDoubleBufferWriter_512_16_16_run_din_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .run_wen(run_wen),
      .din_rsci_oswt(reg_din_rsci_irdy_run_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsci_1 InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst
      (
      .dout_rsci_addr_d(dout_rsci_addr_d_reg),
      .dout_rsci_addr_d_run(nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_addr_d_run[11:0]),
      .dout_rsci_web_d_pff(dout_rsci_web_d_iff),
      .dout_rsci_iswt0_pff(nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff[0:0]),
      .run_wten_pff(nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff[0:0])
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_inst
      (
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(reg_dout_rsc_rls_obj_ld_run_psct_cse)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(reg_dout_rsc_req_obj_iswt0_cse),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferWriter_512_16_16_run_staller InputDoubleBufferWriter_512_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferWriter_512_16_16_run_run_fsm InputDoubleBufferWriter_512_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_5_tr0(exit_while_sva_mx0),
      .while_while_C_1_tr0(or_dcpl_26),
      .while_while_C_2_tr0(nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0[0:0]),
      .while_while_for_for_C_0_tr0(nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0[0:0]),
      .while_while_for_C_1_tr0(operator_32_false_1_slc_33_svs),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign while_while_for_column_value_and_cse = run_wen & (or_dcpl_12 | or_dcpl_11);
  assign while_while_for_column_value_and_1_cse = run_wen & (or_dcpl_15 | or_dcpl_14);
  assign while_while_for_column_value_and_2_cse = run_wen & (or_dcpl_12 | or_dcpl_17);
  assign while_while_for_column_value_and_3_cse = run_wen & (or_dcpl_15 | or_dcpl_17);
  assign while_while_for_column_value_and_4_cse = run_wen & (or_dcpl_12 | or_dcpl_14);
  assign while_while_for_column_value_and_5_cse = run_wen & (or_dcpl_15 | or_dcpl_11);
  assign while_while_for_column_value_and_6_cse = run_wen & (or_dcpl_12 | (while_while_for_for_acc_1_tmp[1:0]!=2'b11));
  assign nl_while_while_for_idx_sva_2 = operator_16_false_1_acc_itm + 9'b000000001;
  assign while_while_for_idx_sva_2 = nl_while_while_for_idx_sva_2[8:0];
  assign total_blocks_sva_1 = conv_u2u_32_32((paramsIn_crt_sva_136_0[31:16]) * (paramsIn_crt_sva_136_0[15:0]));
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ operator_32_false_1_slc_33_svs), (~
      operator_32_false_1_acc_1_itm_32_1), fsm_output[15]);
  assign nl_while_while_for_for_acc_1_tmp = conv_u2s_3_4(while_while_for_for_ic0_idx_3_0_sva_2_0)
      + 4'b0001;
  assign while_while_for_for_acc_1_tmp = nl_while_while_for_for_acc_1_tmp[3:0];
  assign nl_operator_32_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_1_acc_1_nl = nl_operator_32_false_1_acc_1_nl[32:0];
  assign operator_32_false_1_acc_1_itm_32_1 = readslicef_33_1_32((operator_32_false_1_acc_1_nl));
  assign or_dcpl_11 = (while_while_for_for_acc_1_tmp[1:0]!=2'b00);
  assign or_dcpl_12 = (while_while_for_for_acc_1_tmp[3:2]!=2'b00);
  assign or_dcpl_14 = (while_while_for_for_acc_1_tmp[1:0]!=2'b10);
  assign or_dcpl_15 = (while_while_for_for_acc_1_tmp[3:2]!=2'b01);
  assign or_dcpl_17 = (while_while_for_for_acc_1_tmp[1:0]!=2'b01);
  assign nl_while_while_aelse_acc_nl = conv_u2u_9_10(operator_16_false_1_acc_itm)
      + 10'b1100000001;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[9:0];
  assign or_dcpl_26 = (~ operator_32_false_1_slc_33_svs) | (readslicef_10_1_9((while_while_aelse_acc_nl)));
  assign or_dcpl_27 = (fsm_output[15]) | (fsm_output[6]);
  assign and_dcpl_11 = ~((fsm_output[1:0]!=2'b00));
  assign or_dcpl_34 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b00);
  assign or_dcpl_35 = or_dcpl_34 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_36 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b10);
  assign or_dcpl_37 = or_dcpl_36 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_38 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b01);
  assign or_dcpl_39 = or_dcpl_38 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_40 = or_dcpl_38 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_41 = or_dcpl_36 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_42 = or_dcpl_34 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_44 = (while_while_for_for_ic0_idx_3_0_sva_2_0!=3'b011);
  assign nl_while_while_for_acc_2_nl = ({1'b1 , (~ block_size_acc_1_itm)}) + 10'b0000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[9:0];
  assign while_while_for_acc_2_itm_9_1 = readslicef_10_1_9((while_while_for_acc_2_nl));
  assign dout_rsci_web_d_pff = dout_rsci_web_d_iff;
  assign dout_rsci_addr_d = dout_rsci_addr_d_reg;
  assign dout_rsci_din_d = {while_while_for_for_tmp_value_sva , while_while_for_column_value_13_sva
      , while_while_for_column_value_12_sva , while_while_for_column_value_11_sva
      , while_while_for_column_value_10_sva , while_while_for_column_value_9_sva
      , while_while_for_column_value_8_sva , while_while_for_column_value_7_sva ,
      while_while_for_column_value_6_sva , while_while_for_column_value_5_sva , while_while_for_column_value_4_sva
      , while_while_for_column_value_3_sva , while_while_for_column_value_2_sva ,
      while_while_for_column_value_1_sva , while_while_for_column_value_0_sva};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_din_rsci_irdy_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      operator_16_false_1_acc_itm <= 9'b000000000;
      block_size_mul_1_itm <= 9'b000000000;
      operator_32_false_1_slc_33_svs <= 1'b0;
      while_while_for_for_ic0_idx_3_0_sva_2_0 <= 3'b000;
    end
    else if ( run_wen ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= (~ exit_while_sva_mx0) & or_dcpl_27;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_26 & (fsm_output[9]);
      reg_din_rsci_irdy_run_psct_cse <= ((~ (while_while_for_for_acc_1_tmp[3])) &
          (fsm_output[11])) | ((~ operator_32_false_1_slc_33_svs) & (fsm_output[13]))
          | (while_while_for_acc_2_itm_9_1 & (fsm_output[10]));
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~(exit_while_sva_mx0 | (fsm_output[0])))
          | (~((fsm_output[0]) | (fsm_output[15]) | (fsm_output[6]))));
      operator_16_false_1_acc_itm <= MUX_v_9_2_2(9'b000000000, (operator_16_false_1_mux1h_4_nl),
          (not_nl));
      block_size_mul_1_itm <= MUX_v_9_2_2(9'b000000000, (block_size_mux1h_4_nl),
          (nor_9_nl));
      operator_32_false_1_slc_33_svs <= MUX1HOT_s_1_3_2((readslicef_33_1_32((operator_32_false_acc_1_nl))),
          operator_32_false_1_acc_1_itm_32_1, (~ (readslicef_10_1_9((while_while_for_acc_3_nl)))),
          {(fsm_output[5]) , (fsm_output[8]) , (fsm_output[12])});
      while_while_for_for_ic0_idx_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (while_while_for_for_acc_1_tmp[2:0]),
          (fsm_output[11]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_sva_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      paramsIn_crt_sva_136_0 <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_acc_1_itm <= 9'b000000000;
    end
    else if ( run_wen & ((~ and_dcpl_11) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[2])
        | (fsm_output[6])) ) begin
      block_size_acc_1_itm <= MUX1HOT_v_9_3_2((block_size_acc_nl), (block_size_acc_1_nl),
          (block_size_mul_nl), {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[6])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & ((~ and_dcpl_11) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[2])
        | (fsm_output[14]) | (fsm_output[5])) ) begin
      total_blocks_lpi_3 <= MUX_v_32_2_2(total_blocks_sva_1, (while_while_acc_nl),
          fsm_output[14]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_1_sva <= 8'b00000000;
      while_while_for_column_value_0_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_cse ) begin
      while_while_for_column_value_1_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_1_sva, or_dcpl_35);
      while_while_for_column_value_0_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_0_sva, or_dcpl_35);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_13_sva <= 8'b00000000;
      while_while_for_column_value_12_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_1_cse ) begin
      while_while_for_column_value_13_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_13_sva, or_dcpl_37);
      while_while_for_column_value_12_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_12_sva, or_dcpl_37);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_3_sva <= 8'b00000000;
      while_while_for_column_value_2_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_2_cse ) begin
      while_while_for_column_value_3_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_3_sva, or_dcpl_39);
      while_while_for_column_value_2_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_2_sva, or_dcpl_39);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_11_sva <= 8'b00000000;
      while_while_for_column_value_10_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_3_cse ) begin
      while_while_for_column_value_11_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_11_sva, or_dcpl_40);
      while_while_for_column_value_10_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_10_sva, or_dcpl_40);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_5_sva <= 8'b00000000;
      while_while_for_column_value_4_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_4_cse ) begin
      while_while_for_column_value_5_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_5_sva, or_dcpl_41);
      while_while_for_column_value_4_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_4_sva, or_dcpl_41);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_9_sva <= 8'b00000000;
      while_while_for_column_value_8_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_5_cse ) begin
      while_while_for_column_value_9_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_9_sva, or_dcpl_42);
      while_while_for_column_value_8_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_8_sva, or_dcpl_42);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_7_sva <= 8'b00000000;
      while_while_for_column_value_6_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_6_cse ) begin
      while_while_for_column_value_7_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_7_sva, or_dcpl_44);
      while_while_for_column_value_6_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_6_sva, or_dcpl_44);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_tmp_value_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (while_while_for_for_acc_1_tmp[3]) ) begin
      while_while_for_for_tmp_value_sva <= din_rsci_idat_mxwt;
    end
  end
  assign nl_operator_16_false_1_acc_nl = (paramsIn_rsci_idat_mxwt[40:32]) + 9'b111111111;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[8:0];
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_9_10(~ block_size_mul_1_itm) +
      conv_u2u_9_10(~ block_size_acc_1_itm);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[9:0];
  assign or_59_nl = (fsm_output[3]) | (fsm_output[13]) | (fsm_output[11]) | (fsm_output[2]);
  assign operator_16_false_1_mux1h_4_nl = MUX1HOT_v_9_4_2((operator_16_false_1_acc_nl),
      (readslicef_10_9_1((while_while_aelse_acc_1_nl))), while_while_for_idx_sva_2,
      operator_16_false_1_acc_itm, {(fsm_output[1]) , (fsm_output[8]) , (fsm_output[12])
      , (or_59_nl)});
  assign not_nl = ~ (fsm_output[10]);
  assign nl_block_size_mul_1_nl = $signed(conv_u2s_9_10(paramsIn_crt_sva_136_0[88:80]))
      * $signed(block_size_acc_1_itm);
  assign block_size_mul_1_nl = nl_block_size_mul_1_nl[8:0];
  assign nl_while_while_acc_1_nl = block_size_mul_1_itm + block_size_acc_1_itm;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[8:0];
  assign nor_5_nl = ~((~ and_dcpl_11) | (fsm_output[7]) | (fsm_output[2]) | (fsm_output[14])
      | (fsm_output[15]) | (fsm_output[6]));
  assign block_size_mux1h_4_nl = MUX1HOT_v_9_3_2((block_size_mul_1_nl), block_size_mul_1_itm,
      (while_while_acc_1_nl), {(fsm_output[2]) , (nor_5_nl) , (fsm_output[14])});
  assign nor_9_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[7]) | or_dcpl_27);
  assign nl_operator_32_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_acc_1_nl = nl_operator_32_false_acc_1_nl[32:0];
  assign nl_while_while_for_acc_3_nl = ({1'b1 , while_while_for_idx_sva_2}) + conv_u2u_9_10(~
      block_size_acc_1_itm) + 10'b0000000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[9:0];
  assign nl_operator_16_false_acc_nl = (paramsIn_rsci_idat_mxwt[56:48]) + 9'b111111111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[8:0];
  assign nl_block_size_mul_2_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[136:128]))
      * $signed((operator_16_false_acc_nl));
  assign block_size_mul_2_nl = nl_block_size_mul_2_nl[8:0];
  assign nl_block_size_acc_nl = (block_size_mul_2_nl) + (paramsIn_rsci_idat_mxwt[104:96]);
  assign block_size_acc_nl = nl_block_size_acc_nl[8:0];
  assign nl_block_size_mul_3_nl = $signed(conv_u2s_9_10(paramsIn_crt_sva_136_0[136:128]))
      * $signed(operator_16_false_1_acc_itm);
  assign block_size_mul_3_nl = nl_block_size_mul_3_nl[8:0];
  assign nl_block_size_acc_1_nl = (block_size_mul_3_nl) + (paramsIn_crt_sva_136_0[120:112]);
  assign block_size_acc_1_nl = nl_block_size_acc_1_nl[8:0];
  assign nl_block_size_mul_nl = $signed(block_size_mul_1_itm) * $signed(block_size_acc_1_itm);
  assign block_size_mul_nl = nl_block_size_mul_nl[8:0];
  assign nl_while_while_acc_nl = total_blocks_lpi_3 + 32'b11111111111111111111111111111111;
  assign while_while_acc_nl = nl_while_while_acc_nl[31:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_req_vz,
      din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, din_rsci_addr_d,
      din_rsci_dout_d, din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  output [11:0] din_rsci_addr_d;
  input [127:0] din_rsci_dout_d;
  output din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [136:0] paramsIn_rsci_idat_mxwt;
  wire [127:0] din_rsci_dout_d_mxwt;
  wire dout_rsci_wen_comp;
  reg [127:0] dout_rsci_idat;
  wire din_rsc_req_obj_wen_comp;
  wire [8:0] fsm_output;
  wire nor_tmp;
  wire or_dcpl_1;
  wire or_dcpl_8;
  wire nor_tmp_6;
  wire nor_tmp_7;
  wire or_tmp_22;
  wire and_dcpl_25;
  wire and_dcpl_32;
  wire or_dcpl_24;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_39;
  wire or_tmp_36;
  wire or_tmp_55;
  wire exit_while_sva_mx0;
  reg lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7;
  reg exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4;
  reg lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6;
  reg exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4;
  reg lfst_exitL_exit_while_while_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7;
  reg exitL_exitL_exit_while_while_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3;
  reg lfst_exitL_exit_while_while_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6;
  reg exitL_exitL_exit_while_while_for_for_for_lpi_2;
  reg exitL_exit_while_while_for_for_sva;
  reg lfst_exit_while_while_for_for_lpi_2;
  wire exit_while_while_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire exit_while_while_for_lpi_4_dfm_1;
  wire exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  reg while_while_for_for_asn_sft_lpi_4;
  reg while_while_for_stage_0_2;
  reg exit_while_while_for_lpi_4_dfm_st_1;
  reg while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_for_for_for_for_not_mdf_sva_st_1;
  reg while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_for_for_for_asn_sft_lpi_4;
  reg while_while_for_for_for_for_asn_sft_lpi_4;
  reg while_while_for_for_for_asn_sft_lpi_4;
  wire lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0;
  wire and_57_m1c;
  wire while_while_for_for_and_9_tmp;
  reg reg_din_rsc_req_obj_iswt0_cse;
  reg reg_din_rsc_rls_obj_ld_run_psct_cse;
  reg reg_dout_rsci_ivld_run_psct_cse;
  reg reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire while_while_for_for_for_and_cse;
  reg reg_while_while_for_stage_0_cse;
  wire while_while_for_for_for_for_for_for_y_idx_and_cse;
  wire or_1_cse;
  wire or_34_cse;
  wire while_while_for_for_for_and_7_cse;
  wire while_while_for_for_for_for_and_3_cse;
  wire while_while_for_for_for_for_for_and_2_cse;
  wire while_while_aelse_while_while_aelse_and_cse;
  wire [11:0] din_rsci_addr_d_reg;
  wire and_69_rmff;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  reg [136:0] paramsIn_crt_sva_136_0;
  wire [15:0] while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7;
  wire [15:0] while_while_for_for_for_for_wy_idx_lpi_4_dfm_6;
  reg [8:0] while_block_count_8_0_sva;
  reg [8:0] block_size_sva;
  wire [15:0] while_while_for_for_co_idx_lpi_4_dfm_1_mx0;
  reg [8:0] block_size_acc_cse_sva;
  reg [8:0] block_size_acc_1_cse_sva;
  wire [15:0] while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7;
  wire [15:0] while_while_for_for_for_wx_idx_lpi_4_dfm_5;
  reg [31:0] total_blocks_lpi_3;
  reg [8:0] while_current_buffer_size_sva;
  reg [15:0] while_while_for_for_co_idx_lpi_4;
  reg [15:0] while_while_for_for_for_wx_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_wy_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_for_x_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_for_for_y_idx_lpi_4;
  wire [16:0] nl_while_while_for_for_for_for_for_for_y_idx_lpi_4;
  reg [15:0] while_while_for_koo_idx_sva;
  wire lfst_exit_while_while_for_for_lpi_2_mx0c1;
  wire [8:0] block_size_acc_cse_sva_mx0w0;
  wire [9:0] nl_block_size_acc_cse_sva_mx0w0;
  wire [8:0] block_size_acc_1_cse_sva_mx0w0;
  wire [9:0] nl_block_size_acc_1_cse_sva_mx0w0;
  wire [31:0] total_blocks_sva_1;
  wire exit_while_while_for_for_lpi_4_dfm_mx1w0;
  wire exit_while_while_for_for_for_lpi_4_dfm_1;
  wire lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5;
  wire exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
  wire exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_for_not_62;
  wire or_47_tmp;
  wire while_while_for_for_for_wx_idx_and_2_cse;
  wire while_while_for_for_for_for_for_for_acc_2_itm_16_1;
  wire while_while_for_for_for_for_for_acc_2_itm_16_1;
  wire while_while_for_for_for_for_acc_2_itm_16_1;
  wire while_while_for_for_for_acc_2_itm_16_1;
  wire while_while_for_for_acc_3_itm_16_1;
  wire while_while_for_acc_3_itm_16_1;
  wire operator_32_false_1_acc_1_itm_32_1;

  wire[0:0] mux_22_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_9_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_10_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_120_nl;
  wire[0:0] and_143_nl;
  wire[0:0] and_144_nl;
  wire[0:0] nor_11_nl;
  wire[0:0] or_35_nl;
  wire[0:0] and_145_nl;
  wire[0:0] and_146_nl;
  wire[8:0] block_size_mul_nl;
  wire signed [17:0] nl_block_size_mul_nl;
  wire[8:0] block_size_mul_1_nl;
  wire signed [18:0] nl_block_size_mul_1_nl;
  wire[31:0] while_while_acc_1_nl;
  wire[32:0] nl_while_while_acc_1_nl;
  wire[8:0] while_while_acc_2_nl;
  wire[9:0] nl_while_while_acc_2_nl;
  wire[0:0] while_current_buffer_size_not_1_nl;
  wire[8:0] while_block_count_mux_nl;
  wire[8:0] while_while_acc_nl;
  wire[9:0] nl_while_while_acc_nl;
  wire[0:0] while_block_count_not_nl;
  wire[15:0] while_while_for_koo_idx_mux1h_3_nl;
  wire[9:0] while_while_aelse_acc_1_nl;
  wire[10:0] nl_while_while_aelse_acc_1_nl;
  wire[15:0] while_while_for_acc_2_nl;
  wire[16:0] nl_while_while_for_acc_2_nl;
  wire[0:0] while_while_for_koo_idx_and_1_nl;
  wire[0:0] while_while_for_koo_idx_and_2_nl;
  wire[0:0] not_135_nl;
  wire[0:0] while_while_for_mux_3_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] nand_4_nl;
  wire[15:0] while_while_for_for_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_for_and_5_nl;
  wire[15:0] while_while_for_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_and_7_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] and_149_nl;
  wire[0:0] and_150_nl;
  wire[15:0] while_while_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_for_wx_idx_and_nl;
  wire[0:0] while_while_for_for_for_wx_idx_and_1_nl;
  wire[0:0] while_while_for_for_for_mux_35_nl;
  wire[15:0] while_while_for_for_acc_2_nl;
  wire[16:0] nl_while_while_for_for_acc_2_nl;
  wire[0:0] and_53_nl;
  wire[0:0] while_while_for_for_nand_nl;
  wire[0:0] while_while_for_for_and_10_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_13_nl;
  wire[8:0] block_size_mul_2_nl;
  wire signed [18:0] nl_block_size_mul_2_nl;
  wire[8:0] operator_16_false_acc_nl;
  wire[9:0] nl_operator_16_false_acc_nl;
  wire[8:0] block_size_mul_3_nl;
  wire signed [18:0] nl_block_size_mul_3_nl;
  wire[8:0] operator_16_false_1_acc_nl;
  wire[9:0] nl_operator_16_false_1_acc_nl;
  wire[32:0] operator_32_false_acc_1_nl;
  wire[33:0] nl_operator_32_false_acc_1_nl;
  wire[16:0] while_while_for_for_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_for_for_acc_2_nl;
  wire[0:0] or_60_nl;
  wire[0:0] or_69_nl;
  wire[0:0] or_71_nl;
  wire[0:0] or_73_nl;
  wire[16:0] while_while_for_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_acc_3_nl;
  wire[18:0] nl_while_while_for_for_acc_3_nl;
  wire[0:0] while_while_for_for_mux_60_nl;
  wire[16:0] while_while_for_acc_3_nl;
  wire[18:0] nl_while_while_for_acc_3_nl;
  wire[32:0] operator_32_false_1_acc_1_nl;
  wire[33:0] nl_operator_32_false_1_acc_1_nl;
  wire[9:0] while_while_aelse_acc_nl;
  wire[10:0] nl_while_while_aelse_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_10_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_10_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_8_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_8_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_8_nl;
  wire[17:0] nl_while_while_for_for_for_for_for_for_address_mul_8_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_nl;
  wire[17:0] nl_while_while_for_for_for_for_for_for_address_mul_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_9_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_9_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_1_nl;
  wire signed [17:0] nl_while_while_for_for_for_for_for_for_address_mul_1_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_2_nl;
  wire signed [18:0] nl_while_while_for_for_for_for_for_for_address_mul_2_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_5_nl;
  wire signed [18:0] nl_while_while_for_for_for_for_for_for_address_mul_5_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_6_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_6_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_6_nl;
  wire[17:0] nl_while_while_for_for_for_for_for_for_address_mul_6_nl;
  wire [11:0] nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run;
  assign nl_while_while_for_for_for_for_for_for_address_mul_8_nl = (paramsIn_crt_sva_136_0[136:128])
      * (while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7[8:0]);
  assign while_while_for_for_for_for_for_for_address_mul_8_nl = nl_while_while_for_for_for_for_for_for_address_mul_8_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_8_nl = (while_while_for_for_for_for_for_for_address_mul_8_nl)
      + (while_while_for_for_for_for_wy_idx_lpi_4_dfm_6[8:0]);
  assign while_while_for_for_for_for_for_for_address_acc_8_nl = nl_while_while_for_for_for_for_for_for_address_acc_8_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_nl = while_block_count_8_0_sva
      * block_size_sva;
  assign while_while_for_for_for_for_for_for_address_mul_nl = nl_while_while_for_for_for_for_for_for_address_mul_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_10_nl = (while_while_for_for_for_for_for_for_address_acc_8_nl)
      + (while_while_for_for_for_for_for_for_address_mul_nl);
  assign while_while_for_for_for_for_for_for_address_acc_10_nl = nl_while_while_for_for_for_for_for_for_address_acc_10_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_2_nl = $signed(conv_u2s_9_10(while_while_for_for_co_idx_lpi_4_dfm_1_mx0[8:0]))
      * $signed(block_size_acc_cse_sva);
  assign while_while_for_for_for_for_for_for_address_mul_2_nl = nl_while_while_for_for_for_for_for_for_address_mul_2_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_1_nl = $signed((while_while_for_for_for_for_for_for_address_mul_2_nl))
      * $signed(block_size_acc_1_cse_sva);
  assign while_while_for_for_for_for_for_for_address_mul_1_nl = nl_while_while_for_for_for_for_for_for_address_mul_1_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_6_nl = (paramsIn_crt_sva_136_0[136:128])
      * (while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7[8:0]);
  assign while_while_for_for_for_for_for_for_address_mul_6_nl = nl_while_while_for_for_for_for_for_for_address_mul_6_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_6_nl = (while_while_for_for_for_for_for_for_address_mul_6_nl)
      + (while_while_for_for_for_wx_idx_lpi_4_dfm_5[8:0]);
  assign while_while_for_for_for_for_for_for_address_acc_6_nl = nl_while_while_for_for_for_for_for_for_address_acc_6_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_5_nl = $signed(conv_u2s_9_10(while_while_for_for_for_for_for_for_address_acc_6_nl))
      * $signed(block_size_acc_cse_sva);
  assign while_while_for_for_for_for_for_for_address_mul_5_nl = nl_while_while_for_for_for_for_for_for_address_mul_5_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_9_nl = (while_while_for_for_for_for_for_for_address_mul_1_nl)
      + (while_while_for_for_for_for_for_for_address_mul_5_nl);
  assign while_while_for_for_for_for_for_for_address_acc_9_nl = nl_while_while_for_for_for_for_for_for_address_acc_9_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_nl = (while_while_for_for_for_for_for_for_address_acc_10_nl)
      + (while_while_for_for_for_for_for_for_address_acc_9_nl);
  assign while_while_for_for_for_for_for_for_address_acc_nl = nl_while_while_for_for_for_for_for_for_address_acc_nl[8:0];
  assign nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run
      = {3'b0, while_while_for_for_for_for_for_for_address_acc_nl};
  wire [0:0] nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0;
  assign nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0
      = ~(reg_while_while_for_stage_0_cse | while_while_for_stage_0_2);
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsci_1 InputDoubleBufferReader_512_16_16_run_din_rsci_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_addr_d(din_rsci_addr_d_reg),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .din_rsci_addr_d_run(nl_InputDoubleBufferReader_512_16_16_run_din_rsci_1_inst_din_rsci_addr_d_run[11:0]),
      .din_rsci_dout_d_mxwt(din_rsci_dout_d_mxwt),
      .din_rsci_oswt_pff(and_69_rmff)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci InputDoubleBufferReader_512_16_16_run_dout_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .run_wen(run_wen),
      .dout_rsci_oswt(reg_dout_rsci_ivld_run_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_inst
      (
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(reg_din_rsc_rls_obj_ld_run_psct_cse)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_vz(din_rsc_req_vz),
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(reg_din_rsc_req_obj_iswt0_cse),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferReader_512_16_16_run_staller InputDoubleBufferReader_512_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferReader_512_16_16_run_run_fsm InputDoubleBufferReader_512_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_1_tr0(exit_while_sva_mx0),
      .while_while_C_1_tr0(or_dcpl_8),
      .while_while_for_C_0_tr0(nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0[0:0]),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign or_120_nl = while_while_for_for_for_for_for_acc_2_itm_16_1 | (~ or_tmp_22);
  assign and_143_nl = while_while_for_for_for_for_for_acc_2_itm_16_1 & or_tmp_22;
  assign and_144_nl = while_while_for_for_for_for_for_asn_sft_lpi_4 & lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2;
  assign mux_15_nl = MUX_s_1_2_2((or_120_nl), (and_143_nl), and_144_nl);
  assign nor_11_nl = ~((~ while_while_for_for_for_for_for_acc_2_itm_16_1) | lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2);
  assign mux_16_nl = MUX_s_1_2_2((mux_15_nl), (nor_11_nl), while_while_for_for_for_for_asn_sft_lpi_4);
  assign or_35_nl = (~ lfst_exit_while_while_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  assign mux_17_nl = MUX_s_1_2_2((mux_16_nl), nor_tmp_7, or_35_nl);
  assign nor_10_nl = ~(while_while_for_for_for_asn_sft_lpi_4 | (~ (mux_17_nl)));
  assign mux_18_nl = MUX_s_1_2_2(nor_tmp_7, (nor_10_nl), lfst_exitL_exit_while_while_for_for_for_for_lpi_2);
  assign mux_19_nl = MUX_s_1_2_2((mux_18_nl), nor_tmp_6, or_34_cse);
  assign nor_9_nl = ~(while_while_for_for_asn_sft_lpi_4 | (~ (mux_19_nl)));
  assign mux_20_nl = MUX_s_1_2_2(nor_tmp_6, (nor_9_nl), lfst_exitL_exit_while_while_for_for_for_lpi_2);
  assign and_145_nl = while_while_for_for_acc_3_itm_16_1 & while_while_for_for_for_acc_2_itm_16_1
      & while_while_for_for_for_for_acc_2_itm_16_1 & while_while_for_for_for_for_for_acc_2_itm_16_1;
  assign mux_21_nl = MUX_s_1_2_2((mux_20_nl), (and_145_nl), or_1_cse);
  assign and_146_nl = while_while_for_acc_3_itm_16_1 & while_while_for_for_acc_3_itm_16_1
      & while_while_for_for_for_acc_2_itm_16_1 & while_while_for_for_for_for_acc_2_itm_16_1
      & while_while_for_for_for_for_for_acc_2_itm_16_1;
  assign mux_22_nl = MUX_s_1_2_2((mux_21_nl), (and_146_nl), exitL_exit_while_while_for_for_sva);
  assign and_69_rmff = (mux_22_nl) & reg_while_while_for_stage_0_cse & while_while_for_for_for_for_for_for_acc_2_itm_16_1
      & (fsm_output[6]);
  assign while_while_for_for_for_and_cse = run_wen & (~ or_tmp_36);
  assign while_while_for_for_for_and_7_cse = run_wen & (~(while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | or_tmp_36));
  assign while_while_for_for_for_for_and_3_cse = run_wen & (~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | or_tmp_36));
  assign while_while_for_for_for_for_for_and_2_cse = run_wen & (~(while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | or_tmp_36));
  assign or_47_tmp = and_dcpl_32 | while_while_for_for_acc_3_itm_16_1 | (~ reg_while_while_for_stage_0_cse);
  assign while_while_aelse_while_while_aelse_and_cse = reg_while_while_for_stage_0_cse
      & or_dcpl_1;
  assign or_1_cse = (~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2;
  assign while_while_for_for_for_for_for_for_y_idx_and_cse = run_wen & reg_while_while_for_stage_0_cse;
  assign while_while_for_for_and_9_tmp = exit_while_while_for_for_for_for_lpi_4_dfm_1
      & (~ while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & while_while_for_for_not_62;
  assign nor_18_nl = ~(while_while_for_for_asn_sft_lpi_4 | (~((~((~ lfst_exit_while_while_for_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_for_lpi_2)) | while_while_for_for_for_acc_2_itm_16_1)));
  assign mux_8_nl = MUX_s_1_2_2(while_while_for_for_for_acc_2_itm_16_1, (nor_18_nl),
      lfst_exitL_exit_while_while_for_for_for_lpi_2);
  assign and_149_nl = while_while_for_for_acc_3_itm_16_1 & while_while_for_for_for_acc_2_itm_16_1;
  assign mux_9_nl = MUX_s_1_2_2((mux_8_nl), (and_149_nl), or_1_cse);
  assign and_150_nl = while_while_for_acc_3_itm_16_1 & while_while_for_for_acc_3_itm_16_1
      & while_while_for_for_for_acc_2_itm_16_1;
  assign mux_10_nl = MUX_s_1_2_2((mux_9_nl), (and_150_nl), exitL_exit_while_while_for_for_sva);
  assign while_while_for_for_for_wx_idx_and_2_cse = run_wen & (mux_10_nl) & reg_while_while_for_stage_0_cse;
  assign and_57_m1c = (((((~ exitL_exitL_exit_while_while_for_for_for_for_lpi_2)
      & lfst_exit_while_while_for_for_for_lpi_2) | while_while_for_for_asn_sft_lpi_4)
      & lfst_exitL_exit_while_while_for_for_for_lpi_2 & and_dcpl_32) | while_while_for_for_for_acc_2_itm_16_1)
      & reg_while_while_for_stage_0_cse;
  assign or_34_cse = (~ lfst_exit_while_while_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_lpi_2;
  assign nl_operator_16_false_acc_nl = (paramsIn_rsci_idat_mxwt[56:48]) + 9'b111111111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[8:0];
  assign nl_block_size_mul_2_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[136:128]))
      * $signed((operator_16_false_acc_nl));
  assign block_size_mul_2_nl = nl_block_size_mul_2_nl[8:0];
  assign nl_block_size_acc_cse_sva_mx0w0 = (block_size_mul_2_nl) + (paramsIn_rsci_idat_mxwt[104:96]);
  assign block_size_acc_cse_sva_mx0w0 = nl_block_size_acc_cse_sva_mx0w0[8:0];
  assign nl_operator_16_false_1_acc_nl = (paramsIn_rsci_idat_mxwt[40:32]) + 9'b111111111;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[8:0];
  assign nl_block_size_mul_3_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[136:128]))
      * $signed((operator_16_false_1_acc_nl));
  assign block_size_mul_3_nl = nl_block_size_mul_3_nl[8:0];
  assign nl_block_size_acc_1_cse_sva_mx0w0 = (block_size_mul_3_nl) + (paramsIn_rsci_idat_mxwt[120:112]);
  assign block_size_acc_1_cse_sva_mx0w0 = nl_block_size_acc_1_cse_sva_mx0w0[8:0];
  assign nl_operator_32_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_acc_1_nl = nl_operator_32_false_acc_1_nl[32:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ (readslicef_33_1_32((operator_32_false_acc_1_nl)))),
      (~ operator_32_false_1_acc_1_itm_32_1), fsm_output[8]);
  assign total_blocks_sva_1 = conv_u2u_32_32((paramsIn_crt_sva_136_0[31:16]) * (paramsIn_crt_sva_136_0[15:0]));
  assign exit_while_while_for_lpi_4_dfm_1 = (~ while_while_for_acc_3_itm_16_1) &
      exitL_exit_while_while_for_for_sva;
  assign exit_while_while_for_for_lpi_4_dfm_mx1w0 = (~ while_while_for_for_acc_3_itm_16_1)
      & exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6;
  assign nl_while_while_for_for_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7})
      + conv_u2u_16_17(~ (paramsIn_crt_sva_136_0[63:48])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_for_for_acc_2_itm_16_1 = readslicef_17_1_16((while_while_for_for_for_for_for_for_acc_2_nl));
  assign or_60_nl = (~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2))
      | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 | (~ lfst_exit_while_while_for_for_for_for_lpi_2)
      | (~ lfst_exitL_exit_while_while_for_for_for_for_lpi_2) | or_34_cse | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2)
      | or_dcpl_24;
  assign while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_for_for_lpi_4_dfm_1, or_60_nl);
  assign or_69_nl = (~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2
      | (~ lfst_exit_while_while_for_for_for_for_lpi_2) | or_dcpl_39 | or_dcpl_36
      | exitL_exitL_exit_while_while_for_for_for_lpi_2 | or_dcpl_35;
  assign while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_for_lpi_4_dfm_1, or_69_nl);
  assign or_71_nl = or_dcpl_39 | or_dcpl_36 | or_dcpl_24;
  assign while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_lpi_4_dfm_1, or_71_nl);
  assign or_73_nl = (~ lfst_exitL_exit_while_while_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2
      | or_dcpl_35;
  assign while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_lpi_4_dfm_mx1w0, or_73_nl);
  assign exit_while_while_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_acc_2_itm_16_1)
      & exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7;
  assign while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_for_for_for_y_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5);
  assign while_while_for_for_for_for_wy_idx_lpi_4_dfm_6 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_for_wy_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4);
  assign while_while_for_for_co_idx_lpi_4_dfm_1_mx0 = MUX_v_16_2_2(while_while_for_for_co_idx_lpi_4,
      (signext_16_1(~ while_while_for_acc_3_itm_16_1)), exitL_exit_while_while_for_for_sva);
  assign while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_for_for_x_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4);
  assign while_while_for_for_for_wx_idx_lpi_4_dfm_5 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_wx_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3);
  assign lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5 = lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7);
  assign nl_while_while_for_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7})
      + conv_u2u_16_17(~ (paramsIn_crt_sva_136_0[47:32])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_for_acc_2_itm_16_1 = readslicef_17_1_16((while_while_for_for_for_for_for_acc_2_nl));
  assign exit_while_while_for_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_for_acc_2_itm_16_1)
      & exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7;
  assign exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7 = exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4));
  assign lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4 = lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6);
  assign nl_while_while_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_wy_idx_lpi_4_dfm_6})
      + conv_u2u_16_17(~ (paramsIn_crt_sva_136_0[127:112])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_acc_2_itm_16_1 = readslicef_17_1_16((while_while_for_for_for_for_acc_2_nl));
  assign exit_while_while_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_acc_2_itm_16_1)
      & exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6;
  assign exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6 = exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4));
  assign lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4 = lfst_exitL_exit_while_while_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7);
  assign nl_while_while_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_wx_idx_lpi_4_dfm_5})
      + conv_u2u_16_17(~ (paramsIn_crt_sva_136_0[111:96])) + 17'b00000000000000001;
  assign while_while_for_for_for_acc_2_nl = nl_while_while_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_acc_2_itm_16_1 = readslicef_17_1_16((while_while_for_for_for_acc_2_nl));
  assign exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7 = exitL_exitL_exit_while_while_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3));
  assign lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3 = lfst_exitL_exit_while_while_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6);
  assign nl_while_while_for_for_acc_3_nl = ({1'b1 , while_while_for_for_co_idx_lpi_4_dfm_1_mx0})
      + conv_u2u_16_17(~ (paramsIn_crt_sva_136_0[95:80])) + 17'b00000000000000001;
  assign while_while_for_for_acc_3_nl = nl_while_while_for_for_acc_3_nl[16:0];
  assign while_while_for_for_acc_3_itm_16_1 = readslicef_17_1_16((while_while_for_for_acc_3_nl));
  assign while_while_for_for_mux_60_nl = MUX_s_1_2_2(lfst_exit_while_while_for_for_lpi_2,
      lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0, exitL_exit_while_while_for_for_sva);
  assign exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6 = exitL_exitL_exit_while_while_for_for_for_lpi_2
      | (~ (while_while_for_for_mux_60_nl));
  assign lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0 = lfst_exit_while_while_for_for_lpi_2
      & (~ while_while_for_acc_3_itm_16_1);
  assign nl_while_while_for_acc_3_nl = ({1'b1 , while_while_for_koo_idx_sva}) + conv_u2u_16_17(~
      (paramsIn_crt_sva_136_0[79:64])) + 17'b00000000000000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[16:0];
  assign while_while_for_acc_3_itm_16_1 = readslicef_17_1_16((while_while_for_acc_3_nl));
  assign exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_for_for_acc_2_itm_16_1)
      | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  assign exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1 = exit_while_while_for_for_for_for_for_lpi_4_dfm_1
      | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  assign while_while_for_for_not_62 = ~(while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | exit_while_while_for_lpi_4_dfm_1);
  assign nl_operator_32_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_1_acc_1_nl = nl_operator_32_false_1_acc_1_nl[32:0];
  assign operator_32_false_1_acc_1_itm_32_1 = readslicef_33_1_32((operator_32_false_1_acc_1_nl));
  assign nor_tmp = while_while_for_acc_3_itm_16_1 & while_while_for_for_acc_3_itm_16_1;
  assign or_dcpl_1 = while_while_for_acc_3_itm_16_1 | (~ exitL_exit_while_while_for_for_sva);
  assign nl_while_while_aelse_acc_nl = conv_u2u_9_10(while_while_for_koo_idx_sva[8:0])
      + 10'b1100000001;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[9:0];
  assign or_dcpl_8 = ~(exit_while_while_for_lpi_4_dfm_st_1 & (~ (readslicef_10_1_9((while_while_aelse_acc_nl)))));
  assign nor_tmp_6 = while_while_for_for_for_acc_2_itm_16_1 & while_while_for_for_for_for_acc_2_itm_16_1
      & while_while_for_for_for_for_for_acc_2_itm_16_1;
  assign nor_tmp_7 = while_while_for_for_for_for_acc_2_itm_16_1 & while_while_for_for_for_for_for_acc_2_itm_16_1;
  assign or_tmp_22 = (~ lfst_exit_while_while_for_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2);
  assign and_dcpl_25 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_32 = (~ exitL_exitL_exit_while_while_for_for_for_lpi_2) & lfst_exit_while_while_for_for_lpi_2
      & (~ exitL_exit_while_while_for_for_sva);
  assign or_dcpl_24 = exitL_exitL_exit_while_while_for_for_for_lpi_2 | (~ lfst_exit_while_while_for_for_lpi_2)
      | exitL_exit_while_while_for_for_sva;
  assign or_dcpl_35 = (~ lfst_exit_while_while_for_for_lpi_2) | exitL_exit_while_while_for_for_sva;
  assign or_dcpl_36 = ~(lfst_exit_while_while_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_lpi_2);
  assign or_dcpl_39 = (~ lfst_exitL_exit_while_while_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_lpi_2;
  assign or_tmp_36 = (~ (fsm_output[6])) | exit_while_while_for_lpi_4_dfm_1 | (~
      reg_while_while_for_stage_0_cse);
  assign or_tmp_55 = ~((fsm_output[7:4]!=4'b0000));
  assign lfst_exit_while_while_for_for_lpi_2_mx0c1 = exit_while_while_for_lpi_4_dfm_1
      & reg_while_while_for_stage_0_cse & (fsm_output[6]);
  assign din_rsci_addr_d = din_rsci_addr_d_reg;
  assign din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d = din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_din_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_din_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_dout_rsci_ivld_run_psct_cse <= 1'b0;
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      block_size_sva <= 9'b000000000;
      paramsIn_crt_sva_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      block_size_acc_cse_sva <= 9'b000000000;
      block_size_acc_1_cse_sva <= 9'b000000000;
      while_block_count_8_0_sva <= 9'b000000000;
      exit_while_while_for_lpi_4_dfm_st_1 <= 1'b0;
      while_while_for_koo_idx_sva <= 16'b0000000000000000;
      reg_while_while_for_stage_0_cse <= 1'b0;
      exitL_exit_while_while_for_for_sva <= 1'b0;
      while_while_for_stage_0_2 <= 1'b0;
      while_while_for_for_for_for_for_for_not_mdf_sva_st_1 <= 1'b0;
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_din_rsc_req_obj_iswt0_cse <= ~(exit_while_sva_mx0 | (~((fsm_output[2])
          | (fsm_output[8]))));
      reg_din_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_8 & (fsm_output[5]);
      reg_dout_rsci_ivld_run_psct_cse <= (~ exit_while_while_for_lpi_4_dfm_st_1)
          & while_while_for_stage_0_2 & (~(while_while_for_for_for_for_for_for_not_mdf_sva_st_1
          | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1)) & (~(while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1
          | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_asn_sft_lpi_4_dfm_st_1))
          & (fsm_output[6]);
      reg_din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d_run_psct_cse <= and_69_rmff;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[0]) | (fsm_output[2])
          | (fsm_output[8]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      block_size_sva <= MUX_v_9_2_2((block_size_mul_nl), block_size_sva, and_dcpl_25);
      paramsIn_crt_sva_136_0 <= MUX_v_137_2_2(paramsIn_rsci_idat_mxwt, paramsIn_crt_sva_136_0,
          and_dcpl_25);
      block_size_acc_cse_sva <= MUX_v_9_2_2(block_size_acc_cse_sva_mx0w0, block_size_acc_cse_sva,
          and_dcpl_25);
      block_size_acc_1_cse_sva <= MUX_v_9_2_2(block_size_acc_1_cse_sva_mx0w0, block_size_acc_1_cse_sva,
          and_dcpl_25);
      while_block_count_8_0_sva <= MUX_v_9_2_2(9'b000000000, (while_block_count_mux_nl),
          (while_block_count_not_nl));
      exit_while_while_for_lpi_4_dfm_st_1 <= MUX_s_1_2_2(operator_32_false_1_acc_1_itm_32_1,
          exit_while_while_for_lpi_4_dfm_1, fsm_output[6]);
      while_while_for_koo_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, (while_while_for_koo_idx_mux1h_3_nl),
          (not_135_nl));
      reg_while_while_for_stage_0_cse <= while_while_aelse_while_while_aelse_and_cse
          | (~ (fsm_output[6]));
      exitL_exit_while_while_for_for_sva <= (while_while_for_mux_3_nl) | (~ (fsm_output[6]));
      while_while_for_stage_0_2 <= reg_while_while_for_stage_0_cse & (fsm_output[6]);
      while_while_for_for_for_for_for_for_not_mdf_sva_st_1 <= ~ while_while_for_for_for_for_for_for_acc_2_itm_16_1;
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_idat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ (fsm_output[6])) | exit_while_while_for_lpi_4_dfm_st_1
        | (~ while_while_for_stage_0_2) | while_while_for_for_for_for_for_for_not_mdf_sva_st_1
        | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1
        | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_asn_sft_lpi_4_dfm_st_1))
        ) begin
      dout_rsci_idat <= din_rsci_dout_d_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_lpi_2 <= 1'b0;
    end
    else if ( run_wen & ((or_dcpl_1 & reg_while_while_for_stage_0_cse & (fsm_output[6]))
        | lfst_exit_while_while_for_for_lpi_2_mx0c1) ) begin
      lfst_exit_while_while_for_for_lpi_2 <= MUX_s_1_2_2((~ exit_while_while_for_for_lpi_4_dfm_mx1w0),
          lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0, lfst_exit_while_while_for_for_lpi_2_mx0c1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exitL_exit_while_while_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_and_cse ) begin
      exitL_exitL_exit_while_while_for_for_for_lpi_2 <= exit_while_while_for_for_for_lpi_4_dfm_1
          | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      lfst_exitL_exit_while_while_for_for_for_lpi_2 <= ~(exit_while_while_for_for_for_lpi_4_dfm_1
          | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_and_7_cse ) begin
      lfst_exit_while_while_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_lpi_2 <= exit_while_while_for_for_for_for_lpi_4_dfm_1
          | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      lfst_exitL_exit_while_while_for_for_for_for_lpi_2 <= ~(exit_while_while_for_for_for_for_lpi_4_dfm_1
          | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_for_and_3_cse ) begin
      lfst_exit_while_while_for_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
      lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= ~ exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_for_for_and_2_cse ) begin
      lfst_exit_while_while_for_for_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
      lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= ~ exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & ((~ and_dcpl_25) | (fsm_output[2]) | (fsm_output[7])) ) begin
      total_blocks_lpi_3 <= MUX_v_32_2_2(total_blocks_sva_1, (while_while_acc_1_nl),
          fsm_output[7]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_current_buffer_size_sva <= 9'b000000000;
    end
    else if ( (fsm_output[6:4]==3'b000) & run_wen ) begin
      while_current_buffer_size_sva <= MUX_v_9_2_2(9'b000000000, (while_while_acc_2_nl),
          (while_current_buffer_size_not_1_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen & (mux_7_nl) & reg_while_while_for_stage_0_cse ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen & while_while_aelse_while_while_aelse_and_cse ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_for_y_idx_lpi_4 <= 16'b0000000000000000;
      while_while_for_for_for_for_for_x_idx_lpi_4 <= 16'b0000000000000000;
      while_while_for_for_for_for_wy_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( while_while_for_for_for_for_for_for_y_idx_and_cse ) begin
      while_while_for_for_for_for_for_for_y_idx_lpi_4 <= nl_while_while_for_for_for_for_for_for_y_idx_lpi_4[15:0];
      while_while_for_for_for_for_for_x_idx_lpi_4 <= MUX_v_16_2_2(while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7,
          (while_while_for_for_for_for_for_acc_1_nl), while_while_for_for_for_and_5_nl);
      while_while_for_for_for_for_wy_idx_lpi_4 <= MUX_v_16_2_2(while_while_for_for_for_for_wy_idx_lpi_4_dfm_6,
          (while_while_for_for_for_for_acc_1_nl), while_while_for_for_and_7_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5)
        | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
        | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & reg_while_while_for_stage_0_cse
        ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4)
        | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0)
        & reg_while_while_for_stage_0_cse ) begin
      while_while_for_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4)
        | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & reg_while_while_for_stage_0_cse
        ) begin
      while_while_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_wx_idx_lpi_4 <= 16'b0000000000000000;
      while_while_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( while_while_for_for_for_wx_idx_and_2_cse ) begin
      while_while_for_for_for_wx_idx_lpi_4 <= MUX1HOT_v_16_3_2(while_while_for_for_for_wx_idx_lpi_4,
          while_while_for_for_for_wx_idx_lpi_4_dfm_5, (while_while_for_for_for_acc_1_nl),
          {(~ reg_while_while_for_stage_0_cse) , (while_while_for_for_for_wx_idx_and_nl)
          , (while_while_for_for_for_wx_idx_and_1_nl)});
      while_while_for_for_asn_sft_lpi_4 <= MUX_s_1_2_2(while_while_for_for_asn_sft_lpi_4,
          (while_while_for_for_for_mux_35_nl), reg_while_while_for_stage_0_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_co_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( run_wen & (mux_13_nl) & reg_while_while_for_stage_0_cse ) begin
      while_while_for_for_co_idx_lpi_4 <= MUX1HOT_v_16_3_2((while_while_for_for_acc_2_nl),
          while_while_for_for_co_idx_lpi_4, (signext_16_1(~ while_while_for_acc_3_itm_16_1)),
          {(and_53_nl) , (while_while_for_for_nand_nl) , (while_while_for_for_and_10_nl)});
    end
  end
  assign nl_block_size_mul_1_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[88:80]))
      * $signed(block_size_acc_cse_sva_mx0w0);
  assign block_size_mul_1_nl = nl_block_size_mul_1_nl[8:0];
  assign nl_block_size_mul_nl = $signed((block_size_mul_1_nl)) * $signed(block_size_acc_1_cse_sva_mx0w0);
  assign block_size_mul_nl = nl_block_size_mul_nl[8:0];
  assign nl_while_while_acc_nl = while_block_count_8_0_sva + 9'b000000001;
  assign while_while_acc_nl = nl_while_while_acc_nl[8:0];
  assign while_block_count_mux_nl = MUX_v_9_2_2(while_block_count_8_0_sva, (while_while_acc_nl),
      fsm_output[7]);
  assign while_block_count_not_nl = ~ or_tmp_55;
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_9_10(~ while_current_buffer_size_sva)
      + conv_u2u_9_10(~ block_size_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[9:0];
  assign nl_while_while_for_acc_2_nl = while_while_for_koo_idx_sva + 16'b0000000000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[15:0];
  assign while_while_for_koo_idx_and_1_nl = (~ or_47_tmp) & (fsm_output[6]);
  assign while_while_for_koo_idx_and_2_nl = or_47_tmp & (fsm_output[6]);
  assign while_while_for_koo_idx_mux1h_3_nl = MUX1HOT_v_16_3_2(({7'b0000000 , (readslicef_10_9_1((while_while_aelse_acc_1_nl)))}),
      (while_while_for_acc_2_nl), while_while_for_koo_idx_sva, {(fsm_output[4]) ,
      (while_while_for_koo_idx_and_1_nl) , (while_while_for_koo_idx_and_2_nl)});
  assign not_135_nl = ~ (fsm_output[5]);
  assign while_while_for_mux_3_nl = MUX_s_1_2_2(exitL_exit_while_while_for_for_sva,
      exit_while_while_for_for_lpi_4_dfm_mx1w0, reg_while_while_for_stage_0_cse);
  assign nl_while_while_acc_1_nl = total_blocks_lpi_3 + 32'b11111111111111111111111111111111;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[31:0];
  assign nl_while_while_acc_2_nl = while_current_buffer_size_sva + block_size_sva;
  assign while_while_acc_2_nl = nl_while_while_acc_2_nl[8:0];
  assign while_current_buffer_size_not_1_nl = ~ or_tmp_55;
  assign nand_4_nl = ~(lfst_exitL_exit_while_while_for_for_for_lpi_2 & while_while_for_for_asn_sft_lpi_4);
  assign mux_6_nl = MUX_s_1_2_2((nand_4_nl), while_while_for_for_acc_3_itm_16_1,
      or_1_cse);
  assign mux_7_nl = MUX_s_1_2_2((mux_6_nl), nor_tmp, exitL_exit_while_while_for_for_sva);
  assign nl_while_while_for_for_for_for_for_for_y_idx_lpi_4  = while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7
      + 16'b0000000000000001;
  assign nl_while_while_for_for_for_for_for_acc_1_nl = while_while_for_for_for_for_for_x_idx_lpi_4_dfm_7
      + 16'b0000000000000001;
  assign while_while_for_for_for_for_for_acc_1_nl = nl_while_while_for_for_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_for_and_5_nl = (~(while_while_for_for_for_for_for_for_acc_2_itm_16_1
      | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0)) & (~(while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0)) & while_while_for_for_not_62;
  assign nl_while_while_for_for_for_for_acc_1_nl = while_while_for_for_for_for_wy_idx_lpi_4_dfm_6
      + 16'b0000000000000001;
  assign while_while_for_for_for_for_acc_1_nl = nl_while_while_for_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_and_7_nl = exit_while_while_for_for_for_for_for_lpi_4_dfm_1
      & (~ while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & (~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0)) & (~ exit_while_while_for_lpi_4_dfm_1);
  assign nl_while_while_for_for_for_acc_1_nl = while_while_for_for_for_wx_idx_lpi_4_dfm_5
      + 16'b0000000000000001;
  assign while_while_for_for_for_acc_1_nl = nl_while_while_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_for_wx_idx_and_nl = (~ while_while_for_for_and_9_tmp)
      & reg_while_while_for_stage_0_cse;
  assign while_while_for_for_for_wx_idx_and_1_nl = while_while_for_for_and_9_tmp
      & reg_while_while_for_stage_0_cse;
  assign while_while_for_for_for_mux_35_nl = MUX_s_1_2_2(exit_while_while_for_for_lpi_4_dfm_mx1w0,
      while_while_for_for_asn_sft_lpi_4, lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3);
  assign nl_while_while_for_for_acc_2_nl = while_while_for_for_co_idx_lpi_4_dfm_1_mx0
      + 16'b0000000000000001;
  assign while_while_for_for_acc_2_nl = nl_while_while_for_for_acc_2_nl[15:0];
  assign and_53_nl = ((~((~(or_34_cse & (~ while_while_for_for_asn_sft_lpi_4))) &
      lfst_exitL_exit_while_while_for_for_for_lpi_2)) | or_dcpl_24) & (~ while_while_for_for_for_acc_2_itm_16_1)
      & reg_while_while_for_stage_0_cse;
  assign while_while_for_for_nand_nl = ~((~((~ exitL_exit_while_while_for_for_sva)
      & and_57_m1c)) & reg_while_while_for_stage_0_cse);
  assign while_while_for_for_and_10_nl = exitL_exit_while_while_for_for_sva & and_57_m1c;
  assign or_13_nl = (~((~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2))
      | while_while_for_for_acc_3_itm_16_1;
  assign mux_13_nl = MUX_s_1_2_2((or_13_nl), nor_tmp, exitL_exit_while_while_for_for_sva);

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [136:0] MUX_v_137_2_2;
    input [136:0] input_0;
    input [136:0] input_1;
    input [0:0] sel;
    reg [136:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_137_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input [0:0] vector;
  begin
    signext_16_1= {{15{vector[0]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, inputDoubleBufferWriterParams_cns_dat,
      inputDoubleBufferWriterParams_cns_vld, inputDoubleBufferWriterParams_cns_rdy,
      inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;



  // Interconnect Declarations for Component Instantiations 
  InputDoubleBuffer_512_16_16_run_run InputDoubleBuffer_512_16_16_run_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld),
      .inputDoubleBufferReaderParams_cns_rdy(inputDoubleBufferReaderParams_cns_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_csb, dout_rsc_web, dout_rsc_addr, dout_rsc_din,
      dout_rsc_dout, dout_rsc_req_vz, dout_rsc_rls_lz
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output dout_rsc_csb;
  output dout_rsc_web;
  output [11:0] dout_rsc_addr;
  output [127:0] dout_rsc_din;
  input [127:0] dout_rsc_dout;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;


  // Interconnect Declarations
  wire [11:0] dout_rsci_addr_d;
  wire [127:0] dout_rsci_din_d;
  wire [127:0] dout_rsci_dout_d;
  wire dout_rsci_web_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d;
  assign nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d = ~ dout_rsci_web_d_iff;
  InputDoubleBufferWriter_512_16_16_sram_512_128_sram_512_128_rwport_3_128_12_512_128_gen
      dout_rsci (
      .dout(dout_rsc_dout),
      .din(dout_rsc_din),
      .addr(dout_rsc_addr),
      .web(dout_rsc_web),
      .csb(dout_rsc_csb),
      .web_d(dout_rsci_web_d_iff),
      .addr_d(dout_rsci_addr_d),
      .din_d(dout_rsci_din_d),
      .dout_d(dout_rsci_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(1'b0),
      .port_0_rw_ram_ir_internal_WMASK_B_d(nl_dout_rsci_port_0_rw_ram_ir_internal_WMASK_B_d[0:0])
    );
  InputDoubleBufferWriter_512_16_16_run InputDoubleBufferWriter_512_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .dout_rsci_addr_d(dout_rsci_addr_d),
      .dout_rsci_din_d(dout_rsci_din_d),
      .dout_rsci_web_d_pff(dout_rsci_web_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_csb,
      din_rsc_web, din_rsc_addr, din_rsc_din, din_rsc_dout, din_rsc_req_vz, din_rsc_rls_lz,
      dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output din_rsc_csb;
  output din_rsc_web;
  output [11:0] din_rsc_addr;
  output [127:0] din_rsc_din;
  input [127:0] din_rsc_dout;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [11:0] din_rsci_addr_d;
  wire [127:0] din_rsci_dout_d;
  wire din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferReader_512_16_16_sram_512_128_sram_512_128_rwport_8_128_12_512_128_gen
      din_rsci (
      .dout(din_rsc_dout),
      .din(din_rsc_din),
      .addr(din_rsc_addr),
      .web(din_rsc_web),
      .csb(din_rsc_csb),
      .web_d(1'b1),
      .addr_d(din_rsci_addr_d),
      .din_d(128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
      .dout_d(din_rsci_dout_d),
      .port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d),
      .port_0_rw_ram_ir_internal_WMASK_B_d(1'b0)
    );
  InputDoubleBufferReader_512_16_16_run InputDoubleBufferReader_512_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_req_vz(din_rsc_req_vz),
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .din_rsci_addr_d(din_rsci_addr_d),
      .din_rsci_dout_d(din_rsci_dout_d),
      .din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d(din_rsci_port_0_rw_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_struct
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_struct (
  clk, arst_n, inputs_in_rsc_dat_value, inputs_in_rsc_vld, inputs_in_rsc_rdy, inputs_out_rsc_dat_value,
      inputs_out_rsc_vld, inputs_out_rsc_rdy, paramsIn_rsc_dat_STRIDE, paramsIn_rsc_dat_FY,
      paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1, paramsIn_rsc_dat_OC1, paramsIn_rsc_dat_OX0,
      paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1, paramsIn_rsc_dat_OY1, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputs_in_rsc_dat_value;
  input inputs_in_rsc_vld;
  output inputs_in_rsc_rdy;
  output [127:0] inputs_out_rsc_dat_value;
  output inputs_out_rsc_vld;
  input inputs_out_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] paramsIn_rsc_dat_ninputDoubleBufferWriter;
  wire paramsIn_rsc_vld_ninputDoubleBufferWriter;
  wire paramsIn_rsc_rdy_ninputDoubleBufferWriter;
  wire din_rsc_rdy_ninputDoubleBufferWriter;
  wire dout_rsc_csb_ninputDoubleBufferWriter;
  wire dout_rsc_web_ninputDoubleBufferWriter;
  wire [11:0] dout_rsc_addr_ninputDoubleBufferWriter;
  wire [127:0] dout_rsc_din_ninputDoubleBufferWriter;
  wire [127:0] dout_rsc_dout_ninputDoubleBufferWriter;
  wire dout_rsc_req_vz_ninputDoubleBufferWriter;
  wire paramsIn_rsc_rdy_ninputDoubleBufferReader;
  wire din_rsc_csb_ninputDoubleBufferReader;
  wire din_rsc_web_ninputDoubleBufferReader;
  wire [11:0] din_rsc_addr_ninputDoubleBufferReader;
  wire [127:0] din_rsc_din_ninputDoubleBufferReader;
  wire [127:0] din_rsc_dout_ninputDoubleBufferReader;
  wire din_rsc_req_vz_ninputDoubleBufferReader;
  wire [127:0] dout_rsc_dat_ninputDoubleBufferReader;
  wire dout_rsc_vld_ninputDoubleBufferReader;
  wire [143:0] inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst;
  wire inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst;
  wire [143:0] inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst;
  wire paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  wire inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire din_rsc_rdy_ninputDoubleBufferWriter_bud;
  wire dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  wire din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  wire inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire dout_rsc_vld_ninputDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire inputDoubleBufferWriterParams_unc_2;
  wire inputDoubleBufferWriterParams_idle;
  wire mem_cns_R0;
  wire mem_cns_R1;
  wire mem_cns_csb_shi0;
  wire mem_cns_csb_shi1;
  wire mem_cns_web_shi0;
  wire mem_cns_web_shi1;
  wire [11:0] mem_cns_addr_shi0;
  wire [11:0] mem_cns_addr_shi1;
  wire [127:0] mem_cns_din_shi0;
  wire [127:0] mem_cns_din_shi1;
  wire [127:0] mem_cns_dout_sho0;
  wire [127:0] mem_cns_dout_sho1;
  wire mem_cns_S1_iff;
  wire mem_cns_S0_iff;
  wire mem_cns_S0_dmo;
  wire mem_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat = {paramsIn_rsc_dat_STRIDE
      , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1 , paramsIn_rsc_dat_OC1
      , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1 , paramsIn_rsc_dat_OY1};
  ccs_pipe_v5 #(.rscid(32'sd15),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) inputDoubleBufferWriterParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst),
      .din_vld(inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .din(inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_ninputDoubleBufferWriter),
      .dout_vld(paramsIn_rsc_vld_ninputDoubleBufferWriter),
      .dout(paramsIn_rsc_dat_ninputDoubleBufferWriter),
      .sz(inputDoubleBufferWriterParams_unc_2),
      .sz_req(1'b0),
      .is_idle(inputDoubleBufferWriterParams_idle)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd128),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) mem_cns_comp (
      .clk(clk),
      .csb(mem_cns_csb_shi0),
      .web(mem_cns_web_shi0),
      .addr(mem_cns_addr_shi0),
      .din(mem_cns_din_shi0),
      .dout(mem_cns_dout_sho0)
    );
  sram_512_128 #(.WRAPPER_DEPTH(32'sd4096),
  .WRAPPER_WIDTH(32'sd128),
  .WRAPPER_ADDR_BITS(32'sd12),
  .SRAM_DEPTH(32'sd256),
  .SRAM_WIDTH(32'sd32),
  .SRAM_ADDR_BITS(32'sd8),
  .num_inst_depth(32'sd16),
  .num_inst_width(32'sd4)) mem_cns_comp_1 (
      .clk(clk),
      .csb(mem_cns_csb_shi1),
      .web(mem_cns_web_shi1),
      .addr(mem_cns_addr_shi1),
      .din(mem_cns_din_shi1),
      .dout(mem_cns_dout_sho1)
    );
  InputDoubleBufferWriter_512_16_16 inputDoubleBufferWriter (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_ninputDoubleBufferWriter),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_ninputDoubleBufferWriter),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud),
      .din_rsc_dat(inputs_in_rsc_dat_value),
      .din_rsc_vld(inputs_in_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy_ninputDoubleBufferWriter_bud),
      .dout_rsc_csb(dout_rsc_csb_ninputDoubleBufferWriter),
      .dout_rsc_web(dout_rsc_web_ninputDoubleBufferWriter),
      .dout_rsc_addr(dout_rsc_addr_ninputDoubleBufferWriter),
      .dout_rsc_din(dout_rsc_din_ninputDoubleBufferWriter),
      .dout_rsc_dout(dout_rsc_dout_ninputDoubleBufferWriter),
      .dout_rsc_req_vz(dout_rsc_req_vz_ninputDoubleBufferWriter),
      .dout_rsc_rls_lz(dout_rsc_rls_lz_ninputDoubleBufferWriter_bud)
    );
  InputDoubleBufferReader_512_16_16 inputDoubleBufferReader (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .paramsIn_rsc_vld(inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBufferReader_bud),
      .din_rsc_csb(din_rsc_csb_ninputDoubleBufferReader),
      .din_rsc_web(din_rsc_web_ninputDoubleBufferReader),
      .din_rsc_addr(din_rsc_addr_ninputDoubleBufferReader),
      .din_rsc_din(din_rsc_din_ninputDoubleBufferReader),
      .din_rsc_dout(din_rsc_dout_ninputDoubleBufferReader),
      .din_rsc_req_vz(din_rsc_req_vz_ninputDoubleBufferReader),
      .din_rsc_rls_lz(din_rsc_rls_lz_ninputDoubleBufferReader_bud),
      .dout_rsc_dat(dout_rsc_dat_ninputDoubleBufferReader),
      .dout_rsc_vld(dout_rsc_vld_ninputDoubleBufferReader_bud),
      .dout_rsc_rdy(inputs_out_rsc_rdy)
    );
  InputDoubleBuffer_512_16_16_run InputDoubleBuffer_512_16_16_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferReaderParams_cns_rdy(paramsIn_rsc_rdy_ninputDoubleBufferReader)
    );
  unreg_hier unreg (
      .in_0(mem_cns_S0_iff),
      .out_0(mem_cns_R0)
    );
  unreg_hier unreg_1 (
      .in_0(mem_cns_S1_iff),
      .out_0(mem_cns_R1)
    );
  InputDoubleBDjtfoem_cns_bctl InputDoubleBDjtfoem_cns_bctl_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_rdy_ninputDoubleBufferWriter(paramsIn_rsc_rdy_ninputDoubleBufferWriter),
      .din_rsc_rdy_ninputDoubleBufferWriter(din_rsc_rdy_ninputDoubleBufferWriter),
      .dout_rsc_csb_ninputDoubleBufferWriter(dout_rsc_csb_ninputDoubleBufferWriter),
      .dout_rsc_web_ninputDoubleBufferWriter(dout_rsc_web_ninputDoubleBufferWriter),
      .dout_rsc_addr_ninputDoubleBufferWriter(dout_rsc_addr_ninputDoubleBufferWriter),
      .dout_rsc_din_ninputDoubleBufferWriter(dout_rsc_din_ninputDoubleBufferWriter),
      .dout_rsc_dout_ninputDoubleBufferWriter(dout_rsc_dout_ninputDoubleBufferWriter),
      .dout_rsc_req_vz_ninputDoubleBufferWriter(dout_rsc_req_vz_ninputDoubleBufferWriter),
      .paramsIn_rsc_rdy_ninputDoubleBufferReader(paramsIn_rsc_rdy_ninputDoubleBufferReader),
      .din_rsc_csb_ninputDoubleBufferReader(din_rsc_csb_ninputDoubleBufferReader),
      .din_rsc_web_ninputDoubleBufferReader(din_rsc_web_ninputDoubleBufferReader),
      .din_rsc_addr_ninputDoubleBufferReader(din_rsc_addr_ninputDoubleBufferReader),
      .din_rsc_din_ninputDoubleBufferReader(din_rsc_din_ninputDoubleBufferReader),
      .din_rsc_dout_ninputDoubleBufferReader(din_rsc_dout_ninputDoubleBufferReader),
      .din_rsc_req_vz_ninputDoubleBufferReader(din_rsc_req_vz_ninputDoubleBufferReader),
      .dout_rsc_vld_ninputDoubleBufferReader(dout_rsc_vld_ninputDoubleBufferReader),
      .paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud(paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud),
      .din_rsc_rdy_ninputDoubleBufferWriter_bud(din_rsc_rdy_ninputDoubleBufferWriter_bud),
      .dout_rsc_rls_lz_ninputDoubleBufferWriter_bud(dout_rsc_rls_lz_ninputDoubleBufferWriter_bud),
      .din_rsc_rls_lz_ninputDoubleBufferReader_bud(din_rsc_rls_lz_ninputDoubleBufferReader_bud),
      .paramsIn_rsc_rdy_ninputDoubleBufferReader_bud(paramsIn_rsc_rdy_ninputDoubleBufferReader_bud),
      .dout_rsc_vld_ninputDoubleBufferReader_bud(dout_rsc_vld_ninputDoubleBufferReader_bud),
      .mem_cns_S0(mem_cns_S0_dmo),
      .mem_cns_R0(mem_cns_R0),
      .mem_cns_S1(mem_cns_S1_dmo),
      .mem_cns_R1(mem_cns_R1),
      .mem_cns_csb_shi0(mem_cns_csb_shi0),
      .mem_cns_csb_shi1(mem_cns_csb_shi1),
      .mem_cns_web_shi0(mem_cns_web_shi0),
      .mem_cns_web_shi1(mem_cns_web_shi1),
      .mem_cns_addr_shi0(mem_cns_addr_shi0),
      .mem_cns_addr_shi1(mem_cns_addr_shi1),
      .mem_cns_din_shi0(mem_cns_din_shi0),
      .mem_cns_din_shi1(mem_cns_din_shi1),
      .mem_cns_dout_sho0(mem_cns_dout_sho0),
      .mem_cns_dout_sho1(mem_cns_dout_sho1),
      .mem_cns_S1_pff(mem_cns_S1_iff),
      .mem_cns_S0_pff(mem_cns_S0_iff)
    );
  assign inputs_out_rsc_dat_value = dout_rsc_dat_ninputDoubleBufferReader;
  assign inputs_in_rsc_rdy = din_rsc_rdy_ninputDoubleBufferWriter;
  assign inputs_out_rsc_vld = dout_rsc_vld_ninputDoubleBufferReader;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16 (
  clk, arst_n, inputs_in_rsc_dat, inputs_in_rsc_vld, inputs_in_rsc_rdy, inputs_out_rsc_dat,
      inputs_out_rsc_vld, inputs_out_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputs_in_rsc_dat;
  input inputs_in_rsc_vld;
  output inputs_in_rsc_rdy;
  output [127:0] inputs_out_rsc_dat;
  output inputs_out_rsc_vld;
  input inputs_out_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [127:0] inputs_out_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1 = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1 = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0 = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0 = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1 = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1 = paramsIn_rsc_dat[15:0];
  InputDoubleBuffer_512_16_16_struct InputDoubleBuffer_512_16_16_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputs_in_rsc_dat_value(inputs_in_rsc_dat),
      .inputs_in_rsc_vld(inputs_in_rsc_vld),
      .inputs_in_rsc_rdy(inputs_in_rsc_rdy),
      .inputs_out_rsc_dat_value(inputs_out_rsc_dat_value),
      .inputs_out_rsc_vld(inputs_out_rsc_vld),
      .inputs_out_rsc_rdy(inputs_out_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy)
    );
  assign inputs_out_rsc_dat = inputs_out_rsc_dat_value;
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy07
//  Generated date: Sun Feb 23 19:47:57 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ParamsDeserializer_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;


  // FSM State Type Declaration for ParamsDeserializer_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8,
    main_C_8 = 4'd9,
    main_C_9 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ParamsDeserializer_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 11'b00000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_staller
// ------------------------------------------------------------------


module ParamsDeserializer_run_staller (
  run_wen, inputChannel_rsci_wen_comp, outputChannel1_rsci_wen_comp, outputChannel2_rsci_wen_comp,
      outputChannel3_rsci_wen_comp
);
  output run_wen;
  input inputChannel_rsci_wen_comp;
  input outputChannel1_rsci_wen_comp;
  input outputChannel2_rsci_wen_comp;
  input outputChannel3_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = inputChannel_rsci_wen_comp & outputChannel1_rsci_wen_comp & outputChannel2_rsci_wen_comp
      & outputChannel3_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp (
  clk, arst_n, outputChannel3_rsci_oswt, outputChannel3_rsci_wen_comp, outputChannel3_rsci_biwt,
      outputChannel3_rsci_bdwt, outputChannel3_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel3_rsci_oswt;
  output outputChannel3_rsci_wen_comp;
  input outputChannel3_rsci_biwt;
  input outputChannel3_rsci_bdwt;
  output outputChannel3_rsci_bcwt;
  reg outputChannel3_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel3_rsci_wen_comp = (~ outputChannel3_rsci_oswt) | outputChannel3_rsci_biwt
      | outputChannel3_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel3_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel3_rsci_bcwt <= ~((~(outputChannel3_rsci_bcwt | outputChannel3_rsci_biwt))
          | outputChannel3_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl (
  run_wen, outputChannel3_rsci_oswt, outputChannel3_rsci_irdy, outputChannel3_rsci_biwt,
      outputChannel3_rsci_bdwt, outputChannel3_rsci_bcwt, outputChannel3_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel3_rsci_oswt;
  input outputChannel3_rsci_irdy;
  output outputChannel3_rsci_biwt;
  output outputChannel3_rsci_bdwt;
  input outputChannel3_rsci_bcwt;
  output outputChannel3_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel3_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel3_rsci_bdwt = outputChannel3_rsci_oswt & run_wen;
  assign outputChannel3_rsci_biwt = outputChannel3_rsci_ogwt & outputChannel3_rsci_irdy;
  assign outputChannel3_rsci_ogwt = outputChannel3_rsci_oswt & (~ outputChannel3_rsci_bcwt);
  assign outputChannel3_rsci_ivld_run_sct = outputChannel3_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp (
  clk, arst_n, outputChannel2_rsci_oswt, outputChannel2_rsci_wen_comp, outputChannel2_rsci_biwt,
      outputChannel2_rsci_bdwt, outputChannel2_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel2_rsci_oswt;
  output outputChannel2_rsci_wen_comp;
  input outputChannel2_rsci_biwt;
  input outputChannel2_rsci_bdwt;
  output outputChannel2_rsci_bcwt;
  reg outputChannel2_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel2_rsci_wen_comp = (~ outputChannel2_rsci_oswt) | outputChannel2_rsci_biwt
      | outputChannel2_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel2_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel2_rsci_bcwt <= ~((~(outputChannel2_rsci_bcwt | outputChannel2_rsci_biwt))
          | outputChannel2_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl (
  run_wen, outputChannel2_rsci_oswt, outputChannel2_rsci_irdy, outputChannel2_rsci_biwt,
      outputChannel2_rsci_bdwt, outputChannel2_rsci_bcwt, outputChannel2_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel2_rsci_oswt;
  input outputChannel2_rsci_irdy;
  output outputChannel2_rsci_biwt;
  output outputChannel2_rsci_bdwt;
  input outputChannel2_rsci_bcwt;
  output outputChannel2_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel2_rsci_bdwt = outputChannel2_rsci_oswt & run_wen;
  assign outputChannel2_rsci_biwt = outputChannel2_rsci_ogwt & outputChannel2_rsci_irdy;
  assign outputChannel2_rsci_ogwt = outputChannel2_rsci_oswt & (~ outputChannel2_rsci_bcwt);
  assign outputChannel2_rsci_ivld_run_sct = outputChannel2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp (
  clk, arst_n, outputChannel1_rsci_oswt, outputChannel1_rsci_wen_comp, outputChannel1_rsci_biwt,
      outputChannel1_rsci_bdwt, outputChannel1_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel1_rsci_oswt;
  output outputChannel1_rsci_wen_comp;
  input outputChannel1_rsci_biwt;
  input outputChannel1_rsci_bdwt;
  output outputChannel1_rsci_bcwt;
  reg outputChannel1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel1_rsci_wen_comp = (~ outputChannel1_rsci_oswt) | outputChannel1_rsci_biwt
      | outputChannel1_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel1_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel1_rsci_bcwt <= ~((~(outputChannel1_rsci_bcwt | outputChannel1_rsci_biwt))
          | outputChannel1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl (
  run_wen, outputChannel1_rsci_oswt, outputChannel1_rsci_irdy, outputChannel1_rsci_biwt,
      outputChannel1_rsci_bdwt, outputChannel1_rsci_bcwt, outputChannel1_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel1_rsci_oswt;
  input outputChannel1_rsci_irdy;
  output outputChannel1_rsci_biwt;
  output outputChannel1_rsci_bdwt;
  input outputChannel1_rsci_bcwt;
  output outputChannel1_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel1_rsci_bdwt = outputChannel1_rsci_oswt & run_wen;
  assign outputChannel1_rsci_biwt = outputChannel1_rsci_ogwt & outputChannel1_rsci_irdy;
  assign outputChannel1_rsci_ogwt = outputChannel1_rsci_oswt & (~ outputChannel1_rsci_bcwt);
  assign outputChannel1_rsci_ivld_run_sct = outputChannel1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp (
  clk, arst_n, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt,
      inputChannel_rsci_biwt, inputChannel_rsci_bdwt, inputChannel_rsci_bcwt, inputChannel_rsci_idat
);
  input clk;
  input arst_n;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [15:0] inputChannel_rsci_idat_mxwt;
  input inputChannel_rsci_biwt;
  input inputChannel_rsci_bdwt;
  output inputChannel_rsci_bcwt;
  reg inputChannel_rsci_bcwt;
  input [15:0] inputChannel_rsci_idat;


  // Interconnect Declarations
  reg [15:0] inputChannel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_wen_comp = (~ inputChannel_rsci_oswt) | inputChannel_rsci_biwt
      | inputChannel_rsci_bcwt;
  assign inputChannel_rsci_idat_mxwt = MUX_v_16_2_2(inputChannel_rsci_idat, inputChannel_rsci_idat_bfwt,
      inputChannel_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      inputChannel_rsci_bcwt <= ~((~(inputChannel_rsci_bcwt | inputChannel_rsci_biwt))
          | inputChannel_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ inputChannel_rsci_bcwt ) begin
      inputChannel_rsci_idat_bfwt <= inputChannel_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl (
  run_wen, inputChannel_rsci_oswt, inputChannel_rsci_biwt, inputChannel_rsci_bdwt,
      inputChannel_rsci_bcwt, inputChannel_rsci_irdy_run_sct, inputChannel_rsci_ivld
);
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_biwt;
  output inputChannel_rsci_bdwt;
  input inputChannel_rsci_bcwt;
  output inputChannel_rsci_irdy_run_sct;
  input inputChannel_rsci_ivld;


  // Interconnect Declarations
  wire inputChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_bdwt = inputChannel_rsci_oswt & run_wen;
  assign inputChannel_rsci_biwt = inputChannel_rsci_ogwt & inputChannel_rsci_ivld;
  assign inputChannel_rsci_ogwt = inputChannel_rsci_oswt & (~ inputChannel_rsci_bcwt);
  assign inputChannel_rsci_irdy_run_sct = inputChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller (
  run_wen, inputChannel_rsci_wen_comp, serialOutChannel_rsci_wen_comp
);
  output run_wen;
  input inputChannel_rsci_wen_comp;
  input serialOutChannel_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = inputChannel_rsci_wen_comp & serialOutChannel_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
    (
  clk, arst_n, serialOutChannel_rsci_oswt, serialOutChannel_rsci_wen_comp, serialOutChannel_rsci_biwt,
      serialOutChannel_rsci_bdwt, serialOutChannel_rsci_bcwt
);
  input clk;
  input arst_n;
  input serialOutChannel_rsci_oswt;
  output serialOutChannel_rsci_wen_comp;
  input serialOutChannel_rsci_biwt;
  input serialOutChannel_rsci_bdwt;
  output serialOutChannel_rsci_bcwt;
  reg serialOutChannel_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign serialOutChannel_rsci_wen_comp = (~ serialOutChannel_rsci_oswt) | serialOutChannel_rsci_biwt
      | serialOutChannel_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      serialOutChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      serialOutChannel_rsci_bcwt <= ~((~(serialOutChannel_rsci_bcwt | serialOutChannel_rsci_biwt))
          | serialOutChannel_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
    (
  run_wen, serialOutChannel_rsci_oswt, serialOutChannel_rsci_irdy, serialOutChannel_rsci_biwt,
      serialOutChannel_rsci_bdwt, serialOutChannel_rsci_bcwt, serialOutChannel_rsci_ivld_run_sct
);
  input run_wen;
  input serialOutChannel_rsci_oswt;
  input serialOutChannel_rsci_irdy;
  output serialOutChannel_rsci_biwt;
  output serialOutChannel_rsci_bdwt;
  input serialOutChannel_rsci_bcwt;
  output serialOutChannel_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire serialOutChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign serialOutChannel_rsci_bdwt = serialOutChannel_rsci_oswt & run_wen;
  assign serialOutChannel_rsci_biwt = serialOutChannel_rsci_ogwt & serialOutChannel_rsci_irdy;
  assign serialOutChannel_rsci_ogwt = serialOutChannel_rsci_oswt & (~ serialOutChannel_rsci_bcwt);
  assign serialOutChannel_rsci_ivld_run_sct = serialOutChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
    (
  clk, arst_n, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt,
      inputChannel_rsci_biwt, inputChannel_rsci_bdwt, inputChannel_rsci_bcwt, inputChannel_rsci_idat
);
  input clk;
  input arst_n;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [255:0] inputChannel_rsci_idat_mxwt;
  input inputChannel_rsci_biwt;
  input inputChannel_rsci_bdwt;
  output inputChannel_rsci_bcwt;
  reg inputChannel_rsci_bcwt;
  input [255:0] inputChannel_rsci_idat;


  // Interconnect Declarations
  reg [255:0] inputChannel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_wen_comp = (~ inputChannel_rsci_oswt) | inputChannel_rsci_biwt
      | inputChannel_rsci_bcwt;
  assign inputChannel_rsci_idat_mxwt = MUX_v_256_2_2(inputChannel_rsci_idat, inputChannel_rsci_idat_bfwt,
      inputChannel_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      inputChannel_rsci_bcwt <= ~((~(inputChannel_rsci_bcwt | inputChannel_rsci_biwt))
          | inputChannel_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_idat_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ inputChannel_rsci_bcwt ) begin
      inputChannel_rsci_idat_bfwt <= inputChannel_rsci_idat_mxwt;
    end
  end

  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
    (
  run_wen, inputChannel_rsci_oswt, inputChannel_rsci_biwt, inputChannel_rsci_bdwt,
      inputChannel_rsci_bcwt, inputChannel_rsci_irdy_run_sct, inputChannel_rsci_ivld
);
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_biwt;
  output inputChannel_rsci_bdwt;
  input inputChannel_rsci_bcwt;
  output inputChannel_rsci_irdy_run_sct;
  input inputChannel_rsci_ivld;


  // Interconnect Declarations
  wire inputChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_bdwt = inputChannel_rsci_oswt & run_wen;
  assign inputChannel_rsci_biwt = inputChannel_rsci_ogwt & inputChannel_rsci_ivld;
  assign inputChannel_rsci_ogwt = inputChannel_rsci_oswt & (~ inputChannel_rsci_bcwt);
  assign inputChannel_rsci_irdy_run_sct = inputChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module SystolicArrayLooper_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_0_tr0, xy_o_C_0_tr0, OC2_C_0_tr0, co_C_0_tr0,
      winx_C_0_tr0, winy_C_0_tr0, winx_C_1_tr0, co_C_1_tr0, OC2_C_1_tr0, xy_o_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input main_C_0_tr0;
  input xy_o_C_0_tr0;
  input OC2_C_0_tr0;
  input co_C_0_tr0;
  input winx_C_0_tr0;
  input winy_C_0_tr0;
  input winx_C_1_tr0;
  input co_C_1_tr0;
  input OC2_C_1_tr0;
  input xy_o_C_1_tr0;


  // FSM State Type Declaration for SystolicArrayLooper_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    xy_o_C_0 = 4'd2,
    OC2_C_0 = 4'd3,
    co_C_0 = 4'd4,
    winx_C_0 = 4'd5,
    winy_C_0 = 4'd6,
    winx_C_1 = 4'd7,
    co_C_1 = 4'd8,
    OC2_C_1 = 4'd9,
    xy_o_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SystolicArrayLooper_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 11'b00000000010;
        if ( main_C_0_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = xy_o_C_0;
        end
      end
      xy_o_C_0 : begin
        fsm_output = 11'b00000000100;
        if ( xy_o_C_0_tr0 ) begin
          state_var_NS = xy_o_C_1;
        end
        else begin
          state_var_NS = OC2_C_0;
        end
      end
      OC2_C_0 : begin
        fsm_output = 11'b00000001000;
        if ( OC2_C_0_tr0 ) begin
          state_var_NS = OC2_C_1;
        end
        else begin
          state_var_NS = co_C_0;
        end
      end
      co_C_0 : begin
        fsm_output = 11'b00000010000;
        if ( co_C_0_tr0 ) begin
          state_var_NS = co_C_1;
        end
        else begin
          state_var_NS = winx_C_0;
        end
      end
      winx_C_0 : begin
        fsm_output = 11'b00000100000;
        if ( winx_C_0_tr0 ) begin
          state_var_NS = winx_C_1;
        end
        else begin
          state_var_NS = winy_C_0;
        end
      end
      winy_C_0 : begin
        fsm_output = 11'b00001000000;
        if ( winy_C_0_tr0 ) begin
          state_var_NS = winx_C_1;
        end
        else begin
          state_var_NS = winy_C_0;
        end
      end
      winx_C_1 : begin
        fsm_output = 11'b00010000000;
        if ( winx_C_1_tr0 ) begin
          state_var_NS = co_C_1;
        end
        else begin
          state_var_NS = winx_C_0;
        end
      end
      co_C_1 : begin
        fsm_output = 11'b00100000000;
        if ( co_C_1_tr0 ) begin
          state_var_NS = OC2_C_1;
        end
        else begin
          state_var_NS = co_C_0;
        end
      end
      OC2_C_1 : begin
        fsm_output = 11'b01000000000;
        if ( OC2_C_1_tr0 ) begin
          state_var_NS = xy_o_C_1;
        end
        else begin
          state_var_NS = OC2_C_0;
        end
      end
      xy_o_C_1 : begin
        fsm_output = 11'b10000000000;
        if ( xy_o_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = xy_o_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_staller
// ------------------------------------------------------------------


module SystolicArrayLooper_run_staller (
  run_wen, paramsIn_rsci_wen_comp, paramsOut_rsci_wen_comp, loopIndicesOut_rsci_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input paramsOut_rsci_wen_comp;
  input loopIndicesOut_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & paramsOut_rsci_wen_comp & loopIndicesOut_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp (
  clk, arst_n, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input loopIndicesOut_rsci_biwt;
  input loopIndicesOut_rsci_bdwt;
  output loopIndicesOut_rsci_bcwt;
  reg loopIndicesOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_wen_comp = (~ loopIndicesOut_rsci_oswt) | loopIndicesOut_rsci_biwt
      | loopIndicesOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_bcwt <= 1'b0;
    end
    else begin
      loopIndicesOut_rsci_bcwt <= ~((~(loopIndicesOut_rsci_bcwt | loopIndicesOut_rsci_biwt))
          | loopIndicesOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl (
  run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_irdy, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt, loopIndicesOut_rsci_ivld_run_sct
);
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  input loopIndicesOut_rsci_irdy;
  output loopIndicesOut_rsci_biwt;
  output loopIndicesOut_rsci_bdwt;
  input loopIndicesOut_rsci_bcwt;
  output loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_bdwt = loopIndicesOut_rsci_oswt & run_wen;
  assign loopIndicesOut_rsci_biwt = loopIndicesOut_rsci_ogwt & loopIndicesOut_rsci_irdy;
  assign loopIndicesOut_rsci_ogwt = loopIndicesOut_rsci_oswt & (~ loopIndicesOut_rsci_bcwt);
  assign loopIndicesOut_rsci_ivld_run_sct = loopIndicesOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp (
  clk, arst_n, paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_biwt,
      paramsOut_rsci_bdwt, paramsOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input paramsOut_rsci_biwt;
  input paramsOut_rsci_bdwt;
  output paramsOut_rsci_bcwt;
  reg paramsOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_wen_comp = (~ paramsOut_rsci_oswt) | paramsOut_rsci_biwt
      | paramsOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsOut_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsOut_rsci_bcwt <= ~((~(paramsOut_rsci_bcwt | paramsOut_rsci_biwt)) | paramsOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl (
  run_wen, paramsOut_rsci_oswt, paramsOut_rsci_irdy, paramsOut_rsci_biwt, paramsOut_rsci_bdwt,
      paramsOut_rsci_bcwt, paramsOut_rsci_ivld_run_sct
);
  input run_wen;
  input paramsOut_rsci_oswt;
  input paramsOut_rsci_irdy;
  output paramsOut_rsci_biwt;
  output paramsOut_rsci_bdwt;
  input paramsOut_rsci_bcwt;
  output paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire paramsOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_bdwt = paramsOut_rsci_oswt & run_wen;
  assign paramsOut_rsci_biwt = paramsOut_rsci_ogwt & paramsOut_rsci_irdy;
  assign paramsOut_rsci_ogwt = paramsOut_rsci_oswt & (~ paramsOut_rsci_bcwt);
  assign paramsOut_rsci_ivld_run_sct = paramsOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci (
  clk, arst_n, outputChannel3_rsc_dat, outputChannel3_rsc_vld, outputChannel3_rsc_rdy,
      run_wen, outputChannel3_rsci_oswt, outputChannel3_rsci_wen_comp, outputChannel3_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;
  input run_wen;
  input outputChannel3_rsci_oswt;
  output outputChannel3_rsci_wen_comp;
  input [143:0] outputChannel3_rsci_idat;


  // Interconnect Declarations
  wire outputChannel3_rsci_irdy;
  wire outputChannel3_rsci_biwt;
  wire outputChannel3_rsci_bdwt;
  wire outputChannel3_rsci_bcwt;
  wire outputChannel3_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd144)) outputChannel3_rsci (
      .irdy(outputChannel3_rsci_irdy),
      .ivld(outputChannel3_rsci_ivld_run_sct),
      .idat(outputChannel3_rsci_idat),
      .rdy(outputChannel3_rsc_rdy),
      .vld(outputChannel3_rsc_vld),
      .dat(outputChannel3_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel3_rsci_oswt(outputChannel3_rsci_oswt),
      .outputChannel3_rsci_irdy(outputChannel3_rsci_irdy),
      .outputChannel3_rsci_biwt(outputChannel3_rsci_biwt),
      .outputChannel3_rsci_bdwt(outputChannel3_rsci_bdwt),
      .outputChannel3_rsci_bcwt(outputChannel3_rsci_bcwt),
      .outputChannel3_rsci_ivld_run_sct(outputChannel3_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel3_rsci_oswt(outputChannel3_rsci_oswt),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp),
      .outputChannel3_rsci_biwt(outputChannel3_rsci_biwt),
      .outputChannel3_rsci_bdwt(outputChannel3_rsci_bdwt),
      .outputChannel3_rsci_bcwt(outputChannel3_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci (
  clk, arst_n, outputChannel2_rsc_dat, outputChannel2_rsc_vld, outputChannel2_rsc_rdy,
      run_wen, outputChannel2_rsci_oswt, outputChannel2_rsci_wen_comp, outputChannel2_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  input run_wen;
  input outputChannel2_rsci_oswt;
  output outputChannel2_rsci_wen_comp;
  input [143:0] outputChannel2_rsci_idat;


  // Interconnect Declarations
  wire outputChannel2_rsci_irdy;
  wire outputChannel2_rsci_biwt;
  wire outputChannel2_rsci_bdwt;
  wire outputChannel2_rsci_bcwt;
  wire outputChannel2_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd144)) outputChannel2_rsci (
      .irdy(outputChannel2_rsci_irdy),
      .ivld(outputChannel2_rsci_ivld_run_sct),
      .idat(outputChannel2_rsci_idat),
      .rdy(outputChannel2_rsc_rdy),
      .vld(outputChannel2_rsc_vld),
      .dat(outputChannel2_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel2_rsci_oswt(outputChannel2_rsci_oswt),
      .outputChannel2_rsci_irdy(outputChannel2_rsci_irdy),
      .outputChannel2_rsci_biwt(outputChannel2_rsci_biwt),
      .outputChannel2_rsci_bdwt(outputChannel2_rsci_bdwt),
      .outputChannel2_rsci_bcwt(outputChannel2_rsci_bcwt),
      .outputChannel2_rsci_ivld_run_sct(outputChannel2_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel2_rsci_oswt(outputChannel2_rsci_oswt),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel2_rsci_biwt(outputChannel2_rsci_biwt),
      .outputChannel2_rsci_bdwt(outputChannel2_rsci_bdwt),
      .outputChannel2_rsci_bcwt(outputChannel2_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci (
  clk, arst_n, outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy,
      run_wen, outputChannel1_rsci_oswt, outputChannel1_rsci_wen_comp, outputChannel1_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  input run_wen;
  input outputChannel1_rsci_oswt;
  output outputChannel1_rsci_wen_comp;
  input [143:0] outputChannel1_rsci_idat;


  // Interconnect Declarations
  wire outputChannel1_rsci_irdy;
  wire outputChannel1_rsci_biwt;
  wire outputChannel1_rsci_bdwt;
  wire outputChannel1_rsci_bcwt;
  wire outputChannel1_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd144)) outputChannel1_rsci (
      .irdy(outputChannel1_rsci_irdy),
      .ivld(outputChannel1_rsci_ivld_run_sct),
      .idat(outputChannel1_rsci_idat),
      .rdy(outputChannel1_rsc_rdy),
      .vld(outputChannel1_rsc_vld),
      .dat(outputChannel1_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel1_rsci_oswt(outputChannel1_rsci_oswt),
      .outputChannel1_rsci_irdy(outputChannel1_rsci_irdy),
      .outputChannel1_rsci_biwt(outputChannel1_rsci_biwt),
      .outputChannel1_rsci_bdwt(outputChannel1_rsci_bdwt),
      .outputChannel1_rsci_bcwt(outputChannel1_rsci_bcwt),
      .outputChannel1_rsci_ivld_run_sct(outputChannel1_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel1_rsci_oswt(outputChannel1_rsci_oswt),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel1_rsci_biwt(outputChannel1_rsci_biwt),
      .outputChannel1_rsci_bdwt(outputChannel1_rsci_bdwt),
      .outputChannel1_rsci_bcwt(outputChannel1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      run_wen, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [15:0] inputChannel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire inputChannel_rsci_biwt;
  wire inputChannel_rsci_bdwt;
  wire inputChannel_rsci_bcwt;
  wire inputChannel_rsci_irdy_run_sct;
  wire inputChannel_rsci_ivld;
  wire [15:0] inputChannel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd16)) inputChannel_rsci (
      .rdy(inputChannel_rsc_rdy),
      .vld(inputChannel_rsc_vld),
      .dat(inputChannel_rsc_dat),
      .irdy(inputChannel_rsci_irdy_run_sct),
      .ivld(inputChannel_rsci_ivld),
      .idat(inputChannel_rsci_idat)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_irdy_run_sct(inputChannel_rsci_irdy_run_sct),
      .inputChannel_rsci_ivld(inputChannel_rsci_ivld)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_idat(inputChannel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci (
  clk, arst_n, serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy,
      run_wen, serialOutChannel_rsci_oswt, serialOutChannel_rsci_wen_comp, serialOutChannel_rsci_idat
);
  input clk;
  input arst_n;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;
  input run_wen;
  input serialOutChannel_rsci_oswt;
  output serialOutChannel_rsci_wen_comp;
  input [15:0] serialOutChannel_rsci_idat;


  // Interconnect Declarations
  wire serialOutChannel_rsci_irdy;
  wire serialOutChannel_rsci_biwt;
  wire serialOutChannel_rsci_bdwt;
  wire serialOutChannel_rsci_bcwt;
  wire serialOutChannel_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd6),
  .width(32'sd16)) serialOutChannel_rsci (
      .irdy(serialOutChannel_rsci_irdy),
      .ivld(serialOutChannel_rsci_ivld_run_sct),
      .idat(serialOutChannel_rsci_idat),
      .rdy(serialOutChannel_rsc_rdy),
      .vld(serialOutChannel_rsc_vld),
      .dat(serialOutChannel_rsc_dat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .serialOutChannel_rsci_oswt(serialOutChannel_rsci_oswt),
      .serialOutChannel_rsci_irdy(serialOutChannel_rsci_irdy),
      .serialOutChannel_rsci_biwt(serialOutChannel_rsci_biwt),
      .serialOutChannel_rsci_bdwt(serialOutChannel_rsci_bdwt),
      .serialOutChannel_rsci_bcwt(serialOutChannel_rsci_bcwt),
      .serialOutChannel_rsci_ivld_run_sct(serialOutChannel_rsci_ivld_run_sct)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .serialOutChannel_rsci_oswt(serialOutChannel_rsci_oswt),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp),
      .serialOutChannel_rsci_biwt(serialOutChannel_rsci_biwt),
      .serialOutChannel_rsci_bdwt(serialOutChannel_rsci_bdwt),
      .serialOutChannel_rsci_bcwt(serialOutChannel_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      run_wen, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [255:0] inputChannel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire inputChannel_rsci_biwt;
  wire inputChannel_rsci_bdwt;
  wire inputChannel_rsci_bcwt;
  wire inputChannel_rsci_irdy_run_sct;
  wire inputChannel_rsci_ivld;
  wire [255:0] inputChannel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd256)) inputChannel_rsci (
      .rdy(inputChannel_rsc_rdy),
      .vld(inputChannel_rsc_vld),
      .dat(inputChannel_rsc_dat),
      .irdy(inputChannel_rsci_irdy_run_sct),
      .ivld(inputChannel_rsci_ivld),
      .idat(inputChannel_rsci_idat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_irdy_run_sct(inputChannel_rsci_irdy_run_sct),
      .inputChannel_rsci_ivld(inputChannel_rsci_ivld)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_idat(inputChannel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci (
  clk, arst_n, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld, loopIndicesOut_rsc_rdy,
      run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_idat
);
  input clk;
  input arst_n;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input [47:0] loopIndicesOut_rsci_idat;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_irdy;
  wire loopIndicesOut_rsci_biwt;
  wire loopIndicesOut_rsci_bdwt;
  wire loopIndicesOut_rsci_bcwt;
  wire loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd158),
  .width(32'sd48)) loopIndicesOut_rsci (
      .irdy(loopIndicesOut_rsci_irdy),
      .ivld(loopIndicesOut_rsci_ivld_run_sct),
      .idat(loopIndicesOut_rsci_idat),
      .rdy(loopIndicesOut_rsc_rdy),
      .vld(loopIndicesOut_rsc_vld),
      .dat(loopIndicesOut_rsc_dat)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_irdy(loopIndicesOut_rsci_irdy),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt),
      .loopIndicesOut_rsci_ivld_run_sct(loopIndicesOut_rsci_ivld_run_sct)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci (
  clk, arst_n, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy, run_wen,
      paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  input run_wen;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input [143:0] paramsOut_rsci_idat;


  // Interconnect Declarations
  wire paramsOut_rsci_irdy;
  wire paramsOut_rsci_biwt;
  wire paramsOut_rsci_bdwt;
  wire paramsOut_rsci_bcwt;
  wire paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd157),
  .width(32'sd144)) paramsOut_rsci (
      .irdy(paramsOut_rsci_irdy),
      .ivld(paramsOut_rsci_ivld_run_sct),
      .idat(paramsOut_rsci_idat),
      .rdy(paramsOut_rsc_rdy),
      .vld(paramsOut_rsc_vld),
      .dat(paramsOut_rsc_dat)
    );
  SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_irdy(paramsOut_rsci_irdy),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt),
      .paramsOut_rsci_ivld_run_sct(paramsOut_rsci_ivld_run_sct)
    );
  SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd156),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run
// ------------------------------------------------------------------


module ParamsDeserializer_run (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy, outputChannel2_rsc_dat,
      outputChannel2_rsc_vld, outputChannel2_rsc_rdy, outputChannel3_rsc_dat, outputChannel3_rsc_vld,
      outputChannel3_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire inputChannel_rsci_wen_comp;
  wire [15:0] inputChannel_rsci_idat_mxwt;
  wire outputChannel1_rsci_wen_comp;
  wire outputChannel2_rsci_wen_comp;
  wire outputChannel3_rsci_wen_comp;
  wire [10:0] fsm_output;
  wire outputChannel3_and_cse;
  reg reg_outputChannel3_rsci_ivld_run_psct_cse;
  reg reg_inputChannel_rsci_irdy_run_psct_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_15_0_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_31_16_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_47_32_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_63_48_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_79_64_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_95_80_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_111_96_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_127_112_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_143_128_cse;
  reg [15:0] params_OY1_sva;
  reg [15:0] params_OX1_sva;
  reg [15:0] params_OY0_sva;
  reg [15:0] params_OX0_sva;
  reg [15:0] params_OC1_sva;
  reg [15:0] params_IC1_sva;
  reg [15:0] params_FX_sva;
  reg [15:0] params_FY_sva;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  wire [143:0] nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  wire [143:0] nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  ParamsDeserializer_run_inputChannel_rsci ParamsDeserializer_run_inputChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(reg_inputChannel_rsci_irdy_run_psct_cse),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt)
    );
  ParamsDeserializer_run_outputChannel1_rsci ParamsDeserializer_run_outputChannel1_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel1_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel1_rsci_idat(nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat[143:0])
    );
  ParamsDeserializer_run_outputChannel2_rsci ParamsDeserializer_run_outputChannel2_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel2_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel2_rsci_idat(nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat[143:0])
    );
  ParamsDeserializer_run_outputChannel3_rsci ParamsDeserializer_run_outputChannel3_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel3_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp),
      .outputChannel3_rsci_idat(nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat[143:0])
    );
  ParamsDeserializer_run_staller ParamsDeserializer_run_staller_inst (
      .run_wen(run_wen),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp)
    );
  ParamsDeserializer_run_run_fsm ParamsDeserializer_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign outputChannel3_and_cse = run_wen & (fsm_output[9]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_outputChannel3_rsci_idat_15_0_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_31_16_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_47_32_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_63_48_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_79_64_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_95_80_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_111_96_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_127_112_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_143_128_cse <= 16'b0000000000000000;
    end
    else if ( outputChannel3_and_cse ) begin
      reg_outputChannel3_rsci_idat_15_0_cse <= params_OY1_sva;
      reg_outputChannel3_rsci_idat_31_16_cse <= params_OX1_sva;
      reg_outputChannel3_rsci_idat_47_32_cse <= params_OY0_sva;
      reg_outputChannel3_rsci_idat_63_48_cse <= params_OX0_sva;
      reg_outputChannel3_rsci_idat_79_64_cse <= params_OC1_sva;
      reg_outputChannel3_rsci_idat_95_80_cse <= params_IC1_sva;
      reg_outputChannel3_rsci_idat_111_96_cse <= params_FX_sva;
      reg_outputChannel3_rsci_idat_127_112_cse <= params_FY_sva;
      reg_outputChannel3_rsci_idat_143_128_cse <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_outputChannel3_rsci_ivld_run_psct_cse <= 1'b0;
      reg_inputChannel_rsci_irdy_run_psct_cse <= 1'b0;
      params_FY_sva <= 16'b0000000000000000;
    end
    else if ( run_wen ) begin
      reg_outputChannel3_rsci_ivld_run_psct_cse <= fsm_output[9];
      reg_inputChannel_rsci_irdy_run_psct_cse <= ~ (fsm_output[9]);
      params_FY_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OY1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      params_OY1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OX1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      params_OX1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OY0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[3]) ) begin
      params_OY0_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OX0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[4]) ) begin
      params_OX0_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OC1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[5]) ) begin
      params_OC1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_IC1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[6]) ) begin
      params_IC1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_FX_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[7]) ) begin
      params_FX_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire inputChannel_rsci_wen_comp;
  wire [255:0] inputChannel_rsci_idat_mxwt;
  wire serialOutChannel_rsci_wen_comp;
  reg [15:0] serialOutChannel_rsci_idat;
  wire [1:0] fsm_output;
  reg exitL_exit_for_sva;
  wire [4:0] for_i_4_0_sva_3;
  wire [5:0] nl_for_i_4_0_sva_3;
  reg reg_inputChannel_rsci_oswt_cse;
  reg reg_serialOutChannel_rsci_ivld_run_psct_cse;
  wire serialOutChannel_and_cse;
  reg [255:0] input_value_lpi_1_dfm;
  wire [255:0] input_value_lpi_1_dfm_mx0;
  wire [3:0] for_i_4_0_lpi_1_dfm_3_0_1;
  reg [3:0] for_i_4_0_sva_1_3_0;

  wire[0:0] for_not_nl;

  // Interconnect Declarations for Component Instantiations 
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(reg_inputChannel_rsci_oswt_cse),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld),
      .serialOutChannel_rsc_rdy(serialOutChannel_rsc_rdy),
      .run_wen(run_wen),
      .serialOutChannel_rsci_oswt(reg_serialOutChannel_rsci_ivld_run_psct_cse),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp),
      .serialOutChannel_rsci_idat(serialOutChannel_rsci_idat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign serialOutChannel_and_cse = run_wen & (~ (fsm_output[0]));
  assign input_value_lpi_1_dfm_mx0 = MUX_v_256_2_2(input_value_lpi_1_dfm, inputChannel_rsci_idat_mxwt,
      exitL_exit_for_sva);
  assign nl_for_i_4_0_sva_3 = conv_u2s_4_5(for_i_4_0_lpi_1_dfm_3_0_1) + 5'b00001;
  assign for_i_4_0_sva_3 = nl_for_i_4_0_sva_3[4:0];
  assign for_not_nl = ~ exitL_exit_for_sva;
  assign for_i_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, for_i_4_0_sva_1_3_0, (for_not_nl));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputChannel_rsci_oswt_cse <= 1'b0;
      reg_serialOutChannel_rsci_ivld_run_psct_cse <= 1'b0;
      for_i_4_0_sva_1_3_0 <= 4'b0000;
    end
    else if ( run_wen ) begin
      reg_inputChannel_rsci_oswt_cse <= ~((~ (for_i_4_0_sva_3[4])) & (fsm_output[1]));
      reg_serialOutChannel_rsci_ivld_run_psct_cse <= fsm_output[1];
      for_i_4_0_sva_1_3_0 <= for_i_4_0_sva_3[3:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      serialOutChannel_rsci_idat <= 16'b0000000000000000;
      exitL_exit_for_sva <= 1'b1;
    end
    else if ( serialOutChannel_and_cse ) begin
      serialOutChannel_rsci_idat <= MUX_v_16_16_2((input_value_lpi_1_dfm_mx0[15:0]),
          (input_value_lpi_1_dfm_mx0[31:16]), (input_value_lpi_1_dfm_mx0[47:32]),
          (input_value_lpi_1_dfm_mx0[63:48]), (input_value_lpi_1_dfm_mx0[79:64]),
          (input_value_lpi_1_dfm_mx0[95:80]), (input_value_lpi_1_dfm_mx0[111:96]),
          (input_value_lpi_1_dfm_mx0[127:112]), (input_value_lpi_1_dfm_mx0[143:128]),
          (input_value_lpi_1_dfm_mx0[159:144]), (input_value_lpi_1_dfm_mx0[175:160]),
          (input_value_lpi_1_dfm_mx0[191:176]), (input_value_lpi_1_dfm_mx0[207:192]),
          (input_value_lpi_1_dfm_mx0[223:208]), (input_value_lpi_1_dfm_mx0[239:224]),
          (input_value_lpi_1_dfm_mx0[255:240]), for_i_4_0_lpi_1_dfm_3_0_1);
      exitL_exit_for_sva <= for_i_4_0_sva_3[4];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_value_lpi_1_dfm <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (~ (for_i_4_0_sva_3[4])) & run_wen & exitL_exit_for_sva ) begin
      input_value_lpi_1_dfm <= input_value_lpi_1_dfm_mx0;
    end
  end

  function automatic [15:0] MUX_v_16_16_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run
// ------------------------------------------------------------------


module SystolicArrayLooper_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat,
      paramsOut_rsc_vld, paramsOut_rsc_rdy, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld,
      loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire paramsOut_rsci_wen_comp;
  reg [143:0] paramsOut_rsci_idat;
  wire loopIndicesOut_rsci_wen_comp;
  reg [15:0] loopIndicesOut_rsci_idat_47_32;
  reg [15:0] loopIndicesOut_rsci_idat_31_16;
  reg [15:0] loopIndicesOut_rsci_idat_15_0;
  wire [10:0] fsm_output;
  wire and_dcpl_3;
  wire loopIndicesOut_and_cse;
  reg reg_loopIndicesOut_rsci_ivld_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
  wire [15:0] z_out_1;
  wire [16:0] nl_z_out_1;
  reg [143:0] paramsIn_crt_sva;
  reg [15:0] xy_o_p_sva;
  reg [15:0] OC2_koo_idx_sva;
  reg [15:0] co_c_idx_sva;
  reg [15:0] winx_wx_idx_sva;
  reg [31:0] xy_o_mul_1_cse;
  wire loopIndicesOut_rsci_idat_47_32_mx0c0;
  wire [31:0] xy_o_mul_1_cse_1;
  wire xy_o_and_cse;
  wire [16:0] z_out_32_16;

  wire[0:0] loopIndicesOut_not_1_nl;
  wire[33:0] acc_nl;
  wire[34:0] nl_acc_nl;
  wire[0:0] xy_o_xy_o_or_16_nl;
  wire[0:0] xy_o_xy_o_or_17_nl;
  wire[0:0] xy_o_xy_o_or_18_nl;
  wire[0:0] xy_o_xy_o_or_19_nl;
  wire[0:0] xy_o_xy_o_or_20_nl;
  wire[0:0] xy_o_xy_o_or_21_nl;
  wire[0:0] xy_o_xy_o_or_22_nl;
  wire[0:0] xy_o_xy_o_or_23_nl;
  wire[0:0] xy_o_xy_o_or_24_nl;
  wire[0:0] xy_o_xy_o_or_25_nl;
  wire[0:0] xy_o_xy_o_or_26_nl;
  wire[0:0] xy_o_xy_o_or_27_nl;
  wire[0:0] xy_o_xy_o_or_28_nl;
  wire[0:0] xy_o_xy_o_or_29_nl;
  wire[0:0] xy_o_xy_o_or_30_nl;
  wire[0:0] xy_o_xy_o_or_31_nl;
  wire[15:0] xy_o_mux1h_5_nl;
  wire[0:0] xy_o_or_3_nl;
  wire[0:0] xy_o_or_4_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_16_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_17_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_18_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_19_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_20_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_21_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_22_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_23_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_24_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_25_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_26_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_27_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_28_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_29_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_30_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_31_nl;
  wire[15:0] xy_o_mux1h_6_nl;
  wire[0:0] xy_o_or_5_nl;
  wire[15:0] winy_mux1h_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat;
  assign nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat
      = {loopIndicesOut_rsci_idat_47_32 , loopIndicesOut_rsci_idat_31_16 , loopIndicesOut_rsci_idat_15_0};
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_main_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_main_C_0_tr0 = ~ (z_out_32_16[16]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0 = ~ (z_out_32_16[16]);
  SystolicArrayLooper_run_paramsIn_rsci SystolicArrayLooper_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  SystolicArrayLooper_run_paramsOut_rsci SystolicArrayLooper_run_paramsOut_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_idat(paramsOut_rsci_idat)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci SystolicArrayLooper_run_loopIndicesOut_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_idat(nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat[47:0])
    );
  SystolicArrayLooper_run_staller SystolicArrayLooper_run_staller_inst (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp)
    );
  SystolicArrayLooper_run_run_fsm SystolicArrayLooper_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_main_C_0_tr0[0:0]),
      .xy_o_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0[0:0]),
      .OC2_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0[0:0]),
      .co_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0[0:0]),
      .winx_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0[0:0]),
      .winy_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0[0:0]),
      .winx_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0[0:0]),
      .co_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0[0:0]),
      .OC2_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0[0:0]),
      .xy_o_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0[0:0])
    );
  assign reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm = ((fsm_output[6:5]!=2'b00))
      & (z_out_32_16[0]);
  assign loopIndicesOut_and_cse = run_wen & reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
  assign xy_o_and_cse = run_wen & (~ and_dcpl_3);
  assign xy_o_mul_1_cse_1 = conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16]) * (paramsIn_rsci_idat_mxwt[15:0]));
  assign and_dcpl_3 = ~((fsm_output[1:0]!=2'b00));
  assign loopIndicesOut_rsci_idat_47_32_mx0c0 = (z_out_32_16[0]) & (fsm_output[5]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_15_0 <= 16'b0000000000000000;
      loopIndicesOut_rsci_idat_31_16 <= 16'b0000000000000000;
      paramsOut_rsci_idat <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( loopIndicesOut_and_cse ) begin
      loopIndicesOut_rsci_idat_15_0 <= co_c_idx_sva;
      loopIndicesOut_rsci_idat_31_16 <= winx_wx_idx_sva;
      paramsOut_rsci_idat <= paramsIn_crt_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( run_wen & (loopIndicesOut_rsci_idat_47_32_mx0c0 | ((z_out_32_16[0])
        & (fsm_output[6]))) ) begin
      loopIndicesOut_rsci_idat_47_32 <= MUX_v_16_2_2(16'b0000000000000000, z_out_1,
          (loopIndicesOut_not_1_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((and_dcpl_3 & (~ (fsm_output[10])))
          | (~((~ (z_out_32_16[16])) | (fsm_output[0]))));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      xy_o_mul_1_cse <= 32'b00000000000000000000000000000000;
      paramsIn_crt_sva <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( xy_o_and_cse ) begin
      xy_o_mul_1_cse <= xy_o_mul_1_cse_1;
      paramsIn_crt_sva <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      xy_o_p_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[10]) | (fsm_output[1])) ) begin
      xy_o_p_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[10]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      OC2_koo_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[9]) | (fsm_output[2])) ) begin
      OC2_koo_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[9]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      co_c_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[8]) | (fsm_output[3])) ) begin
      co_c_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[8]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      winx_wx_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[7]) | (fsm_output[4])) ) begin
      winx_wx_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[7]));
    end
  end
  assign loopIndicesOut_not_1_nl = ~ loopIndicesOut_rsci_idat_47_32_mx0c0;
  assign xy_o_xy_o_or_16_nl = (~((xy_o_mul_1_cse_1[31]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_17_nl = (~((xy_o_mul_1_cse_1[30]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_18_nl = (~((xy_o_mul_1_cse_1[29]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_19_nl = (~((xy_o_mul_1_cse_1[28]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_20_nl = (~((xy_o_mul_1_cse_1[27]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_21_nl = (~((xy_o_mul_1_cse_1[26]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_22_nl = (~((xy_o_mul_1_cse_1[25]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_23_nl = (~((xy_o_mul_1_cse_1[24]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_24_nl = (~((xy_o_mul_1_cse_1[23]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_25_nl = (~((xy_o_mul_1_cse_1[22]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_26_nl = (~((xy_o_mul_1_cse_1[21]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_27_nl = (~((xy_o_mul_1_cse_1[20]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_28_nl = (~((xy_o_mul_1_cse_1[19]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_29_nl = (~((xy_o_mul_1_cse_1[18]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_30_nl = (~((xy_o_mul_1_cse_1[17]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_xy_o_or_31_nl = (~((xy_o_mul_1_cse_1[16]) | (fsm_output[10]))) | (fsm_output[9:2]!=8'b00000000);
  assign xy_o_or_3_nl = (fsm_output[10:6]!=5'b00000);
  assign xy_o_mux1h_5_nl = MUX1HOT_v_16_6_2((~ (xy_o_mul_1_cse_1[15:0])), z_out_1,
      (~ (paramsIn_crt_sva[79:64])), (~ (paramsIn_crt_sva[95:80])), (~ (paramsIn_crt_sva[111:96])),
      (~ (paramsIn_crt_sva[127:112])), {(fsm_output[1]) , (xy_o_or_3_nl) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign xy_o_or_4_nl = (~((fsm_output[5:1]!=5'b00000))) | (fsm_output[10:6]!=5'b00000);
  assign xy_o_xy_o_xy_o_nor_16_nl = ~((xy_o_mul_1_cse[31]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_17_nl = ~((xy_o_mul_1_cse[30]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_18_nl = ~((xy_o_mul_1_cse[29]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_19_nl = ~((xy_o_mul_1_cse[28]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_20_nl = ~((xy_o_mul_1_cse[27]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_21_nl = ~((xy_o_mul_1_cse[26]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_22_nl = ~((xy_o_mul_1_cse[25]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_23_nl = ~((xy_o_mul_1_cse[24]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_24_nl = ~((xy_o_mul_1_cse[23]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_25_nl = ~((xy_o_mul_1_cse[22]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_26_nl = ~((xy_o_mul_1_cse[21]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_27_nl = ~((xy_o_mul_1_cse[20]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_28_nl = ~((xy_o_mul_1_cse[19]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_29_nl = ~((xy_o_mul_1_cse[18]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_30_nl = ~((xy_o_mul_1_cse[17]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_31_nl = ~((xy_o_mul_1_cse[16]) | (fsm_output[9:1]!=9'b000000000));
  assign xy_o_or_5_nl = (fsm_output[5:1]!=5'b00000);
  assign xy_o_mux1h_6_nl = MUX1HOT_v_16_6_2(16'b0000000000000001, (~ (xy_o_mul_1_cse[15:0])),
      (~ (paramsIn_crt_sva[79:64])), (~ (paramsIn_crt_sva[95:80])), (~ (paramsIn_crt_sva[111:96])),
      (~ (paramsIn_crt_sva[127:112])), {(xy_o_or_5_nl) , (fsm_output[10]) , (fsm_output[9])
      , (fsm_output[8]) , (fsm_output[7]) , (fsm_output[6])});
  assign nl_acc_nl = ({1'b1 , (xy_o_xy_o_or_16_nl) , (xy_o_xy_o_or_17_nl) , (xy_o_xy_o_or_18_nl)
      , (xy_o_xy_o_or_19_nl) , (xy_o_xy_o_or_20_nl) , (xy_o_xy_o_or_21_nl) , (xy_o_xy_o_or_22_nl)
      , (xy_o_xy_o_or_23_nl) , (xy_o_xy_o_or_24_nl) , (xy_o_xy_o_or_25_nl) , (xy_o_xy_o_or_26_nl)
      , (xy_o_xy_o_or_27_nl) , (xy_o_xy_o_or_28_nl) , (xy_o_xy_o_or_29_nl) , (xy_o_xy_o_or_30_nl)
      , (xy_o_xy_o_or_31_nl) , (xy_o_mux1h_5_nl) , (xy_o_or_4_nl)}) + conv_u2u_33_34({(xy_o_xy_o_xy_o_nor_16_nl)
      , (xy_o_xy_o_xy_o_nor_17_nl) , (xy_o_xy_o_xy_o_nor_18_nl) , (xy_o_xy_o_xy_o_nor_19_nl)
      , (xy_o_xy_o_xy_o_nor_20_nl) , (xy_o_xy_o_xy_o_nor_21_nl) , (xy_o_xy_o_xy_o_nor_22_nl)
      , (xy_o_xy_o_xy_o_nor_23_nl) , (xy_o_xy_o_xy_o_nor_24_nl) , (xy_o_xy_o_xy_o_nor_25_nl)
      , (xy_o_xy_o_xy_o_nor_26_nl) , (xy_o_xy_o_xy_o_nor_27_nl) , (xy_o_xy_o_xy_o_nor_28_nl)
      , (xy_o_xy_o_xy_o_nor_29_nl) , (xy_o_xy_o_xy_o_nor_30_nl) , (xy_o_xy_o_xy_o_nor_31_nl)
      , (xy_o_mux1h_6_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[33:0];
  assign z_out_32_16 = readslicef_34_17_17((acc_nl));
  assign winy_mux1h_1_nl = MUX1HOT_v_16_5_2(loopIndicesOut_rsci_idat_47_32, xy_o_p_sva,
      OC2_koo_idx_sva, co_c_idx_sva, winx_wx_idx_sva, {(fsm_output[6]) , (fsm_output[10])
      , (fsm_output[9]) , (fsm_output[8]) , (fsm_output[7])});
  assign nl_z_out_1 = (winy_mux1h_1_nl) + 16'b0000000000000001;
  assign z_out_1 = nl_z_out_1[15:0];

  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [16:0] readslicef_34_17_17;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 17;
    readslicef_34_17_17 = tmp[16:0];
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer
// ------------------------------------------------------------------


module ParamsDeserializer (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy, outputChannel2_rsc_dat,
      outputChannel2_rsc_vld, outputChannel2_rsc_rdy, outputChannel3_rsc_dat, outputChannel3_rsc_vld,
      outputChannel3_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ParamsDeserializer_run ParamsDeserializer_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16 (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld),
      .serialOutChannel_rsc_rdy(serialOutChannel_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper
// ------------------------------------------------------------------


module SystolicArrayLooper (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat,
      paramsOut_rsc_vld, paramsOut_rsc_rdy, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld,
      loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  SystolicArrayLooper_run SystolicArrayLooper_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16
// ------------------------------------------------------------------


module SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16 (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [255:0] output_rsc_dat_nsystolicArrayCore;
  wire [143:0] paramsIn_rsc_dat_nsystolicArrayCore;
  wire paramsIn_rsc_vld_nsystolicArrayCore;
  wire [47:0] loopIndicesIn_rsc_dat_nsystolicArrayCore;
  wire loopIndicesIn_rsc_vld_nsystolicArrayCore;
  wire [143:0] paramsOut_rsc_dat_nsystolicArrayLooper;
  wire paramsOut_rsc_rdy_nsystolicArrayLooper;
  wire [47:0] loopIndicesOut_rsc_dat_nsystolicArrayLooper;
  wire loopIndicesOut_rsc_rdy_nsystolicArrayLooper;
  wire input_rsc_rdy_nsystolicArrayCore_bud;
  wire weight_rsc_rdy_nsystolicArrayCore_bud;
  wire output_rsc_vld_nsystolicArrayCore_bud;
  wire paramsIn_rsc_rdy_nsystolicArrayCore_bud;
  wire paramsOut_rsc_vld_nsystolicArrayLooper_bud;
  wire loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud;
  wire loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud;
  wire paramsIn_rsc_rdy_nsystolicArrayLooper_bud;
  wire paramsChannel_unc_2;
  wire paramsChannel_idle;
  wire loopIndicesChannel_unc_2;
  wire loopIndicesChannel_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd163),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) paramsChannel_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(paramsOut_rsc_rdy_nsystolicArrayLooper),
      .din_vld(paramsOut_rsc_vld_nsystolicArrayLooper_bud),
      .din(paramsOut_rsc_dat_nsystolicArrayLooper),
      .dout_rdy(paramsIn_rsc_rdy_nsystolicArrayCore_bud),
      .dout_vld(paramsIn_rsc_vld_nsystolicArrayCore),
      .dout(paramsIn_rsc_dat_nsystolicArrayCore),
      .sz(paramsChannel_unc_2),
      .sz_req(1'b0),
      .is_idle(paramsChannel_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd164),
  .width(32'sd48),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) loopIndicesChannel_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(loopIndicesOut_rsc_rdy_nsystolicArrayLooper),
      .din_vld(loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud),
      .din(loopIndicesOut_rsc_dat_nsystolicArrayLooper),
      .dout_rdy(loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud),
      .dout_vld(loopIndicesIn_rsc_vld_nsystolicArrayCore),
      .dout(loopIndicesIn_rsc_dat_nsystolicArrayCore),
      .sz(loopIndicesChannel_unc_2),
      .sz_req(1'b0),
      .is_idle(loopIndicesChannel_idle)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16 systolicArrayCore (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy_nsystolicArrayCore_bud),
      .weight_rsc_dat(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy_nsystolicArrayCore_bud),
      .output_rsc_dat(output_rsc_dat_nsystolicArrayCore),
      .output_rsc_vld(output_rsc_vld_nsystolicArrayCore_bud),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nsystolicArrayCore),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nsystolicArrayCore),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArrayCore_bud),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat_nsystolicArrayCore),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld_nsystolicArrayCore),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud)
    );
  SystolicArrayLooper systolicArrayLooper_1 (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArrayLooper_bud),
      .paramsOut_rsc_dat(paramsOut_rsc_dat_nsystolicArrayLooper),
      .paramsOut_rsc_vld(paramsOut_rsc_vld_nsystolicArrayLooper_bud),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy_nsystolicArrayLooper),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat_nsystolicArrayLooper),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy_nsystolicArrayLooper)
    );
  assign input_rsc_rdy = input_rsc_rdy_nsystolicArrayCore_bud;
  assign weight_rsc_rdy = weight_rsc_rdy_nsystolicArrayCore_bud;
  assign output_rsc_vld = output_rsc_vld_nsystolicArrayCore_bud;
  assign output_rsc_dat = output_rsc_dat_nsystolicArrayCore;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nsystolicArrayLooper_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Conv
// ------------------------------------------------------------------


module Conv (
  clk, arst_n, input_serial_rsc_dat, input_serial_rsc_vld, input_serial_rsc_rdy,
      weight_serial_rsc_dat, weight_serial_rsc_vld, weight_serial_rsc_rdy, output_serial_rsc_dat,
      output_serial_rsc_vld, output_serial_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] input_serial_rsc_dat;
  input input_serial_rsc_vld;
  output input_serial_rsc_rdy;
  input [15:0] weight_serial_rsc_dat;
  input weight_serial_rsc_vld;
  output weight_serial_rsc_rdy;
  output [15:0] output_serial_rsc_dat;
  output output_serial_rsc_vld;
  input output_serial_rsc_rdy;
  input [15:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] outputChannel1_rsc_dat_nparamsDeserializer;
  wire outputChannel1_rsc_rdy_nparamsDeserializer;
  wire [143:0] outputChannel2_rsc_dat_nparamsDeserializer;
  wire outputChannel2_rsc_rdy_nparamsDeserializer;
  wire [143:0] outputChannel3_rsc_dat_nparamsDeserializer;
  wire outputChannel3_rsc_rdy_nparamsDeserializer;
  wire [255:0] inputChannel_rsc_dat_noutputSerializer;
  wire inputChannel_rsc_vld_noutputSerializer;
  wire [15:0] serialOutChannel_rsc_dat_noutputSerializer;
  wire [127:0] inputs_out_rsc_dat_ninputDoubleBuffer;
  wire inputs_out_rsc_rdy_ninputDoubleBuffer;
  wire [143:0] paramsIn_rsc_dat_ninputDoubleBuffer;
  wire paramsIn_rsc_vld_ninputDoubleBuffer;
  wire [127:0] weights_out_rsc_dat_nweightDoubleBuffer;
  wire weights_out_rsc_rdy_nweightDoubleBuffer;
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBuffer;
  wire paramsIn_rsc_vld_nweightDoubleBuffer;
  wire [127:0] input_rsc_dat_nsystolicArray;
  wire input_rsc_vld_nsystolicArray;
  wire [127:0] weight_rsc_dat_nsystolicArray;
  wire weight_rsc_vld_nsystolicArray;
  wire [255:0] output_rsc_dat_nsystolicArray;
  wire output_rsc_rdy_nsystolicArray;
  wire [143:0] paramsIn_rsc_dat_nsystolicArray;
  wire paramsIn_rsc_vld_nsystolicArray;
  wire inputChannel_rsc_rdy_nparamsDeserializer_bud;
  wire outputChannel1_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_ninputDoubleBuffer_bud;
  wire outputChannel2_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_nweightDoubleBuffer_bud;
  wire outputChannel3_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_nsystolicArray_bud;
  wire inputChannel_rsc_rdy_noutputSerializer_bud;
  wire output_rsc_vld_nsystolicArray_bud;
  wire serialOutChannel_rsc_vld_noutputSerializer_bud;
  wire inputs_in_rsc_rdy_ninputDoubleBuffer_bud;
  wire inputs_out_rsc_vld_ninputDoubleBuffer_bud;
  wire input_rsc_rdy_nsystolicArray_bud;
  wire weights_in_rsc_rdy_nweightDoubleBuffer_bud;
  wire weights_out_rsc_vld_nweightDoubleBuffer_bud;
  wire weight_rsc_rdy_nsystolicArray_bud;
  wire inputDoubleBufferParams_unc_2;
  wire inputDoubleBufferParams_idle;
  wire weightDoubleBufferParams_unc_2;
  wire weightDoubleBufferParams_idle;
  wire systolicArrayParams_unc_2;
  wire systolicArrayParams_idle;
  wire output_unc_2;
  wire output_idle;
  wire input_out_unc_2;
  wire input_out_idle;
  wire weight_out_unc_2;
  wire weight_out_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd169),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) inputDoubleBufferParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel1_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel1_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel1_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_ninputDoubleBuffer_bud),
      .dout_vld(paramsIn_rsc_vld_ninputDoubleBuffer),
      .dout(paramsIn_rsc_dat_ninputDoubleBuffer),
      .sz(inputDoubleBufferParams_unc_2),
      .sz_req(1'b0),
      .is_idle(inputDoubleBufferParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd170),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel2_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel2_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel2_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBuffer_bud),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBuffer),
      .dout(paramsIn_rsc_dat_nweightDoubleBuffer),
      .sz(weightDoubleBufferParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd174),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) systolicArrayParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel3_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel3_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel3_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_nsystolicArray_bud),
      .dout_vld(paramsIn_rsc_vld_nsystolicArray),
      .dout(paramsIn_rsc_dat_nsystolicArray),
      .sz(systolicArrayParams_unc_2),
      .sz_req(1'b0),
      .is_idle(systolicArrayParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd173),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) output_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(output_rsc_rdy_nsystolicArray),
      .din_vld(output_rsc_vld_nsystolicArray_bud),
      .din(output_rsc_dat_nsystolicArray),
      .dout_rdy(inputChannel_rsc_rdy_noutputSerializer_bud),
      .dout_vld(inputChannel_rsc_vld_noutputSerializer),
      .dout(inputChannel_rsc_dat_noutputSerializer),
      .sz(output_unc_2),
      .sz_req(1'b0),
      .is_idle(output_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd171),
  .width(32'sd128),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) input_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(inputs_out_rsc_rdy_ninputDoubleBuffer),
      .din_vld(inputs_out_rsc_vld_ninputDoubleBuffer_bud),
      .din(inputs_out_rsc_dat_ninputDoubleBuffer),
      .dout_rdy(input_rsc_rdy_nsystolicArray_bud),
      .dout_vld(input_rsc_vld_nsystolicArray),
      .dout(input_rsc_dat_nsystolicArray),
      .sz(input_out_unc_2),
      .sz_req(1'b0),
      .is_idle(input_out_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd172),
  .width(32'sd128),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weight_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weights_out_rsc_rdy_nweightDoubleBuffer),
      .din_vld(weights_out_rsc_vld_nweightDoubleBuffer_bud),
      .din(weights_out_rsc_dat_nweightDoubleBuffer),
      .dout_rdy(weight_rsc_rdy_nsystolicArray_bud),
      .dout_vld(weight_rsc_vld_nsystolicArray),
      .dout(weight_rsc_dat_nsystolicArray),
      .sz(weight_out_unc_2),
      .sz_req(1'b0),
      .is_idle(weight_out_idle)
    );
  ParamsDeserializer paramsDeserializer_1 (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(paramsIn_rsc_dat),
      .inputChannel_rsc_vld(paramsIn_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy_nparamsDeserializer_bud),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat_nparamsDeserializer),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld_nparamsDeserializer_bud),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy_nparamsDeserializer),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat_nparamsDeserializer),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld_nparamsDeserializer_bud),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy_nparamsDeserializer),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat_nparamsDeserializer),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld_nparamsDeserializer_bud),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy_nparamsDeserializer)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16 outputSerializer (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat_noutputSerializer),
      .inputChannel_rsc_vld(inputChannel_rsc_vld_noutputSerializer),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy_noutputSerializer_bud),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat_noutputSerializer),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld_noutputSerializer_bud),
      .serialOutChannel_rsc_rdy(output_serial_rsc_rdy)
    );
  InputDoubleBuffer_512_16_16 inputDoubleBuffer (
      .clk(clk),
      .arst_n(arst_n),
      .inputs_in_rsc_dat(input_serial_rsc_dat),
      .inputs_in_rsc_vld(input_serial_rsc_vld),
      .inputs_in_rsc_rdy(inputs_in_rsc_rdy_ninputDoubleBuffer_bud),
      .inputs_out_rsc_dat(inputs_out_rsc_dat_ninputDoubleBuffer),
      .inputs_out_rsc_vld(inputs_out_rsc_vld_ninputDoubleBuffer_bud),
      .inputs_out_rsc_rdy(inputs_out_rsc_rdy_ninputDoubleBuffer),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_ninputDoubleBuffer),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_ninputDoubleBuffer),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBuffer_bud)
    );
  WeightDoubleBuffer_384_16_16 weightDoubleBuffer (
      .clk(clk),
      .arst_n(arst_n),
      .weights_in_rsc_dat(weight_serial_rsc_dat),
      .weights_in_rsc_vld(weight_serial_rsc_vld),
      .weights_in_rsc_rdy(weights_in_rsc_rdy_nweightDoubleBuffer_bud),
      .weights_out_rsc_dat(weights_out_rsc_dat_nweightDoubleBuffer),
      .weights_out_rsc_vld(weights_out_rsc_vld_nweightDoubleBuffer_bud),
      .weights_out_rsc_rdy(weights_out_rsc_rdy_nweightDoubleBuffer),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBuffer),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBuffer),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBuffer_bud)
    );
  SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16 systolicArray (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat_nsystolicArray),
      .input_rsc_vld(input_rsc_vld_nsystolicArray),
      .input_rsc_rdy(input_rsc_rdy_nsystolicArray_bud),
      .weight_rsc_dat(weight_rsc_dat_nsystolicArray),
      .weight_rsc_vld(weight_rsc_vld_nsystolicArray),
      .weight_rsc_rdy(weight_rsc_rdy_nsystolicArray_bud),
      .output_rsc_dat(output_rsc_dat_nsystolicArray),
      .output_rsc_vld(output_rsc_vld_nsystolicArray_bud),
      .output_rsc_rdy(output_rsc_rdy_nsystolicArray),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nsystolicArray),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nsystolicArray),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArray_bud)
    );
  assign paramsIn_rsc_rdy = inputChannel_rsc_rdy_nparamsDeserializer_bud;
  assign output_serial_rsc_vld = serialOutChannel_rsc_vld_noutputSerializer_bud;
  assign output_serial_rsc_dat = serialOutChannel_rsc_dat_noutputSerializer;
  assign input_serial_rsc_rdy = inputs_in_rsc_rdy_ninputDoubleBuffer_bud;
  assign weight_serial_rsc_rdy = weights_in_rsc_rdy_nweightDoubleBuffer_bud;
endmodule



