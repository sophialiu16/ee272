
//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/Fifo_ODTYPE_16__221b3917049bbc5c28349b3242b352d67c53_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:07:21 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_16_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_16_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;
  reg [15:0] regs_13_sva_dfm;
  reg [15:0] regs_14_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd97),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd98),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd117),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_14_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_14_sva_dfm <= 16'b0000000000000000;
      regs_13_sva_dfm <= 16'b0000000000000000;
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_14_sva_dfm <= regs_13_sva_dfm;
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_16
// ------------------------------------------------------------------


module Fifo_ODTYPE_16 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_16_run Fifo_ODTYPE_16_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_15__0588a2793143081c26ab62d19350374879f4_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:07:29 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_15_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_15_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;
  reg [15:0] regs_13_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd94),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd95),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd118),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_13_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_13_sva_dfm <= 16'b0000000000000000;
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_15
// ------------------------------------------------------------------


module Fifo_ODTYPE_15 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_15_run Fifo_ODTYPE_15_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_14__45e500b517c70224a67c6e90729192d87795_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:07:37 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_14_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_14_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;
  reg [15:0] regs_12_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd91),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd92),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd119),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_12_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_12_sva_dfm <= 16'b0000000000000000;
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_14
// ------------------------------------------------------------------


module Fifo_ODTYPE_14 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_14_run Fifo_ODTYPE_14_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_13__cfc4e6d714c299c88f1ea11a4aa19dcd7536_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:07:45 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_13_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_13_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;
  reg [15:0] regs_11_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd88),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd89),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd120),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_11_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_11_sva_dfm <= 16'b0000000000000000;
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_13
// ------------------------------------------------------------------


module Fifo_ODTYPE_13 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_13_run Fifo_ODTYPE_13_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_12__20588fe682fdeb9113d6793626c8c22872d7_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:07:53 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_12_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_12_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;
  reg [15:0] regs_10_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd85),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd86),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd121),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_10_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_10_sva_dfm <= 16'b0000000000000000;
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_12
// ------------------------------------------------------------------


module Fifo_ODTYPE_12 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_12_run Fifo_ODTYPE_12_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_11__917724a8fd2b9046ed510e9c8c2f6e0c7078_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:01 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_11_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_11_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;
  reg [15:0] regs_9_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd82),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd83),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd122),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_9_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_9_sva_dfm <= 16'b0000000000000000;
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_11
// ------------------------------------------------------------------


module Fifo_ODTYPE_11 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_11_run Fifo_ODTYPE_11_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_10__98cb450ab203be4fbf6a1bbccd8ea7be6e1a_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:10 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_10_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_10_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;
  reg [15:0] regs_8_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd79),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd80),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd123),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_8_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_8_sva_dfm <= 16'b0000000000000000;
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_10
// ------------------------------------------------------------------


module Fifo_ODTYPE_10 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_10_run Fifo_ODTYPE_10_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_9__59d17ff0eccb20043113c483bd4832ad6bb0_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:18 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_9_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_9_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;
  reg [15:0] regs_7_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd76),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd77),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd124),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_7_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_7_sva_dfm <= 16'b0000000000000000;
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_9
// ------------------------------------------------------------------


module Fifo_ODTYPE_9 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_9_run Fifo_ODTYPE_9_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_8__fe12db0fc7a2f935da96abaa8a4058ea6952_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:26 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_8_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_8_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;
  reg [15:0] regs_6_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd73),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd74),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd125),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_6_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_6_sva_dfm <= 16'b0000000000000000;
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_8
// ------------------------------------------------------------------


module Fifo_ODTYPE_8 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_8_run Fifo_ODTYPE_8_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_7__d003a84803bb8a29bae7687df0b778f666f4_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:34 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_7_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_7_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;
  reg [15:0] regs_5_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd70),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd71),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd126),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_5_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_5_sva_dfm <= 16'b0000000000000000;
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_7
// ------------------------------------------------------------------


module Fifo_ODTYPE_7 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_7_run Fifo_ODTYPE_7_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_6__ef9cbbb510dc9b7e23fbd9ad2a0b75166496_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:42 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_6_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_6_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;
  reg [15:0] regs_4_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd67),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd68),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd127),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_4_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_4_sva_dfm <= 16'b0000000000000000;
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_6
// ------------------------------------------------------------------


module Fifo_ODTYPE_6 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_6_run Fifo_ODTYPE_6_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_5__3e4e6554e1972e837dfae32d6649bb6d6238_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:51 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_5_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_5_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;
  reg [15:0] regs_3_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd64),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd65),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd128),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_3_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_3_sva_dfm <= 16'b0000000000000000;
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_5
// ------------------------------------------------------------------


module Fifo_ODTYPE_5 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_5_run Fifo_ODTYPE_5_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_4__156db601d575e3447c254544adc35f885fda_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:08:59 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_4_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_4_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;
  reg [15:0] regs_2_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd61),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd62),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd129),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_2_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_2_sva_dfm <= 16'b0000000000000000;
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_4
// ------------------------------------------------------------------


module Fifo_ODTYPE_4 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_4_run Fifo_ODTYPE_4_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_3__7b12ca58716272e54ee61060556848705d7c_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:07 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_3_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_3_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [15:0] regs_0_sva;
  reg [15:0] regs_1_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd58),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd59),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd130),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_1_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_1_sva_dfm <= 16'b0000000000000000;
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( regs_and_cse ) begin
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_3
// ------------------------------------------------------------------


module Fifo_ODTYPE_3 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_3_run Fifo_ODTYPE_3_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_2__d9255459d1985bba09ce948bd73b39735b1e_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:15 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_2_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_2_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [15:0] regs_0_sva;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd55),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd56),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd131),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_0_sva;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_0_sva <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_2
// ------------------------------------------------------------------


module Fifo_ODTYPE_2 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_2_run Fifo_ODTYPE_2_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_16__d38d5c3f7f7d770ed3944fd5fef6db0b7c26_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:32 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_16_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_16_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;
  reg [7:0] regs_13_sva_dfm;
  reg [7:0] regs_14_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd50),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd51),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd133),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_14_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_14_sva_dfm <= 8'b00000000;
      regs_13_sva_dfm <= 8'b00000000;
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_14_sva_dfm <= regs_13_sva_dfm;
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_16
// ------------------------------------------------------------------


module Fifo_IDTYPE_16 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_16_run Fifo_IDTYPE_16_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_15__a3693e6df94c682291b73c0533bd535379c8_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:41 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_15_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_15_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;
  reg [7:0] regs_13_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd47),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd48),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd134),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_13_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_13_sva_dfm <= 8'b00000000;
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_13_sva_dfm <= regs_12_sva_dfm;
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_15
// ------------------------------------------------------------------


module Fifo_IDTYPE_15 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_15_run Fifo_IDTYPE_15_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_14__6ed558445f9b0ba26813510e683ff2e6776a_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:49 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_14_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_14_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;
  reg [7:0] regs_12_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd45),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd135),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_12_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_12_sva_dfm <= 8'b00000000;
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_12_sva_dfm <= regs_11_sva_dfm;
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_14
// ------------------------------------------------------------------


module Fifo_IDTYPE_14 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_14_run Fifo_IDTYPE_14_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_13__3ab39e6656c571656f9f918808a98c90750c_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:58 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_13_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_13_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;
  reg [7:0] regs_11_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd41),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd42),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd136),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_11_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_11_sva_dfm <= 8'b00000000;
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_11_sva_dfm <= regs_10_sva_dfm;
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_13
// ------------------------------------------------------------------


module Fifo_IDTYPE_13 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_13_run Fifo_IDTYPE_13_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_12__41334737f9db89f3401ddbdb180284a372ae_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:07 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_12_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_12_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;
  reg [7:0] regs_10_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd38),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd39),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd137),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_10_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_10_sva_dfm <= 8'b00000000;
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_10_sva_dfm <= regs_9_sva_dfm;
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_12
// ------------------------------------------------------------------


module Fifo_IDTYPE_12 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_12_run Fifo_IDTYPE_12_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_11__b143065b8a794d7c3150cb2396006f267050_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:16 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_11_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_11_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;
  reg [7:0] regs_9_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd35),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd36),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd138),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_9_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_9_sva_dfm <= 8'b00000000;
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_9_sva_dfm <= regs_8_sva_dfm;
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_11
// ------------------------------------------------------------------


module Fifo_IDTYPE_11 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_11_run Fifo_IDTYPE_11_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_10__2ffa16ce99a732e8d71a5f721f0f2d316df3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:25 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_10_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_10_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;
  reg [7:0] regs_8_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd32),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd33),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd139),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_8_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_8_sva_dfm <= 8'b00000000;
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_8_sva_dfm <= regs_7_sva_dfm;
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_10
// ------------------------------------------------------------------


module Fifo_IDTYPE_10 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_10_run Fifo_IDTYPE_10_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_9__3850d4c5a858cb636c57c5c7832e8f086b8a_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:33 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_9_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_9_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;
  reg [7:0] regs_7_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd29),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd30),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd140),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_7_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_7_sva_dfm <= 8'b00000000;
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_7_sva_dfm <= regs_6_sva_dfm;
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_9
// ------------------------------------------------------------------


module Fifo_IDTYPE_9 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_9_run Fifo_IDTYPE_9_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_8__088804bffe2cbc7474b0591ee11c8c42692d_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:42 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_8_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_8_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;
  reg [7:0] regs_6_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd26),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd27),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd141),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_6_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_6_sva_dfm <= 8'b00000000;
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_6_sva_dfm <= regs_5_sva_dfm;
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_8
// ------------------------------------------------------------------


module Fifo_IDTYPE_8 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_8_run Fifo_IDTYPE_8_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_7__219aaa96b5533f6efa14178ba0ae3f9266d0_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:51 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_7_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_7_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;
  reg [7:0] regs_5_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd23),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd24),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd142),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_5_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_5_sva_dfm <= 8'b00000000;
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_5_sva_dfm <= regs_4_sva_dfm;
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_7
// ------------------------------------------------------------------


module Fifo_IDTYPE_7 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_7_run Fifo_IDTYPE_7_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_6__4caa842e06e3cce2ef6eb0925cfd318a6473_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:10:59 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_6_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_6_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;
  reg [7:0] regs_4_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd20),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd21),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd143),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_4_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_4_sva_dfm <= 8'b00000000;
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_4_sva_dfm <= regs_3_sva_dfm;
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_6
// ------------------------------------------------------------------


module Fifo_IDTYPE_6 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_6_run Fifo_IDTYPE_6_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_5__74b9abe40f59f3bac195e723964a8a776216_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:11:08 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_5_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_5_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;
  reg [7:0] regs_3_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd17),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd18),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd144),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_3_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_3_sva_dfm <= 8'b00000000;
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_3_sva_dfm <= regs_2_sva_dfm;
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_5
// ------------------------------------------------------------------


module Fifo_IDTYPE_5 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_5_run Fifo_IDTYPE_5_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_4__99dd0c69a5e527ded4c3d01075afb99b5fb9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:11:17 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_4_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_4_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;
  reg [7:0] regs_2_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd14),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd15),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd145),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_2_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_2_sva_dfm <= 8'b00000000;
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_2_sva_dfm <= regs_1_sva_dfm;
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_4
// ------------------------------------------------------------------


module Fifo_IDTYPE_4 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_4_run Fifo_IDTYPE_4_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_3__9ab5ce9495ab244439c9135630c9d9035d5c_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:11:25 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_3_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_3_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  wire regs_and_cse;
  reg [7:0] regs_0_sva;
  reg [7:0] regs_1_sva_dfm;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd12),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd146),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign regs_and_cse = ccs_ccore_en & ccs_ccore_start_rsci_idat;
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_1_sva_dfm;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_1_sva_dfm <= 8'b00000000;
      regs_0_sva <= 8'b00000000;
    end
    else if ( regs_and_cse ) begin
      regs_1_sva_dfm <= regs_0_sva;
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_3
// ------------------------------------------------------------------


module Fifo_IDTYPE_3 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_3_run Fifo_IDTYPE_3_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_2__e3a3a79fd6d2b9552fe00c731f1f97345afd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:11:34 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_2_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_2_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [7:0] regs_0_sva;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd147),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= regs_0_sva;
    end
  end
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      regs_0_sva <= 8'b00000000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      regs_0_sva <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_2
// ------------------------------------------------------------------


module Fifo_IDTYPE_2 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_2_run Fifo_IDTYPE_2_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../ProcessingElementless_IDTYPEcomma_ODTYPEgreater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:05:20 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ProcessingElement_IDTYPE_ODTYPE_run
// ------------------------------------------------------------------


module ProcessingElement_IDTYPE_ODTYPE_run (
  clk, arst_n, input_in_rsc_dat, psum_in_rsc_dat, weight_rsc_dat, input_out_rsc_z,
      psum_out_rsc_z, ccs_ccore_en
);
  input clk;
  input arst_n;
  input [7:0] input_in_rsc_dat;
  input [15:0] psum_in_rsc_dat;
  input [7:0] weight_rsc_dat;
  output [7:0] input_out_rsc_z;
  output [15:0] psum_out_rsc_z;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_in_rsci_idat;
  wire [15:0] psum_in_rsci_idat;
  wire [7:0] weight_rsci_idat;
  reg [7:0] input_out_rsci_d;
  reg [15:0] psum_out_rsci_d;
  wire [16:0] nl_psum_out_rsci_d;

  wire[15:0] mul_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd8)) input_in_rsci (
      .dat(input_in_rsc_dat),
      .idat(input_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd16)) psum_in_rsci (
      .dat(psum_in_rsc_dat),
      .idat(psum_in_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd8)) weight_rsci (
      .dat(weight_rsc_dat),
      .idat(weight_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd8)) input_out_rsci (
      .d(input_out_rsci_d),
      .z(input_out_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd5),
  .width(32'sd16)) psum_out_rsci (
      .d(psum_out_rsci_d),
      .z(psum_out_rsc_z)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_out_rsci_d <= 8'b00000000;
      psum_out_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      input_out_rsci_d <= input_in_rsci_idat;
      psum_out_rsci_d <= nl_psum_out_rsci_d[15:0];
    end
  end
  assign mul_nl = conv_s2u_16_16($signed((input_in_rsci_idat)) * $signed((weight_rsci_idat)));
  assign nl_psum_out_rsci_d  = (mul_nl) + psum_in_rsci_idat;

  function automatic [15:0] conv_s2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_16 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ProcessingElement_IDTYPE_ODTYPE
// ------------------------------------------------------------------


module ProcessingElement_IDTYPE_ODTYPE (
  clk, arst_n, input_in_rsc_dat, psum_in_rsc_dat, weight_rsc_dat, input_out_rsc_z,
      psum_out_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_en
);
  input clk;
  input arst_n;
  input [7:0] input_in_rsc_dat;
  input [15:0] psum_in_rsc_dat;
  input [7:0] weight_rsc_dat;
  output [7:0] input_out_rsc_z;
  output [15:0] psum_out_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  ProcessingElement_IDTYPE_ODTYPE_run ProcessingElement_IDTYPE_ODTYPE_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .input_in_rsc_dat(input_in_rsc_dat),
      .psum_in_rsc_dat(psum_in_rsc_dat),
      .weight_rsc_dat(weight_rsc_dat),
      .input_out_rsc_z(input_out_rsc_z),
      .psum_out_rsc_z(psum_out_rsc_z),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_ODTYPE_1__9c4a99f532013522e5120280b322b342544e_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:09:23 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_1_run
// ------------------------------------------------------------------


module Fifo_ODTYPE_1_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_clk, ccs_ccore_arst, ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [15:0] input_rsci_idat;
  reg [15:0] output_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd53),
  .width(32'sd16)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd54),
  .width(32'sd16)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 16'b0000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_ODTYPE_1
// ------------------------------------------------------------------


module Fifo_ODTYPE_1 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [15:0] input_rsc_dat;
  output [15:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_ODTYPE_1_run Fifo_ODTYPE_1_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/Fifo_IDTYPE_1__93d204e0bede44f1c5761a5d5c8023bb542f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:11:42 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_1_run
// ------------------------------------------------------------------


module Fifo_IDTYPE_1_run (
  input_rsc_dat, output_rsc_z, ccs_ccore_clk, ccs_ccore_arst, ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [7:0] input_rsci_idat;
  reg [7:0] output_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd8)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd8)) output_rsci (
      .d(output_rsci_d),
      .z(output_rsc_z)
    );
  always @(posedge ccs_ccore_clk or negedge ccs_ccore_arst) begin
    if ( ~ ccs_ccore_arst ) begin
      output_rsci_d <= 8'b00000000;
    end
    else if ( ccs_ccore_en ) begin
      output_rsci_d <= input_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Fifo_IDTYPE_1
// ------------------------------------------------------------------


module Fifo_IDTYPE_1 (
  input_rsc_dat, output_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_arst,
      ccs_ccore_en
);
  input [7:0] input_rsc_dat;
  output [7:0] output_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_arst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  Fifo_IDTYPE_1_run Fifo_IDTYPE_1_run_inst (
      .input_rsc_dat(input_rsc_dat),
      .output_rsc_z(output_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_arst(ccs_ccore_arst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_ram_sync_1R1W.v 
module ccs_ram_sync_1R1W
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

   // synopsys translate_off
	reg [data_width-1:0] q;

	reg [data_width-1:0] mem [depth-1:0];
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end
   // synopsys translate_on

endmodule

//------> ../SystolicArrayCoreless_IDTYPEcomma_WDTYPEcomma_ODTYPEcomma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:17:20 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_164_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_164_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_163_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_163_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_162_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_162_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_161_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_161_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_160_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_160_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_159_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_159_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_158_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_158_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_157_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_157_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_156_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_156_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_155_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_155_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_154_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_154_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_153_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_153_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_152_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_152_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_151_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_151_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_150_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_150_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_149_16_8_256_256_16_5_gen
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_149_16_8_256_256_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [7:0] wadr;
  input [15:0] q;
  output re;
  output [7:0] radr;
  input [7:0] radr_d;
  input [7:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, input_rsci_wen_comp, weight_rsci_wen_comp, output_rsci_wen_comp,
      paramsIn_rsci_wen_comp, loopIndicesIn_rsci_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input input_rsci_wen_comp;
  input weight_rsci_wen_comp;
  input output_rsci_wen_comp;
  input paramsIn_rsci_wen_comp;
  input loopIndicesIn_rsci_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = input_rsci_wen_comp & weight_rsci_wen_comp & output_rsci_wen_comp
      & paramsIn_rsci_wen_comp & loopIndicesIn_rsci_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp (
  ensig_cgo_iro, ensig_cgo_iro_1, run_wen, ensig_cgo, accum_fifo_15_rsci_ccs_ccore_en,
      ensig_cgo_1, output_fifo_0_rsci_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo_iro_1;
  input run_wen;
  input ensig_cgo;
  output accum_fifo_15_rsci_ccs_ccore_en;
  input ensig_cgo_1;
  output output_fifo_0_rsci_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign accum_fifo_15_rsci_ccs_ccore_en = run_wen & (ensig_cgo | ensig_cgo_iro);
  assign output_fifo_0_rsci_ccs_ccore_en = run_wen & (ensig_cgo_1 | ensig_cgo_iro_1);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    CGHpart
// ------------------------------------------------------------------


module CGHpart (
  CGHpart_isig
);
  input CGHpart_isig;



  // Interconnect Declarations for Component Instantiations 
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_15_i_radr_d, accumulation_buffer_rsc_0_15_i_wadr_d,
      accumulation_buffer_rsc_0_15_i_q_d, accumulation_buffer_rsc_0_15_i_radr_d_run,
      accumulation_buffer_rsc_0_15_i_wadr_d_run, accumulation_buffer_rsc_0_15_i_q_d_mxwt,
      accumulation_buffer_rsc_0_15_i_biwt, accumulation_buffer_rsc_0_15_i_bdwt, accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_15_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_15_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_15_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_15_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_15_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_15_i_biwt;
  input accumulation_buffer_rsc_0_15_i_bdwt;
  input accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_15_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_15_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_15_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_15_i_q_d,
      accumulation_buffer_rsc_0_15_i_q_d_bfwt, accumulation_buffer_rsc_0_15_i_bcwt);
  assign accumulation_buffer_rsc_0_15_i_radr_d = {(~ accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_15_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_15_i_wadr_d = {(~ accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_15_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_15_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_15_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_15_i_bcwt <= ~((~(accumulation_buffer_rsc_0_15_i_bcwt
          | accumulation_buffer_rsc_0_15_i_biwt)) | accumulation_buffer_rsc_0_15_i_bdwt);
      accumulation_buffer_rsc_0_15_i_q_d_bfwt <= accumulation_buffer_rsc_0_15_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_15_i_oswt, accumulation_buffer_rsc_0_15_i_biwt,
      accumulation_buffer_rsc_0_15_i_bdwt, accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_15_i_oswt_pff, accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_15_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_15_i_oswt;
  output accumulation_buffer_rsc_0_15_i_biwt;
  output accumulation_buffer_rsc_0_15_i_bdwt;
  output accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_15_i_oswt_pff;
  output accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_15_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_15_i_bdwt = accumulation_buffer_rsc_0_15_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_15_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_15_i_oswt;
  assign accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_15_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_15_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_14_i_radr_d, accumulation_buffer_rsc_0_14_i_wadr_d,
      accumulation_buffer_rsc_0_14_i_q_d, accumulation_buffer_rsc_0_14_i_radr_d_run,
      accumulation_buffer_rsc_0_14_i_wadr_d_run, accumulation_buffer_rsc_0_14_i_q_d_mxwt,
      accumulation_buffer_rsc_0_14_i_biwt, accumulation_buffer_rsc_0_14_i_bdwt, accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_14_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_14_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_14_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_14_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_14_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_14_i_biwt;
  input accumulation_buffer_rsc_0_14_i_bdwt;
  input accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_14_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_14_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_14_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_14_i_q_d,
      accumulation_buffer_rsc_0_14_i_q_d_bfwt, accumulation_buffer_rsc_0_14_i_bcwt);
  assign accumulation_buffer_rsc_0_14_i_radr_d = {(~ accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_14_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_14_i_wadr_d = {(~ accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_14_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_14_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_14_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_14_i_bcwt <= ~((~(accumulation_buffer_rsc_0_14_i_bcwt
          | accumulation_buffer_rsc_0_14_i_biwt)) | accumulation_buffer_rsc_0_14_i_bdwt);
      accumulation_buffer_rsc_0_14_i_q_d_bfwt <= accumulation_buffer_rsc_0_14_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_14_i_oswt, accumulation_buffer_rsc_0_14_i_biwt,
      accumulation_buffer_rsc_0_14_i_bdwt, accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_14_i_oswt_pff, accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_14_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_14_i_oswt;
  output accumulation_buffer_rsc_0_14_i_biwt;
  output accumulation_buffer_rsc_0_14_i_bdwt;
  output accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_14_i_oswt_pff;
  output accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_14_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_14_i_bdwt = accumulation_buffer_rsc_0_14_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_14_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_14_i_oswt;
  assign accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_14_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_14_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_13_i_radr_d, accumulation_buffer_rsc_0_13_i_wadr_d,
      accumulation_buffer_rsc_0_13_i_q_d, accumulation_buffer_rsc_0_13_i_radr_d_run,
      accumulation_buffer_rsc_0_13_i_wadr_d_run, accumulation_buffer_rsc_0_13_i_q_d_mxwt,
      accumulation_buffer_rsc_0_13_i_biwt, accumulation_buffer_rsc_0_13_i_bdwt, accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_13_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_13_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_13_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_13_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_13_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_13_i_biwt;
  input accumulation_buffer_rsc_0_13_i_bdwt;
  input accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_13_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_13_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_13_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_13_i_q_d,
      accumulation_buffer_rsc_0_13_i_q_d_bfwt, accumulation_buffer_rsc_0_13_i_bcwt);
  assign accumulation_buffer_rsc_0_13_i_radr_d = {(~ accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_13_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_13_i_wadr_d = {(~ accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_13_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_13_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_13_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_13_i_bcwt <= ~((~(accumulation_buffer_rsc_0_13_i_bcwt
          | accumulation_buffer_rsc_0_13_i_biwt)) | accumulation_buffer_rsc_0_13_i_bdwt);
      accumulation_buffer_rsc_0_13_i_q_d_bfwt <= accumulation_buffer_rsc_0_13_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_13_i_oswt, accumulation_buffer_rsc_0_13_i_biwt,
      accumulation_buffer_rsc_0_13_i_bdwt, accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_13_i_oswt_pff, accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_13_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_13_i_oswt;
  output accumulation_buffer_rsc_0_13_i_biwt;
  output accumulation_buffer_rsc_0_13_i_bdwt;
  output accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_13_i_oswt_pff;
  output accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_13_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_13_i_bdwt = accumulation_buffer_rsc_0_13_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_13_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_13_i_oswt;
  assign accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_13_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_13_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_12_i_radr_d, accumulation_buffer_rsc_0_12_i_wadr_d,
      accumulation_buffer_rsc_0_12_i_q_d, accumulation_buffer_rsc_0_12_i_radr_d_run,
      accumulation_buffer_rsc_0_12_i_wadr_d_run, accumulation_buffer_rsc_0_12_i_q_d_mxwt,
      accumulation_buffer_rsc_0_12_i_biwt, accumulation_buffer_rsc_0_12_i_bdwt, accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_12_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_12_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_12_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_12_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_12_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_12_i_biwt;
  input accumulation_buffer_rsc_0_12_i_bdwt;
  input accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_12_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_12_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_12_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_12_i_q_d,
      accumulation_buffer_rsc_0_12_i_q_d_bfwt, accumulation_buffer_rsc_0_12_i_bcwt);
  assign accumulation_buffer_rsc_0_12_i_radr_d = {(~ accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_12_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_12_i_wadr_d = {(~ accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_12_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_12_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_12_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_12_i_bcwt <= ~((~(accumulation_buffer_rsc_0_12_i_bcwt
          | accumulation_buffer_rsc_0_12_i_biwt)) | accumulation_buffer_rsc_0_12_i_bdwt);
      accumulation_buffer_rsc_0_12_i_q_d_bfwt <= accumulation_buffer_rsc_0_12_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_12_i_oswt, accumulation_buffer_rsc_0_12_i_biwt,
      accumulation_buffer_rsc_0_12_i_bdwt, accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_12_i_oswt_pff, accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_12_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_12_i_oswt;
  output accumulation_buffer_rsc_0_12_i_biwt;
  output accumulation_buffer_rsc_0_12_i_bdwt;
  output accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_12_i_oswt_pff;
  output accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_12_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_12_i_bdwt = accumulation_buffer_rsc_0_12_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_12_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_12_i_oswt;
  assign accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_12_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_12_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_11_i_radr_d, accumulation_buffer_rsc_0_11_i_wadr_d,
      accumulation_buffer_rsc_0_11_i_q_d, accumulation_buffer_rsc_0_11_i_radr_d_run,
      accumulation_buffer_rsc_0_11_i_wadr_d_run, accumulation_buffer_rsc_0_11_i_q_d_mxwt,
      accumulation_buffer_rsc_0_11_i_biwt, accumulation_buffer_rsc_0_11_i_bdwt, accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_11_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_11_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_11_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_11_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_11_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_11_i_biwt;
  input accumulation_buffer_rsc_0_11_i_bdwt;
  input accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_11_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_11_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_11_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_11_i_q_d,
      accumulation_buffer_rsc_0_11_i_q_d_bfwt, accumulation_buffer_rsc_0_11_i_bcwt);
  assign accumulation_buffer_rsc_0_11_i_radr_d = {(~ accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_11_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_11_i_wadr_d = {(~ accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_11_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_11_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_11_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_11_i_bcwt <= ~((~(accumulation_buffer_rsc_0_11_i_bcwt
          | accumulation_buffer_rsc_0_11_i_biwt)) | accumulation_buffer_rsc_0_11_i_bdwt);
      accumulation_buffer_rsc_0_11_i_q_d_bfwt <= accumulation_buffer_rsc_0_11_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_11_i_oswt, accumulation_buffer_rsc_0_11_i_biwt,
      accumulation_buffer_rsc_0_11_i_bdwt, accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_11_i_oswt_pff, accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_11_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_11_i_oswt;
  output accumulation_buffer_rsc_0_11_i_biwt;
  output accumulation_buffer_rsc_0_11_i_bdwt;
  output accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_11_i_oswt_pff;
  output accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_11_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_11_i_bdwt = accumulation_buffer_rsc_0_11_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_11_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_11_i_oswt;
  assign accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_11_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_11_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_10_i_radr_d, accumulation_buffer_rsc_0_10_i_wadr_d,
      accumulation_buffer_rsc_0_10_i_q_d, accumulation_buffer_rsc_0_10_i_radr_d_run,
      accumulation_buffer_rsc_0_10_i_wadr_d_run, accumulation_buffer_rsc_0_10_i_q_d_mxwt,
      accumulation_buffer_rsc_0_10_i_biwt, accumulation_buffer_rsc_0_10_i_bdwt, accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_10_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_10_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_10_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_10_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_10_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_10_i_biwt;
  input accumulation_buffer_rsc_0_10_i_bdwt;
  input accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_10_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_10_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_10_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_10_i_q_d,
      accumulation_buffer_rsc_0_10_i_q_d_bfwt, accumulation_buffer_rsc_0_10_i_bcwt);
  assign accumulation_buffer_rsc_0_10_i_radr_d = {(~ accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_10_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_10_i_wadr_d = {(~ accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_10_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_10_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_10_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_10_i_bcwt <= ~((~(accumulation_buffer_rsc_0_10_i_bcwt
          | accumulation_buffer_rsc_0_10_i_biwt)) | accumulation_buffer_rsc_0_10_i_bdwt);
      accumulation_buffer_rsc_0_10_i_q_d_bfwt <= accumulation_buffer_rsc_0_10_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_10_i_oswt, accumulation_buffer_rsc_0_10_i_biwt,
      accumulation_buffer_rsc_0_10_i_bdwt, accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_10_i_oswt_pff, accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_10_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_10_i_oswt;
  output accumulation_buffer_rsc_0_10_i_biwt;
  output accumulation_buffer_rsc_0_10_i_bdwt;
  output accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_10_i_oswt_pff;
  output accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_10_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_10_i_bdwt = accumulation_buffer_rsc_0_10_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_10_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_10_i_oswt;
  assign accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_10_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_10_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_9_i_radr_d, accumulation_buffer_rsc_0_9_i_wadr_d,
      accumulation_buffer_rsc_0_9_i_q_d, accumulation_buffer_rsc_0_9_i_radr_d_run,
      accumulation_buffer_rsc_0_9_i_wadr_d_run, accumulation_buffer_rsc_0_9_i_q_d_mxwt,
      accumulation_buffer_rsc_0_9_i_biwt, accumulation_buffer_rsc_0_9_i_bdwt, accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_9_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_9_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_9_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_9_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_9_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_9_i_biwt;
  input accumulation_buffer_rsc_0_9_i_bdwt;
  input accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_9_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_9_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_9_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_9_i_q_d,
      accumulation_buffer_rsc_0_9_i_q_d_bfwt, accumulation_buffer_rsc_0_9_i_bcwt);
  assign accumulation_buffer_rsc_0_9_i_radr_d = {(~ accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_9_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_9_i_wadr_d = {(~ accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_9_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_9_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_9_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_9_i_bcwt <= ~((~(accumulation_buffer_rsc_0_9_i_bcwt
          | accumulation_buffer_rsc_0_9_i_biwt)) | accumulation_buffer_rsc_0_9_i_bdwt);
      accumulation_buffer_rsc_0_9_i_q_d_bfwt <= accumulation_buffer_rsc_0_9_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_9_i_oswt, accumulation_buffer_rsc_0_9_i_biwt,
      accumulation_buffer_rsc_0_9_i_bdwt, accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_9_i_oswt_pff, accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_9_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_9_i_oswt;
  output accumulation_buffer_rsc_0_9_i_biwt;
  output accumulation_buffer_rsc_0_9_i_bdwt;
  output accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_9_i_oswt_pff;
  output accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_9_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_9_i_bdwt = accumulation_buffer_rsc_0_9_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_9_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_9_i_oswt;
  assign accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_9_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_9_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_8_i_radr_d, accumulation_buffer_rsc_0_8_i_wadr_d,
      accumulation_buffer_rsc_0_8_i_q_d, accumulation_buffer_rsc_0_8_i_radr_d_run,
      accumulation_buffer_rsc_0_8_i_wadr_d_run, accumulation_buffer_rsc_0_8_i_q_d_mxwt,
      accumulation_buffer_rsc_0_8_i_biwt, accumulation_buffer_rsc_0_8_i_bdwt, accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_8_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_8_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_8_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_8_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_8_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_8_i_biwt;
  input accumulation_buffer_rsc_0_8_i_bdwt;
  input accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_8_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_8_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_8_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_8_i_q_d,
      accumulation_buffer_rsc_0_8_i_q_d_bfwt, accumulation_buffer_rsc_0_8_i_bcwt);
  assign accumulation_buffer_rsc_0_8_i_radr_d = {(~ accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_8_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_8_i_wadr_d = {(~ accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_8_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_8_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_8_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_8_i_bcwt <= ~((~(accumulation_buffer_rsc_0_8_i_bcwt
          | accumulation_buffer_rsc_0_8_i_biwt)) | accumulation_buffer_rsc_0_8_i_bdwt);
      accumulation_buffer_rsc_0_8_i_q_d_bfwt <= accumulation_buffer_rsc_0_8_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_8_i_oswt, accumulation_buffer_rsc_0_8_i_biwt,
      accumulation_buffer_rsc_0_8_i_bdwt, accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_8_i_oswt_pff, accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_8_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_8_i_oswt;
  output accumulation_buffer_rsc_0_8_i_biwt;
  output accumulation_buffer_rsc_0_8_i_bdwt;
  output accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_8_i_oswt_pff;
  output accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_8_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_8_i_bdwt = accumulation_buffer_rsc_0_8_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_8_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_8_i_oswt;
  assign accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_8_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_8_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_7_i_radr_d, accumulation_buffer_rsc_0_7_i_wadr_d,
      accumulation_buffer_rsc_0_7_i_q_d, accumulation_buffer_rsc_0_7_i_radr_d_run,
      accumulation_buffer_rsc_0_7_i_wadr_d_run, accumulation_buffer_rsc_0_7_i_q_d_mxwt,
      accumulation_buffer_rsc_0_7_i_biwt, accumulation_buffer_rsc_0_7_i_bdwt, accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_7_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_7_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_7_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_7_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_7_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_7_i_biwt;
  input accumulation_buffer_rsc_0_7_i_bdwt;
  input accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_7_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_7_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_7_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_7_i_q_d,
      accumulation_buffer_rsc_0_7_i_q_d_bfwt, accumulation_buffer_rsc_0_7_i_bcwt);
  assign accumulation_buffer_rsc_0_7_i_radr_d = {(~ accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_7_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_7_i_wadr_d = {(~ accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_7_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_7_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_7_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_7_i_bcwt <= ~((~(accumulation_buffer_rsc_0_7_i_bcwt
          | accumulation_buffer_rsc_0_7_i_biwt)) | accumulation_buffer_rsc_0_7_i_bdwt);
      accumulation_buffer_rsc_0_7_i_q_d_bfwt <= accumulation_buffer_rsc_0_7_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_7_i_oswt, accumulation_buffer_rsc_0_7_i_biwt,
      accumulation_buffer_rsc_0_7_i_bdwt, accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_7_i_oswt_pff, accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_7_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_7_i_oswt;
  output accumulation_buffer_rsc_0_7_i_biwt;
  output accumulation_buffer_rsc_0_7_i_bdwt;
  output accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_7_i_oswt_pff;
  output accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_7_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_7_i_bdwt = accumulation_buffer_rsc_0_7_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_7_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_7_i_oswt;
  assign accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_7_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_7_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_6_i_radr_d, accumulation_buffer_rsc_0_6_i_wadr_d,
      accumulation_buffer_rsc_0_6_i_q_d, accumulation_buffer_rsc_0_6_i_radr_d_run,
      accumulation_buffer_rsc_0_6_i_wadr_d_run, accumulation_buffer_rsc_0_6_i_q_d_mxwt,
      accumulation_buffer_rsc_0_6_i_biwt, accumulation_buffer_rsc_0_6_i_bdwt, accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_6_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_6_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_6_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_6_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_6_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_6_i_biwt;
  input accumulation_buffer_rsc_0_6_i_bdwt;
  input accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_6_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_6_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_6_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_6_i_q_d,
      accumulation_buffer_rsc_0_6_i_q_d_bfwt, accumulation_buffer_rsc_0_6_i_bcwt);
  assign accumulation_buffer_rsc_0_6_i_radr_d = {(~ accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_6_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_6_i_wadr_d = {(~ accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_6_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_6_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_6_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_6_i_bcwt <= ~((~(accumulation_buffer_rsc_0_6_i_bcwt
          | accumulation_buffer_rsc_0_6_i_biwt)) | accumulation_buffer_rsc_0_6_i_bdwt);
      accumulation_buffer_rsc_0_6_i_q_d_bfwt <= accumulation_buffer_rsc_0_6_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_6_i_oswt, accumulation_buffer_rsc_0_6_i_biwt,
      accumulation_buffer_rsc_0_6_i_bdwt, accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_6_i_oswt_pff, accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_6_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_6_i_oswt;
  output accumulation_buffer_rsc_0_6_i_biwt;
  output accumulation_buffer_rsc_0_6_i_bdwt;
  output accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_6_i_oswt_pff;
  output accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_6_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_6_i_bdwt = accumulation_buffer_rsc_0_6_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_6_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_6_i_oswt;
  assign accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_6_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_6_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_5_i_radr_d, accumulation_buffer_rsc_0_5_i_wadr_d,
      accumulation_buffer_rsc_0_5_i_q_d, accumulation_buffer_rsc_0_5_i_radr_d_run,
      accumulation_buffer_rsc_0_5_i_wadr_d_run, accumulation_buffer_rsc_0_5_i_q_d_mxwt,
      accumulation_buffer_rsc_0_5_i_biwt, accumulation_buffer_rsc_0_5_i_bdwt, accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_5_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_5_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_5_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_5_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_5_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_5_i_biwt;
  input accumulation_buffer_rsc_0_5_i_bdwt;
  input accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_5_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_5_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_5_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_5_i_q_d,
      accumulation_buffer_rsc_0_5_i_q_d_bfwt, accumulation_buffer_rsc_0_5_i_bcwt);
  assign accumulation_buffer_rsc_0_5_i_radr_d = {(~ accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_5_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_5_i_wadr_d = {(~ accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_5_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_5_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_5_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_5_i_bcwt <= ~((~(accumulation_buffer_rsc_0_5_i_bcwt
          | accumulation_buffer_rsc_0_5_i_biwt)) | accumulation_buffer_rsc_0_5_i_bdwt);
      accumulation_buffer_rsc_0_5_i_q_d_bfwt <= accumulation_buffer_rsc_0_5_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_5_i_oswt, accumulation_buffer_rsc_0_5_i_biwt,
      accumulation_buffer_rsc_0_5_i_bdwt, accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_5_i_oswt_pff, accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_5_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_5_i_oswt;
  output accumulation_buffer_rsc_0_5_i_biwt;
  output accumulation_buffer_rsc_0_5_i_bdwt;
  output accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_5_i_oswt_pff;
  output accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_5_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_5_i_bdwt = accumulation_buffer_rsc_0_5_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_5_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_5_i_oswt;
  assign accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_5_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_5_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_4_i_radr_d, accumulation_buffer_rsc_0_4_i_wadr_d,
      accumulation_buffer_rsc_0_4_i_q_d, accumulation_buffer_rsc_0_4_i_radr_d_run,
      accumulation_buffer_rsc_0_4_i_wadr_d_run, accumulation_buffer_rsc_0_4_i_q_d_mxwt,
      accumulation_buffer_rsc_0_4_i_biwt, accumulation_buffer_rsc_0_4_i_bdwt, accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_4_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_4_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_4_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_4_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_4_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_4_i_biwt;
  input accumulation_buffer_rsc_0_4_i_bdwt;
  input accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_4_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_4_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_4_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_4_i_q_d,
      accumulation_buffer_rsc_0_4_i_q_d_bfwt, accumulation_buffer_rsc_0_4_i_bcwt);
  assign accumulation_buffer_rsc_0_4_i_radr_d = {(~ accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_4_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_4_i_wadr_d = {(~ accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_4_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_4_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_4_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_4_i_bcwt <= ~((~(accumulation_buffer_rsc_0_4_i_bcwt
          | accumulation_buffer_rsc_0_4_i_biwt)) | accumulation_buffer_rsc_0_4_i_bdwt);
      accumulation_buffer_rsc_0_4_i_q_d_bfwt <= accumulation_buffer_rsc_0_4_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_4_i_oswt, accumulation_buffer_rsc_0_4_i_biwt,
      accumulation_buffer_rsc_0_4_i_bdwt, accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_4_i_oswt_pff, accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_4_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_4_i_oswt;
  output accumulation_buffer_rsc_0_4_i_biwt;
  output accumulation_buffer_rsc_0_4_i_bdwt;
  output accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_4_i_oswt_pff;
  output accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_4_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_4_i_bdwt = accumulation_buffer_rsc_0_4_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_4_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_4_i_oswt;
  assign accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_4_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_4_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_3_i_radr_d, accumulation_buffer_rsc_0_3_i_wadr_d,
      accumulation_buffer_rsc_0_3_i_q_d, accumulation_buffer_rsc_0_3_i_radr_d_run,
      accumulation_buffer_rsc_0_3_i_wadr_d_run, accumulation_buffer_rsc_0_3_i_q_d_mxwt,
      accumulation_buffer_rsc_0_3_i_biwt, accumulation_buffer_rsc_0_3_i_bdwt, accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_3_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_3_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_3_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_3_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_3_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_3_i_biwt;
  input accumulation_buffer_rsc_0_3_i_bdwt;
  input accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_3_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_3_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_3_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_3_i_q_d,
      accumulation_buffer_rsc_0_3_i_q_d_bfwt, accumulation_buffer_rsc_0_3_i_bcwt);
  assign accumulation_buffer_rsc_0_3_i_radr_d = {(~ accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_3_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_3_i_wadr_d = {(~ accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_3_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_3_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_3_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_3_i_bcwt <= ~((~(accumulation_buffer_rsc_0_3_i_bcwt
          | accumulation_buffer_rsc_0_3_i_biwt)) | accumulation_buffer_rsc_0_3_i_bdwt);
      accumulation_buffer_rsc_0_3_i_q_d_bfwt <= accumulation_buffer_rsc_0_3_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_3_i_oswt, accumulation_buffer_rsc_0_3_i_biwt,
      accumulation_buffer_rsc_0_3_i_bdwt, accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_3_i_oswt_pff, accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_3_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_3_i_oswt;
  output accumulation_buffer_rsc_0_3_i_biwt;
  output accumulation_buffer_rsc_0_3_i_bdwt;
  output accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_3_i_oswt_pff;
  output accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_3_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_3_i_bdwt = accumulation_buffer_rsc_0_3_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_3_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_3_i_oswt;
  assign accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_3_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_3_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_2_i_radr_d, accumulation_buffer_rsc_0_2_i_wadr_d,
      accumulation_buffer_rsc_0_2_i_q_d, accumulation_buffer_rsc_0_2_i_radr_d_run,
      accumulation_buffer_rsc_0_2_i_wadr_d_run, accumulation_buffer_rsc_0_2_i_q_d_mxwt,
      accumulation_buffer_rsc_0_2_i_biwt, accumulation_buffer_rsc_0_2_i_bdwt, accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_2_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_2_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_2_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_2_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_2_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_2_i_biwt;
  input accumulation_buffer_rsc_0_2_i_bdwt;
  input accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_2_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_2_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_2_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_2_i_q_d,
      accumulation_buffer_rsc_0_2_i_q_d_bfwt, accumulation_buffer_rsc_0_2_i_bcwt);
  assign accumulation_buffer_rsc_0_2_i_radr_d = {(~ accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_2_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_2_i_wadr_d = {(~ accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_2_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_2_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_2_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_2_i_bcwt <= ~((~(accumulation_buffer_rsc_0_2_i_bcwt
          | accumulation_buffer_rsc_0_2_i_biwt)) | accumulation_buffer_rsc_0_2_i_bdwt);
      accumulation_buffer_rsc_0_2_i_q_d_bfwt <= accumulation_buffer_rsc_0_2_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_2_i_oswt, accumulation_buffer_rsc_0_2_i_biwt,
      accumulation_buffer_rsc_0_2_i_bdwt, accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_2_i_oswt_pff, accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_2_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_2_i_oswt;
  output accumulation_buffer_rsc_0_2_i_biwt;
  output accumulation_buffer_rsc_0_2_i_bdwt;
  output accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_2_i_oswt_pff;
  output accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_2_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_2_i_bdwt = accumulation_buffer_rsc_0_2_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_2_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_2_i_oswt;
  assign accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_2_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_2_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_1_i_radr_d, accumulation_buffer_rsc_0_1_i_wadr_d,
      accumulation_buffer_rsc_0_1_i_q_d, accumulation_buffer_rsc_0_1_i_radr_d_run,
      accumulation_buffer_rsc_0_1_i_wadr_d_run, accumulation_buffer_rsc_0_1_i_q_d_mxwt,
      accumulation_buffer_rsc_0_1_i_biwt, accumulation_buffer_rsc_0_1_i_bdwt, accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_1_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_1_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_1_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_1_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_1_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_1_i_biwt;
  input accumulation_buffer_rsc_0_1_i_bdwt;
  input accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_1_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_1_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_1_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_1_i_q_d,
      accumulation_buffer_rsc_0_1_i_q_d_bfwt, accumulation_buffer_rsc_0_1_i_bcwt);
  assign accumulation_buffer_rsc_0_1_i_radr_d = {(~ accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_1_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_1_i_wadr_d = {(~ accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_1_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_1_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_1_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_1_i_bcwt <= ~((~(accumulation_buffer_rsc_0_1_i_bcwt
          | accumulation_buffer_rsc_0_1_i_biwt)) | accumulation_buffer_rsc_0_1_i_bdwt);
      accumulation_buffer_rsc_0_1_i_q_d_bfwt <= accumulation_buffer_rsc_0_1_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_1_i_oswt, accumulation_buffer_rsc_0_1_i_biwt,
      accumulation_buffer_rsc_0_1_i_bdwt, accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_1_i_oswt_pff, accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_1_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_1_i_oswt;
  output accumulation_buffer_rsc_0_1_i_biwt;
  output accumulation_buffer_rsc_0_1_i_bdwt;
  output accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_1_i_oswt_pff;
  output accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_1_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_1_i_bdwt = accumulation_buffer_rsc_0_1_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_1_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_1_i_oswt;
  assign accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_1_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_1_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
    (
  clk, arst_n, accumulation_buffer_rsc_0_0_i_radr_d, accumulation_buffer_rsc_0_0_i_wadr_d,
      accumulation_buffer_rsc_0_0_i_q_d, accumulation_buffer_rsc_0_0_i_radr_d_run,
      accumulation_buffer_rsc_0_0_i_wadr_d_run, accumulation_buffer_rsc_0_0_i_q_d_mxwt,
      accumulation_buffer_rsc_0_0_i_biwt, accumulation_buffer_rsc_0_0_i_bdwt, accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_0_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_0_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_q_d;
  input [7:0] accumulation_buffer_rsc_0_0_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_0_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_0_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_0_i_biwt;
  input accumulation_buffer_rsc_0_0_i_bdwt;
  input accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff;


  // Interconnect Declarations
  reg accumulation_buffer_rsc_0_0_i_bcwt;
  reg [15:0] accumulation_buffer_rsc_0_0_i_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_0_i_q_d_mxwt = MUX_v_16_2_2(accumulation_buffer_rsc_0_0_i_q_d,
      accumulation_buffer_rsc_0_0_i_q_d_bfwt, accumulation_buffer_rsc_0_0_i_bcwt);
  assign accumulation_buffer_rsc_0_0_i_radr_d = {(~ accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff) , (accumulation_buffer_rsc_0_0_i_radr_d_run[5:0])};
  assign accumulation_buffer_rsc_0_0_i_wadr_d = {(~ accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff)
      , (~ accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff) , (accumulation_buffer_rsc_0_0_i_wadr_d_run[5:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulation_buffer_rsc_0_0_i_bcwt <= 1'b0;
      accumulation_buffer_rsc_0_0_i_q_d_bfwt <= 16'b0000000000000000;
    end
    else begin
      accumulation_buffer_rsc_0_0_i_bcwt <= ~((~(accumulation_buffer_rsc_0_0_i_bcwt
          | accumulation_buffer_rsc_0_0_i_biwt)) | accumulation_buffer_rsc_0_0_i_bdwt);
      accumulation_buffer_rsc_0_0_i_q_d_bfwt <= accumulation_buffer_rsc_0_0_i_q_d_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
    (
  run_wen, run_wten, accumulation_buffer_rsc_0_0_i_oswt, accumulation_buffer_rsc_0_0_i_biwt,
      accumulation_buffer_rsc_0_0_i_bdwt, accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff,
      accumulation_buffer_rsc_0_0_i_oswt_pff, accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff,
      accumulation_buffer_rsc_0_0_i_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_0_i_oswt;
  output accumulation_buffer_rsc_0_0_i_biwt;
  output accumulation_buffer_rsc_0_0_i_bdwt;
  output accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_0_i_oswt_pff;
  output accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff;
  input accumulation_buffer_rsc_0_0_i_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accumulation_buffer_rsc_0_0_i_bdwt = accumulation_buffer_rsc_0_0_i_oswt
      & run_wen;
  assign accumulation_buffer_rsc_0_0_i_biwt = (~ run_wten) & accumulation_buffer_rsc_0_0_i_oswt;
  assign accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff = accumulation_buffer_rsc_0_0_i_oswt_pff
      & run_wen;
  assign accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff = accumulation_buffer_rsc_0_0_i_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
    (
  clk, arst_n, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt,
      loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt, loopIndicesIn_rsci_bcwt,
      loopIndicesIn_rsci_idat
);
  input clk;
  input arst_n;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [47:0] loopIndicesIn_rsci_idat_mxwt;
  input loopIndicesIn_rsci_biwt;
  input loopIndicesIn_rsci_bdwt;
  output loopIndicesIn_rsci_bcwt;
  reg loopIndicesIn_rsci_bcwt;
  input [47:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations
  reg [47:0] loopIndicesIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_wen_comp = (~ loopIndicesIn_rsci_oswt) | loopIndicesIn_rsci_biwt
      | loopIndicesIn_rsci_bcwt;
  assign loopIndicesIn_rsci_idat_mxwt = MUX_v_48_2_2(loopIndicesIn_rsci_idat, loopIndicesIn_rsci_idat_bfwt,
      loopIndicesIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_rsci_bcwt <= 1'b0;
      loopIndicesIn_rsci_idat_bfwt <= 48'b000000000000000000000000000000000000000000000000;
    end
    else begin
      loopIndicesIn_rsci_bcwt <= ~((~(loopIndicesIn_rsci_bcwt | loopIndicesIn_rsci_biwt))
          | loopIndicesIn_rsci_bdwt);
      loopIndicesIn_rsci_idat_bfwt <= loopIndicesIn_rsci_idat_mxwt;
    end
  end

  function automatic [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
    (
  run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt,
      loopIndicesIn_rsci_bcwt, loopIndicesIn_rsci_irdy_run_sct, loopIndicesIn_rsci_ivld
);
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_biwt;
  output loopIndicesIn_rsci_bdwt;
  input loopIndicesIn_rsci_bcwt;
  output loopIndicesIn_rsci_irdy_run_sct;
  input loopIndicesIn_rsci_ivld;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_bdwt = loopIndicesIn_rsci_oswt & run_wen;
  assign loopIndicesIn_rsci_biwt = loopIndicesIn_rsci_ogwt & loopIndicesIn_rsci_ivld;
  assign loopIndicesIn_rsci_ogwt = loopIndicesIn_rsci_oswt & (~ loopIndicesIn_rsci_bcwt);
  assign loopIndicesIn_rsci_irdy_run_sct = loopIndicesIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
    (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [79:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [47:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [31:0] reg_paramsIn_rsci_idat_bfwt_ftd_17;
  wire [47:0] paramsIn_rsci_idat_mxwt_opt_127_80;
  wire [31:0] paramsIn_rsci_idat_mxwt_opt_63_32;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_127_80 = MUX_v_48_2_2((paramsIn_rsci_idat[127:80]),
      reg_paramsIn_rsci_idat_bfwt_ftd, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_63_32 = MUX_v_32_2_2((paramsIn_rsci_idat[63:32]),
      reg_paramsIn_rsci_idat_bfwt_ftd_17, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {paramsIn_rsci_idat_mxwt_opt_127_80 , paramsIn_rsci_idat_mxwt_opt_63_32};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
      reg_paramsIn_rsci_idat_bfwt_ftd <= 48'b000000000000000000000000000000000000000000000000;
      reg_paramsIn_rsci_idat_bfwt_ftd_17 <= 32'b00000000000000000000000000000000;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_opt_127_80;
      reg_paramsIn_rsci_idat_bfwt_ftd_17 <= paramsIn_rsci_idat_mxwt_opt_63_32;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
    (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp
    (
  clk, arst_n, output_rsci_oswt, output_rsci_wen_comp, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_bcwt
);
  input clk;
  input arst_n;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input output_rsci_biwt;
  input output_rsci_bdwt;
  output output_rsci_bcwt;
  reg output_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_wen_comp = (~ output_rsci_oswt) | output_rsci_biwt | output_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_rsci_bcwt <= 1'b0;
    end
    else begin
      output_rsci_bcwt <= ~((~(output_rsci_bcwt | output_rsci_biwt)) | output_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl
    (
  run_wen, output_rsci_oswt, output_rsci_irdy, output_rsci_biwt, output_rsci_bdwt,
      output_rsci_bcwt, output_rsci_ivld_run_sct
);
  input run_wen;
  input output_rsci_oswt;
  input output_rsci_irdy;
  output output_rsci_biwt;
  output output_rsci_bdwt;
  input output_rsci_bcwt;
  output output_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire output_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_rsci_bdwt = output_rsci_oswt & run_wen;
  assign output_rsci_biwt = output_rsci_ogwt & output_rsci_irdy;
  assign output_rsci_ogwt = output_rsci_oswt & (~ output_rsci_bcwt);
  assign output_rsci_ivld_run_sct = output_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp
    (
  clk, arst_n, weight_rsci_oswt, weight_rsci_wen_comp, weight_rsci_idat_mxwt, weight_rsci_biwt,
      weight_rsci_bdwt, weight_rsci_bcwt, weight_rsci_idat
);
  input clk;
  input arst_n;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [127:0] weight_rsci_idat_mxwt;
  input weight_rsci_biwt;
  input weight_rsci_bdwt;
  output weight_rsci_bcwt;
  reg weight_rsci_bcwt;
  input [127:0] weight_rsci_idat;


  // Interconnect Declarations
  reg [127:0] weight_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_wen_comp = (~ weight_rsci_oswt) | weight_rsci_biwt | weight_rsci_bcwt;
  assign weight_rsci_idat_mxwt = MUX_v_128_2_2(weight_rsci_idat, weight_rsci_idat_bfwt,
      weight_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_rsci_bcwt <= 1'b0;
    end
    else begin
      weight_rsci_bcwt <= ~((~(weight_rsci_bcwt | weight_rsci_biwt)) | weight_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_rsci_idat_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ weight_rsci_bcwt ) begin
      weight_rsci_idat_bfwt <= weight_rsci_idat_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl
    (
  run_wen, weight_rsci_oswt, weight_rsci_biwt, weight_rsci_bdwt, weight_rsci_bcwt,
      weight_rsci_irdy_run_sct, weight_rsci_ivld
);
  input run_wen;
  input weight_rsci_oswt;
  output weight_rsci_biwt;
  output weight_rsci_bdwt;
  input weight_rsci_bcwt;
  output weight_rsci_irdy_run_sct;
  input weight_rsci_ivld;


  // Interconnect Declarations
  wire weight_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_rsci_bdwt = weight_rsci_oswt & run_wen;
  assign weight_rsci_biwt = weight_rsci_ogwt & weight_rsci_ivld;
  assign weight_rsci_ogwt = weight_rsci_oswt & (~ weight_rsci_bcwt);
  assign weight_rsci_irdy_run_sct = weight_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp
    (
  clk, arst_n, input_rsci_oswt, input_rsci_wen_comp, input_rsci_idat_mxwt, input_rsci_biwt,
      input_rsci_bdwt, input_rsci_bcwt, input_rsci_idat
);
  input clk;
  input arst_n;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [127:0] input_rsci_idat_mxwt;
  input input_rsci_biwt;
  input input_rsci_bdwt;
  output input_rsci_bcwt;
  reg input_rsci_bcwt;
  input [127:0] input_rsci_idat;


  // Interconnect Declarations
  reg [127:0] input_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_wen_comp = (~ input_rsci_oswt) | input_rsci_biwt | input_rsci_bcwt;
  assign input_rsci_idat_mxwt = MUX_v_128_2_2(input_rsci_idat, input_rsci_idat_bfwt,
      input_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_rsci_bcwt <= 1'b0;
      input_rsci_idat_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      input_rsci_bcwt <= ~((~(input_rsci_bcwt | input_rsci_biwt)) | input_rsci_bdwt);
      input_rsci_idat_bfwt <= input_rsci_idat_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl
    (
  run_wen, input_rsci_oswt, input_rsci_biwt, input_rsci_bdwt, input_rsci_bcwt, input_rsci_irdy_run_sct,
      input_rsci_ivld
);
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_biwt;
  output input_rsci_bdwt;
  input input_rsci_bcwt;
  output input_rsci_irdy_run_sct;
  input input_rsci_ivld;


  // Interconnect Declarations
  wire input_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_rsci_bdwt = input_rsci_oswt & run_wen;
  assign input_rsci_biwt = input_rsci_ogwt & input_rsci_ivld;
  assign input_rsci_ogwt = input_rsci_oswt & (~ input_rsci_bcwt);
  assign input_rsci_irdy_run_sct = input_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_15_i_radr_d, accumulation_buffer_rsc_0_15_i_wadr_d,
      accumulation_buffer_rsc_0_15_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_15_i_oswt,
      accumulation_buffer_rsc_0_15_i_radr_d_run, accumulation_buffer_rsc_0_15_i_wadr_d_run,
      accumulation_buffer_rsc_0_15_i_q_d_mxwt, accumulation_buffer_rsc_0_15_i_oswt_pff,
      accumulation_buffer_rsc_0_15_i_iswt0_1_pff, accumulation_buffer_rsc_0_15_i_we_d_pff,
      accumulation_buffer_rsc_0_15_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_15_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_15_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_15_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_15_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_15_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_15_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_15_i_oswt_pff;
  input accumulation_buffer_rsc_0_15_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_15_i_we_d_pff;
  output accumulation_buffer_rsc_0_15_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_15_i_biwt;
  wire accumulation_buffer_rsc_0_15_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_15_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_15_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_15_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_15_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_15_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_15_i_oswt(accumulation_buffer_rsc_0_15_i_oswt),
      .accumulation_buffer_rsc_0_15_i_biwt(accumulation_buffer_rsc_0_15_i_biwt),
      .accumulation_buffer_rsc_0_15_i_bdwt(accumulation_buffer_rsc_0_15_i_bdwt),
      .accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_15_i_oswt_pff(accumulation_buffer_rsc_0_15_i_oswt_pff),
      .accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_15_i_iswt0_1_pff(accumulation_buffer_rsc_0_15_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_15_i_radr_d(accumulation_buffer_rsc_0_15_i_radr_d_reg),
      .accumulation_buffer_rsc_0_15_i_wadr_d(accumulation_buffer_rsc_0_15_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_15_i_q_d(accumulation_buffer_rsc_0_15_i_q_d),
      .accumulation_buffer_rsc_0_15_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_15_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_accumulation_buffer_rsc_0_15_wait_dp_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_15_i_q_d_mxwt(accumulation_buffer_rsc_0_15_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_15_i_biwt(accumulation_buffer_rsc_0_15_i_biwt),
      .accumulation_buffer_rsc_0_15_i_bdwt(accumulation_buffer_rsc_0_15_i_bdwt),
      .accumulation_buffer_rsc_0_15_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_15_i_radr_d = accumulation_buffer_rsc_0_15_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_wadr_d = accumulation_buffer_rsc_0_15_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_we_d_pff = accumulation_buffer_rsc_0_15_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_15_i_re_d_pff = accumulation_buffer_rsc_0_15_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_14_i_radr_d, accumulation_buffer_rsc_0_14_i_wadr_d,
      accumulation_buffer_rsc_0_14_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_14_i_oswt,
      accumulation_buffer_rsc_0_14_i_radr_d_run, accumulation_buffer_rsc_0_14_i_wadr_d_run,
      accumulation_buffer_rsc_0_14_i_q_d_mxwt, accumulation_buffer_rsc_0_14_i_oswt_pff,
      accumulation_buffer_rsc_0_14_i_iswt0_1_pff, accumulation_buffer_rsc_0_14_i_we_d_pff,
      accumulation_buffer_rsc_0_14_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_14_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_14_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_14_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_14_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_14_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_14_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_14_i_oswt_pff;
  input accumulation_buffer_rsc_0_14_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_14_i_we_d_pff;
  output accumulation_buffer_rsc_0_14_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_14_i_biwt;
  wire accumulation_buffer_rsc_0_14_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_14_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_14_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_14_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_14_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_14_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_14_i_oswt(accumulation_buffer_rsc_0_14_i_oswt),
      .accumulation_buffer_rsc_0_14_i_biwt(accumulation_buffer_rsc_0_14_i_biwt),
      .accumulation_buffer_rsc_0_14_i_bdwt(accumulation_buffer_rsc_0_14_i_bdwt),
      .accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_14_i_oswt_pff(accumulation_buffer_rsc_0_14_i_oswt_pff),
      .accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_14_i_iswt0_1_pff(accumulation_buffer_rsc_0_14_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_14_i_radr_d(accumulation_buffer_rsc_0_14_i_radr_d_reg),
      .accumulation_buffer_rsc_0_14_i_wadr_d(accumulation_buffer_rsc_0_14_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_14_i_q_d(accumulation_buffer_rsc_0_14_i_q_d),
      .accumulation_buffer_rsc_0_14_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_14_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_accumulation_buffer_rsc_0_14_wait_dp_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_14_i_q_d_mxwt(accumulation_buffer_rsc_0_14_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_14_i_biwt(accumulation_buffer_rsc_0_14_i_biwt),
      .accumulation_buffer_rsc_0_14_i_bdwt(accumulation_buffer_rsc_0_14_i_bdwt),
      .accumulation_buffer_rsc_0_14_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_14_i_radr_d = accumulation_buffer_rsc_0_14_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_wadr_d = accumulation_buffer_rsc_0_14_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_we_d_pff = accumulation_buffer_rsc_0_14_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_14_i_re_d_pff = accumulation_buffer_rsc_0_14_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_13_i_radr_d, accumulation_buffer_rsc_0_13_i_wadr_d,
      accumulation_buffer_rsc_0_13_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_13_i_oswt,
      accumulation_buffer_rsc_0_13_i_radr_d_run, accumulation_buffer_rsc_0_13_i_wadr_d_run,
      accumulation_buffer_rsc_0_13_i_q_d_mxwt, accumulation_buffer_rsc_0_13_i_oswt_pff,
      accumulation_buffer_rsc_0_13_i_iswt0_1_pff, accumulation_buffer_rsc_0_13_i_we_d_pff,
      accumulation_buffer_rsc_0_13_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_13_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_13_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_13_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_13_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_13_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_13_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_13_i_oswt_pff;
  input accumulation_buffer_rsc_0_13_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_13_i_we_d_pff;
  output accumulation_buffer_rsc_0_13_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_13_i_biwt;
  wire accumulation_buffer_rsc_0_13_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_13_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_13_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_13_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_13_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_13_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_13_i_oswt(accumulation_buffer_rsc_0_13_i_oswt),
      .accumulation_buffer_rsc_0_13_i_biwt(accumulation_buffer_rsc_0_13_i_biwt),
      .accumulation_buffer_rsc_0_13_i_bdwt(accumulation_buffer_rsc_0_13_i_bdwt),
      .accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_13_i_oswt_pff(accumulation_buffer_rsc_0_13_i_oswt_pff),
      .accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_13_i_iswt0_1_pff(accumulation_buffer_rsc_0_13_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_13_i_radr_d(accumulation_buffer_rsc_0_13_i_radr_d_reg),
      .accumulation_buffer_rsc_0_13_i_wadr_d(accumulation_buffer_rsc_0_13_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_13_i_q_d(accumulation_buffer_rsc_0_13_i_q_d),
      .accumulation_buffer_rsc_0_13_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_13_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_accumulation_buffer_rsc_0_13_wait_dp_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_13_i_q_d_mxwt(accumulation_buffer_rsc_0_13_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_13_i_biwt(accumulation_buffer_rsc_0_13_i_biwt),
      .accumulation_buffer_rsc_0_13_i_bdwt(accumulation_buffer_rsc_0_13_i_bdwt),
      .accumulation_buffer_rsc_0_13_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_13_i_radr_d = accumulation_buffer_rsc_0_13_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_wadr_d = accumulation_buffer_rsc_0_13_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_we_d_pff = accumulation_buffer_rsc_0_13_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_13_i_re_d_pff = accumulation_buffer_rsc_0_13_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_12_i_radr_d, accumulation_buffer_rsc_0_12_i_wadr_d,
      accumulation_buffer_rsc_0_12_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_12_i_oswt,
      accumulation_buffer_rsc_0_12_i_radr_d_run, accumulation_buffer_rsc_0_12_i_wadr_d_run,
      accumulation_buffer_rsc_0_12_i_q_d_mxwt, accumulation_buffer_rsc_0_12_i_oswt_pff,
      accumulation_buffer_rsc_0_12_i_iswt0_1_pff, accumulation_buffer_rsc_0_12_i_we_d_pff,
      accumulation_buffer_rsc_0_12_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_12_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_12_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_12_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_12_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_12_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_12_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_12_i_oswt_pff;
  input accumulation_buffer_rsc_0_12_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_12_i_we_d_pff;
  output accumulation_buffer_rsc_0_12_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_12_i_biwt;
  wire accumulation_buffer_rsc_0_12_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_12_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_12_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_12_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_12_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_12_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_12_i_oswt(accumulation_buffer_rsc_0_12_i_oswt),
      .accumulation_buffer_rsc_0_12_i_biwt(accumulation_buffer_rsc_0_12_i_biwt),
      .accumulation_buffer_rsc_0_12_i_bdwt(accumulation_buffer_rsc_0_12_i_bdwt),
      .accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_12_i_oswt_pff(accumulation_buffer_rsc_0_12_i_oswt_pff),
      .accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_12_i_iswt0_1_pff(accumulation_buffer_rsc_0_12_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_12_i_radr_d(accumulation_buffer_rsc_0_12_i_radr_d_reg),
      .accumulation_buffer_rsc_0_12_i_wadr_d(accumulation_buffer_rsc_0_12_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_12_i_q_d(accumulation_buffer_rsc_0_12_i_q_d),
      .accumulation_buffer_rsc_0_12_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_12_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_accumulation_buffer_rsc_0_12_wait_dp_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_12_i_q_d_mxwt(accumulation_buffer_rsc_0_12_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_12_i_biwt(accumulation_buffer_rsc_0_12_i_biwt),
      .accumulation_buffer_rsc_0_12_i_bdwt(accumulation_buffer_rsc_0_12_i_bdwt),
      .accumulation_buffer_rsc_0_12_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_12_i_radr_d = accumulation_buffer_rsc_0_12_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_wadr_d = accumulation_buffer_rsc_0_12_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_we_d_pff = accumulation_buffer_rsc_0_12_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_12_i_re_d_pff = accumulation_buffer_rsc_0_12_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_11_i_radr_d, accumulation_buffer_rsc_0_11_i_wadr_d,
      accumulation_buffer_rsc_0_11_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_11_i_oswt,
      accumulation_buffer_rsc_0_11_i_radr_d_run, accumulation_buffer_rsc_0_11_i_wadr_d_run,
      accumulation_buffer_rsc_0_11_i_q_d_mxwt, accumulation_buffer_rsc_0_11_i_oswt_pff,
      accumulation_buffer_rsc_0_11_i_iswt0_1_pff, accumulation_buffer_rsc_0_11_i_we_d_pff,
      accumulation_buffer_rsc_0_11_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_11_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_11_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_11_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_11_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_11_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_11_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_11_i_oswt_pff;
  input accumulation_buffer_rsc_0_11_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_11_i_we_d_pff;
  output accumulation_buffer_rsc_0_11_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_11_i_biwt;
  wire accumulation_buffer_rsc_0_11_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_11_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_11_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_11_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_11_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_11_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_11_i_oswt(accumulation_buffer_rsc_0_11_i_oswt),
      .accumulation_buffer_rsc_0_11_i_biwt(accumulation_buffer_rsc_0_11_i_biwt),
      .accumulation_buffer_rsc_0_11_i_bdwt(accumulation_buffer_rsc_0_11_i_bdwt),
      .accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_11_i_oswt_pff(accumulation_buffer_rsc_0_11_i_oswt_pff),
      .accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_11_i_iswt0_1_pff(accumulation_buffer_rsc_0_11_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_11_i_radr_d(accumulation_buffer_rsc_0_11_i_radr_d_reg),
      .accumulation_buffer_rsc_0_11_i_wadr_d(accumulation_buffer_rsc_0_11_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_11_i_q_d(accumulation_buffer_rsc_0_11_i_q_d),
      .accumulation_buffer_rsc_0_11_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_11_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_accumulation_buffer_rsc_0_11_wait_dp_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_11_i_q_d_mxwt(accumulation_buffer_rsc_0_11_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_11_i_biwt(accumulation_buffer_rsc_0_11_i_biwt),
      .accumulation_buffer_rsc_0_11_i_bdwt(accumulation_buffer_rsc_0_11_i_bdwt),
      .accumulation_buffer_rsc_0_11_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_11_i_radr_d = accumulation_buffer_rsc_0_11_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_wadr_d = accumulation_buffer_rsc_0_11_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_we_d_pff = accumulation_buffer_rsc_0_11_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_11_i_re_d_pff = accumulation_buffer_rsc_0_11_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_10_i_radr_d, accumulation_buffer_rsc_0_10_i_wadr_d,
      accumulation_buffer_rsc_0_10_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_10_i_oswt,
      accumulation_buffer_rsc_0_10_i_radr_d_run, accumulation_buffer_rsc_0_10_i_wadr_d_run,
      accumulation_buffer_rsc_0_10_i_q_d_mxwt, accumulation_buffer_rsc_0_10_i_oswt_pff,
      accumulation_buffer_rsc_0_10_i_iswt0_1_pff, accumulation_buffer_rsc_0_10_i_we_d_pff,
      accumulation_buffer_rsc_0_10_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_10_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_10_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_10_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_10_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_10_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_10_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_10_i_oswt_pff;
  input accumulation_buffer_rsc_0_10_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_10_i_we_d_pff;
  output accumulation_buffer_rsc_0_10_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_10_i_biwt;
  wire accumulation_buffer_rsc_0_10_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_10_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_10_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_10_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_10_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_10_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_10_i_oswt(accumulation_buffer_rsc_0_10_i_oswt),
      .accumulation_buffer_rsc_0_10_i_biwt(accumulation_buffer_rsc_0_10_i_biwt),
      .accumulation_buffer_rsc_0_10_i_bdwt(accumulation_buffer_rsc_0_10_i_bdwt),
      .accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_10_i_oswt_pff(accumulation_buffer_rsc_0_10_i_oswt_pff),
      .accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_10_i_iswt0_1_pff(accumulation_buffer_rsc_0_10_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_10_i_radr_d(accumulation_buffer_rsc_0_10_i_radr_d_reg),
      .accumulation_buffer_rsc_0_10_i_wadr_d(accumulation_buffer_rsc_0_10_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_10_i_q_d(accumulation_buffer_rsc_0_10_i_q_d),
      .accumulation_buffer_rsc_0_10_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_10_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_accumulation_buffer_rsc_0_10_wait_dp_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_10_i_q_d_mxwt(accumulation_buffer_rsc_0_10_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_10_i_biwt(accumulation_buffer_rsc_0_10_i_biwt),
      .accumulation_buffer_rsc_0_10_i_bdwt(accumulation_buffer_rsc_0_10_i_bdwt),
      .accumulation_buffer_rsc_0_10_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_10_i_radr_d = accumulation_buffer_rsc_0_10_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_wadr_d = accumulation_buffer_rsc_0_10_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_we_d_pff = accumulation_buffer_rsc_0_10_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_10_i_re_d_pff = accumulation_buffer_rsc_0_10_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_9_i_radr_d, accumulation_buffer_rsc_0_9_i_wadr_d,
      accumulation_buffer_rsc_0_9_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_9_i_oswt,
      accumulation_buffer_rsc_0_9_i_radr_d_run, accumulation_buffer_rsc_0_9_i_wadr_d_run,
      accumulation_buffer_rsc_0_9_i_q_d_mxwt, accumulation_buffer_rsc_0_9_i_oswt_pff,
      accumulation_buffer_rsc_0_9_i_iswt0_1_pff, accumulation_buffer_rsc_0_9_i_we_d_pff,
      accumulation_buffer_rsc_0_9_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_9_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_9_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_9_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_9_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_9_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_9_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_9_i_oswt_pff;
  input accumulation_buffer_rsc_0_9_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_9_i_we_d_pff;
  output accumulation_buffer_rsc_0_9_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_9_i_biwt;
  wire accumulation_buffer_rsc_0_9_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_9_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_9_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_9_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_9_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_9_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_9_i_oswt(accumulation_buffer_rsc_0_9_i_oswt),
      .accumulation_buffer_rsc_0_9_i_biwt(accumulation_buffer_rsc_0_9_i_biwt),
      .accumulation_buffer_rsc_0_9_i_bdwt(accumulation_buffer_rsc_0_9_i_bdwt),
      .accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_9_i_oswt_pff(accumulation_buffer_rsc_0_9_i_oswt_pff),
      .accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_9_i_iswt0_1_pff(accumulation_buffer_rsc_0_9_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_9_i_radr_d(accumulation_buffer_rsc_0_9_i_radr_d_reg),
      .accumulation_buffer_rsc_0_9_i_wadr_d(accumulation_buffer_rsc_0_9_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_9_i_q_d(accumulation_buffer_rsc_0_9_i_q_d),
      .accumulation_buffer_rsc_0_9_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_9_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_accumulation_buffer_rsc_0_9_wait_dp_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_9_i_q_d_mxwt(accumulation_buffer_rsc_0_9_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_9_i_biwt(accumulation_buffer_rsc_0_9_i_biwt),
      .accumulation_buffer_rsc_0_9_i_bdwt(accumulation_buffer_rsc_0_9_i_bdwt),
      .accumulation_buffer_rsc_0_9_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_9_i_radr_d = accumulation_buffer_rsc_0_9_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_wadr_d = accumulation_buffer_rsc_0_9_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_we_d_pff = accumulation_buffer_rsc_0_9_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_9_i_re_d_pff = accumulation_buffer_rsc_0_9_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_8_i_radr_d, accumulation_buffer_rsc_0_8_i_wadr_d,
      accumulation_buffer_rsc_0_8_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_8_i_oswt,
      accumulation_buffer_rsc_0_8_i_radr_d_run, accumulation_buffer_rsc_0_8_i_wadr_d_run,
      accumulation_buffer_rsc_0_8_i_q_d_mxwt, accumulation_buffer_rsc_0_8_i_oswt_pff,
      accumulation_buffer_rsc_0_8_i_iswt0_1_pff, accumulation_buffer_rsc_0_8_i_we_d_pff,
      accumulation_buffer_rsc_0_8_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_8_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_8_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_8_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_8_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_8_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_8_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_8_i_oswt_pff;
  input accumulation_buffer_rsc_0_8_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_8_i_we_d_pff;
  output accumulation_buffer_rsc_0_8_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_8_i_biwt;
  wire accumulation_buffer_rsc_0_8_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_8_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_8_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_8_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_8_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_8_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_8_i_oswt(accumulation_buffer_rsc_0_8_i_oswt),
      .accumulation_buffer_rsc_0_8_i_biwt(accumulation_buffer_rsc_0_8_i_biwt),
      .accumulation_buffer_rsc_0_8_i_bdwt(accumulation_buffer_rsc_0_8_i_bdwt),
      .accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_8_i_oswt_pff(accumulation_buffer_rsc_0_8_i_oswt_pff),
      .accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_8_i_iswt0_1_pff(accumulation_buffer_rsc_0_8_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_8_i_radr_d(accumulation_buffer_rsc_0_8_i_radr_d_reg),
      .accumulation_buffer_rsc_0_8_i_wadr_d(accumulation_buffer_rsc_0_8_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_8_i_q_d(accumulation_buffer_rsc_0_8_i_q_d),
      .accumulation_buffer_rsc_0_8_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_8_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_accumulation_buffer_rsc_0_8_wait_dp_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_8_i_q_d_mxwt(accumulation_buffer_rsc_0_8_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_8_i_biwt(accumulation_buffer_rsc_0_8_i_biwt),
      .accumulation_buffer_rsc_0_8_i_bdwt(accumulation_buffer_rsc_0_8_i_bdwt),
      .accumulation_buffer_rsc_0_8_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_8_i_radr_d = accumulation_buffer_rsc_0_8_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_wadr_d = accumulation_buffer_rsc_0_8_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_we_d_pff = accumulation_buffer_rsc_0_8_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_8_i_re_d_pff = accumulation_buffer_rsc_0_8_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_7_i_radr_d, accumulation_buffer_rsc_0_7_i_wadr_d,
      accumulation_buffer_rsc_0_7_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_7_i_oswt,
      accumulation_buffer_rsc_0_7_i_radr_d_run, accumulation_buffer_rsc_0_7_i_wadr_d_run,
      accumulation_buffer_rsc_0_7_i_q_d_mxwt, accumulation_buffer_rsc_0_7_i_oswt_pff,
      accumulation_buffer_rsc_0_7_i_iswt0_1_pff, accumulation_buffer_rsc_0_7_i_we_d_pff,
      accumulation_buffer_rsc_0_7_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_7_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_7_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_7_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_7_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_7_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_7_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_7_i_oswt_pff;
  input accumulation_buffer_rsc_0_7_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_7_i_we_d_pff;
  output accumulation_buffer_rsc_0_7_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_7_i_biwt;
  wire accumulation_buffer_rsc_0_7_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_7_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_7_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_7_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_7_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_7_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_7_i_oswt(accumulation_buffer_rsc_0_7_i_oswt),
      .accumulation_buffer_rsc_0_7_i_biwt(accumulation_buffer_rsc_0_7_i_biwt),
      .accumulation_buffer_rsc_0_7_i_bdwt(accumulation_buffer_rsc_0_7_i_bdwt),
      .accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_7_i_oswt_pff(accumulation_buffer_rsc_0_7_i_oswt_pff),
      .accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_7_i_iswt0_1_pff(accumulation_buffer_rsc_0_7_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_7_i_radr_d(accumulation_buffer_rsc_0_7_i_radr_d_reg),
      .accumulation_buffer_rsc_0_7_i_wadr_d(accumulation_buffer_rsc_0_7_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_7_i_q_d(accumulation_buffer_rsc_0_7_i_q_d),
      .accumulation_buffer_rsc_0_7_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_7_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_accumulation_buffer_rsc_0_7_wait_dp_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_7_i_q_d_mxwt(accumulation_buffer_rsc_0_7_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_7_i_biwt(accumulation_buffer_rsc_0_7_i_biwt),
      .accumulation_buffer_rsc_0_7_i_bdwt(accumulation_buffer_rsc_0_7_i_bdwt),
      .accumulation_buffer_rsc_0_7_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_7_i_radr_d = accumulation_buffer_rsc_0_7_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_wadr_d = accumulation_buffer_rsc_0_7_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_we_d_pff = accumulation_buffer_rsc_0_7_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_7_i_re_d_pff = accumulation_buffer_rsc_0_7_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_6_i_radr_d, accumulation_buffer_rsc_0_6_i_wadr_d,
      accumulation_buffer_rsc_0_6_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_6_i_oswt,
      accumulation_buffer_rsc_0_6_i_radr_d_run, accumulation_buffer_rsc_0_6_i_wadr_d_run,
      accumulation_buffer_rsc_0_6_i_q_d_mxwt, accumulation_buffer_rsc_0_6_i_oswt_pff,
      accumulation_buffer_rsc_0_6_i_iswt0_1_pff, accumulation_buffer_rsc_0_6_i_we_d_pff,
      accumulation_buffer_rsc_0_6_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_6_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_6_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_6_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_6_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_6_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_6_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_6_i_oswt_pff;
  input accumulation_buffer_rsc_0_6_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_6_i_we_d_pff;
  output accumulation_buffer_rsc_0_6_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_6_i_biwt;
  wire accumulation_buffer_rsc_0_6_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_6_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_6_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_6_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_6_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_6_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_6_i_oswt(accumulation_buffer_rsc_0_6_i_oswt),
      .accumulation_buffer_rsc_0_6_i_biwt(accumulation_buffer_rsc_0_6_i_biwt),
      .accumulation_buffer_rsc_0_6_i_bdwt(accumulation_buffer_rsc_0_6_i_bdwt),
      .accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_6_i_oswt_pff(accumulation_buffer_rsc_0_6_i_oswt_pff),
      .accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_6_i_iswt0_1_pff(accumulation_buffer_rsc_0_6_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_6_i_radr_d(accumulation_buffer_rsc_0_6_i_radr_d_reg),
      .accumulation_buffer_rsc_0_6_i_wadr_d(accumulation_buffer_rsc_0_6_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_6_i_q_d(accumulation_buffer_rsc_0_6_i_q_d),
      .accumulation_buffer_rsc_0_6_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_6_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_accumulation_buffer_rsc_0_6_wait_dp_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_6_i_q_d_mxwt(accumulation_buffer_rsc_0_6_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_6_i_biwt(accumulation_buffer_rsc_0_6_i_biwt),
      .accumulation_buffer_rsc_0_6_i_bdwt(accumulation_buffer_rsc_0_6_i_bdwt),
      .accumulation_buffer_rsc_0_6_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_6_i_radr_d = accumulation_buffer_rsc_0_6_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_wadr_d = accumulation_buffer_rsc_0_6_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_we_d_pff = accumulation_buffer_rsc_0_6_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_6_i_re_d_pff = accumulation_buffer_rsc_0_6_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_5_i_radr_d, accumulation_buffer_rsc_0_5_i_wadr_d,
      accumulation_buffer_rsc_0_5_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_5_i_oswt,
      accumulation_buffer_rsc_0_5_i_radr_d_run, accumulation_buffer_rsc_0_5_i_wadr_d_run,
      accumulation_buffer_rsc_0_5_i_q_d_mxwt, accumulation_buffer_rsc_0_5_i_oswt_pff,
      accumulation_buffer_rsc_0_5_i_iswt0_1_pff, accumulation_buffer_rsc_0_5_i_we_d_pff,
      accumulation_buffer_rsc_0_5_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_5_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_5_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_5_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_5_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_5_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_5_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_5_i_oswt_pff;
  input accumulation_buffer_rsc_0_5_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_5_i_we_d_pff;
  output accumulation_buffer_rsc_0_5_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_5_i_biwt;
  wire accumulation_buffer_rsc_0_5_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_5_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_5_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_5_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_5_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_5_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_5_i_oswt(accumulation_buffer_rsc_0_5_i_oswt),
      .accumulation_buffer_rsc_0_5_i_biwt(accumulation_buffer_rsc_0_5_i_biwt),
      .accumulation_buffer_rsc_0_5_i_bdwt(accumulation_buffer_rsc_0_5_i_bdwt),
      .accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_5_i_oswt_pff(accumulation_buffer_rsc_0_5_i_oswt_pff),
      .accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_5_i_iswt0_1_pff(accumulation_buffer_rsc_0_5_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_5_i_radr_d(accumulation_buffer_rsc_0_5_i_radr_d_reg),
      .accumulation_buffer_rsc_0_5_i_wadr_d(accumulation_buffer_rsc_0_5_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_5_i_q_d(accumulation_buffer_rsc_0_5_i_q_d),
      .accumulation_buffer_rsc_0_5_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_5_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_accumulation_buffer_rsc_0_5_wait_dp_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_5_i_q_d_mxwt(accumulation_buffer_rsc_0_5_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_5_i_biwt(accumulation_buffer_rsc_0_5_i_biwt),
      .accumulation_buffer_rsc_0_5_i_bdwt(accumulation_buffer_rsc_0_5_i_bdwt),
      .accumulation_buffer_rsc_0_5_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_5_i_radr_d = accumulation_buffer_rsc_0_5_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_wadr_d = accumulation_buffer_rsc_0_5_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_we_d_pff = accumulation_buffer_rsc_0_5_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_5_i_re_d_pff = accumulation_buffer_rsc_0_5_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_4_i_radr_d, accumulation_buffer_rsc_0_4_i_wadr_d,
      accumulation_buffer_rsc_0_4_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_4_i_oswt,
      accumulation_buffer_rsc_0_4_i_radr_d_run, accumulation_buffer_rsc_0_4_i_wadr_d_run,
      accumulation_buffer_rsc_0_4_i_q_d_mxwt, accumulation_buffer_rsc_0_4_i_oswt_pff,
      accumulation_buffer_rsc_0_4_i_iswt0_1_pff, accumulation_buffer_rsc_0_4_i_we_d_pff,
      accumulation_buffer_rsc_0_4_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_4_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_4_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_4_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_4_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_4_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_4_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_4_i_oswt_pff;
  input accumulation_buffer_rsc_0_4_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_4_i_we_d_pff;
  output accumulation_buffer_rsc_0_4_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_4_i_biwt;
  wire accumulation_buffer_rsc_0_4_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_4_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_4_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_4_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_4_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_4_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_4_i_oswt(accumulation_buffer_rsc_0_4_i_oswt),
      .accumulation_buffer_rsc_0_4_i_biwt(accumulation_buffer_rsc_0_4_i_biwt),
      .accumulation_buffer_rsc_0_4_i_bdwt(accumulation_buffer_rsc_0_4_i_bdwt),
      .accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_4_i_oswt_pff(accumulation_buffer_rsc_0_4_i_oswt_pff),
      .accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_4_i_iswt0_1_pff(accumulation_buffer_rsc_0_4_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_4_i_radr_d(accumulation_buffer_rsc_0_4_i_radr_d_reg),
      .accumulation_buffer_rsc_0_4_i_wadr_d(accumulation_buffer_rsc_0_4_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_4_i_q_d(accumulation_buffer_rsc_0_4_i_q_d),
      .accumulation_buffer_rsc_0_4_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_4_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_accumulation_buffer_rsc_0_4_wait_dp_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_4_i_q_d_mxwt(accumulation_buffer_rsc_0_4_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_4_i_biwt(accumulation_buffer_rsc_0_4_i_biwt),
      .accumulation_buffer_rsc_0_4_i_bdwt(accumulation_buffer_rsc_0_4_i_bdwt),
      .accumulation_buffer_rsc_0_4_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_4_i_radr_d = accumulation_buffer_rsc_0_4_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_wadr_d = accumulation_buffer_rsc_0_4_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_we_d_pff = accumulation_buffer_rsc_0_4_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_4_i_re_d_pff = accumulation_buffer_rsc_0_4_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_3_i_radr_d, accumulation_buffer_rsc_0_3_i_wadr_d,
      accumulation_buffer_rsc_0_3_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_3_i_oswt,
      accumulation_buffer_rsc_0_3_i_radr_d_run, accumulation_buffer_rsc_0_3_i_wadr_d_run,
      accumulation_buffer_rsc_0_3_i_q_d_mxwt, accumulation_buffer_rsc_0_3_i_oswt_pff,
      accumulation_buffer_rsc_0_3_i_iswt0_1_pff, accumulation_buffer_rsc_0_3_i_we_d_pff,
      accumulation_buffer_rsc_0_3_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_3_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_3_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_3_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_3_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_3_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_3_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_3_i_oswt_pff;
  input accumulation_buffer_rsc_0_3_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_3_i_we_d_pff;
  output accumulation_buffer_rsc_0_3_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_3_i_biwt;
  wire accumulation_buffer_rsc_0_3_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_3_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_3_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_3_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_3_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_3_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_3_i_oswt(accumulation_buffer_rsc_0_3_i_oswt),
      .accumulation_buffer_rsc_0_3_i_biwt(accumulation_buffer_rsc_0_3_i_biwt),
      .accumulation_buffer_rsc_0_3_i_bdwt(accumulation_buffer_rsc_0_3_i_bdwt),
      .accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_3_i_oswt_pff(accumulation_buffer_rsc_0_3_i_oswt_pff),
      .accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_3_i_iswt0_1_pff(accumulation_buffer_rsc_0_3_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_3_i_radr_d(accumulation_buffer_rsc_0_3_i_radr_d_reg),
      .accumulation_buffer_rsc_0_3_i_wadr_d(accumulation_buffer_rsc_0_3_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_3_i_q_d(accumulation_buffer_rsc_0_3_i_q_d),
      .accumulation_buffer_rsc_0_3_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_3_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_accumulation_buffer_rsc_0_3_wait_dp_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_3_i_q_d_mxwt(accumulation_buffer_rsc_0_3_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_3_i_biwt(accumulation_buffer_rsc_0_3_i_biwt),
      .accumulation_buffer_rsc_0_3_i_bdwt(accumulation_buffer_rsc_0_3_i_bdwt),
      .accumulation_buffer_rsc_0_3_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_3_i_radr_d = accumulation_buffer_rsc_0_3_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_wadr_d = accumulation_buffer_rsc_0_3_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_we_d_pff = accumulation_buffer_rsc_0_3_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_3_i_re_d_pff = accumulation_buffer_rsc_0_3_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_2_i_radr_d, accumulation_buffer_rsc_0_2_i_wadr_d,
      accumulation_buffer_rsc_0_2_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_2_i_oswt,
      accumulation_buffer_rsc_0_2_i_radr_d_run, accumulation_buffer_rsc_0_2_i_wadr_d_run,
      accumulation_buffer_rsc_0_2_i_q_d_mxwt, accumulation_buffer_rsc_0_2_i_oswt_pff,
      accumulation_buffer_rsc_0_2_i_iswt0_1_pff, accumulation_buffer_rsc_0_2_i_we_d_pff,
      accumulation_buffer_rsc_0_2_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_2_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_2_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_2_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_2_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_2_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_2_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_2_i_oswt_pff;
  input accumulation_buffer_rsc_0_2_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_2_i_we_d_pff;
  output accumulation_buffer_rsc_0_2_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_2_i_biwt;
  wire accumulation_buffer_rsc_0_2_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_2_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_2_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_2_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_2_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_2_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_2_i_oswt(accumulation_buffer_rsc_0_2_i_oswt),
      .accumulation_buffer_rsc_0_2_i_biwt(accumulation_buffer_rsc_0_2_i_biwt),
      .accumulation_buffer_rsc_0_2_i_bdwt(accumulation_buffer_rsc_0_2_i_bdwt),
      .accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_2_i_oswt_pff(accumulation_buffer_rsc_0_2_i_oswt_pff),
      .accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_2_i_iswt0_1_pff(accumulation_buffer_rsc_0_2_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_2_i_radr_d(accumulation_buffer_rsc_0_2_i_radr_d_reg),
      .accumulation_buffer_rsc_0_2_i_wadr_d(accumulation_buffer_rsc_0_2_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_2_i_q_d(accumulation_buffer_rsc_0_2_i_q_d),
      .accumulation_buffer_rsc_0_2_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_2_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_accumulation_buffer_rsc_0_2_wait_dp_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_2_i_q_d_mxwt(accumulation_buffer_rsc_0_2_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_2_i_biwt(accumulation_buffer_rsc_0_2_i_biwt),
      .accumulation_buffer_rsc_0_2_i_bdwt(accumulation_buffer_rsc_0_2_i_bdwt),
      .accumulation_buffer_rsc_0_2_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_2_i_radr_d = accumulation_buffer_rsc_0_2_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_wadr_d = accumulation_buffer_rsc_0_2_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_we_d_pff = accumulation_buffer_rsc_0_2_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_2_i_re_d_pff = accumulation_buffer_rsc_0_2_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_1_i_radr_d, accumulation_buffer_rsc_0_1_i_wadr_d,
      accumulation_buffer_rsc_0_1_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_1_i_oswt,
      accumulation_buffer_rsc_0_1_i_radr_d_run, accumulation_buffer_rsc_0_1_i_wadr_d_run,
      accumulation_buffer_rsc_0_1_i_q_d_mxwt, accumulation_buffer_rsc_0_1_i_oswt_pff,
      accumulation_buffer_rsc_0_1_i_iswt0_1_pff, accumulation_buffer_rsc_0_1_i_we_d_pff,
      accumulation_buffer_rsc_0_1_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_1_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_1_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_1_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_1_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_1_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_1_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_1_i_oswt_pff;
  input accumulation_buffer_rsc_0_1_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_1_i_we_d_pff;
  output accumulation_buffer_rsc_0_1_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_1_i_biwt;
  wire accumulation_buffer_rsc_0_1_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_1_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_1_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_1_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_1_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_1_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_1_i_oswt(accumulation_buffer_rsc_0_1_i_oswt),
      .accumulation_buffer_rsc_0_1_i_biwt(accumulation_buffer_rsc_0_1_i_biwt),
      .accumulation_buffer_rsc_0_1_i_bdwt(accumulation_buffer_rsc_0_1_i_bdwt),
      .accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_1_i_oswt_pff(accumulation_buffer_rsc_0_1_i_oswt_pff),
      .accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_1_i_iswt0_1_pff(accumulation_buffer_rsc_0_1_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_1_i_radr_d(accumulation_buffer_rsc_0_1_i_radr_d_reg),
      .accumulation_buffer_rsc_0_1_i_wadr_d(accumulation_buffer_rsc_0_1_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_1_i_q_d(accumulation_buffer_rsc_0_1_i_q_d),
      .accumulation_buffer_rsc_0_1_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_1_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_accumulation_buffer_rsc_0_1_wait_dp_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_1_i_q_d_mxwt(accumulation_buffer_rsc_0_1_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_1_i_biwt(accumulation_buffer_rsc_0_1_i_biwt),
      .accumulation_buffer_rsc_0_1_i_bdwt(accumulation_buffer_rsc_0_1_i_bdwt),
      .accumulation_buffer_rsc_0_1_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_1_i_radr_d = accumulation_buffer_rsc_0_1_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_wadr_d = accumulation_buffer_rsc_0_1_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_we_d_pff = accumulation_buffer_rsc_0_1_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_1_i_re_d_pff = accumulation_buffer_rsc_0_1_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
    (
  clk, arst_n, accumulation_buffer_rsc_0_0_i_radr_d, accumulation_buffer_rsc_0_0_i_wadr_d,
      accumulation_buffer_rsc_0_0_i_q_d, run_wen, run_wten, accumulation_buffer_rsc_0_0_i_oswt,
      accumulation_buffer_rsc_0_0_i_radr_d_run, accumulation_buffer_rsc_0_0_i_wadr_d_run,
      accumulation_buffer_rsc_0_0_i_q_d_mxwt, accumulation_buffer_rsc_0_0_i_oswt_pff,
      accumulation_buffer_rsc_0_0_i_iswt0_1_pff, accumulation_buffer_rsc_0_0_i_we_d_pff,
      accumulation_buffer_rsc_0_0_i_re_d_pff
);
  input clk;
  input arst_n;
  output [7:0] accumulation_buffer_rsc_0_0_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_0_i_wadr_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_q_d;
  input run_wen;
  input run_wten;
  input accumulation_buffer_rsc_0_0_i_oswt;
  input [7:0] accumulation_buffer_rsc_0_0_i_radr_d_run;
  input [7:0] accumulation_buffer_rsc_0_0_i_wadr_d_run;
  output [15:0] accumulation_buffer_rsc_0_0_i_q_d_mxwt;
  input accumulation_buffer_rsc_0_0_i_oswt_pff;
  input accumulation_buffer_rsc_0_0_i_iswt0_1_pff;
  output accumulation_buffer_rsc_0_0_i_we_d_pff;
  output accumulation_buffer_rsc_0_0_i_re_d_pff;


  // Interconnect Declarations
  wire accumulation_buffer_rsc_0_0_i_biwt;
  wire accumulation_buffer_rsc_0_0_i_bdwt;
  wire [7:0] accumulation_buffer_rsc_0_0_i_radr_d_reg;
  wire accumulation_buffer_rsc_0_0_i_radr_d_run_sct_iff;
  wire [7:0] accumulation_buffer_rsc_0_0_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_radr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_0_i_radr_d_run[5:0])};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run
      = {2'b00 , (accumulation_buffer_rsc_0_0_i_wadr_d_run[5:0])};
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_0_i_oswt(accumulation_buffer_rsc_0_0_i_oswt),
      .accumulation_buffer_rsc_0_0_i_biwt(accumulation_buffer_rsc_0_0_i_biwt),
      .accumulation_buffer_rsc_0_0_i_bdwt(accumulation_buffer_rsc_0_0_i_bdwt),
      .accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_0_i_oswt_pff(accumulation_buffer_rsc_0_0_i_oswt_pff),
      .accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_0_i_iswt0_1_pff(accumulation_buffer_rsc_0_0_i_iswt0_1_pff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_0_i_radr_d(accumulation_buffer_rsc_0_0_i_radr_d_reg),
      .accumulation_buffer_rsc_0_0_i_wadr_d(accumulation_buffer_rsc_0_0_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_0_i_q_d(accumulation_buffer_rsc_0_0_i_q_d),
      .accumulation_buffer_rsc_0_0_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_0_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_accumulation_buffer_rsc_0_0_wait_dp_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_0_i_q_d_mxwt(accumulation_buffer_rsc_0_0_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_0_i_biwt(accumulation_buffer_rsc_0_0_i_biwt),
      .accumulation_buffer_rsc_0_0_i_bdwt(accumulation_buffer_rsc_0_0_i_bdwt),
      .accumulation_buffer_rsc_0_0_i_radr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_radr_d_run_sct_iff),
      .accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_pff(accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_iff)
    );
  assign accumulation_buffer_rsc_0_0_i_radr_d = accumulation_buffer_rsc_0_0_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_wadr_d = accumulation_buffer_rsc_0_0_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_we_d_pff = accumulation_buffer_rsc_0_0_i_wadr_d_run_sct_iff;
  assign accumulation_buffer_rsc_0_0_i_re_d_pff = accumulation_buffer_rsc_0_0_i_radr_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci (
  clk, arst_n, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld, loopIndicesIn_rsc_rdy,
      run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [47:0] loopIndicesIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_biwt;
  wire loopIndicesIn_rsci_bdwt;
  wire loopIndicesIn_rsci_bcwt;
  wire loopIndicesIn_rsci_irdy_run_sct;
  wire loopIndicesIn_rsci_ivld;
  wire [47:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd104),
  .width(32'sd48)) loopIndicesIn_rsci (
      .rdy(loopIndicesIn_rsc_rdy),
      .vld(loopIndicesIn_rsc_vld),
      .dat(loopIndicesIn_rsc_dat),
      .irdy(loopIndicesIn_rsci_irdy_run_sct),
      .ivld(loopIndicesIn_rsci_ivld),
      .idat(loopIndicesIn_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_irdy_run_sct(loopIndicesIn_rsci_irdy_run_sct),
      .loopIndicesIn_rsci_ivld(loopIndicesIn_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_idat(loopIndicesIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [79:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [79:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd103),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci (
  clk, arst_n, output_rsc_dat, output_rsc_vld, output_rsc_rdy, run_wen, output_rsci_oswt,
      output_rsci_wen_comp, output_rsci_idat
);
  input clk;
  input arst_n;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input run_wen;
  input output_rsci_oswt;
  output output_rsci_wen_comp;
  input [255:0] output_rsci_idat;


  // Interconnect Declarations
  wire output_rsci_irdy;
  wire output_rsci_biwt;
  wire output_rsci_bdwt;
  wire output_rsci_bcwt;
  wire output_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd102),
  .width(32'sd256)) output_rsci (
      .irdy(output_rsci_irdy),
      .ivld(output_rsci_ivld_run_sct),
      .idat(output_rsci_idat),
      .rdy(output_rsc_rdy),
      .vld(output_rsc_vld),
      .dat(output_rsc_dat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_irdy(output_rsci_irdy),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt),
      .output_rsci_ivld_run_sct(output_rsci_ivld_run_sct)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_output_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_rsci_oswt(output_rsci_oswt),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_biwt(output_rsci_biwt),
      .output_rsci_bdwt(output_rsci_bdwt),
      .output_rsci_bcwt(output_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci (
  clk, arst_n, weight_rsc_dat, weight_rsc_vld, weight_rsc_rdy, run_wen, weight_rsci_oswt,
      weight_rsci_wen_comp, weight_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  input run_wen;
  input weight_rsci_oswt;
  output weight_rsci_wen_comp;
  output [127:0] weight_rsci_idat_mxwt;


  // Interconnect Declarations
  wire weight_rsci_biwt;
  wire weight_rsci_bdwt;
  wire weight_rsci_bcwt;
  wire weight_rsci_irdy_run_sct;
  wire weight_rsci_ivld;
  wire [127:0] weight_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd101),
  .width(32'sd128)) weight_rsci (
      .rdy(weight_rsc_rdy),
      .vld(weight_rsc_vld),
      .dat(weight_rsc_dat),
      .irdy(weight_rsci_irdy_run_sct),
      .ivld(weight_rsci_ivld),
      .idat(weight_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_bcwt(weight_rsci_bcwt),
      .weight_rsci_irdy_run_sct(weight_rsci_irdy_run_sct),
      .weight_rsci_ivld(weight_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_weight_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weight_rsci_oswt(weight_rsci_oswt),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_idat_mxwt(weight_rsci_idat_mxwt),
      .weight_rsci_biwt(weight_rsci_biwt),
      .weight_rsci_bdwt(weight_rsci_bdwt),
      .weight_rsci_bcwt(weight_rsci_bcwt),
      .weight_rsci_idat(weight_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, run_wen, input_rsci_oswt,
      input_rsci_wen_comp, input_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input run_wen;
  input input_rsci_oswt;
  output input_rsci_wen_comp;
  output [127:0] input_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_rsci_biwt;
  wire input_rsci_bdwt;
  wire input_rsci_bcwt;
  wire input_rsci_irdy_run_sct;
  wire input_rsci_ivld;
  wire [127:0] input_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd100),
  .width(32'sd128)) input_rsci (
      .rdy(input_rsc_rdy),
      .vld(input_rsc_vld),
      .dat(input_rsc_dat),
      .irdy(input_rsci_irdy_run_sct),
      .ivld(input_rsci_ivld),
      .idat(input_rsci_idat)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_irdy_run_sct(input_rsci_irdy_run_sct),
      .input_rsci_ivld(input_rsci_ivld)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_input_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsci_oswt(input_rsci_oswt),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt),
      .input_rsci_biwt(input_rsci_biwt),
      .input_rsci_bdwt(input_rsci_bdwt),
      .input_rsci_bcwt(input_rsci_bcwt),
      .input_rsci_idat(input_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy, accumulation_buffer_rsc_0_0_i_radr_d, accumulation_buffer_rsc_0_0_i_wadr_d,
      accumulation_buffer_rsc_0_0_i_d_d, accumulation_buffer_rsc_0_0_i_q_d, accumulation_buffer_rsc_0_1_i_radr_d,
      accumulation_buffer_rsc_0_1_i_wadr_d, accumulation_buffer_rsc_0_1_i_d_d, accumulation_buffer_rsc_0_1_i_q_d,
      accumulation_buffer_rsc_0_2_i_radr_d, accumulation_buffer_rsc_0_2_i_wadr_d,
      accumulation_buffer_rsc_0_2_i_d_d, accumulation_buffer_rsc_0_2_i_q_d, accumulation_buffer_rsc_0_3_i_radr_d,
      accumulation_buffer_rsc_0_3_i_wadr_d, accumulation_buffer_rsc_0_3_i_d_d, accumulation_buffer_rsc_0_3_i_q_d,
      accumulation_buffer_rsc_0_4_i_radr_d, accumulation_buffer_rsc_0_4_i_wadr_d,
      accumulation_buffer_rsc_0_4_i_d_d, accumulation_buffer_rsc_0_4_i_q_d, accumulation_buffer_rsc_0_5_i_radr_d,
      accumulation_buffer_rsc_0_5_i_wadr_d, accumulation_buffer_rsc_0_5_i_d_d, accumulation_buffer_rsc_0_5_i_q_d,
      accumulation_buffer_rsc_0_6_i_radr_d, accumulation_buffer_rsc_0_6_i_wadr_d,
      accumulation_buffer_rsc_0_6_i_d_d, accumulation_buffer_rsc_0_6_i_q_d, accumulation_buffer_rsc_0_7_i_radr_d,
      accumulation_buffer_rsc_0_7_i_wadr_d, accumulation_buffer_rsc_0_7_i_d_d, accumulation_buffer_rsc_0_7_i_q_d,
      accumulation_buffer_rsc_0_8_i_radr_d, accumulation_buffer_rsc_0_8_i_wadr_d,
      accumulation_buffer_rsc_0_8_i_d_d, accumulation_buffer_rsc_0_8_i_q_d, accumulation_buffer_rsc_0_9_i_radr_d,
      accumulation_buffer_rsc_0_9_i_wadr_d, accumulation_buffer_rsc_0_9_i_d_d, accumulation_buffer_rsc_0_9_i_q_d,
      accumulation_buffer_rsc_0_10_i_radr_d, accumulation_buffer_rsc_0_10_i_wadr_d,
      accumulation_buffer_rsc_0_10_i_d_d, accumulation_buffer_rsc_0_10_i_q_d, accumulation_buffer_rsc_0_11_i_radr_d,
      accumulation_buffer_rsc_0_11_i_wadr_d, accumulation_buffer_rsc_0_11_i_d_d,
      accumulation_buffer_rsc_0_11_i_q_d, accumulation_buffer_rsc_0_12_i_radr_d,
      accumulation_buffer_rsc_0_12_i_wadr_d, accumulation_buffer_rsc_0_12_i_d_d,
      accumulation_buffer_rsc_0_12_i_q_d, accumulation_buffer_rsc_0_13_i_radr_d,
      accumulation_buffer_rsc_0_13_i_wadr_d, accumulation_buffer_rsc_0_13_i_d_d,
      accumulation_buffer_rsc_0_13_i_q_d, accumulation_buffer_rsc_0_14_i_radr_d,
      accumulation_buffer_rsc_0_14_i_wadr_d, accumulation_buffer_rsc_0_14_i_d_d,
      accumulation_buffer_rsc_0_14_i_q_d, accumulation_buffer_rsc_0_15_i_radr_d,
      accumulation_buffer_rsc_0_15_i_wadr_d, accumulation_buffer_rsc_0_15_i_d_d,
      accumulation_buffer_rsc_0_15_i_q_d, accumulation_buffer_rsc_0_0_i_we_d_pff,
      accumulation_buffer_rsc_0_0_i_re_d_pff, accumulation_buffer_rsc_0_1_i_we_d_pff,
      accumulation_buffer_rsc_0_1_i_re_d_pff, accumulation_buffer_rsc_0_2_i_we_d_pff,
      accumulation_buffer_rsc_0_2_i_re_d_pff, accumulation_buffer_rsc_0_3_i_we_d_pff,
      accumulation_buffer_rsc_0_3_i_re_d_pff, accumulation_buffer_rsc_0_4_i_we_d_pff,
      accumulation_buffer_rsc_0_4_i_re_d_pff, accumulation_buffer_rsc_0_5_i_we_d_pff,
      accumulation_buffer_rsc_0_5_i_re_d_pff, accumulation_buffer_rsc_0_6_i_we_d_pff,
      accumulation_buffer_rsc_0_6_i_re_d_pff, accumulation_buffer_rsc_0_7_i_we_d_pff,
      accumulation_buffer_rsc_0_7_i_re_d_pff, accumulation_buffer_rsc_0_8_i_we_d_pff,
      accumulation_buffer_rsc_0_8_i_re_d_pff, accumulation_buffer_rsc_0_9_i_we_d_pff,
      accumulation_buffer_rsc_0_9_i_re_d_pff, accumulation_buffer_rsc_0_10_i_we_d_pff,
      accumulation_buffer_rsc_0_10_i_re_d_pff, accumulation_buffer_rsc_0_11_i_we_d_pff,
      accumulation_buffer_rsc_0_11_i_re_d_pff, accumulation_buffer_rsc_0_12_i_we_d_pff,
      accumulation_buffer_rsc_0_12_i_re_d_pff, accumulation_buffer_rsc_0_13_i_we_d_pff,
      accumulation_buffer_rsc_0_13_i_re_d_pff, accumulation_buffer_rsc_0_14_i_we_d_pff,
      accumulation_buffer_rsc_0_14_i_re_d_pff, accumulation_buffer_rsc_0_15_i_we_d_pff,
      accumulation_buffer_rsc_0_15_i_re_d_pff
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  output [7:0] accumulation_buffer_rsc_0_0_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_0_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_0_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_0_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_1_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_1_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_1_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_1_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_2_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_2_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_2_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_2_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_3_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_3_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_3_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_3_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_4_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_4_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_4_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_4_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_5_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_5_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_5_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_5_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_6_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_6_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_6_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_6_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_7_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_7_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_7_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_7_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_8_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_8_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_8_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_8_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_9_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_9_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_9_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_9_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_10_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_10_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_10_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_10_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_11_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_11_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_11_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_11_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_12_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_12_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_12_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_12_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_13_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_13_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_13_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_13_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_14_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_14_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_14_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_14_i_q_d;
  output [7:0] accumulation_buffer_rsc_0_15_i_radr_d;
  output [7:0] accumulation_buffer_rsc_0_15_i_wadr_d;
  output [15:0] accumulation_buffer_rsc_0_15_i_d_d;
  input [15:0] accumulation_buffer_rsc_0_15_i_q_d;
  output accumulation_buffer_rsc_0_0_i_we_d_pff;
  output accumulation_buffer_rsc_0_0_i_re_d_pff;
  output accumulation_buffer_rsc_0_1_i_we_d_pff;
  output accumulation_buffer_rsc_0_1_i_re_d_pff;
  output accumulation_buffer_rsc_0_2_i_we_d_pff;
  output accumulation_buffer_rsc_0_2_i_re_d_pff;
  output accumulation_buffer_rsc_0_3_i_we_d_pff;
  output accumulation_buffer_rsc_0_3_i_re_d_pff;
  output accumulation_buffer_rsc_0_4_i_we_d_pff;
  output accumulation_buffer_rsc_0_4_i_re_d_pff;
  output accumulation_buffer_rsc_0_5_i_we_d_pff;
  output accumulation_buffer_rsc_0_5_i_re_d_pff;
  output accumulation_buffer_rsc_0_6_i_we_d_pff;
  output accumulation_buffer_rsc_0_6_i_re_d_pff;
  output accumulation_buffer_rsc_0_7_i_we_d_pff;
  output accumulation_buffer_rsc_0_7_i_re_d_pff;
  output accumulation_buffer_rsc_0_8_i_we_d_pff;
  output accumulation_buffer_rsc_0_8_i_re_d_pff;
  output accumulation_buffer_rsc_0_9_i_we_d_pff;
  output accumulation_buffer_rsc_0_9_i_re_d_pff;
  output accumulation_buffer_rsc_0_10_i_we_d_pff;
  output accumulation_buffer_rsc_0_10_i_re_d_pff;
  output accumulation_buffer_rsc_0_11_i_we_d_pff;
  output accumulation_buffer_rsc_0_11_i_re_d_pff;
  output accumulation_buffer_rsc_0_12_i_we_d_pff;
  output accumulation_buffer_rsc_0_12_i_re_d_pff;
  output accumulation_buffer_rsc_0_13_i_we_d_pff;
  output accumulation_buffer_rsc_0_13_i_re_d_pff;
  output accumulation_buffer_rsc_0_14_i_we_d_pff;
  output accumulation_buffer_rsc_0_14_i_re_d_pff;
  output accumulation_buffer_rsc_0_15_i_we_d_pff;
  output accumulation_buffer_rsc_0_15_i_re_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire input_rsci_wen_comp;
  wire [127:0] input_rsci_idat_mxwt;
  wire weight_rsci_wen_comp;
  wire [127:0] weight_rsci_idat_mxwt;
  wire output_rsci_wen_comp;
  wire paramsIn_rsci_wen_comp;
  wire [79:0] paramsIn_rsci_idat_mxwt;
  wire loopIndicesIn_rsci_wen_comp;
  wire [47:0] loopIndicesIn_rsci_idat_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_0_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_1_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_2_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_3_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_4_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_5_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_6_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_7_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_8_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_9_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_10_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_11_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_12_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_13_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_14_i_q_d_mxwt;
  wire [15:0] accumulation_buffer_rsc_0_15_i_q_d_mxwt;
  wire [15:0] accum_fifo_15_rsci_output_rsc_z;
  wire accum_fifo_15_rsci_ccs_ccore_en;
  wire [15:0] output_fifo_0_rsci_output_rsc_z;
  wire output_fifo_0_rsci_ccs_ccore_en;
  wire [15:0] accum_fifo_14_rsci_output_rsc_z;
  wire [15:0] output_fifo_1_rsci_output_rsc_z;
  wire [15:0] accum_fifo_13_rsci_output_rsc_z;
  wire [15:0] output_fifo_2_rsci_output_rsc_z;
  wire [15:0] accum_fifo_12_rsci_output_rsc_z;
  wire [15:0] output_fifo_3_rsci_output_rsc_z;
  wire [15:0] accum_fifo_11_rsci_output_rsc_z;
  wire [15:0] output_fifo_4_rsci_output_rsc_z;
  wire [15:0] accum_fifo_10_rsci_output_rsc_z;
  wire [15:0] output_fifo_5_rsci_output_rsc_z;
  wire [15:0] accum_fifo_9_rsci_output_rsc_z;
  wire [15:0] output_fifo_6_rsci_output_rsc_z;
  wire [15:0] accum_fifo_8_rsci_output_rsc_z;
  wire [15:0] output_fifo_7_rsci_output_rsc_z;
  wire [15:0] accum_fifo_7_rsci_output_rsc_z;
  wire [15:0] output_fifo_8_rsci_output_rsc_z;
  wire [15:0] accum_fifo_6_rsci_output_rsc_z;
  wire [15:0] output_fifo_9_rsci_output_rsc_z;
  wire [15:0] accum_fifo_5_rsci_output_rsc_z;
  wire [15:0] output_fifo_10_rsci_output_rsc_z;
  wire [15:0] accum_fifo_4_rsci_output_rsc_z;
  wire [15:0] output_fifo_11_rsci_output_rsc_z;
  wire [15:0] accum_fifo_3_rsci_output_rsc_z;
  wire [15:0] output_fifo_12_rsci_output_rsc_z;
  wire [15:0] accum_fifo_2_rsci_output_rsc_z;
  wire [15:0] output_fifo_13_rsci_output_rsc_z;
  wire [15:0] accum_fifo_1_rsci_output_rsc_z;
  wire [15:0] output_fifo_14_rsci_output_rsc_z;
  wire [7:0] input_fifo_15_rsci_output_rsc_z;
  wire [7:0] input_fifo_14_rsci_output_rsc_z;
  wire [7:0] input_fifo_13_rsci_output_rsc_z;
  wire [7:0] input_fifo_12_rsci_output_rsc_z;
  wire [7:0] input_fifo_11_rsci_output_rsc_z;
  wire [7:0] input_fifo_10_rsci_output_rsc_z;
  wire [7:0] input_fifo_9_rsci_output_rsc_z;
  wire [7:0] input_fifo_8_rsci_output_rsc_z;
  wire [7:0] input_fifo_7_rsci_output_rsc_z;
  wire [7:0] input_fifo_6_rsci_output_rsc_z;
  wire [7:0] input_fifo_5_rsci_output_rsc_z;
  wire [7:0] input_fifo_4_rsci_output_rsc_z;
  wire [7:0] input_fifo_3_rsci_output_rsc_z;
  wire [7:0] input_fifo_2_rsci_output_rsc_z;
  wire [7:0] input_fifo_1_rsci_output_rsc_z;
  wire [7:0] pe_0_0_run_cmp_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_1_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_1_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_2_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_2_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_3_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_3_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_4_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_4_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_5_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_5_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_6_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_6_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_7_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_7_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_8_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_8_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_9_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_9_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_10_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_10_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_11_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_11_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_12_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_12_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_13_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_13_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_14_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_14_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_15_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_15_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_16_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_16_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_17_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_17_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_18_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_18_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_19_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_19_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_20_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_20_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_21_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_21_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_22_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_22_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_23_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_23_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_24_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_24_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_25_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_25_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_26_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_26_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_27_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_27_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_28_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_28_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_29_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_29_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_30_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_30_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_31_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_31_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_32_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_32_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_33_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_33_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_34_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_34_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_35_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_35_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_36_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_36_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_37_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_37_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_38_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_38_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_39_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_39_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_40_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_40_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_41_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_41_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_42_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_42_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_43_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_43_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_44_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_44_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_45_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_45_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_46_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_46_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_47_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_47_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_48_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_48_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_49_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_49_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_50_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_50_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_51_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_51_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_52_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_52_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_53_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_53_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_54_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_54_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_55_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_55_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_56_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_56_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_57_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_57_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_58_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_58_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_59_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_59_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_60_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_60_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_61_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_61_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_62_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_62_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_63_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_63_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_64_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_64_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_65_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_65_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_66_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_66_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_67_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_67_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_68_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_68_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_69_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_69_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_70_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_70_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_71_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_71_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_72_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_72_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_73_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_73_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_74_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_74_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_75_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_75_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_76_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_76_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_77_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_77_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_78_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_78_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_79_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_79_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_80_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_80_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_81_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_81_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_82_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_82_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_83_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_83_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_84_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_84_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_85_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_85_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_86_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_86_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_87_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_87_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_88_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_88_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_89_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_89_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_90_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_90_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_91_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_91_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_92_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_92_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_93_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_93_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_94_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_94_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_95_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_95_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_96_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_96_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_97_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_97_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_98_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_98_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_99_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_99_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_100_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_100_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_101_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_101_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_102_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_102_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_103_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_103_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_104_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_104_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_105_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_105_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_106_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_106_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_107_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_107_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_108_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_108_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_109_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_109_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_110_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_110_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_111_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_111_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_112_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_112_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_113_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_113_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_114_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_114_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_115_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_115_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_116_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_116_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_117_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_117_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_118_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_118_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_119_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_119_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_120_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_120_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_121_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_121_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_122_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_122_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_123_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_123_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_124_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_124_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_125_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_125_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_126_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_126_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_127_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_127_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_128_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_128_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_129_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_129_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_130_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_130_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_131_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_131_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_132_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_132_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_133_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_133_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_134_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_134_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_135_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_135_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_136_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_136_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_137_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_137_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_138_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_138_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_139_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_139_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_140_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_140_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_141_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_141_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_142_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_142_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_143_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_143_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_144_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_144_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_145_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_145_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_146_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_146_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_147_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_147_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_148_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_148_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_149_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_149_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_150_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_150_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_151_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_151_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_152_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_152_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_153_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_153_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_154_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_154_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_155_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_155_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_156_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_156_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_157_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_157_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_158_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_158_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_159_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_159_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_160_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_160_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_161_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_161_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_162_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_162_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_163_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_163_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_164_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_164_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_165_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_165_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_166_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_166_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_167_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_167_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_168_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_168_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_169_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_169_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_170_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_170_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_171_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_171_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_172_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_172_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_173_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_173_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_174_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_174_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_175_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_175_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_176_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_176_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_177_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_177_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_178_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_178_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_179_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_179_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_180_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_180_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_181_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_181_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_182_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_182_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_183_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_183_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_184_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_184_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_185_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_185_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_186_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_186_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_187_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_187_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_188_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_188_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_189_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_189_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_190_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_190_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_191_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_191_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_192_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_192_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_193_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_193_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_194_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_194_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_195_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_195_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_196_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_196_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_197_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_197_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_198_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_198_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_199_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_199_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_200_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_200_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_201_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_201_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_202_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_202_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_203_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_203_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_204_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_204_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_205_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_205_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_206_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_206_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_207_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_207_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_208_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_208_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_209_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_209_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_210_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_210_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_211_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_211_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_212_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_212_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_213_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_213_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_214_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_214_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_215_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_215_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_216_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_216_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_217_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_217_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_218_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_218_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_219_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_219_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_220_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_220_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_221_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_221_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_222_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_222_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_223_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_223_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_224_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_224_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_225_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_225_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_226_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_226_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_227_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_227_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_228_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_228_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_229_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_229_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_230_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_230_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_231_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_231_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_232_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_232_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_233_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_233_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_234_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_234_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_235_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_235_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_236_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_236_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_237_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_237_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_238_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_238_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_239_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_239_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_240_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_240_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_241_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_241_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_242_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_242_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_243_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_243_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_244_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_244_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_245_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_245_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_246_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_246_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_247_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_247_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_248_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_248_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_249_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_249_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_250_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_250_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_251_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_251_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_252_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_252_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_253_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_253_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_254_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_254_psum_out_rsc_z;
  wire [7:0] pe_0_0_run_cmp_255_input_out_rsc_z;
  wire [15:0] pe_0_0_run_cmp_255_psum_out_rsc_z;
  wire [15:0] accum_fifo_0_run_cmp_output_rsc_z;
  wire [15:0] accum_fifo_0_run_cmp_1_output_rsc_z;
  wire [7:0] input_fifo_0_run_cmp_output_rsc_z;
  reg [15:0] output_rsci_idat_255_240;
  reg [15:0] output_rsci_idat_239_224;
  reg [15:0] output_rsci_idat_223_208;
  reg [15:0] output_rsci_idat_207_192;
  reg [15:0] output_rsci_idat_191_176;
  reg [15:0] output_rsci_idat_175_160;
  reg [15:0] output_rsci_idat_159_144;
  reg [15:0] output_rsci_idat_143_128;
  reg [15:0] output_rsci_idat_127_112;
  reg [15:0] output_rsci_idat_111_96;
  reg [15:0] output_rsci_idat_95_80;
  reg [15:0] output_rsci_idat_79_64;
  reg [15:0] output_rsci_idat_63_48;
  reg [15:0] output_rsci_idat_47_32;
  reg [15:0] output_rsci_idat_31_16;
  reg [15:0] output_rsci_idat_15_0;
  wire [1:0] fsm_output;
  wire step_if_2_if_step_if_2_if_nor_1_tmp;
  wire and_dcpl_1;
  wire and_dcpl_4;
  wire or_dcpl_4;
  wire or_dcpl_7;
  wire or_dcpl_8;
  wire or_dcpl_13;
  wire or_dcpl_14;
  wire or_dcpl_17;
  wire or_dcpl_19;
  wire or_dcpl_20;
  wire or_dcpl_23;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_30;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire and_dcpl_10;
  wire and_dcpl_13;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_49;
  wire or_dcpl_50;
  wire or_dcpl_51;
  wire or_dcpl_52;
  wire or_dcpl_53;
  wire or_dcpl_54;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire or_dcpl_58;
  wire or_dcpl_59;
  wire or_dcpl_60;
  wire or_dcpl_61;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire or_dcpl_64;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire or_dcpl_67;
  wire or_dcpl_68;
  wire or_dcpl_69;
  wire or_dcpl_70;
  wire or_dcpl_71;
  wire or_dcpl_72;
  wire and_dcpl_18;
  wire or_dcpl_74;
  wire or_tmp_3;
  wire not_tmp_36;
  wire or_tmp_39;
  wire not_tmp_251;
  wire or_tmp_47;
  wire step_if_for_and_stg_2_7_sva_mx1;
  reg operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
  wire step_if_for_and_stg_2_6_sva_mx1;
  wire step_if_for_and_stg_2_5_sva_mx1;
  wire step_if_for_and_stg_2_4_sva_mx1;
  wire step_if_for_and_stg_2_3_sva_mx1;
  wire step_if_for_and_stg_2_2_sva_mx1;
  wire step_if_for_and_stg_2_1_sva_mx1;
  wire step_if_for_and_stg_2_0_sva_mx1;
  wire step_if_for_and_stg_1_0_sva_1;
  wire step_if_for_and_stg_1_1_sva_1;
  wire step_if_for_and_stg_1_2_sva_1;
  wire step_if_for_and_stg_1_3_sva_1;
  reg [15:0] step_step_lpi_1;
  wire [16:0] nl_step_step_lpi_1;
  reg exitL_exit_step_sva;
  wire [15:0] step_step_lpi_1_dfm_1;
  reg main_stage_0_3;
  reg step_not_mdf_sva_st_1;
  reg main_stage_0_2;
  reg operator_16_false_slc_operator_16_false_acc_16_itm_2;
  reg step_not_mdf_sva_st_2;
  reg operator_16_false_slc_operator_16_false_acc_16_itm_1;
  reg step_if_3_if_step_if_3_if_and_1_itm_3;
  reg operator_16_false_slc_operator_16_false_acc_16_itm_3;
  reg main_stage_0_4;
  reg [3:0] step_step_lpi_1_dfm_1_3_0;
  reg step_if_1_acc_cse_32;
  reg step_and_10_psp;
  reg step_and_128_psp;
  reg step_and_psp;
  reg step_and_144_psp;
  reg step_and_16_psp;
  reg step_and_160_psp;
  reg step_and_32_psp;
  reg step_and_176_psp;
  reg step_and_48_psp;
  reg step_and_192_psp;
  reg step_and_64_psp;
  reg step_and_208_psp;
  reg step_and_80_psp;
  reg step_and_100_psp;
  reg step_and_224_psp;
  reg step_and_96_psp;
  reg step_and_240_psp;
  reg step_and_112_psp;
  wire [47:0] loopIndicesIn_crt_lpi_1_dfm_mx0;
  wire [16:0] operator_16_false_2_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_2_acc_psp_sva_1;
  wire [16:0] operator_16_false_1_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_1_acc_psp_sva_1;
  wire [16:0] operator_16_false_3_acc_psp_sva_1;
  wire [17:0] nl_operator_16_false_3_acc_psp_sva_1;
  reg reg_loopIndicesIn_rsci_oswt_cse;
  wire output_and_cse;
  reg reg_ensig_cgo_303_cse;
  reg reg_ensig_cgo_302_cse;
  reg reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse;
  reg reg_output_rsci_ivld_run_psct_cse;
  reg reg_weight_rsci_irdy_run_psct_cse;
  reg reg_input_rsci_irdy_run_psct_cse;
  wire step_and_241_cse;
  wire [7:0] accumulation_buffer_rsc_0_0_i_radr_d_reg;
  wire and_1019_rmff;
  wire [7:0] accumulation_buffer_rsc_0_0_i_wadr_d_reg;
  wire and_12_rmff;
  wire accumulation_buffer_rsc_0_0_i_we_d_iff;
  wire accumulation_buffer_rsc_0_0_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_1_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_1_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_1_i_we_d_iff;
  wire accumulation_buffer_rsc_0_1_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_2_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_2_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_2_i_we_d_iff;
  wire accumulation_buffer_rsc_0_2_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_3_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_3_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_3_i_we_d_iff;
  wire accumulation_buffer_rsc_0_3_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_4_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_4_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_4_i_we_d_iff;
  wire accumulation_buffer_rsc_0_4_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_5_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_5_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_5_i_we_d_iff;
  wire accumulation_buffer_rsc_0_5_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_6_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_6_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_6_i_we_d_iff;
  wire accumulation_buffer_rsc_0_6_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_7_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_7_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_7_i_we_d_iff;
  wire accumulation_buffer_rsc_0_7_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_8_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_8_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_8_i_we_d_iff;
  wire accumulation_buffer_rsc_0_8_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_9_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_9_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_9_i_we_d_iff;
  wire accumulation_buffer_rsc_0_9_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_10_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_10_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_10_i_we_d_iff;
  wire accumulation_buffer_rsc_0_10_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_11_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_11_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_11_i_we_d_iff;
  wire accumulation_buffer_rsc_0_11_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_12_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_12_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_12_i_we_d_iff;
  wire accumulation_buffer_rsc_0_12_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_13_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_13_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_13_i_we_d_iff;
  wire accumulation_buffer_rsc_0_13_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_14_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_14_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_14_i_we_d_iff;
  wire accumulation_buffer_rsc_0_14_i_re_d_iff;
  wire [7:0] accumulation_buffer_rsc_0_15_i_radr_d_reg;
  wire [7:0] accumulation_buffer_rsc_0_15_i_wadr_d_reg;
  wire accumulation_buffer_rsc_0_15_i_we_d_iff;
  wire accumulation_buffer_rsc_0_15_i_re_d_iff;
  wire and_23_rmff;
  wire and_27_rmff;
  reg [15:0] psum_reg_16_1_sva;
  reg [15:0] psum_reg_16_2_sva;
  reg [15:0] psum_reg_16_3_sva;
  reg [15:0] psum_reg_16_4_sva;
  reg [15:0] psum_reg_16_5_sva;
  reg [15:0] psum_reg_16_6_sva;
  reg [15:0] psum_reg_16_7_sva;
  reg [15:0] psum_reg_16_8_sva;
  reg [15:0] psum_reg_16_9_sva;
  reg [15:0] psum_reg_16_10_sva;
  reg [15:0] psum_reg_16_11_sva;
  reg [15:0] psum_reg_16_12_sva;
  reg [15:0] psum_reg_16_13_sva;
  reg [15:0] psum_reg_16_14_sva;
  reg [15:0] psum_reg_16_15_sva;
  wire [127:0] step_in_col_value_lpi_1_dfm_mx0;
  reg [7:0] step_mux_4_itm_1;
  reg [7:0] input_reg_16_15_sva;
  reg [15:0] psum_reg_15_16_sva;
  reg [7:0] step_mux_259_itm_1;
  reg [7:0] input_reg_15_15_sva;
  reg [15:0] psum_reg_14_16_sva;
  reg [7:0] step_mux_243_itm_1;
  reg [7:0] input_reg_14_15_sva;
  reg [15:0] psum_reg_13_16_sva;
  reg [7:0] step_mux_227_itm_1;
  reg [7:0] input_reg_13_15_sva;
  reg [15:0] psum_reg_12_16_sva;
  reg [7:0] step_mux_211_itm_1;
  reg [7:0] input_reg_12_15_sva;
  reg [15:0] psum_reg_11_16_sva;
  reg [7:0] step_mux_195_itm_1;
  reg [7:0] input_reg_11_15_sva;
  reg [15:0] psum_reg_10_16_sva;
  reg [7:0] step_mux_179_itm_1;
  reg [7:0] input_reg_10_15_sva;
  reg [15:0] psum_reg_9_16_sva;
  reg [7:0] step_mux_163_itm_1;
  reg [7:0] input_reg_9_15_sva;
  reg [15:0] psum_reg_8_16_sva;
  reg [7:0] step_mux_147_itm_1;
  reg [7:0] input_reg_8_15_sva;
  reg [15:0] psum_reg_7_16_sva;
  reg [7:0] step_mux_131_itm_1;
  reg [7:0] input_reg_7_15_sva;
  reg [15:0] psum_reg_6_16_sva;
  reg [7:0] step_mux_115_itm_1;
  reg [7:0] input_reg_6_15_sva;
  reg [15:0] psum_reg_5_16_sva;
  reg [7:0] step_mux_99_itm_1;
  reg [7:0] input_reg_5_15_sva;
  reg [15:0] psum_reg_4_16_sva;
  reg [7:0] step_mux_83_itm_1;
  reg [7:0] input_reg_4_15_sva;
  reg [15:0] psum_reg_3_16_sva;
  reg [7:0] step_mux_67_itm_1;
  reg [7:0] input_reg_3_15_sva;
  reg [15:0] psum_reg_2_16_sva;
  reg [7:0] step_mux_51_itm_1;
  reg [7:0] input_reg_2_15_sva;
  reg [15:0] psum_reg_1_16_sva;
  reg [7:0] step_mux_35_itm_1;
  reg [7:0] input_reg_1_15_sva;
  reg [7:0] step_mux_19_itm_1;
  reg [7:0] input_reg_16_14_sva;
  reg [15:0] psum_reg_15_15_sva;
  reg [7:0] step_mux_258_itm_1;
  reg [7:0] input_reg_15_14_sva;
  reg [15:0] psum_reg_14_15_sva;
  reg [7:0] step_mux_242_itm_1;
  reg [7:0] input_reg_14_14_sva;
  reg [15:0] psum_reg_13_15_sva;
  reg [7:0] step_mux_226_itm_1;
  reg [7:0] input_reg_13_14_sva;
  reg [15:0] psum_reg_12_15_sva;
  reg [7:0] step_mux_210_itm_1;
  reg [7:0] input_reg_12_14_sva;
  reg [15:0] psum_reg_11_15_sva;
  reg [7:0] step_mux_194_itm_1;
  reg [7:0] input_reg_11_14_sva;
  reg [15:0] psum_reg_10_15_sva;
  reg [7:0] step_mux_178_itm_1;
  reg [7:0] input_reg_10_14_sva;
  reg [15:0] psum_reg_9_15_sva;
  reg [7:0] step_mux_162_itm_1;
  reg [7:0] input_reg_9_14_sva;
  reg [15:0] psum_reg_8_15_sva;
  reg [7:0] step_mux_146_itm_1;
  reg [7:0] input_reg_8_14_sva;
  reg [15:0] psum_reg_7_15_sva;
  reg [7:0] step_mux_130_itm_1;
  reg [7:0] input_reg_7_14_sva;
  reg [15:0] psum_reg_6_15_sva;
  reg [7:0] step_mux_114_itm_1;
  reg [7:0] input_reg_6_14_sva;
  reg [15:0] psum_reg_5_15_sva;
  reg [7:0] step_mux_98_itm_1;
  reg [7:0] input_reg_5_14_sva;
  reg [15:0] psum_reg_4_15_sva;
  reg [7:0] step_mux_82_itm_1;
  reg [7:0] input_reg_4_14_sva;
  reg [15:0] psum_reg_3_15_sva;
  reg [7:0] step_mux_66_itm_1;
  reg [7:0] input_reg_3_14_sva;
  reg [15:0] psum_reg_2_15_sva;
  reg [7:0] step_mux_50_itm_1;
  reg [7:0] input_reg_2_14_sva;
  reg [15:0] psum_reg_1_15_sva;
  reg [7:0] step_mux_34_itm_1;
  reg [7:0] input_reg_1_14_sva;
  reg [7:0] step_mux_18_itm_1;
  reg [7:0] input_reg_16_13_sva;
  reg [15:0] psum_reg_15_14_sva;
  reg [7:0] step_mux_257_itm_1;
  reg [7:0] input_reg_15_13_sva;
  reg [15:0] psum_reg_14_14_sva;
  reg [7:0] step_mux_241_itm_1;
  reg [7:0] input_reg_14_13_sva;
  reg [15:0] psum_reg_13_14_sva;
  reg [7:0] step_mux_225_itm_1;
  reg [7:0] input_reg_13_13_sva;
  reg [15:0] psum_reg_12_14_sva;
  reg [7:0] step_mux_209_itm_1;
  reg [7:0] input_reg_12_13_sva;
  reg [15:0] psum_reg_11_14_sva;
  reg [7:0] step_mux_193_itm_1;
  reg [7:0] input_reg_11_13_sva;
  reg [15:0] psum_reg_10_14_sva;
  reg [7:0] step_mux_177_itm_1;
  reg [7:0] input_reg_10_13_sva;
  reg [15:0] psum_reg_9_14_sva;
  reg [7:0] step_mux_161_itm_1;
  reg [7:0] input_reg_9_13_sva;
  reg [15:0] psum_reg_8_14_sva;
  reg [7:0] step_mux_145_itm_1;
  reg [7:0] input_reg_8_13_sva;
  reg [15:0] psum_reg_7_14_sva;
  reg [7:0] step_mux_129_itm_1;
  reg [7:0] input_reg_7_13_sva;
  reg [15:0] psum_reg_6_14_sva;
  reg [7:0] step_mux_113_itm_1;
  reg [7:0] input_reg_6_13_sva;
  reg [15:0] psum_reg_5_14_sva;
  reg [7:0] step_mux_97_itm_1;
  reg [7:0] input_reg_5_13_sva;
  reg [15:0] psum_reg_4_14_sva;
  reg [7:0] step_mux_81_itm_1;
  reg [7:0] input_reg_4_13_sva;
  reg [15:0] psum_reg_3_14_sva;
  reg [7:0] step_mux_65_itm_1;
  reg [7:0] input_reg_3_13_sva;
  reg [15:0] psum_reg_2_14_sva;
  reg [7:0] step_mux_49_itm_1;
  reg [7:0] input_reg_2_13_sva;
  reg [15:0] psum_reg_1_14_sva;
  reg [7:0] step_mux_33_itm_1;
  reg [7:0] input_reg_1_13_sva;
  reg [7:0] step_mux_17_itm_1;
  reg [7:0] input_reg_16_12_sva;
  reg [15:0] psum_reg_15_13_sva;
  reg [7:0] step_mux_256_itm_1;
  reg [7:0] input_reg_15_12_sva;
  reg [15:0] psum_reg_14_13_sva;
  reg [7:0] step_mux_240_itm_1;
  reg [7:0] input_reg_14_12_sva;
  reg [15:0] psum_reg_13_13_sva;
  reg [7:0] step_mux_224_itm_1;
  reg [7:0] input_reg_13_12_sva;
  reg [15:0] psum_reg_12_13_sva;
  reg [7:0] step_mux_208_itm_1;
  reg [7:0] input_reg_12_12_sva;
  reg [15:0] psum_reg_11_13_sva;
  reg [7:0] step_mux_192_itm_1;
  reg [7:0] input_reg_11_12_sva;
  reg [15:0] psum_reg_10_13_sva;
  reg [7:0] step_mux_176_itm_1;
  reg [7:0] input_reg_10_12_sva;
  reg [15:0] psum_reg_9_13_sva;
  reg [7:0] step_mux_160_itm_1;
  reg [7:0] input_reg_9_12_sva;
  reg [15:0] psum_reg_8_13_sva;
  reg [7:0] step_mux_144_itm_1;
  reg [7:0] input_reg_8_12_sva;
  reg [15:0] psum_reg_7_13_sva;
  reg [7:0] step_mux_128_itm_1;
  reg [7:0] input_reg_7_12_sva;
  reg [15:0] psum_reg_6_13_sva;
  reg [7:0] step_mux_112_itm_1;
  reg [7:0] input_reg_6_12_sva;
  reg [15:0] psum_reg_5_13_sva;
  reg [7:0] step_mux_96_itm_1;
  reg [7:0] input_reg_5_12_sva;
  reg [15:0] psum_reg_4_13_sva;
  reg [7:0] step_mux_80_itm_1;
  reg [7:0] input_reg_4_12_sva;
  reg [15:0] psum_reg_3_13_sva;
  reg [7:0] step_mux_64_itm_1;
  reg [7:0] input_reg_3_12_sva;
  reg [15:0] psum_reg_2_13_sva;
  reg [7:0] step_mux_48_itm_1;
  reg [7:0] input_reg_2_12_sva;
  reg [15:0] psum_reg_1_13_sva;
  reg [7:0] step_mux_32_itm_1;
  reg [7:0] input_reg_1_12_sva;
  reg [7:0] step_mux_16_itm_1;
  reg [7:0] input_reg_16_11_sva;
  reg [15:0] psum_reg_15_12_sva;
  reg [7:0] step_mux_255_itm_1;
  reg [7:0] input_reg_15_11_sva;
  reg [15:0] psum_reg_14_12_sva;
  reg [7:0] step_mux_239_itm_1;
  reg [7:0] input_reg_14_11_sva;
  reg [15:0] psum_reg_13_12_sva;
  reg [7:0] step_mux_223_itm_1;
  reg [7:0] input_reg_13_11_sva;
  reg [15:0] psum_reg_12_12_sva;
  reg [7:0] step_mux_207_itm_1;
  reg [7:0] input_reg_12_11_sva;
  reg [15:0] psum_reg_11_12_sva;
  reg [7:0] step_mux_191_itm_1;
  reg [7:0] input_reg_11_11_sva;
  reg [15:0] psum_reg_10_12_sva;
  reg [7:0] step_mux_175_itm_1;
  reg [7:0] input_reg_10_11_sva;
  reg [15:0] psum_reg_9_12_sva;
  reg [7:0] step_mux_159_itm_1;
  reg [7:0] input_reg_9_11_sva;
  reg [15:0] psum_reg_8_12_sva;
  reg [7:0] step_mux_143_itm_1;
  reg [7:0] input_reg_8_11_sva;
  reg [15:0] psum_reg_7_12_sva;
  reg [7:0] step_mux_127_itm_1;
  reg [7:0] input_reg_7_11_sva;
  reg [15:0] psum_reg_6_12_sva;
  reg [7:0] step_mux_111_itm_1;
  reg [7:0] input_reg_6_11_sva;
  reg [15:0] psum_reg_5_12_sva;
  reg [7:0] step_mux_95_itm_1;
  reg [7:0] input_reg_5_11_sva;
  reg [15:0] psum_reg_4_12_sva;
  reg [7:0] step_mux_79_itm_1;
  reg [7:0] input_reg_4_11_sva;
  reg [15:0] psum_reg_3_12_sva;
  reg [7:0] step_mux_63_itm_1;
  reg [7:0] input_reg_3_11_sva;
  reg [15:0] psum_reg_2_12_sva;
  reg [7:0] step_mux_47_itm_1;
  reg [7:0] input_reg_2_11_sva;
  reg [15:0] psum_reg_1_12_sva;
  reg [7:0] step_mux_31_itm_1;
  reg [7:0] input_reg_1_11_sva;
  reg [7:0] step_mux_15_itm_1;
  reg [7:0] input_reg_16_10_sva;
  reg [15:0] psum_reg_15_11_sva;
  reg [7:0] step_mux_254_itm_1;
  reg [7:0] input_reg_15_10_sva;
  reg [15:0] psum_reg_14_11_sva;
  reg [7:0] step_mux_238_itm_1;
  reg [7:0] input_reg_14_10_sva;
  reg [15:0] psum_reg_13_11_sva;
  reg [7:0] step_mux_222_itm_1;
  reg [7:0] input_reg_13_10_sva;
  reg [15:0] psum_reg_12_11_sva;
  reg [7:0] step_mux_206_itm_1;
  reg [7:0] input_reg_12_10_sva;
  reg [15:0] psum_reg_11_11_sva;
  reg [7:0] step_mux_190_itm_1;
  reg [7:0] input_reg_11_10_sva;
  reg [15:0] psum_reg_10_11_sva;
  reg [7:0] step_mux_174_itm_1;
  reg [7:0] input_reg_10_10_sva;
  reg [15:0] psum_reg_9_11_sva;
  reg [7:0] step_mux_158_itm_1;
  reg [7:0] input_reg_9_10_sva;
  reg [15:0] psum_reg_8_11_sva;
  reg [7:0] step_mux_142_itm_1;
  reg [7:0] input_reg_8_10_sva;
  reg [15:0] psum_reg_7_11_sva;
  reg [7:0] step_mux_126_itm_1;
  reg [7:0] input_reg_7_10_sva;
  reg [15:0] psum_reg_6_11_sva;
  reg [7:0] step_mux_110_itm_1;
  reg [7:0] input_reg_6_10_sva;
  reg [15:0] psum_reg_5_11_sva;
  reg [7:0] step_mux_94_itm_1;
  reg [7:0] input_reg_5_10_sva;
  reg [15:0] psum_reg_4_11_sva;
  reg [7:0] step_mux_78_itm_1;
  reg [7:0] input_reg_4_10_sva;
  reg [15:0] psum_reg_3_11_sva;
  reg [7:0] step_mux_62_itm_1;
  reg [7:0] input_reg_3_10_sva;
  reg [15:0] psum_reg_2_11_sva;
  reg [7:0] step_mux_46_itm_1;
  reg [7:0] input_reg_2_10_sva;
  reg [15:0] psum_reg_1_11_sva;
  reg [7:0] step_mux_30_itm_1;
  reg [7:0] input_reg_1_10_sva;
  reg [7:0] step_mux_14_itm_1;
  reg [7:0] input_reg_16_9_sva;
  reg [15:0] psum_reg_15_10_sva;
  reg [7:0] step_mux_253_itm_1;
  reg [7:0] input_reg_15_9_sva;
  reg [15:0] psum_reg_14_10_sva;
  reg [7:0] step_mux_237_itm_1;
  reg [7:0] input_reg_14_9_sva;
  reg [15:0] psum_reg_13_10_sva;
  reg [7:0] step_mux_221_itm_1;
  reg [7:0] input_reg_13_9_sva;
  reg [15:0] psum_reg_12_10_sva;
  reg [7:0] step_mux_205_itm_1;
  reg [7:0] input_reg_12_9_sva;
  reg [15:0] psum_reg_11_10_sva;
  reg [7:0] step_mux_189_itm_1;
  reg [7:0] input_reg_11_9_sva;
  reg [15:0] psum_reg_10_10_sva;
  reg [7:0] step_mux_173_itm_1;
  reg [7:0] input_reg_10_9_sva;
  reg [15:0] psum_reg_9_10_sva;
  reg [7:0] step_mux_157_itm_1;
  reg [7:0] input_reg_9_9_sva;
  reg [15:0] psum_reg_8_10_sva;
  reg [7:0] step_mux_141_itm_1;
  reg [7:0] input_reg_8_9_sva;
  reg [15:0] psum_reg_7_10_sva;
  reg [7:0] step_mux_125_itm_1;
  reg [7:0] input_reg_7_9_sva;
  reg [15:0] psum_reg_6_10_sva;
  reg [7:0] step_mux_109_itm_1;
  reg [7:0] input_reg_6_9_sva;
  reg [15:0] psum_reg_5_10_sva;
  reg [7:0] step_mux_93_itm_1;
  reg [7:0] input_reg_5_9_sva;
  reg [15:0] psum_reg_4_10_sva;
  reg [7:0] step_mux_77_itm_1;
  reg [7:0] input_reg_4_9_sva;
  reg [15:0] psum_reg_3_10_sva;
  reg [7:0] step_mux_61_itm_1;
  reg [7:0] input_reg_3_9_sva;
  reg [15:0] psum_reg_2_10_sva;
  reg [7:0] step_mux_45_itm_1;
  reg [7:0] input_reg_2_9_sva;
  reg [15:0] psum_reg_1_10_sva;
  reg [7:0] step_mux_29_itm_1;
  reg [7:0] input_reg_1_9_sva;
  reg [7:0] step_mux_13_itm_1;
  reg [7:0] input_reg_16_8_sva;
  reg [15:0] psum_reg_15_9_sva;
  reg [7:0] step_mux_252_itm_1;
  reg [7:0] input_reg_15_8_sva;
  reg [15:0] psum_reg_14_9_sva;
  reg [7:0] step_mux_236_itm_1;
  reg [7:0] input_reg_14_8_sva;
  reg [15:0] psum_reg_13_9_sva;
  reg [7:0] step_mux_220_itm_1;
  reg [7:0] input_reg_13_8_sva;
  reg [15:0] psum_reg_12_9_sva;
  reg [7:0] step_mux_204_itm_1;
  reg [7:0] input_reg_12_8_sva;
  reg [15:0] psum_reg_11_9_sva;
  reg [7:0] step_mux_188_itm_1;
  reg [7:0] input_reg_11_8_sva;
  reg [15:0] psum_reg_10_9_sva;
  reg [7:0] step_mux_172_itm_1;
  reg [7:0] input_reg_10_8_sva;
  reg [15:0] psum_reg_9_9_sva;
  reg [7:0] step_mux_156_itm_1;
  reg [7:0] input_reg_9_8_sva;
  reg [15:0] psum_reg_8_9_sva;
  reg [7:0] step_mux_140_itm_1;
  reg [7:0] input_reg_8_8_sva;
  reg [15:0] psum_reg_7_9_sva;
  reg [7:0] step_mux_124_itm_1;
  reg [7:0] input_reg_7_8_sva;
  reg [15:0] psum_reg_6_9_sva;
  reg [7:0] step_mux_108_itm_1;
  reg [7:0] input_reg_6_8_sva;
  reg [15:0] psum_reg_5_9_sva;
  reg [7:0] step_mux_92_itm_1;
  reg [7:0] input_reg_5_8_sva;
  reg [15:0] psum_reg_4_9_sva;
  reg [7:0] step_mux_76_itm_1;
  reg [7:0] input_reg_4_8_sva;
  reg [15:0] psum_reg_3_9_sva;
  reg [7:0] step_mux_60_itm_1;
  reg [7:0] input_reg_3_8_sva;
  reg [15:0] psum_reg_2_9_sva;
  reg [7:0] step_mux_44_itm_1;
  reg [7:0] input_reg_2_8_sva;
  reg [15:0] psum_reg_1_9_sva;
  reg [7:0] step_mux_28_itm_1;
  reg [7:0] input_reg_1_8_sva;
  reg [7:0] step_mux_12_itm_1;
  reg [7:0] input_reg_16_7_sva;
  reg [15:0] psum_reg_15_8_sva;
  reg [7:0] step_mux_251_itm_1;
  reg [7:0] input_reg_15_7_sva;
  reg [15:0] psum_reg_14_8_sva;
  reg [7:0] step_mux_235_itm_1;
  reg [7:0] input_reg_14_7_sva;
  reg [15:0] psum_reg_13_8_sva;
  reg [7:0] step_mux_219_itm_1;
  reg [7:0] input_reg_13_7_sva;
  reg [15:0] psum_reg_12_8_sva;
  reg [7:0] step_mux_203_itm_1;
  reg [7:0] input_reg_12_7_sva;
  reg [15:0] psum_reg_11_8_sva;
  reg [7:0] step_mux_187_itm_1;
  reg [7:0] input_reg_11_7_sva;
  reg [15:0] psum_reg_10_8_sva;
  reg [7:0] step_mux_171_itm_1;
  reg [7:0] input_reg_10_7_sva;
  reg [15:0] psum_reg_9_8_sva;
  reg [7:0] step_mux_155_itm_1;
  reg [7:0] input_reg_9_7_sva;
  reg [15:0] psum_reg_8_8_sva;
  reg [7:0] step_mux_139_itm_1;
  reg [7:0] input_reg_8_7_sva;
  reg [15:0] psum_reg_7_8_sva;
  reg [7:0] step_mux_123_itm_1;
  reg [7:0] input_reg_7_7_sva;
  reg [15:0] psum_reg_6_8_sva;
  reg [7:0] step_mux_107_itm_1;
  reg [7:0] input_reg_6_7_sva;
  reg [15:0] psum_reg_5_8_sva;
  reg [7:0] step_mux_91_itm_1;
  reg [7:0] input_reg_5_7_sva;
  reg [15:0] psum_reg_4_8_sva;
  reg [7:0] step_mux_75_itm_1;
  reg [7:0] input_reg_4_7_sva;
  reg [15:0] psum_reg_3_8_sva;
  reg [7:0] step_mux_59_itm_1;
  reg [7:0] input_reg_3_7_sva;
  reg [15:0] psum_reg_2_8_sva;
  reg [7:0] step_mux_43_itm_1;
  reg [7:0] input_reg_2_7_sva;
  reg [15:0] psum_reg_1_8_sva;
  reg [7:0] step_mux_27_itm_1;
  reg [7:0] input_reg_1_7_sva;
  reg [7:0] step_mux_11_itm_1;
  reg [7:0] input_reg_16_6_sva;
  reg [15:0] psum_reg_15_7_sva;
  reg [7:0] step_mux_250_itm_1;
  reg [7:0] input_reg_15_6_sva;
  reg [15:0] psum_reg_14_7_sva;
  reg [7:0] step_mux_234_itm_1;
  reg [7:0] input_reg_14_6_sva;
  reg [15:0] psum_reg_13_7_sva;
  reg [7:0] step_mux_218_itm_1;
  reg [7:0] input_reg_13_6_sva;
  reg [15:0] psum_reg_12_7_sva;
  reg [7:0] step_mux_202_itm_1;
  reg [7:0] input_reg_12_6_sva;
  reg [15:0] psum_reg_11_7_sva;
  reg [7:0] step_mux_186_itm_1;
  reg [7:0] input_reg_11_6_sva;
  reg [15:0] psum_reg_10_7_sva;
  reg [7:0] step_mux_170_itm_1;
  reg [7:0] input_reg_10_6_sva;
  reg [15:0] psum_reg_9_7_sva;
  reg [7:0] step_mux_154_itm_1;
  reg [7:0] input_reg_9_6_sva;
  reg [15:0] psum_reg_8_7_sva;
  reg [7:0] step_mux_138_itm_1;
  reg [7:0] input_reg_8_6_sva;
  reg [15:0] psum_reg_7_7_sva;
  reg [7:0] step_mux_122_itm_1;
  reg [7:0] input_reg_7_6_sva;
  reg [15:0] psum_reg_6_7_sva;
  reg [7:0] step_mux_106_itm_1;
  reg [7:0] input_reg_6_6_sva;
  reg [15:0] psum_reg_5_7_sva;
  reg [7:0] step_mux_90_itm_1;
  reg [7:0] input_reg_5_6_sva;
  reg [15:0] psum_reg_4_7_sva;
  reg [7:0] step_mux_74_itm_1;
  reg [7:0] input_reg_4_6_sva;
  reg [15:0] psum_reg_3_7_sva;
  reg [7:0] step_mux_58_itm_1;
  reg [7:0] input_reg_3_6_sva;
  reg [15:0] psum_reg_2_7_sva;
  reg [7:0] step_mux_42_itm_1;
  reg [7:0] input_reg_2_6_sva;
  reg [15:0] psum_reg_1_7_sva;
  reg [7:0] step_mux_26_itm_1;
  reg [7:0] input_reg_1_6_sva;
  reg [7:0] step_mux_10_itm_1;
  reg [7:0] input_reg_16_5_sva;
  reg [15:0] psum_reg_15_6_sva;
  reg [7:0] step_mux_249_itm_1;
  reg [7:0] input_reg_15_5_sva;
  reg [15:0] psum_reg_14_6_sva;
  reg [7:0] step_mux_233_itm_1;
  reg [7:0] input_reg_14_5_sva;
  reg [15:0] psum_reg_13_6_sva;
  reg [7:0] step_mux_217_itm_1;
  reg [7:0] input_reg_13_5_sva;
  reg [15:0] psum_reg_12_6_sva;
  reg [7:0] step_mux_201_itm_1;
  reg [7:0] input_reg_12_5_sva;
  reg [15:0] psum_reg_11_6_sva;
  reg [7:0] step_mux_185_itm_1;
  reg [7:0] input_reg_11_5_sva;
  reg [15:0] psum_reg_10_6_sva;
  reg [7:0] step_mux_169_itm_1;
  reg [7:0] input_reg_10_5_sva;
  reg [15:0] psum_reg_9_6_sva;
  reg [7:0] step_mux_153_itm_1;
  reg [7:0] input_reg_9_5_sva;
  reg [15:0] psum_reg_8_6_sva;
  reg [7:0] step_mux_137_itm_1;
  reg [7:0] input_reg_8_5_sva;
  reg [15:0] psum_reg_7_6_sva;
  reg [7:0] step_mux_121_itm_1;
  reg [7:0] input_reg_7_5_sva;
  reg [15:0] psum_reg_6_6_sva;
  reg [7:0] step_mux_105_itm_1;
  reg [7:0] input_reg_6_5_sva;
  reg [15:0] psum_reg_5_6_sva;
  reg [7:0] step_mux_89_itm_1;
  reg [7:0] input_reg_5_5_sva;
  reg [15:0] psum_reg_4_6_sva;
  reg [7:0] step_mux_73_itm_1;
  reg [7:0] input_reg_4_5_sva;
  reg [15:0] psum_reg_3_6_sva;
  reg [7:0] step_mux_57_itm_1;
  reg [7:0] input_reg_3_5_sva;
  reg [15:0] psum_reg_2_6_sva;
  reg [7:0] step_mux_41_itm_1;
  reg [7:0] input_reg_2_5_sva;
  reg [15:0] psum_reg_1_6_sva;
  reg [7:0] step_mux_25_itm_1;
  reg [7:0] input_reg_1_5_sva;
  reg [7:0] step_mux_9_itm_1;
  reg [7:0] input_reg_16_4_sva;
  reg [15:0] psum_reg_15_5_sva;
  reg [7:0] step_mux_248_itm_1;
  reg [7:0] input_reg_15_4_sva;
  reg [15:0] psum_reg_14_5_sva;
  reg [7:0] step_mux_232_itm_1;
  reg [7:0] input_reg_14_4_sva;
  reg [15:0] psum_reg_13_5_sva;
  reg [7:0] step_mux_216_itm_1;
  reg [7:0] input_reg_13_4_sva;
  reg [15:0] psum_reg_12_5_sva;
  reg [7:0] step_mux_200_itm_1;
  reg [7:0] input_reg_12_4_sva;
  reg [15:0] psum_reg_11_5_sva;
  reg [7:0] step_mux_184_itm_1;
  reg [7:0] input_reg_11_4_sva;
  reg [15:0] psum_reg_10_5_sva;
  reg [7:0] step_mux_168_itm_1;
  reg [7:0] input_reg_10_4_sva;
  reg [15:0] psum_reg_9_5_sva;
  reg [7:0] step_mux_152_itm_1;
  reg [7:0] input_reg_9_4_sva;
  reg [15:0] psum_reg_8_5_sva;
  reg [7:0] step_mux_136_itm_1;
  reg [7:0] input_reg_8_4_sva;
  reg [15:0] psum_reg_7_5_sva;
  reg [7:0] step_mux_120_itm_1;
  reg [7:0] input_reg_7_4_sva;
  reg [15:0] psum_reg_6_5_sva;
  reg [7:0] step_mux_104_itm_1;
  reg [7:0] input_reg_6_4_sva;
  reg [15:0] psum_reg_5_5_sva;
  reg [7:0] step_mux_88_itm_1;
  reg [7:0] input_reg_5_4_sva;
  reg [15:0] psum_reg_4_5_sva;
  reg [7:0] step_mux_72_itm_1;
  reg [7:0] input_reg_4_4_sva;
  reg [15:0] psum_reg_3_5_sva;
  reg [7:0] step_mux_56_itm_1;
  reg [7:0] input_reg_3_4_sva;
  reg [15:0] psum_reg_2_5_sva;
  reg [7:0] step_mux_40_itm_1;
  reg [7:0] input_reg_2_4_sva;
  reg [15:0] psum_reg_1_5_sva;
  reg [7:0] step_mux_24_itm_1;
  reg [7:0] input_reg_1_4_sva;
  reg [7:0] step_mux_8_itm_1;
  reg [7:0] input_reg_16_3_sva;
  reg [15:0] psum_reg_15_4_sva;
  reg [7:0] step_mux_247_itm_1;
  reg [7:0] input_reg_15_3_sva;
  reg [15:0] psum_reg_14_4_sva;
  reg [7:0] step_mux_231_itm_1;
  reg [7:0] input_reg_14_3_sva;
  reg [15:0] psum_reg_13_4_sva;
  reg [7:0] step_mux_215_itm_1;
  reg [7:0] input_reg_13_3_sva;
  reg [15:0] psum_reg_12_4_sva;
  reg [7:0] step_mux_199_itm_1;
  reg [7:0] input_reg_12_3_sva;
  reg [15:0] psum_reg_11_4_sva;
  reg [7:0] step_mux_183_itm_1;
  reg [7:0] input_reg_11_3_sva;
  reg [15:0] psum_reg_10_4_sva;
  reg [7:0] step_mux_167_itm_1;
  reg [7:0] input_reg_10_3_sva;
  reg [15:0] psum_reg_9_4_sva;
  reg [7:0] step_mux_151_itm_1;
  reg [7:0] input_reg_9_3_sva;
  reg [15:0] psum_reg_8_4_sva;
  reg [7:0] step_mux_135_itm_1;
  reg [7:0] input_reg_8_3_sva;
  reg [15:0] psum_reg_7_4_sva;
  reg [7:0] step_mux_119_itm_1;
  reg [7:0] input_reg_7_3_sva;
  reg [15:0] psum_reg_6_4_sva;
  reg [7:0] step_mux_103_itm_1;
  reg [7:0] input_reg_6_3_sva;
  reg [15:0] psum_reg_5_4_sva;
  reg [7:0] step_mux_87_itm_1;
  reg [7:0] input_reg_5_3_sva;
  reg [15:0] psum_reg_4_4_sva;
  reg [7:0] step_mux_71_itm_1;
  reg [7:0] input_reg_4_3_sva;
  reg [15:0] psum_reg_3_4_sva;
  reg [7:0] step_mux_55_itm_1;
  reg [7:0] input_reg_3_3_sva;
  reg [15:0] psum_reg_2_4_sva;
  reg [7:0] step_mux_39_itm_1;
  reg [7:0] input_reg_2_3_sva;
  reg [15:0] psum_reg_1_4_sva;
  reg [7:0] step_mux_23_itm_1;
  reg [7:0] input_reg_1_3_sva;
  reg [7:0] step_mux_7_itm_1;
  reg [7:0] input_reg_16_2_sva;
  reg [15:0] psum_reg_15_3_sva;
  reg [7:0] step_mux_246_itm_1;
  reg [7:0] input_reg_15_2_sva;
  reg [15:0] psum_reg_14_3_sva;
  reg [7:0] step_mux_230_itm_1;
  reg [7:0] input_reg_14_2_sva;
  reg [15:0] psum_reg_13_3_sva;
  reg [7:0] step_mux_214_itm_1;
  reg [7:0] input_reg_13_2_sva;
  reg [15:0] psum_reg_12_3_sva;
  reg [7:0] step_mux_198_itm_1;
  reg [7:0] input_reg_12_2_sva;
  reg [15:0] psum_reg_11_3_sva;
  reg [7:0] step_mux_182_itm_1;
  reg [7:0] input_reg_11_2_sva;
  reg [15:0] psum_reg_10_3_sva;
  reg [7:0] step_mux_166_itm_1;
  reg [7:0] input_reg_10_2_sva;
  reg [15:0] psum_reg_9_3_sva;
  reg [7:0] step_mux_150_itm_1;
  reg [7:0] input_reg_9_2_sva;
  reg [15:0] psum_reg_8_3_sva;
  reg [7:0] step_mux_134_itm_1;
  reg [7:0] input_reg_8_2_sva;
  reg [15:0] psum_reg_7_3_sva;
  reg [7:0] step_mux_118_itm_1;
  reg [7:0] input_reg_7_2_sva;
  reg [15:0] psum_reg_6_3_sva;
  reg [7:0] step_mux_102_itm_1;
  reg [7:0] input_reg_6_2_sva;
  reg [15:0] psum_reg_5_3_sva;
  reg [7:0] step_mux_86_itm_1;
  reg [7:0] input_reg_5_2_sva;
  reg [15:0] psum_reg_4_3_sva;
  reg [7:0] step_mux_70_itm_1;
  reg [7:0] input_reg_4_2_sva;
  reg [15:0] psum_reg_3_3_sva;
  reg [7:0] step_mux_54_itm_1;
  reg [7:0] input_reg_3_2_sva;
  reg [15:0] psum_reg_2_3_sva;
  reg [7:0] step_mux_38_itm_1;
  reg [7:0] input_reg_2_2_sva;
  reg [15:0] psum_reg_1_3_sva;
  reg [7:0] step_mux_22_itm_1;
  reg [7:0] input_reg_1_2_sva;
  reg [7:0] step_mux_6_itm_1;
  reg [7:0] input_reg_16_1_sva;
  reg [15:0] psum_reg_15_2_sva;
  reg [7:0] step_mux_245_itm_1;
  reg [7:0] input_reg_15_1_sva;
  reg [15:0] psum_reg_14_2_sva;
  reg [7:0] step_mux_229_itm_1;
  reg [7:0] input_reg_14_1_sva;
  reg [15:0] psum_reg_13_2_sva;
  reg [7:0] step_mux_213_itm_1;
  reg [7:0] input_reg_13_1_sva;
  reg [15:0] psum_reg_12_2_sva;
  reg [7:0] step_mux_197_itm_1;
  reg [7:0] input_reg_12_1_sva;
  reg [15:0] psum_reg_11_2_sva;
  reg [7:0] step_mux_181_itm_1;
  reg [7:0] input_reg_11_1_sva;
  reg [15:0] psum_reg_10_2_sva;
  reg [7:0] step_mux_165_itm_1;
  reg [7:0] input_reg_10_1_sva;
  reg [15:0] psum_reg_9_2_sva;
  reg [7:0] step_mux_149_itm_1;
  reg [7:0] input_reg_9_1_sva;
  reg [15:0] psum_reg_8_2_sva;
  reg [7:0] step_mux_133_itm_1;
  reg [7:0] input_reg_8_1_sva;
  reg [15:0] psum_reg_7_2_sva;
  reg [7:0] step_mux_117_itm_1;
  reg [7:0] input_reg_7_1_sva;
  reg [15:0] psum_reg_6_2_sva;
  reg [7:0] step_mux_101_itm_1;
  reg [7:0] input_reg_6_1_sva;
  reg [15:0] psum_reg_5_2_sva;
  reg [7:0] step_mux_85_itm_1;
  reg [7:0] input_reg_5_1_sva;
  reg [15:0] psum_reg_4_2_sva;
  reg [7:0] step_mux_69_itm_1;
  reg [7:0] input_reg_4_1_sva;
  reg [15:0] psum_reg_3_2_sva;
  reg [7:0] step_mux_53_itm_1;
  reg [7:0] input_reg_3_1_sva;
  reg [15:0] psum_reg_2_2_sva;
  reg [7:0] step_mux_37_itm_1;
  reg [7:0] input_reg_2_1_sva;
  reg [15:0] psum_reg_1_2_sva;
  reg [7:0] step_mux_21_itm_1;
  reg [7:0] input_reg_1_1_sva;
  reg [7:0] step_mux_5_itm_1;
  reg [15:0] psum_reg_15_1_sva;
  reg [7:0] step_mux_244_itm_1;
  reg [15:0] psum_reg_14_1_sva;
  reg [7:0] step_mux_228_itm_1;
  reg [15:0] psum_reg_13_1_sva;
  reg [7:0] step_mux_212_itm_1;
  reg [15:0] psum_reg_12_1_sva;
  reg [7:0] step_mux_196_itm_1;
  reg [15:0] psum_reg_11_1_sva;
  reg [7:0] step_mux_180_itm_1;
  reg [15:0] psum_reg_10_1_sva;
  reg [7:0] step_mux_164_itm_1;
  reg [15:0] psum_reg_9_1_sva;
  reg [7:0] step_mux_148_itm_1;
  reg [15:0] psum_reg_8_1_sva;
  reg [7:0] step_mux_132_itm_1;
  reg [15:0] psum_reg_7_1_sva;
  reg [7:0] step_mux_116_itm_1;
  reg [15:0] psum_reg_6_1_sva;
  reg [7:0] step_mux_100_itm_1;
  reg [15:0] psum_reg_5_1_sva;
  reg [7:0] step_mux_84_itm_1;
  reg [15:0] psum_reg_4_1_sva;
  reg [7:0] step_mux_68_itm_1;
  reg [15:0] psum_reg_3_1_sva;
  reg [7:0] step_mux_52_itm_1;
  reg [15:0] psum_reg_2_1_sva;
  reg [7:0] step_mux_36_itm_1;
  reg [15:0] psum_reg_1_1_sva;
  reg [7:0] step_mux_20_itm_1;
  reg [15:0] psum_reg_16_16_sva;
  reg [5:0] step_if_3_for_1_operator_16_false_acc_cse_sva_3;
  reg [127:0] step_in_col_value_lpi_1;
  reg [7:0] weight_reg_7_15_sva;
  reg [7:0] weight_reg_8_0_sva;
  reg [7:0] weight_reg_7_14_sva;
  reg [7:0] weight_reg_8_1_sva;
  reg [7:0] weight_reg_7_13_sva;
  reg [7:0] weight_reg_8_2_sva;
  reg [7:0] weight_reg_7_12_sva;
  reg [7:0] weight_reg_8_3_sva;
  reg [7:0] weight_reg_7_11_sva;
  reg [7:0] weight_reg_8_4_sva;
  reg [7:0] weight_reg_7_10_sva;
  reg [7:0] weight_reg_8_5_sva;
  reg [7:0] weight_reg_7_9_sva;
  reg [7:0] weight_reg_8_6_sva;
  reg [7:0] weight_reg_7_8_sva;
  reg [7:0] weight_reg_8_7_sva;
  reg [7:0] weight_reg_7_7_sva;
  reg [7:0] weight_reg_8_8_sva;
  reg [7:0] weight_reg_7_6_sva;
  reg [7:0] weight_reg_8_9_sva;
  reg [7:0] weight_reg_7_5_sva;
  reg [7:0] weight_reg_8_10_sva;
  reg [7:0] weight_reg_7_4_sva;
  reg [7:0] weight_reg_8_11_sva;
  reg [7:0] weight_reg_7_3_sva;
  reg [7:0] weight_reg_8_12_sva;
  reg [7:0] weight_reg_7_2_sva;
  reg [7:0] weight_reg_8_13_sva;
  reg [7:0] weight_reg_7_1_sva;
  reg [7:0] weight_reg_8_14_sva;
  reg [7:0] weight_reg_7_0_sva;
  reg [7:0] weight_reg_8_15_sva;
  reg [7:0] weight_reg_6_15_sva;
  reg [7:0] weight_reg_9_0_sva;
  reg [7:0] weight_reg_6_14_sva;
  reg [7:0] weight_reg_9_1_sva;
  reg [7:0] weight_reg_6_13_sva;
  reg [7:0] weight_reg_9_2_sva;
  reg [7:0] weight_reg_6_12_sva;
  reg [7:0] weight_reg_9_3_sva;
  reg [7:0] weight_reg_6_11_sva;
  reg [7:0] weight_reg_9_4_sva;
  reg [7:0] weight_reg_6_10_sva;
  reg [7:0] weight_reg_9_5_sva;
  reg [7:0] weight_reg_6_9_sva;
  reg [7:0] weight_reg_9_6_sva;
  reg [7:0] weight_reg_6_8_sva;
  reg [7:0] weight_reg_9_7_sva;
  reg [7:0] weight_reg_6_7_sva;
  reg [7:0] weight_reg_9_8_sva;
  reg [7:0] weight_reg_6_6_sva;
  reg [7:0] weight_reg_9_9_sva;
  reg [7:0] weight_reg_6_5_sva;
  reg [7:0] weight_reg_9_10_sva;
  reg [7:0] weight_reg_6_4_sva;
  reg [7:0] weight_reg_9_11_sva;
  reg [7:0] weight_reg_6_3_sva;
  reg [7:0] weight_reg_9_12_sva;
  reg [7:0] weight_reg_6_2_sva;
  reg [7:0] weight_reg_9_13_sva;
  reg [7:0] weight_reg_6_1_sva;
  reg [7:0] weight_reg_9_14_sva;
  reg [7:0] weight_reg_6_0_sva;
  reg [7:0] weight_reg_9_15_sva;
  reg [7:0] weight_reg_5_15_sva;
  reg [7:0] weight_reg_10_0_sva;
  reg [7:0] weight_reg_5_14_sva;
  reg [7:0] weight_reg_10_1_sva;
  reg [7:0] weight_reg_5_13_sva;
  reg [7:0] weight_reg_10_2_sva;
  reg [7:0] weight_reg_5_12_sva;
  reg [7:0] weight_reg_10_3_sva;
  reg [7:0] weight_reg_5_11_sva;
  reg [7:0] weight_reg_10_4_sva;
  reg [7:0] weight_reg_5_10_sva;
  reg [7:0] weight_reg_10_5_sva;
  reg [7:0] weight_reg_5_9_sva;
  reg [7:0] weight_reg_10_6_sva;
  reg [7:0] weight_reg_5_8_sva;
  reg [7:0] weight_reg_10_7_sva;
  reg [7:0] weight_reg_5_7_sva;
  reg [7:0] weight_reg_10_8_sva;
  reg [7:0] weight_reg_5_6_sva;
  reg [7:0] weight_reg_10_9_sva;
  reg [7:0] weight_reg_5_5_sva;
  reg [7:0] weight_reg_10_10_sva;
  reg [7:0] weight_reg_5_4_sva;
  reg [7:0] weight_reg_10_11_sva;
  reg [7:0] weight_reg_5_3_sva;
  reg [7:0] weight_reg_10_12_sva;
  reg [7:0] weight_reg_5_2_sva;
  reg [7:0] weight_reg_10_13_sva;
  reg [7:0] weight_reg_5_1_sva;
  reg [7:0] weight_reg_10_14_sva;
  reg [7:0] weight_reg_5_0_sva;
  reg [7:0] weight_reg_10_15_sva;
  reg [7:0] weight_reg_4_15_sva;
  reg [7:0] weight_reg_11_0_sva;
  reg [7:0] weight_reg_4_14_sva;
  reg [7:0] weight_reg_11_1_sva;
  reg [7:0] weight_reg_4_13_sva;
  reg [7:0] weight_reg_11_2_sva;
  reg [7:0] weight_reg_4_12_sva;
  reg [7:0] weight_reg_11_3_sva;
  reg [7:0] weight_reg_4_11_sva;
  reg [7:0] weight_reg_11_4_sva;
  reg [7:0] weight_reg_4_10_sva;
  reg [7:0] weight_reg_11_5_sva;
  reg [7:0] weight_reg_4_9_sva;
  reg [7:0] weight_reg_11_6_sva;
  reg [7:0] weight_reg_4_8_sva;
  reg [7:0] weight_reg_11_7_sva;
  reg [7:0] weight_reg_4_7_sva;
  reg [7:0] weight_reg_11_8_sva;
  reg [7:0] weight_reg_4_6_sva;
  reg [7:0] weight_reg_11_9_sva;
  reg [7:0] weight_reg_4_5_sva;
  reg [7:0] weight_reg_11_10_sva;
  reg [7:0] weight_reg_4_4_sva;
  reg [7:0] weight_reg_11_11_sva;
  reg [7:0] weight_reg_4_3_sva;
  reg [7:0] weight_reg_11_12_sva;
  reg [7:0] weight_reg_4_2_sva;
  reg [7:0] weight_reg_11_13_sva;
  reg [7:0] weight_reg_4_1_sva;
  reg [7:0] weight_reg_11_14_sva;
  reg [7:0] weight_reg_4_0_sva;
  reg [7:0] weight_reg_11_15_sva;
  reg [7:0] weight_reg_3_15_sva;
  reg [7:0] weight_reg_12_0_sva;
  reg [7:0] weight_reg_3_14_sva;
  reg [7:0] weight_reg_12_1_sva;
  reg [7:0] weight_reg_3_13_sva;
  reg [7:0] weight_reg_12_2_sva;
  reg [7:0] weight_reg_3_12_sva;
  reg [7:0] weight_reg_12_3_sva;
  reg [7:0] weight_reg_3_11_sva;
  reg [7:0] weight_reg_12_4_sva;
  reg [7:0] weight_reg_3_10_sva;
  reg [7:0] weight_reg_12_5_sva;
  reg [7:0] weight_reg_3_9_sva;
  reg [7:0] weight_reg_12_6_sva;
  reg [7:0] weight_reg_3_8_sva;
  reg [7:0] weight_reg_12_7_sva;
  reg [7:0] weight_reg_3_7_sva;
  reg [7:0] weight_reg_12_8_sva;
  reg [7:0] weight_reg_3_6_sva;
  reg [7:0] weight_reg_12_9_sva;
  reg [7:0] weight_reg_3_5_sva;
  reg [7:0] weight_reg_12_10_sva;
  reg [7:0] weight_reg_3_4_sva;
  reg [7:0] weight_reg_12_11_sva;
  reg [7:0] weight_reg_3_3_sva;
  reg [7:0] weight_reg_12_12_sva;
  reg [7:0] weight_reg_3_2_sva;
  reg [7:0] weight_reg_12_13_sva;
  reg [7:0] weight_reg_3_1_sva;
  reg [7:0] weight_reg_12_14_sva;
  reg [7:0] weight_reg_3_0_sva;
  reg [7:0] weight_reg_12_15_sva;
  reg [7:0] weight_reg_2_15_sva;
  reg [7:0] weight_reg_13_0_sva;
  reg [7:0] weight_reg_2_14_sva;
  reg [7:0] weight_reg_13_1_sva;
  reg [7:0] weight_reg_2_13_sva;
  reg [7:0] weight_reg_13_2_sva;
  reg [7:0] weight_reg_2_12_sva;
  reg [7:0] weight_reg_13_3_sva;
  reg [7:0] weight_reg_2_11_sva;
  reg [7:0] weight_reg_13_4_sva;
  reg [7:0] weight_reg_2_10_sva;
  reg [7:0] weight_reg_13_5_sva;
  reg [7:0] weight_reg_2_9_sva;
  reg [7:0] weight_reg_13_6_sva;
  reg [7:0] weight_reg_2_8_sva;
  reg [7:0] weight_reg_13_7_sva;
  reg [7:0] weight_reg_2_7_sva;
  reg [7:0] weight_reg_13_8_sva;
  reg [7:0] weight_reg_2_6_sva;
  reg [7:0] weight_reg_13_9_sva;
  reg [7:0] weight_reg_2_5_sva;
  reg [7:0] weight_reg_13_10_sva;
  reg [7:0] weight_reg_2_4_sva;
  reg [7:0] weight_reg_13_11_sva;
  reg [7:0] weight_reg_2_3_sva;
  reg [7:0] weight_reg_13_12_sva;
  reg [7:0] weight_reg_2_2_sva;
  reg [7:0] weight_reg_13_13_sva;
  reg [7:0] weight_reg_2_1_sva;
  reg [7:0] weight_reg_13_14_sva;
  reg [7:0] weight_reg_2_0_sva;
  reg [7:0] weight_reg_13_15_sva;
  reg [7:0] weight_reg_1_15_sva;
  reg [7:0] weight_reg_14_0_sva;
  reg [7:0] weight_reg_1_14_sva;
  reg [7:0] weight_reg_14_1_sva;
  reg [7:0] weight_reg_1_13_sva;
  reg [7:0] weight_reg_14_2_sva;
  reg [7:0] weight_reg_1_12_sva;
  reg [7:0] weight_reg_14_3_sva;
  reg [7:0] weight_reg_1_11_sva;
  reg [7:0] weight_reg_14_4_sva;
  reg [7:0] weight_reg_1_10_sva;
  reg [7:0] weight_reg_14_5_sva;
  reg [7:0] weight_reg_1_9_sva;
  reg [7:0] weight_reg_14_6_sva;
  reg [7:0] weight_reg_1_8_sva;
  reg [7:0] weight_reg_14_7_sva;
  reg [7:0] weight_reg_1_7_sva;
  reg [7:0] weight_reg_14_8_sva;
  reg [7:0] weight_reg_1_6_sva;
  reg [7:0] weight_reg_14_9_sva;
  reg [7:0] weight_reg_1_5_sva;
  reg [7:0] weight_reg_14_10_sva;
  reg [7:0] weight_reg_1_4_sva;
  reg [7:0] weight_reg_14_11_sva;
  reg [7:0] weight_reg_1_3_sva;
  reg [7:0] weight_reg_14_12_sva;
  reg [7:0] weight_reg_1_2_sva;
  reg [7:0] weight_reg_14_13_sva;
  reg [7:0] weight_reg_1_1_sva;
  reg [7:0] weight_reg_14_14_sva;
  reg [7:0] weight_reg_1_0_sva;
  reg [7:0] weight_reg_14_15_sva;
  reg [7:0] weight_reg_0_15_sva;
  reg [7:0] weight_reg_15_0_sva;
  reg [7:0] weight_reg_0_14_sva;
  reg [7:0] weight_reg_15_1_sva;
  reg [7:0] weight_reg_0_13_sva;
  reg [7:0] weight_reg_15_2_sva;
  reg [7:0] weight_reg_0_12_sva;
  reg [7:0] weight_reg_15_3_sva;
  reg [7:0] weight_reg_0_11_sva;
  reg [7:0] weight_reg_15_4_sva;
  reg [7:0] weight_reg_0_10_sva;
  reg [7:0] weight_reg_15_5_sva;
  reg [7:0] weight_reg_0_9_sva;
  reg [7:0] weight_reg_15_6_sva;
  reg [7:0] weight_reg_0_8_sva;
  reg [7:0] weight_reg_15_7_sva;
  reg [7:0] weight_reg_0_7_sva;
  reg [7:0] weight_reg_15_8_sva;
  reg [7:0] weight_reg_0_6_sva;
  reg [7:0] weight_reg_15_9_sva;
  reg [7:0] weight_reg_0_5_sva;
  reg [7:0] weight_reg_15_10_sva;
  reg [7:0] weight_reg_0_4_sva;
  reg [7:0] weight_reg_15_11_sva;
  reg [7:0] weight_reg_0_3_sva;
  reg [7:0] weight_reg_15_12_sva;
  reg [7:0] weight_reg_0_2_sva;
  reg [7:0] weight_reg_15_13_sva;
  reg [7:0] weight_reg_0_1_sva;
  reg [7:0] weight_reg_15_14_sva;
  reg [7:0] weight_reg_0_0_sva;
  reg [7:0] weight_reg_15_15_sva;
  reg [47:0] loopIndicesIn_crt_lpi_1_dfm;
  reg step_if_for_and_stg_2_7_sva;
  reg step_if_for_and_stg_2_6_sva;
  reg step_if_for_and_stg_2_5_sva;
  reg step_if_for_and_stg_2_4_sva;
  reg step_if_for_and_stg_2_3_sva;
  reg step_if_for_and_stg_2_2_sva;
  reg step_if_for_and_stg_2_1_sva;
  reg step_if_for_and_stg_2_0_sva;
  reg [5:0] step_if_3_for_1_operator_16_false_acc_cse_sva_1;
  wire [6:0] nl_step_if_3_for_1_operator_16_false_acc_cse_sva_1;
  reg [5:0] step_if_3_for_1_operator_16_false_acc_cse_sva_2;
  reg step_if_3_if_step_if_3_if_and_1_itm_2;
  reg [47:0] paramsIn_crt_lpi_1_dfm_127_80;
  reg [31:0] paramsIn_crt_lpi_1_dfm_63_32;
  wire [47:0] paramsIn_crt_lpi_1_dfm_127_80_mx0;
  wire [31:0] paramsIn_crt_lpi_1_dfm_63_32_mx0;
  wire step_if_for_and_stg_2_0_sva_mx1w0;
  wire step_if_for_and_stg_2_1_sva_mx1w0;
  wire step_if_for_and_stg_2_2_sva_mx1w0;
  wire step_if_for_and_stg_2_3_sva_mx1w0;
  wire step_if_for_and_stg_2_4_sva_mx1w0;
  wire step_if_for_and_stg_2_5_sva_mx1w0;
  wire step_if_for_and_stg_2_6_sva_mx1w0;
  wire step_if_for_and_stg_2_7_sva_mx1w0;
  wire step_and_96_psp_1;
  wire step_and_psp_1;
  wire psum_reg_and_cse;
  wire step_if_3_if_and_cse;
  wire step_and_499_cse;
  wire and_1562_cse;
  wire step_if_3_if_and_1_cse;
  wire step_if_for_and_20_cse;
  wire step_and_757_cse;
  reg reg_step_not_mdf_sva_3_cse;
  wire weight_reg_and_cse;
  wire weight_reg_and_1_cse;
  wire weight_reg_and_32_cse;
  wire weight_reg_and_33_cse;
  wire weight_reg_and_64_cse;
  wire weight_reg_and_65_cse;
  wire weight_reg_and_96_cse;
  wire weight_reg_and_97_cse;
  wire weight_reg_and_128_cse;
  wire weight_reg_and_129_cse;
  wire weight_reg_and_160_cse;
  wire weight_reg_and_161_cse;
  wire weight_reg_and_192_cse;
  wire weight_reg_and_193_cse;
  wire weight_reg_and_224_cse;
  wire weight_reg_and_225_cse;
  wire [31:0] step_mul_itm;
  wire operator_32_false_acc_itm_31;
  wire operator_16_false_acc_itm_12_1;
  wire step_if_1_acc_itm_32_1;
  wire operator_16_false_acc_itm_16_1;

  wire[0:0] or_73_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] or_1168_nl;
  wire[0:0] nor_290_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] or_1167_nl;
  wire[0:0] nor_289_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_1166_nl;
  wire[0:0] nor_288_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] or_1165_nl;
  wire[0:0] nor_287_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] or_1164_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] or_1163_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] mux_107_nl;
  wire[0:0] or_1162_nl;
  wire[0:0] nor_284_nl;
  wire[0:0] mux_138_nl;
  wire[0:0] or_1161_nl;
  wire[0:0] nor_283_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] or_1160_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] or_1159_nl;
  wire[0:0] nor_281_nl;
  wire[0:0] mux_171_nl;
  wire[0:0] or_1158_nl;
  wire[0:0] nor_280_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] or_1157_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] or_1156_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] or_1155_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] step_if_3_if_step_if_3_if_and_1_nl;
  wire[0:0] and_19_nl;
  wire[31:0] operator_32_false_acc_nl;
  wire[32:0] nl_operator_32_false_acc_nl;
  wire[32:0] operator_32_false_acc_1_nl;
  wire[33:0] nl_operator_32_false_acc_1_nl;
  wire[12:0] operator_16_false_acc_nl;
  wire[13:0] nl_operator_16_false_acc_nl;
  wire[32:0] step_if_1_acc_nl;
  wire[34:0] nl_step_if_1_acc_nl;
  wire[16:0] operator_16_false_acc_nl_1;
  wire[17:0] nl_operator_16_false_acc_nl_1;
  wire[0:0] step_not_12_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[0:0] step_if_2_aelse_1_not_18_nl;
  wire [15:0] nl_accum_fifo_15_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_18_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_15_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_15_i_q_d_mxwt, (step_if_2_aelse_1_not_18_nl));
  wire[0:0] psum_reg_and_256_nl;
  wire [15:0] nl_output_fifo_0_rsci_input_rsc_dat;
  assign psum_reg_and_256_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_0_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_1_sva, pe_0_0_run_cmp_241_psum_out_rsc_z,
      psum_reg_and_256_nl);
  wire[0:0] step_if_2_aelse_1_not_19_nl;
  wire [15:0] nl_accum_fifo_14_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_19_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_14_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_14_i_q_d_mxwt, (step_if_2_aelse_1_not_19_nl));
  wire[0:0] psum_reg_and_257_nl;
  wire [15:0] nl_output_fifo_1_rsci_input_rsc_dat;
  assign psum_reg_and_257_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_1_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_2_sva, pe_0_0_run_cmp_225_psum_out_rsc_z,
      psum_reg_and_257_nl);
  wire[0:0] step_if_2_aelse_1_not_20_nl;
  wire [15:0] nl_accum_fifo_13_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_20_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_13_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_13_i_q_d_mxwt, (step_if_2_aelse_1_not_20_nl));
  wire[0:0] psum_reg_and_258_nl;
  wire [15:0] nl_output_fifo_2_rsci_input_rsc_dat;
  assign psum_reg_and_258_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_2_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_3_sva, pe_0_0_run_cmp_209_psum_out_rsc_z,
      psum_reg_and_258_nl);
  wire[0:0] step_if_2_aelse_1_not_21_nl;
  wire [15:0] nl_accum_fifo_12_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_21_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_12_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_12_i_q_d_mxwt, (step_if_2_aelse_1_not_21_nl));
  wire[0:0] psum_reg_and_259_nl;
  wire [15:0] nl_output_fifo_3_rsci_input_rsc_dat;
  assign psum_reg_and_259_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_3_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_4_sva, pe_0_0_run_cmp_193_psum_out_rsc_z,
      psum_reg_and_259_nl);
  wire[0:0] step_if_2_aelse_1_not_22_nl;
  wire [15:0] nl_accum_fifo_11_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_22_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_11_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_11_i_q_d_mxwt, (step_if_2_aelse_1_not_22_nl));
  wire[0:0] psum_reg_and_260_nl;
  wire [15:0] nl_output_fifo_4_rsci_input_rsc_dat;
  assign psum_reg_and_260_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_4_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_5_sva, pe_0_0_run_cmp_177_psum_out_rsc_z,
      psum_reg_and_260_nl);
  wire[0:0] step_if_2_aelse_1_not_23_nl;
  wire [15:0] nl_accum_fifo_10_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_23_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_10_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_10_i_q_d_mxwt, (step_if_2_aelse_1_not_23_nl));
  wire[0:0] psum_reg_and_261_nl;
  wire [15:0] nl_output_fifo_5_rsci_input_rsc_dat;
  assign psum_reg_and_261_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_5_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_6_sva, pe_0_0_run_cmp_161_psum_out_rsc_z,
      psum_reg_and_261_nl);
  wire[0:0] step_if_2_aelse_1_not_24_nl;
  wire [15:0] nl_accum_fifo_9_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_24_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_9_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_9_i_q_d_mxwt, (step_if_2_aelse_1_not_24_nl));
  wire[0:0] psum_reg_and_262_nl;
  wire [15:0] nl_output_fifo_6_rsci_input_rsc_dat;
  assign psum_reg_and_262_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_6_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_7_sva, pe_0_0_run_cmp_145_psum_out_rsc_z,
      psum_reg_and_262_nl);
  wire[0:0] step_if_2_aelse_1_not_25_nl;
  wire [15:0] nl_accum_fifo_8_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_25_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_8_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_8_i_q_d_mxwt, (step_if_2_aelse_1_not_25_nl));
  wire[0:0] psum_reg_and_263_nl;
  wire [15:0] nl_output_fifo_7_rsci_input_rsc_dat;
  assign psum_reg_and_263_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_7_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_8_sva, pe_0_0_run_cmp_129_psum_out_rsc_z,
      psum_reg_and_263_nl);
  wire[0:0] step_if_2_aelse_1_not_26_nl;
  wire [15:0] nl_accum_fifo_7_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_26_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_7_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_7_i_q_d_mxwt, (step_if_2_aelse_1_not_26_nl));
  wire[0:0] psum_reg_and_264_nl;
  wire [15:0] nl_output_fifo_8_rsci_input_rsc_dat;
  assign psum_reg_and_264_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_8_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_9_sva, pe_0_0_run_cmp_113_psum_out_rsc_z,
      psum_reg_and_264_nl);
  wire[0:0] step_if_2_aelse_1_not_27_nl;
  wire [15:0] nl_accum_fifo_6_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_27_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_6_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_6_i_q_d_mxwt, (step_if_2_aelse_1_not_27_nl));
  wire[0:0] psum_reg_and_265_nl;
  wire [15:0] nl_output_fifo_9_rsci_input_rsc_dat;
  assign psum_reg_and_265_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_9_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_10_sva, pe_0_0_run_cmp_97_psum_out_rsc_z,
      psum_reg_and_265_nl);
  wire[0:0] step_if_2_aelse_1_not_28_nl;
  wire [15:0] nl_accum_fifo_5_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_28_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_5_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_5_i_q_d_mxwt, (step_if_2_aelse_1_not_28_nl));
  wire[0:0] psum_reg_and_266_nl;
  wire [15:0] nl_output_fifo_10_rsci_input_rsc_dat;
  assign psum_reg_and_266_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_10_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_11_sva,
      pe_0_0_run_cmp_81_psum_out_rsc_z, psum_reg_and_266_nl);
  wire[0:0] step_if_2_aelse_1_not_29_nl;
  wire [15:0] nl_accum_fifo_4_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_29_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_4_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_4_i_q_d_mxwt, (step_if_2_aelse_1_not_29_nl));
  wire[0:0] psum_reg_and_267_nl;
  wire [15:0] nl_output_fifo_11_rsci_input_rsc_dat;
  assign psum_reg_and_267_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_11_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_12_sva,
      pe_0_0_run_cmp_65_psum_out_rsc_z, psum_reg_and_267_nl);
  wire[0:0] step_if_2_aelse_1_not_30_nl;
  wire [15:0] nl_accum_fifo_3_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_30_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_3_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_3_i_q_d_mxwt, (step_if_2_aelse_1_not_30_nl));
  wire[0:0] psum_reg_and_268_nl;
  wire [15:0] nl_output_fifo_12_rsci_input_rsc_dat;
  assign psum_reg_and_268_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_12_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_13_sva,
      pe_0_0_run_cmp_49_psum_out_rsc_z, psum_reg_and_268_nl);
  wire[0:0] step_if_2_aelse_1_not_31_nl;
  wire [15:0] nl_accum_fifo_2_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_31_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_2_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_2_i_q_d_mxwt, (step_if_2_aelse_1_not_31_nl));
  wire[0:0] psum_reg_and_269_nl;
  wire [15:0] nl_output_fifo_13_rsci_input_rsc_dat;
  assign psum_reg_and_269_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_13_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_14_sva,
      pe_0_0_run_cmp_33_psum_out_rsc_z, psum_reg_and_269_nl);
  wire[0:0] step_if_2_aelse_1_not_32_nl;
  wire [15:0] nl_accum_fifo_1_rsci_input_rsc_dat;
  assign step_if_2_aelse_1_not_32_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_1_rsci_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_1_i_q_d_mxwt, (step_if_2_aelse_1_not_32_nl));
  wire[0:0] psum_reg_and_270_nl;
  wire [15:0] nl_output_fifo_14_rsci_input_rsc_dat;
  assign psum_reg_and_270_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_output_fifo_14_rsci_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_15_sva,
      pe_0_0_run_cmp_17_psum_out_rsc_z, psum_reg_and_270_nl);
  wire [7:0] nl_input_fifo_15_rsci_input_rsc_dat;
  assign nl_input_fifo_15_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[127:120];
  wire [7:0] nl_input_fifo_14_rsci_input_rsc_dat;
  assign nl_input_fifo_14_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[119:112];
  wire [7:0] nl_input_fifo_13_rsci_input_rsc_dat;
  assign nl_input_fifo_13_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[111:104];
  wire [7:0] nl_input_fifo_12_rsci_input_rsc_dat;
  assign nl_input_fifo_12_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[103:96];
  wire [7:0] nl_input_fifo_11_rsci_input_rsc_dat;
  assign nl_input_fifo_11_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[95:88];
  wire [7:0] nl_input_fifo_10_rsci_input_rsc_dat;
  assign nl_input_fifo_10_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[87:80];
  wire [7:0] nl_input_fifo_9_rsci_input_rsc_dat;
  assign nl_input_fifo_9_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[79:72];
  wire [7:0] nl_input_fifo_8_rsci_input_rsc_dat;
  assign nl_input_fifo_8_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[71:64];
  wire [7:0] nl_input_fifo_7_rsci_input_rsc_dat;
  assign nl_input_fifo_7_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[63:56];
  wire [7:0] nl_input_fifo_6_rsci_input_rsc_dat;
  assign nl_input_fifo_6_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[55:48];
  wire [7:0] nl_input_fifo_5_rsci_input_rsc_dat;
  assign nl_input_fifo_5_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[47:40];
  wire [7:0] nl_input_fifo_4_rsci_input_rsc_dat;
  assign nl_input_fifo_4_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[39:32];
  wire [7:0] nl_input_fifo_3_rsci_input_rsc_dat;
  assign nl_input_fifo_3_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[31:24];
  wire [7:0] nl_input_fifo_2_rsci_input_rsc_dat;
  assign nl_input_fifo_2_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[23:16];
  wire [7:0] nl_input_fifo_1_rsci_input_rsc_dat;
  assign nl_input_fifo_1_rsci_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[15:8];
  wire [7:0] nl_pe_0_0_run_cmp_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_weight_rsc_dat = step_mux_4_itm_1;
  wire[0:0] input_reg_and_nl;
  wire [7:0] nl_pe_0_0_run_cmp_1_input_in_rsc_dat;
  assign input_reg_and_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_1_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_15_sva,
      pe_0_0_run_cmp_17_input_out_rsc_z, input_reg_and_nl);
  wire[0:0] psum_reg_and_271_nl;
  wire [15:0] nl_pe_0_0_run_cmp_1_psum_in_rsc_dat;
  assign psum_reg_and_271_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_1_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_16_sva, pe_0_0_run_cmp_2_psum_out_rsc_z,
      psum_reg_and_271_nl);
  wire [7:0] nl_pe_0_0_run_cmp_1_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_1_weight_rsc_dat = step_mux_259_itm_1;
  wire[0:0] input_reg_and_240_nl;
  wire [7:0] nl_pe_0_0_run_cmp_2_input_in_rsc_dat;
  assign input_reg_and_240_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_2_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_15_sva,
      pe_0_0_run_cmp_18_input_out_rsc_z, input_reg_and_240_nl);
  wire[0:0] psum_reg_and_272_nl;
  wire [15:0] nl_pe_0_0_run_cmp_2_psum_in_rsc_dat;
  assign psum_reg_and_272_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_2_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_16_sva, pe_0_0_run_cmp_3_psum_out_rsc_z,
      psum_reg_and_272_nl);
  wire [7:0] nl_pe_0_0_run_cmp_2_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_2_weight_rsc_dat = step_mux_243_itm_1;
  wire[0:0] input_reg_and_241_nl;
  wire [7:0] nl_pe_0_0_run_cmp_3_input_in_rsc_dat;
  assign input_reg_and_241_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_3_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_15_sva,
      pe_0_0_run_cmp_19_input_out_rsc_z, input_reg_and_241_nl);
  wire[0:0] psum_reg_and_273_nl;
  wire [15:0] nl_pe_0_0_run_cmp_3_psum_in_rsc_dat;
  assign psum_reg_and_273_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_3_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_16_sva, pe_0_0_run_cmp_4_psum_out_rsc_z,
      psum_reg_and_273_nl);
  wire [7:0] nl_pe_0_0_run_cmp_3_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_3_weight_rsc_dat = step_mux_227_itm_1;
  wire[0:0] input_reg_and_242_nl;
  wire [7:0] nl_pe_0_0_run_cmp_4_input_in_rsc_dat;
  assign input_reg_and_242_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_4_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_15_sva,
      pe_0_0_run_cmp_20_input_out_rsc_z, input_reg_and_242_nl);
  wire[0:0] psum_reg_and_274_nl;
  wire [15:0] nl_pe_0_0_run_cmp_4_psum_in_rsc_dat;
  assign psum_reg_and_274_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_4_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_16_sva, pe_0_0_run_cmp_5_psum_out_rsc_z,
      psum_reg_and_274_nl);
  wire [7:0] nl_pe_0_0_run_cmp_4_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_4_weight_rsc_dat = step_mux_211_itm_1;
  wire[0:0] input_reg_and_243_nl;
  wire [7:0] nl_pe_0_0_run_cmp_5_input_in_rsc_dat;
  assign input_reg_and_243_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_5_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_15_sva,
      pe_0_0_run_cmp_21_input_out_rsc_z, input_reg_and_243_nl);
  wire[0:0] psum_reg_and_275_nl;
  wire [15:0] nl_pe_0_0_run_cmp_5_psum_in_rsc_dat;
  assign psum_reg_and_275_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_5_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_16_sva, pe_0_0_run_cmp_6_psum_out_rsc_z,
      psum_reg_and_275_nl);
  wire [7:0] nl_pe_0_0_run_cmp_5_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_5_weight_rsc_dat = step_mux_195_itm_1;
  wire[0:0] input_reg_and_244_nl;
  wire [7:0] nl_pe_0_0_run_cmp_6_input_in_rsc_dat;
  assign input_reg_and_244_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_6_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_15_sva,
      pe_0_0_run_cmp_22_input_out_rsc_z, input_reg_and_244_nl);
  wire[0:0] psum_reg_and_276_nl;
  wire [15:0] nl_pe_0_0_run_cmp_6_psum_in_rsc_dat;
  assign psum_reg_and_276_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_6_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_16_sva, pe_0_0_run_cmp_7_psum_out_rsc_z,
      psum_reg_and_276_nl);
  wire [7:0] nl_pe_0_0_run_cmp_6_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_6_weight_rsc_dat = step_mux_179_itm_1;
  wire[0:0] input_reg_and_245_nl;
  wire [7:0] nl_pe_0_0_run_cmp_7_input_in_rsc_dat;
  assign input_reg_and_245_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_7_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_15_sva,
      pe_0_0_run_cmp_23_input_out_rsc_z, input_reg_and_245_nl);
  wire[0:0] psum_reg_and_277_nl;
  wire [15:0] nl_pe_0_0_run_cmp_7_psum_in_rsc_dat;
  assign psum_reg_and_277_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_7_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_16_sva, pe_0_0_run_cmp_8_psum_out_rsc_z,
      psum_reg_and_277_nl);
  wire [7:0] nl_pe_0_0_run_cmp_7_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_7_weight_rsc_dat = step_mux_163_itm_1;
  wire[0:0] input_reg_and_246_nl;
  wire [7:0] nl_pe_0_0_run_cmp_8_input_in_rsc_dat;
  assign input_reg_and_246_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_8_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_15_sva, pe_0_0_run_cmp_24_input_out_rsc_z,
      input_reg_and_246_nl);
  wire[0:0] psum_reg_and_278_nl;
  wire [15:0] nl_pe_0_0_run_cmp_8_psum_in_rsc_dat;
  assign psum_reg_and_278_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_8_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_16_sva, pe_0_0_run_cmp_9_psum_out_rsc_z,
      psum_reg_and_278_nl);
  wire [7:0] nl_pe_0_0_run_cmp_8_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_8_weight_rsc_dat = step_mux_147_itm_1;
  wire[0:0] input_reg_and_247_nl;
  wire [7:0] nl_pe_0_0_run_cmp_9_input_in_rsc_dat;
  assign input_reg_and_247_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_9_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_15_sva, pe_0_0_run_cmp_25_input_out_rsc_z,
      input_reg_and_247_nl);
  wire[0:0] psum_reg_and_279_nl;
  wire [15:0] nl_pe_0_0_run_cmp_9_psum_in_rsc_dat;
  assign psum_reg_and_279_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_9_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_16_sva, pe_0_0_run_cmp_10_psum_out_rsc_z,
      psum_reg_and_279_nl);
  wire [7:0] nl_pe_0_0_run_cmp_9_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_9_weight_rsc_dat = step_mux_131_itm_1;
  wire[0:0] input_reg_and_248_nl;
  wire [7:0] nl_pe_0_0_run_cmp_10_input_in_rsc_dat;
  assign input_reg_and_248_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_10_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_15_sva,
      pe_0_0_run_cmp_26_input_out_rsc_z, input_reg_and_248_nl);
  wire[0:0] psum_reg_and_280_nl;
  wire [15:0] nl_pe_0_0_run_cmp_10_psum_in_rsc_dat;
  assign psum_reg_and_280_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_10_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_16_sva, pe_0_0_run_cmp_11_psum_out_rsc_z,
      psum_reg_and_280_nl);
  wire [7:0] nl_pe_0_0_run_cmp_10_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_10_weight_rsc_dat = step_mux_115_itm_1;
  wire[0:0] input_reg_and_249_nl;
  wire [7:0] nl_pe_0_0_run_cmp_11_input_in_rsc_dat;
  assign input_reg_and_249_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_11_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_15_sva,
      pe_0_0_run_cmp_27_input_out_rsc_z, input_reg_and_249_nl);
  wire[0:0] psum_reg_and_281_nl;
  wire [15:0] nl_pe_0_0_run_cmp_11_psum_in_rsc_dat;
  assign psum_reg_and_281_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_11_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_16_sva, pe_0_0_run_cmp_12_psum_out_rsc_z,
      psum_reg_and_281_nl);
  wire [7:0] nl_pe_0_0_run_cmp_11_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_11_weight_rsc_dat = step_mux_99_itm_1;
  wire[0:0] input_reg_and_250_nl;
  wire [7:0] nl_pe_0_0_run_cmp_12_input_in_rsc_dat;
  assign input_reg_and_250_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_12_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_15_sva,
      pe_0_0_run_cmp_28_input_out_rsc_z, input_reg_and_250_nl);
  wire[0:0] psum_reg_and_282_nl;
  wire [15:0] nl_pe_0_0_run_cmp_12_psum_in_rsc_dat;
  assign psum_reg_and_282_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_12_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_16_sva, pe_0_0_run_cmp_13_psum_out_rsc_z,
      psum_reg_and_282_nl);
  wire [7:0] nl_pe_0_0_run_cmp_12_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_12_weight_rsc_dat = step_mux_83_itm_1;
  wire[0:0] input_reg_and_251_nl;
  wire [7:0] nl_pe_0_0_run_cmp_13_input_in_rsc_dat;
  assign input_reg_and_251_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_13_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_15_sva,
      pe_0_0_run_cmp_29_input_out_rsc_z, input_reg_and_251_nl);
  wire[0:0] psum_reg_and_283_nl;
  wire [15:0] nl_pe_0_0_run_cmp_13_psum_in_rsc_dat;
  assign psum_reg_and_283_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_13_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_16_sva, pe_0_0_run_cmp_14_psum_out_rsc_z,
      psum_reg_and_283_nl);
  wire [7:0] nl_pe_0_0_run_cmp_13_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_13_weight_rsc_dat = step_mux_67_itm_1;
  wire[0:0] input_reg_and_252_nl;
  wire [7:0] nl_pe_0_0_run_cmp_14_input_in_rsc_dat;
  assign input_reg_and_252_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_14_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_15_sva,
      pe_0_0_run_cmp_30_input_out_rsc_z, input_reg_and_252_nl);
  wire[0:0] psum_reg_and_284_nl;
  wire [15:0] nl_pe_0_0_run_cmp_14_psum_in_rsc_dat;
  assign psum_reg_and_284_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_14_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_16_sva, pe_0_0_run_cmp_15_psum_out_rsc_z,
      psum_reg_and_284_nl);
  wire [7:0] nl_pe_0_0_run_cmp_14_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_14_weight_rsc_dat = step_mux_51_itm_1;
  wire[0:0] input_reg_and_253_nl;
  wire [7:0] nl_pe_0_0_run_cmp_15_input_in_rsc_dat;
  assign input_reg_and_253_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_15_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_15_sva,
      pe_0_0_run_cmp_31_input_out_rsc_z, input_reg_and_253_nl);
  wire[0:0] psum_reg_and_285_nl;
  wire [15:0] nl_pe_0_0_run_cmp_15_psum_in_rsc_dat;
  assign psum_reg_and_285_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_15_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_16_sva, pe_0_0_run_cmp_16_psum_out_rsc_z,
      psum_reg_and_285_nl);
  wire [7:0] nl_pe_0_0_run_cmp_15_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_15_weight_rsc_dat = step_mux_35_itm_1;
  wire[0:0] input_reg_and_254_nl;
  wire [7:0] nl_pe_0_0_run_cmp_16_input_in_rsc_dat;
  assign input_reg_and_254_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_16_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_15_sva,
      pe_0_0_run_cmp_32_input_out_rsc_z, input_reg_and_254_nl);
  wire [7:0] nl_pe_0_0_run_cmp_16_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_16_weight_rsc_dat = step_mux_19_itm_1;
  wire[0:0] input_reg_and_255_nl;
  wire [7:0] nl_pe_0_0_run_cmp_17_input_in_rsc_dat;
  assign input_reg_and_255_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_17_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_14_sva,
      pe_0_0_run_cmp_33_input_out_rsc_z, input_reg_and_255_nl);
  wire[0:0] psum_reg_and_286_nl;
  wire [15:0] nl_pe_0_0_run_cmp_17_psum_in_rsc_dat;
  assign psum_reg_and_286_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_17_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_15_sva,
      pe_0_0_run_cmp_18_psum_out_rsc_z, psum_reg_and_286_nl);
  wire [7:0] nl_pe_0_0_run_cmp_17_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_17_weight_rsc_dat = step_mux_258_itm_1;
  wire[0:0] input_reg_and_256_nl;
  wire [7:0] nl_pe_0_0_run_cmp_18_input_in_rsc_dat;
  assign input_reg_and_256_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_18_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_14_sva,
      pe_0_0_run_cmp_34_input_out_rsc_z, input_reg_and_256_nl);
  wire[0:0] psum_reg_and_287_nl;
  wire [15:0] nl_pe_0_0_run_cmp_18_psum_in_rsc_dat;
  assign psum_reg_and_287_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_18_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_15_sva,
      pe_0_0_run_cmp_19_psum_out_rsc_z, psum_reg_and_287_nl);
  wire [7:0] nl_pe_0_0_run_cmp_18_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_18_weight_rsc_dat = step_mux_242_itm_1;
  wire[0:0] input_reg_and_257_nl;
  wire [7:0] nl_pe_0_0_run_cmp_19_input_in_rsc_dat;
  assign input_reg_and_257_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_19_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_14_sva,
      pe_0_0_run_cmp_35_input_out_rsc_z, input_reg_and_257_nl);
  wire[0:0] psum_reg_and_288_nl;
  wire [15:0] nl_pe_0_0_run_cmp_19_psum_in_rsc_dat;
  assign psum_reg_and_288_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_19_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_15_sva,
      pe_0_0_run_cmp_20_psum_out_rsc_z, psum_reg_and_288_nl);
  wire [7:0] nl_pe_0_0_run_cmp_19_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_19_weight_rsc_dat = step_mux_226_itm_1;
  wire[0:0] input_reg_and_258_nl;
  wire [7:0] nl_pe_0_0_run_cmp_20_input_in_rsc_dat;
  assign input_reg_and_258_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_20_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_14_sva,
      pe_0_0_run_cmp_36_input_out_rsc_z, input_reg_and_258_nl);
  wire[0:0] psum_reg_and_289_nl;
  wire [15:0] nl_pe_0_0_run_cmp_20_psum_in_rsc_dat;
  assign psum_reg_and_289_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_20_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_15_sva,
      pe_0_0_run_cmp_21_psum_out_rsc_z, psum_reg_and_289_nl);
  wire [7:0] nl_pe_0_0_run_cmp_20_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_20_weight_rsc_dat = step_mux_210_itm_1;
  wire[0:0] input_reg_and_259_nl;
  wire [7:0] nl_pe_0_0_run_cmp_21_input_in_rsc_dat;
  assign input_reg_and_259_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_21_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_14_sva,
      pe_0_0_run_cmp_37_input_out_rsc_z, input_reg_and_259_nl);
  wire[0:0] psum_reg_and_290_nl;
  wire [15:0] nl_pe_0_0_run_cmp_21_psum_in_rsc_dat;
  assign psum_reg_and_290_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_21_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_15_sva,
      pe_0_0_run_cmp_22_psum_out_rsc_z, psum_reg_and_290_nl);
  wire [7:0] nl_pe_0_0_run_cmp_21_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_21_weight_rsc_dat = step_mux_194_itm_1;
  wire[0:0] input_reg_and_260_nl;
  wire [7:0] nl_pe_0_0_run_cmp_22_input_in_rsc_dat;
  assign input_reg_and_260_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_22_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_14_sva,
      pe_0_0_run_cmp_38_input_out_rsc_z, input_reg_and_260_nl);
  wire[0:0] psum_reg_and_291_nl;
  wire [15:0] nl_pe_0_0_run_cmp_22_psum_in_rsc_dat;
  assign psum_reg_and_291_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_22_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_15_sva,
      pe_0_0_run_cmp_23_psum_out_rsc_z, psum_reg_and_291_nl);
  wire [7:0] nl_pe_0_0_run_cmp_22_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_22_weight_rsc_dat = step_mux_178_itm_1;
  wire[0:0] input_reg_and_261_nl;
  wire [7:0] nl_pe_0_0_run_cmp_23_input_in_rsc_dat;
  assign input_reg_and_261_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_23_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_14_sva,
      pe_0_0_run_cmp_39_input_out_rsc_z, input_reg_and_261_nl);
  wire[0:0] psum_reg_and_292_nl;
  wire [15:0] nl_pe_0_0_run_cmp_23_psum_in_rsc_dat;
  assign psum_reg_and_292_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_23_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_15_sva, pe_0_0_run_cmp_24_psum_out_rsc_z,
      psum_reg_and_292_nl);
  wire [7:0] nl_pe_0_0_run_cmp_23_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_23_weight_rsc_dat = step_mux_162_itm_1;
  wire[0:0] input_reg_and_262_nl;
  wire [7:0] nl_pe_0_0_run_cmp_24_input_in_rsc_dat;
  assign input_reg_and_262_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_24_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_14_sva,
      pe_0_0_run_cmp_40_input_out_rsc_z, input_reg_and_262_nl);
  wire[0:0] psum_reg_and_293_nl;
  wire [15:0] nl_pe_0_0_run_cmp_24_psum_in_rsc_dat;
  assign psum_reg_and_293_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_24_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_15_sva, pe_0_0_run_cmp_25_psum_out_rsc_z,
      psum_reg_and_293_nl);
  wire [7:0] nl_pe_0_0_run_cmp_24_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_24_weight_rsc_dat = step_mux_146_itm_1;
  wire[0:0] input_reg_and_263_nl;
  wire [7:0] nl_pe_0_0_run_cmp_25_input_in_rsc_dat;
  assign input_reg_and_263_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_25_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_14_sva,
      pe_0_0_run_cmp_41_input_out_rsc_z, input_reg_and_263_nl);
  wire[0:0] psum_reg_and_294_nl;
  wire [15:0] nl_pe_0_0_run_cmp_25_psum_in_rsc_dat;
  assign psum_reg_and_294_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_25_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_15_sva, pe_0_0_run_cmp_26_psum_out_rsc_z,
      psum_reg_and_294_nl);
  wire [7:0] nl_pe_0_0_run_cmp_25_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_25_weight_rsc_dat = step_mux_130_itm_1;
  wire[0:0] input_reg_and_264_nl;
  wire [7:0] nl_pe_0_0_run_cmp_26_input_in_rsc_dat;
  assign input_reg_and_264_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_26_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_14_sva,
      pe_0_0_run_cmp_42_input_out_rsc_z, input_reg_and_264_nl);
  wire[0:0] psum_reg_and_295_nl;
  wire [15:0] nl_pe_0_0_run_cmp_26_psum_in_rsc_dat;
  assign psum_reg_and_295_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_26_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_15_sva, pe_0_0_run_cmp_27_psum_out_rsc_z,
      psum_reg_and_295_nl);
  wire [7:0] nl_pe_0_0_run_cmp_26_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_26_weight_rsc_dat = step_mux_114_itm_1;
  wire[0:0] input_reg_and_265_nl;
  wire [7:0] nl_pe_0_0_run_cmp_27_input_in_rsc_dat;
  assign input_reg_and_265_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_27_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_14_sva,
      pe_0_0_run_cmp_43_input_out_rsc_z, input_reg_and_265_nl);
  wire[0:0] psum_reg_and_296_nl;
  wire [15:0] nl_pe_0_0_run_cmp_27_psum_in_rsc_dat;
  assign psum_reg_and_296_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_27_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_15_sva, pe_0_0_run_cmp_28_psum_out_rsc_z,
      psum_reg_and_296_nl);
  wire [7:0] nl_pe_0_0_run_cmp_27_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_27_weight_rsc_dat = step_mux_98_itm_1;
  wire[0:0] input_reg_and_266_nl;
  wire [7:0] nl_pe_0_0_run_cmp_28_input_in_rsc_dat;
  assign input_reg_and_266_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_28_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_14_sva,
      pe_0_0_run_cmp_44_input_out_rsc_z, input_reg_and_266_nl);
  wire[0:0] psum_reg_and_297_nl;
  wire [15:0] nl_pe_0_0_run_cmp_28_psum_in_rsc_dat;
  assign psum_reg_and_297_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_28_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_15_sva, pe_0_0_run_cmp_29_psum_out_rsc_z,
      psum_reg_and_297_nl);
  wire [7:0] nl_pe_0_0_run_cmp_28_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_28_weight_rsc_dat = step_mux_82_itm_1;
  wire[0:0] input_reg_and_267_nl;
  wire [7:0] nl_pe_0_0_run_cmp_29_input_in_rsc_dat;
  assign input_reg_and_267_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_29_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_14_sva,
      pe_0_0_run_cmp_45_input_out_rsc_z, input_reg_and_267_nl);
  wire[0:0] psum_reg_and_298_nl;
  wire [15:0] nl_pe_0_0_run_cmp_29_psum_in_rsc_dat;
  assign psum_reg_and_298_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_29_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_15_sva, pe_0_0_run_cmp_30_psum_out_rsc_z,
      psum_reg_and_298_nl);
  wire [7:0] nl_pe_0_0_run_cmp_29_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_29_weight_rsc_dat = step_mux_66_itm_1;
  wire[0:0] input_reg_and_268_nl;
  wire [7:0] nl_pe_0_0_run_cmp_30_input_in_rsc_dat;
  assign input_reg_and_268_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_30_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_14_sva,
      pe_0_0_run_cmp_46_input_out_rsc_z, input_reg_and_268_nl);
  wire[0:0] psum_reg_and_299_nl;
  wire [15:0] nl_pe_0_0_run_cmp_30_psum_in_rsc_dat;
  assign psum_reg_and_299_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_30_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_15_sva, pe_0_0_run_cmp_31_psum_out_rsc_z,
      psum_reg_and_299_nl);
  wire [7:0] nl_pe_0_0_run_cmp_30_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_30_weight_rsc_dat = step_mux_50_itm_1;
  wire[0:0] input_reg_and_269_nl;
  wire [7:0] nl_pe_0_0_run_cmp_31_input_in_rsc_dat;
  assign input_reg_and_269_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_31_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_14_sva,
      pe_0_0_run_cmp_47_input_out_rsc_z, input_reg_and_269_nl);
  wire[0:0] psum_reg_and_300_nl;
  wire [15:0] nl_pe_0_0_run_cmp_31_psum_in_rsc_dat;
  assign psum_reg_and_300_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_31_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_15_sva, pe_0_0_run_cmp_32_psum_out_rsc_z,
      psum_reg_and_300_nl);
  wire [7:0] nl_pe_0_0_run_cmp_31_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_31_weight_rsc_dat = step_mux_34_itm_1;
  wire[0:0] input_reg_and_270_nl;
  wire [7:0] nl_pe_0_0_run_cmp_32_input_in_rsc_dat;
  assign input_reg_and_270_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_32_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_14_sva,
      pe_0_0_run_cmp_48_input_out_rsc_z, input_reg_and_270_nl);
  wire [7:0] nl_pe_0_0_run_cmp_32_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_32_weight_rsc_dat = step_mux_18_itm_1;
  wire[0:0] input_reg_and_271_nl;
  wire [7:0] nl_pe_0_0_run_cmp_33_input_in_rsc_dat;
  assign input_reg_and_271_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_33_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_13_sva,
      pe_0_0_run_cmp_49_input_out_rsc_z, input_reg_and_271_nl);
  wire[0:0] psum_reg_and_301_nl;
  wire [15:0] nl_pe_0_0_run_cmp_33_psum_in_rsc_dat;
  assign psum_reg_and_301_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_33_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_14_sva,
      pe_0_0_run_cmp_34_psum_out_rsc_z, psum_reg_and_301_nl);
  wire [7:0] nl_pe_0_0_run_cmp_33_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_33_weight_rsc_dat = step_mux_257_itm_1;
  wire[0:0] input_reg_and_272_nl;
  wire [7:0] nl_pe_0_0_run_cmp_34_input_in_rsc_dat;
  assign input_reg_and_272_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_34_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_13_sva,
      pe_0_0_run_cmp_50_input_out_rsc_z, input_reg_and_272_nl);
  wire[0:0] psum_reg_and_302_nl;
  wire [15:0] nl_pe_0_0_run_cmp_34_psum_in_rsc_dat;
  assign psum_reg_and_302_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_34_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_14_sva,
      pe_0_0_run_cmp_35_psum_out_rsc_z, psum_reg_and_302_nl);
  wire [7:0] nl_pe_0_0_run_cmp_34_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_34_weight_rsc_dat = step_mux_241_itm_1;
  wire[0:0] input_reg_and_273_nl;
  wire [7:0] nl_pe_0_0_run_cmp_35_input_in_rsc_dat;
  assign input_reg_and_273_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_35_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_13_sva,
      pe_0_0_run_cmp_51_input_out_rsc_z, input_reg_and_273_nl);
  wire[0:0] psum_reg_and_303_nl;
  wire [15:0] nl_pe_0_0_run_cmp_35_psum_in_rsc_dat;
  assign psum_reg_and_303_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_35_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_14_sva,
      pe_0_0_run_cmp_36_psum_out_rsc_z, psum_reg_and_303_nl);
  wire [7:0] nl_pe_0_0_run_cmp_35_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_35_weight_rsc_dat = step_mux_225_itm_1;
  wire[0:0] input_reg_and_274_nl;
  wire [7:0] nl_pe_0_0_run_cmp_36_input_in_rsc_dat;
  assign input_reg_and_274_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_36_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_13_sva,
      pe_0_0_run_cmp_52_input_out_rsc_z, input_reg_and_274_nl);
  wire[0:0] psum_reg_and_304_nl;
  wire [15:0] nl_pe_0_0_run_cmp_36_psum_in_rsc_dat;
  assign psum_reg_and_304_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_36_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_14_sva,
      pe_0_0_run_cmp_37_psum_out_rsc_z, psum_reg_and_304_nl);
  wire [7:0] nl_pe_0_0_run_cmp_36_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_36_weight_rsc_dat = step_mux_209_itm_1;
  wire[0:0] input_reg_and_275_nl;
  wire [7:0] nl_pe_0_0_run_cmp_37_input_in_rsc_dat;
  assign input_reg_and_275_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_37_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_13_sva,
      pe_0_0_run_cmp_53_input_out_rsc_z, input_reg_and_275_nl);
  wire[0:0] psum_reg_and_305_nl;
  wire [15:0] nl_pe_0_0_run_cmp_37_psum_in_rsc_dat;
  assign psum_reg_and_305_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_37_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_14_sva,
      pe_0_0_run_cmp_38_psum_out_rsc_z, psum_reg_and_305_nl);
  wire [7:0] nl_pe_0_0_run_cmp_37_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_37_weight_rsc_dat = step_mux_193_itm_1;
  wire[0:0] input_reg_and_276_nl;
  wire [7:0] nl_pe_0_0_run_cmp_38_input_in_rsc_dat;
  assign input_reg_and_276_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_38_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_13_sva,
      pe_0_0_run_cmp_54_input_out_rsc_z, input_reg_and_276_nl);
  wire[0:0] psum_reg_and_306_nl;
  wire [15:0] nl_pe_0_0_run_cmp_38_psum_in_rsc_dat;
  assign psum_reg_and_306_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_38_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_14_sva,
      pe_0_0_run_cmp_39_psum_out_rsc_z, psum_reg_and_306_nl);
  wire [7:0] nl_pe_0_0_run_cmp_38_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_38_weight_rsc_dat = step_mux_177_itm_1;
  wire[0:0] input_reg_and_277_nl;
  wire [7:0] nl_pe_0_0_run_cmp_39_input_in_rsc_dat;
  assign input_reg_and_277_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_39_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_13_sva,
      pe_0_0_run_cmp_55_input_out_rsc_z, input_reg_and_277_nl);
  wire[0:0] psum_reg_and_307_nl;
  wire [15:0] nl_pe_0_0_run_cmp_39_psum_in_rsc_dat;
  assign psum_reg_and_307_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_39_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_14_sva, pe_0_0_run_cmp_40_psum_out_rsc_z,
      psum_reg_and_307_nl);
  wire [7:0] nl_pe_0_0_run_cmp_39_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_39_weight_rsc_dat = step_mux_161_itm_1;
  wire[0:0] input_reg_and_278_nl;
  wire [7:0] nl_pe_0_0_run_cmp_40_input_in_rsc_dat;
  assign input_reg_and_278_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_40_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_13_sva,
      pe_0_0_run_cmp_56_input_out_rsc_z, input_reg_and_278_nl);
  wire[0:0] psum_reg_and_308_nl;
  wire [15:0] nl_pe_0_0_run_cmp_40_psum_in_rsc_dat;
  assign psum_reg_and_308_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_40_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_14_sva, pe_0_0_run_cmp_41_psum_out_rsc_z,
      psum_reg_and_308_nl);
  wire [7:0] nl_pe_0_0_run_cmp_40_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_40_weight_rsc_dat = step_mux_145_itm_1;
  wire[0:0] input_reg_and_279_nl;
  wire [7:0] nl_pe_0_0_run_cmp_41_input_in_rsc_dat;
  assign input_reg_and_279_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_41_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_13_sva,
      pe_0_0_run_cmp_57_input_out_rsc_z, input_reg_and_279_nl);
  wire[0:0] psum_reg_and_309_nl;
  wire [15:0] nl_pe_0_0_run_cmp_41_psum_in_rsc_dat;
  assign psum_reg_and_309_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_41_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_14_sva, pe_0_0_run_cmp_42_psum_out_rsc_z,
      psum_reg_and_309_nl);
  wire [7:0] nl_pe_0_0_run_cmp_41_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_41_weight_rsc_dat = step_mux_129_itm_1;
  wire[0:0] input_reg_and_280_nl;
  wire [7:0] nl_pe_0_0_run_cmp_42_input_in_rsc_dat;
  assign input_reg_and_280_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_42_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_13_sva,
      pe_0_0_run_cmp_58_input_out_rsc_z, input_reg_and_280_nl);
  wire[0:0] psum_reg_and_310_nl;
  wire [15:0] nl_pe_0_0_run_cmp_42_psum_in_rsc_dat;
  assign psum_reg_and_310_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_42_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_14_sva, pe_0_0_run_cmp_43_psum_out_rsc_z,
      psum_reg_and_310_nl);
  wire [7:0] nl_pe_0_0_run_cmp_42_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_42_weight_rsc_dat = step_mux_113_itm_1;
  wire[0:0] input_reg_and_281_nl;
  wire [7:0] nl_pe_0_0_run_cmp_43_input_in_rsc_dat;
  assign input_reg_and_281_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_43_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_13_sva,
      pe_0_0_run_cmp_59_input_out_rsc_z, input_reg_and_281_nl);
  wire[0:0] psum_reg_and_311_nl;
  wire [15:0] nl_pe_0_0_run_cmp_43_psum_in_rsc_dat;
  assign psum_reg_and_311_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_43_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_14_sva, pe_0_0_run_cmp_44_psum_out_rsc_z,
      psum_reg_and_311_nl);
  wire [7:0] nl_pe_0_0_run_cmp_43_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_43_weight_rsc_dat = step_mux_97_itm_1;
  wire[0:0] input_reg_and_282_nl;
  wire [7:0] nl_pe_0_0_run_cmp_44_input_in_rsc_dat;
  assign input_reg_and_282_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_44_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_13_sva,
      pe_0_0_run_cmp_60_input_out_rsc_z, input_reg_and_282_nl);
  wire[0:0] psum_reg_and_312_nl;
  wire [15:0] nl_pe_0_0_run_cmp_44_psum_in_rsc_dat;
  assign psum_reg_and_312_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_44_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_14_sva, pe_0_0_run_cmp_45_psum_out_rsc_z,
      psum_reg_and_312_nl);
  wire [7:0] nl_pe_0_0_run_cmp_44_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_44_weight_rsc_dat = step_mux_81_itm_1;
  wire[0:0] input_reg_and_283_nl;
  wire [7:0] nl_pe_0_0_run_cmp_45_input_in_rsc_dat;
  assign input_reg_and_283_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_45_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_13_sva,
      pe_0_0_run_cmp_61_input_out_rsc_z, input_reg_and_283_nl);
  wire[0:0] psum_reg_and_313_nl;
  wire [15:0] nl_pe_0_0_run_cmp_45_psum_in_rsc_dat;
  assign psum_reg_and_313_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_45_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_14_sva, pe_0_0_run_cmp_46_psum_out_rsc_z,
      psum_reg_and_313_nl);
  wire [7:0] nl_pe_0_0_run_cmp_45_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_45_weight_rsc_dat = step_mux_65_itm_1;
  wire[0:0] input_reg_and_284_nl;
  wire [7:0] nl_pe_0_0_run_cmp_46_input_in_rsc_dat;
  assign input_reg_and_284_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_46_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_13_sva,
      pe_0_0_run_cmp_62_input_out_rsc_z, input_reg_and_284_nl);
  wire[0:0] psum_reg_and_314_nl;
  wire [15:0] nl_pe_0_0_run_cmp_46_psum_in_rsc_dat;
  assign psum_reg_and_314_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_46_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_14_sva, pe_0_0_run_cmp_47_psum_out_rsc_z,
      psum_reg_and_314_nl);
  wire [7:0] nl_pe_0_0_run_cmp_46_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_46_weight_rsc_dat = step_mux_49_itm_1;
  wire[0:0] input_reg_and_285_nl;
  wire [7:0] nl_pe_0_0_run_cmp_47_input_in_rsc_dat;
  assign input_reg_and_285_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_47_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_13_sva,
      pe_0_0_run_cmp_63_input_out_rsc_z, input_reg_and_285_nl);
  wire[0:0] psum_reg_and_315_nl;
  wire [15:0] nl_pe_0_0_run_cmp_47_psum_in_rsc_dat;
  assign psum_reg_and_315_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_47_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_14_sva, pe_0_0_run_cmp_48_psum_out_rsc_z,
      psum_reg_and_315_nl);
  wire [7:0] nl_pe_0_0_run_cmp_47_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_47_weight_rsc_dat = step_mux_33_itm_1;
  wire[0:0] input_reg_and_286_nl;
  wire [7:0] nl_pe_0_0_run_cmp_48_input_in_rsc_dat;
  assign input_reg_and_286_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_48_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_13_sva,
      pe_0_0_run_cmp_64_input_out_rsc_z, input_reg_and_286_nl);
  wire [7:0] nl_pe_0_0_run_cmp_48_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_48_weight_rsc_dat = step_mux_17_itm_1;
  wire[0:0] input_reg_and_287_nl;
  wire [7:0] nl_pe_0_0_run_cmp_49_input_in_rsc_dat;
  assign input_reg_and_287_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_49_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_12_sva,
      pe_0_0_run_cmp_65_input_out_rsc_z, input_reg_and_287_nl);
  wire[0:0] psum_reg_and_316_nl;
  wire [15:0] nl_pe_0_0_run_cmp_49_psum_in_rsc_dat;
  assign psum_reg_and_316_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_49_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_13_sva,
      pe_0_0_run_cmp_50_psum_out_rsc_z, psum_reg_and_316_nl);
  wire [7:0] nl_pe_0_0_run_cmp_49_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_49_weight_rsc_dat = step_mux_256_itm_1;
  wire[0:0] input_reg_and_288_nl;
  wire [7:0] nl_pe_0_0_run_cmp_50_input_in_rsc_dat;
  assign input_reg_and_288_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_50_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_12_sva,
      pe_0_0_run_cmp_66_input_out_rsc_z, input_reg_and_288_nl);
  wire[0:0] psum_reg_and_317_nl;
  wire [15:0] nl_pe_0_0_run_cmp_50_psum_in_rsc_dat;
  assign psum_reg_and_317_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_50_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_13_sva,
      pe_0_0_run_cmp_51_psum_out_rsc_z, psum_reg_and_317_nl);
  wire [7:0] nl_pe_0_0_run_cmp_50_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_50_weight_rsc_dat = step_mux_240_itm_1;
  wire[0:0] input_reg_and_289_nl;
  wire [7:0] nl_pe_0_0_run_cmp_51_input_in_rsc_dat;
  assign input_reg_and_289_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_51_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_12_sva,
      pe_0_0_run_cmp_67_input_out_rsc_z, input_reg_and_289_nl);
  wire[0:0] psum_reg_and_318_nl;
  wire [15:0] nl_pe_0_0_run_cmp_51_psum_in_rsc_dat;
  assign psum_reg_and_318_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_51_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_13_sva,
      pe_0_0_run_cmp_52_psum_out_rsc_z, psum_reg_and_318_nl);
  wire [7:0] nl_pe_0_0_run_cmp_51_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_51_weight_rsc_dat = step_mux_224_itm_1;
  wire[0:0] input_reg_and_290_nl;
  wire [7:0] nl_pe_0_0_run_cmp_52_input_in_rsc_dat;
  assign input_reg_and_290_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_52_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_12_sva,
      pe_0_0_run_cmp_68_input_out_rsc_z, input_reg_and_290_nl);
  wire[0:0] psum_reg_and_319_nl;
  wire [15:0] nl_pe_0_0_run_cmp_52_psum_in_rsc_dat;
  assign psum_reg_and_319_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_52_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_13_sva,
      pe_0_0_run_cmp_53_psum_out_rsc_z, psum_reg_and_319_nl);
  wire [7:0] nl_pe_0_0_run_cmp_52_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_52_weight_rsc_dat = step_mux_208_itm_1;
  wire[0:0] input_reg_and_291_nl;
  wire [7:0] nl_pe_0_0_run_cmp_53_input_in_rsc_dat;
  assign input_reg_and_291_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_53_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_12_sva,
      pe_0_0_run_cmp_69_input_out_rsc_z, input_reg_and_291_nl);
  wire[0:0] psum_reg_and_320_nl;
  wire [15:0] nl_pe_0_0_run_cmp_53_psum_in_rsc_dat;
  assign psum_reg_and_320_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_53_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_13_sva,
      pe_0_0_run_cmp_54_psum_out_rsc_z, psum_reg_and_320_nl);
  wire [7:0] nl_pe_0_0_run_cmp_53_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_53_weight_rsc_dat = step_mux_192_itm_1;
  wire[0:0] input_reg_and_292_nl;
  wire [7:0] nl_pe_0_0_run_cmp_54_input_in_rsc_dat;
  assign input_reg_and_292_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_54_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_12_sva,
      pe_0_0_run_cmp_70_input_out_rsc_z, input_reg_and_292_nl);
  wire[0:0] psum_reg_and_321_nl;
  wire [15:0] nl_pe_0_0_run_cmp_54_psum_in_rsc_dat;
  assign psum_reg_and_321_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_54_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_13_sva,
      pe_0_0_run_cmp_55_psum_out_rsc_z, psum_reg_and_321_nl);
  wire [7:0] nl_pe_0_0_run_cmp_54_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_54_weight_rsc_dat = step_mux_176_itm_1;
  wire[0:0] input_reg_and_293_nl;
  wire [7:0] nl_pe_0_0_run_cmp_55_input_in_rsc_dat;
  assign input_reg_and_293_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_55_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_12_sva,
      pe_0_0_run_cmp_71_input_out_rsc_z, input_reg_and_293_nl);
  wire[0:0] psum_reg_and_322_nl;
  wire [15:0] nl_pe_0_0_run_cmp_55_psum_in_rsc_dat;
  assign psum_reg_and_322_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_55_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_13_sva, pe_0_0_run_cmp_56_psum_out_rsc_z,
      psum_reg_and_322_nl);
  wire [7:0] nl_pe_0_0_run_cmp_55_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_55_weight_rsc_dat = step_mux_160_itm_1;
  wire[0:0] input_reg_and_294_nl;
  wire [7:0] nl_pe_0_0_run_cmp_56_input_in_rsc_dat;
  assign input_reg_and_294_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_56_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_12_sva,
      pe_0_0_run_cmp_72_input_out_rsc_z, input_reg_and_294_nl);
  wire[0:0] psum_reg_and_323_nl;
  wire [15:0] nl_pe_0_0_run_cmp_56_psum_in_rsc_dat;
  assign psum_reg_and_323_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_56_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_13_sva, pe_0_0_run_cmp_57_psum_out_rsc_z,
      psum_reg_and_323_nl);
  wire [7:0] nl_pe_0_0_run_cmp_56_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_56_weight_rsc_dat = step_mux_144_itm_1;
  wire[0:0] input_reg_and_295_nl;
  wire [7:0] nl_pe_0_0_run_cmp_57_input_in_rsc_dat;
  assign input_reg_and_295_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_57_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_12_sva,
      pe_0_0_run_cmp_73_input_out_rsc_z, input_reg_and_295_nl);
  wire[0:0] psum_reg_and_324_nl;
  wire [15:0] nl_pe_0_0_run_cmp_57_psum_in_rsc_dat;
  assign psum_reg_and_324_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_57_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_13_sva, pe_0_0_run_cmp_58_psum_out_rsc_z,
      psum_reg_and_324_nl);
  wire [7:0] nl_pe_0_0_run_cmp_57_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_57_weight_rsc_dat = step_mux_128_itm_1;
  wire[0:0] input_reg_and_296_nl;
  wire [7:0] nl_pe_0_0_run_cmp_58_input_in_rsc_dat;
  assign input_reg_and_296_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_58_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_12_sva,
      pe_0_0_run_cmp_74_input_out_rsc_z, input_reg_and_296_nl);
  wire[0:0] psum_reg_and_325_nl;
  wire [15:0] nl_pe_0_0_run_cmp_58_psum_in_rsc_dat;
  assign psum_reg_and_325_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_58_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_13_sva, pe_0_0_run_cmp_59_psum_out_rsc_z,
      psum_reg_and_325_nl);
  wire [7:0] nl_pe_0_0_run_cmp_58_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_58_weight_rsc_dat = step_mux_112_itm_1;
  wire[0:0] input_reg_and_297_nl;
  wire [7:0] nl_pe_0_0_run_cmp_59_input_in_rsc_dat;
  assign input_reg_and_297_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_59_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_12_sva,
      pe_0_0_run_cmp_75_input_out_rsc_z, input_reg_and_297_nl);
  wire[0:0] psum_reg_and_326_nl;
  wire [15:0] nl_pe_0_0_run_cmp_59_psum_in_rsc_dat;
  assign psum_reg_and_326_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_59_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_13_sva, pe_0_0_run_cmp_60_psum_out_rsc_z,
      psum_reg_and_326_nl);
  wire [7:0] nl_pe_0_0_run_cmp_59_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_59_weight_rsc_dat = step_mux_96_itm_1;
  wire[0:0] input_reg_and_298_nl;
  wire [7:0] nl_pe_0_0_run_cmp_60_input_in_rsc_dat;
  assign input_reg_and_298_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_60_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_12_sva,
      pe_0_0_run_cmp_76_input_out_rsc_z, input_reg_and_298_nl);
  wire[0:0] psum_reg_and_327_nl;
  wire [15:0] nl_pe_0_0_run_cmp_60_psum_in_rsc_dat;
  assign psum_reg_and_327_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_60_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_13_sva, pe_0_0_run_cmp_61_psum_out_rsc_z,
      psum_reg_and_327_nl);
  wire [7:0] nl_pe_0_0_run_cmp_60_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_60_weight_rsc_dat = step_mux_80_itm_1;
  wire[0:0] input_reg_and_299_nl;
  wire [7:0] nl_pe_0_0_run_cmp_61_input_in_rsc_dat;
  assign input_reg_and_299_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_61_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_12_sva,
      pe_0_0_run_cmp_77_input_out_rsc_z, input_reg_and_299_nl);
  wire[0:0] psum_reg_and_328_nl;
  wire [15:0] nl_pe_0_0_run_cmp_61_psum_in_rsc_dat;
  assign psum_reg_and_328_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_61_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_13_sva, pe_0_0_run_cmp_62_psum_out_rsc_z,
      psum_reg_and_328_nl);
  wire [7:0] nl_pe_0_0_run_cmp_61_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_61_weight_rsc_dat = step_mux_64_itm_1;
  wire[0:0] input_reg_and_300_nl;
  wire [7:0] nl_pe_0_0_run_cmp_62_input_in_rsc_dat;
  assign input_reg_and_300_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_62_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_12_sva,
      pe_0_0_run_cmp_78_input_out_rsc_z, input_reg_and_300_nl);
  wire[0:0] psum_reg_and_329_nl;
  wire [15:0] nl_pe_0_0_run_cmp_62_psum_in_rsc_dat;
  assign psum_reg_and_329_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_62_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_13_sva, pe_0_0_run_cmp_63_psum_out_rsc_z,
      psum_reg_and_329_nl);
  wire [7:0] nl_pe_0_0_run_cmp_62_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_62_weight_rsc_dat = step_mux_48_itm_1;
  wire[0:0] input_reg_and_301_nl;
  wire [7:0] nl_pe_0_0_run_cmp_63_input_in_rsc_dat;
  assign input_reg_and_301_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_63_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_12_sva,
      pe_0_0_run_cmp_79_input_out_rsc_z, input_reg_and_301_nl);
  wire[0:0] psum_reg_and_330_nl;
  wire [15:0] nl_pe_0_0_run_cmp_63_psum_in_rsc_dat;
  assign psum_reg_and_330_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_63_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_13_sva, pe_0_0_run_cmp_64_psum_out_rsc_z,
      psum_reg_and_330_nl);
  wire [7:0] nl_pe_0_0_run_cmp_63_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_63_weight_rsc_dat = step_mux_32_itm_1;
  wire[0:0] input_reg_and_302_nl;
  wire [7:0] nl_pe_0_0_run_cmp_64_input_in_rsc_dat;
  assign input_reg_and_302_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_64_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_12_sva,
      pe_0_0_run_cmp_80_input_out_rsc_z, input_reg_and_302_nl);
  wire [7:0] nl_pe_0_0_run_cmp_64_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_64_weight_rsc_dat = step_mux_16_itm_1;
  wire[0:0] input_reg_and_303_nl;
  wire [7:0] nl_pe_0_0_run_cmp_65_input_in_rsc_dat;
  assign input_reg_and_303_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_65_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_11_sva,
      pe_0_0_run_cmp_81_input_out_rsc_z, input_reg_and_303_nl);
  wire[0:0] psum_reg_and_331_nl;
  wire [15:0] nl_pe_0_0_run_cmp_65_psum_in_rsc_dat;
  assign psum_reg_and_331_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_65_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_12_sva,
      pe_0_0_run_cmp_66_psum_out_rsc_z, psum_reg_and_331_nl);
  wire [7:0] nl_pe_0_0_run_cmp_65_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_65_weight_rsc_dat = step_mux_255_itm_1;
  wire[0:0] input_reg_and_304_nl;
  wire [7:0] nl_pe_0_0_run_cmp_66_input_in_rsc_dat;
  assign input_reg_and_304_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_66_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_11_sva,
      pe_0_0_run_cmp_82_input_out_rsc_z, input_reg_and_304_nl);
  wire[0:0] psum_reg_and_332_nl;
  wire [15:0] nl_pe_0_0_run_cmp_66_psum_in_rsc_dat;
  assign psum_reg_and_332_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_66_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_12_sva,
      pe_0_0_run_cmp_67_psum_out_rsc_z, psum_reg_and_332_nl);
  wire [7:0] nl_pe_0_0_run_cmp_66_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_66_weight_rsc_dat = step_mux_239_itm_1;
  wire[0:0] input_reg_and_305_nl;
  wire [7:0] nl_pe_0_0_run_cmp_67_input_in_rsc_dat;
  assign input_reg_and_305_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_67_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_11_sva,
      pe_0_0_run_cmp_83_input_out_rsc_z, input_reg_and_305_nl);
  wire[0:0] psum_reg_and_333_nl;
  wire [15:0] nl_pe_0_0_run_cmp_67_psum_in_rsc_dat;
  assign psum_reg_and_333_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_67_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_12_sva,
      pe_0_0_run_cmp_68_psum_out_rsc_z, psum_reg_and_333_nl);
  wire [7:0] nl_pe_0_0_run_cmp_67_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_67_weight_rsc_dat = step_mux_223_itm_1;
  wire[0:0] input_reg_and_306_nl;
  wire [7:0] nl_pe_0_0_run_cmp_68_input_in_rsc_dat;
  assign input_reg_and_306_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_68_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_11_sva,
      pe_0_0_run_cmp_84_input_out_rsc_z, input_reg_and_306_nl);
  wire[0:0] psum_reg_and_334_nl;
  wire [15:0] nl_pe_0_0_run_cmp_68_psum_in_rsc_dat;
  assign psum_reg_and_334_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_68_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_12_sva,
      pe_0_0_run_cmp_69_psum_out_rsc_z, psum_reg_and_334_nl);
  wire [7:0] nl_pe_0_0_run_cmp_68_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_68_weight_rsc_dat = step_mux_207_itm_1;
  wire[0:0] input_reg_and_307_nl;
  wire [7:0] nl_pe_0_0_run_cmp_69_input_in_rsc_dat;
  assign input_reg_and_307_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_69_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_11_sva,
      pe_0_0_run_cmp_85_input_out_rsc_z, input_reg_and_307_nl);
  wire[0:0] psum_reg_and_335_nl;
  wire [15:0] nl_pe_0_0_run_cmp_69_psum_in_rsc_dat;
  assign psum_reg_and_335_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_69_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_12_sva,
      pe_0_0_run_cmp_70_psum_out_rsc_z, psum_reg_and_335_nl);
  wire [7:0] nl_pe_0_0_run_cmp_69_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_69_weight_rsc_dat = step_mux_191_itm_1;
  wire[0:0] input_reg_and_308_nl;
  wire [7:0] nl_pe_0_0_run_cmp_70_input_in_rsc_dat;
  assign input_reg_and_308_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_70_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_11_sva,
      pe_0_0_run_cmp_86_input_out_rsc_z, input_reg_and_308_nl);
  wire[0:0] psum_reg_and_336_nl;
  wire [15:0] nl_pe_0_0_run_cmp_70_psum_in_rsc_dat;
  assign psum_reg_and_336_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_70_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_12_sva,
      pe_0_0_run_cmp_71_psum_out_rsc_z, psum_reg_and_336_nl);
  wire [7:0] nl_pe_0_0_run_cmp_70_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_70_weight_rsc_dat = step_mux_175_itm_1;
  wire[0:0] input_reg_and_309_nl;
  wire [7:0] nl_pe_0_0_run_cmp_71_input_in_rsc_dat;
  assign input_reg_and_309_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_71_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_11_sva,
      pe_0_0_run_cmp_87_input_out_rsc_z, input_reg_and_309_nl);
  wire[0:0] psum_reg_and_337_nl;
  wire [15:0] nl_pe_0_0_run_cmp_71_psum_in_rsc_dat;
  assign psum_reg_and_337_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_71_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_12_sva, pe_0_0_run_cmp_72_psum_out_rsc_z,
      psum_reg_and_337_nl);
  wire [7:0] nl_pe_0_0_run_cmp_71_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_71_weight_rsc_dat = step_mux_159_itm_1;
  wire[0:0] input_reg_and_310_nl;
  wire [7:0] nl_pe_0_0_run_cmp_72_input_in_rsc_dat;
  assign input_reg_and_310_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_72_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_11_sva,
      pe_0_0_run_cmp_88_input_out_rsc_z, input_reg_and_310_nl);
  wire[0:0] psum_reg_and_338_nl;
  wire [15:0] nl_pe_0_0_run_cmp_72_psum_in_rsc_dat;
  assign psum_reg_and_338_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_72_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_12_sva, pe_0_0_run_cmp_73_psum_out_rsc_z,
      psum_reg_and_338_nl);
  wire [7:0] nl_pe_0_0_run_cmp_72_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_72_weight_rsc_dat = step_mux_143_itm_1;
  wire[0:0] input_reg_and_311_nl;
  wire [7:0] nl_pe_0_0_run_cmp_73_input_in_rsc_dat;
  assign input_reg_and_311_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_73_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_11_sva,
      pe_0_0_run_cmp_89_input_out_rsc_z, input_reg_and_311_nl);
  wire[0:0] psum_reg_and_339_nl;
  wire [15:0] nl_pe_0_0_run_cmp_73_psum_in_rsc_dat;
  assign psum_reg_and_339_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_73_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_12_sva, pe_0_0_run_cmp_74_psum_out_rsc_z,
      psum_reg_and_339_nl);
  wire [7:0] nl_pe_0_0_run_cmp_73_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_73_weight_rsc_dat = step_mux_127_itm_1;
  wire[0:0] input_reg_and_312_nl;
  wire [7:0] nl_pe_0_0_run_cmp_74_input_in_rsc_dat;
  assign input_reg_and_312_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_74_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_11_sva,
      pe_0_0_run_cmp_90_input_out_rsc_z, input_reg_and_312_nl);
  wire[0:0] psum_reg_and_340_nl;
  wire [15:0] nl_pe_0_0_run_cmp_74_psum_in_rsc_dat;
  assign psum_reg_and_340_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_74_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_12_sva, pe_0_0_run_cmp_75_psum_out_rsc_z,
      psum_reg_and_340_nl);
  wire [7:0] nl_pe_0_0_run_cmp_74_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_74_weight_rsc_dat = step_mux_111_itm_1;
  wire[0:0] input_reg_and_313_nl;
  wire [7:0] nl_pe_0_0_run_cmp_75_input_in_rsc_dat;
  assign input_reg_and_313_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_75_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_11_sva,
      pe_0_0_run_cmp_91_input_out_rsc_z, input_reg_and_313_nl);
  wire[0:0] psum_reg_and_341_nl;
  wire [15:0] nl_pe_0_0_run_cmp_75_psum_in_rsc_dat;
  assign psum_reg_and_341_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_75_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_12_sva, pe_0_0_run_cmp_76_psum_out_rsc_z,
      psum_reg_and_341_nl);
  wire [7:0] nl_pe_0_0_run_cmp_75_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_75_weight_rsc_dat = step_mux_95_itm_1;
  wire[0:0] input_reg_and_314_nl;
  wire [7:0] nl_pe_0_0_run_cmp_76_input_in_rsc_dat;
  assign input_reg_and_314_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_76_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_11_sva,
      pe_0_0_run_cmp_92_input_out_rsc_z, input_reg_and_314_nl);
  wire[0:0] psum_reg_and_342_nl;
  wire [15:0] nl_pe_0_0_run_cmp_76_psum_in_rsc_dat;
  assign psum_reg_and_342_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_76_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_12_sva, pe_0_0_run_cmp_77_psum_out_rsc_z,
      psum_reg_and_342_nl);
  wire [7:0] nl_pe_0_0_run_cmp_76_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_76_weight_rsc_dat = step_mux_79_itm_1;
  wire[0:0] input_reg_and_315_nl;
  wire [7:0] nl_pe_0_0_run_cmp_77_input_in_rsc_dat;
  assign input_reg_and_315_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_77_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_11_sva,
      pe_0_0_run_cmp_93_input_out_rsc_z, input_reg_and_315_nl);
  wire[0:0] psum_reg_and_343_nl;
  wire [15:0] nl_pe_0_0_run_cmp_77_psum_in_rsc_dat;
  assign psum_reg_and_343_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_77_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_12_sva, pe_0_0_run_cmp_78_psum_out_rsc_z,
      psum_reg_and_343_nl);
  wire [7:0] nl_pe_0_0_run_cmp_77_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_77_weight_rsc_dat = step_mux_63_itm_1;
  wire[0:0] input_reg_and_316_nl;
  wire [7:0] nl_pe_0_0_run_cmp_78_input_in_rsc_dat;
  assign input_reg_and_316_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_78_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_11_sva,
      pe_0_0_run_cmp_94_input_out_rsc_z, input_reg_and_316_nl);
  wire[0:0] psum_reg_and_344_nl;
  wire [15:0] nl_pe_0_0_run_cmp_78_psum_in_rsc_dat;
  assign psum_reg_and_344_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_78_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_12_sva, pe_0_0_run_cmp_79_psum_out_rsc_z,
      psum_reg_and_344_nl);
  wire [7:0] nl_pe_0_0_run_cmp_78_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_78_weight_rsc_dat = step_mux_47_itm_1;
  wire[0:0] input_reg_and_317_nl;
  wire [7:0] nl_pe_0_0_run_cmp_79_input_in_rsc_dat;
  assign input_reg_and_317_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_79_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_11_sva,
      pe_0_0_run_cmp_95_input_out_rsc_z, input_reg_and_317_nl);
  wire[0:0] psum_reg_and_345_nl;
  wire [15:0] nl_pe_0_0_run_cmp_79_psum_in_rsc_dat;
  assign psum_reg_and_345_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_79_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_12_sva, pe_0_0_run_cmp_80_psum_out_rsc_z,
      psum_reg_and_345_nl);
  wire [7:0] nl_pe_0_0_run_cmp_79_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_79_weight_rsc_dat = step_mux_31_itm_1;
  wire[0:0] input_reg_and_318_nl;
  wire [7:0] nl_pe_0_0_run_cmp_80_input_in_rsc_dat;
  assign input_reg_and_318_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_80_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_11_sva,
      pe_0_0_run_cmp_96_input_out_rsc_z, input_reg_and_318_nl);
  wire [7:0] nl_pe_0_0_run_cmp_80_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_80_weight_rsc_dat = step_mux_15_itm_1;
  wire[0:0] input_reg_and_319_nl;
  wire [7:0] nl_pe_0_0_run_cmp_81_input_in_rsc_dat;
  assign input_reg_and_319_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_81_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_10_sva,
      pe_0_0_run_cmp_97_input_out_rsc_z, input_reg_and_319_nl);
  wire[0:0] psum_reg_and_346_nl;
  wire [15:0] nl_pe_0_0_run_cmp_81_psum_in_rsc_dat;
  assign psum_reg_and_346_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_81_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_11_sva,
      pe_0_0_run_cmp_82_psum_out_rsc_z, psum_reg_and_346_nl);
  wire [7:0] nl_pe_0_0_run_cmp_81_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_81_weight_rsc_dat = step_mux_254_itm_1;
  wire[0:0] input_reg_and_320_nl;
  wire [7:0] nl_pe_0_0_run_cmp_82_input_in_rsc_dat;
  assign input_reg_and_320_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_82_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_10_sva,
      pe_0_0_run_cmp_98_input_out_rsc_z, input_reg_and_320_nl);
  wire[0:0] psum_reg_and_347_nl;
  wire [15:0] nl_pe_0_0_run_cmp_82_psum_in_rsc_dat;
  assign psum_reg_and_347_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_82_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_11_sva,
      pe_0_0_run_cmp_83_psum_out_rsc_z, psum_reg_and_347_nl);
  wire [7:0] nl_pe_0_0_run_cmp_82_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_82_weight_rsc_dat = step_mux_238_itm_1;
  wire[0:0] input_reg_and_321_nl;
  wire [7:0] nl_pe_0_0_run_cmp_83_input_in_rsc_dat;
  assign input_reg_and_321_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_83_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_10_sva,
      pe_0_0_run_cmp_99_input_out_rsc_z, input_reg_and_321_nl);
  wire[0:0] psum_reg_and_348_nl;
  wire [15:0] nl_pe_0_0_run_cmp_83_psum_in_rsc_dat;
  assign psum_reg_and_348_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_83_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_11_sva,
      pe_0_0_run_cmp_84_psum_out_rsc_z, psum_reg_and_348_nl);
  wire [7:0] nl_pe_0_0_run_cmp_83_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_83_weight_rsc_dat = step_mux_222_itm_1;
  wire[0:0] input_reg_and_322_nl;
  wire [7:0] nl_pe_0_0_run_cmp_84_input_in_rsc_dat;
  assign input_reg_and_322_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_84_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_10_sva,
      pe_0_0_run_cmp_100_input_out_rsc_z, input_reg_and_322_nl);
  wire[0:0] psum_reg_and_349_nl;
  wire [15:0] nl_pe_0_0_run_cmp_84_psum_in_rsc_dat;
  assign psum_reg_and_349_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_84_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_11_sva,
      pe_0_0_run_cmp_85_psum_out_rsc_z, psum_reg_and_349_nl);
  wire [7:0] nl_pe_0_0_run_cmp_84_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_84_weight_rsc_dat = step_mux_206_itm_1;
  wire[0:0] input_reg_and_323_nl;
  wire [7:0] nl_pe_0_0_run_cmp_85_input_in_rsc_dat;
  assign input_reg_and_323_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_85_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_10_sva,
      pe_0_0_run_cmp_101_input_out_rsc_z, input_reg_and_323_nl);
  wire[0:0] psum_reg_and_350_nl;
  wire [15:0] nl_pe_0_0_run_cmp_85_psum_in_rsc_dat;
  assign psum_reg_and_350_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_85_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_11_sva,
      pe_0_0_run_cmp_86_psum_out_rsc_z, psum_reg_and_350_nl);
  wire [7:0] nl_pe_0_0_run_cmp_85_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_85_weight_rsc_dat = step_mux_190_itm_1;
  wire[0:0] input_reg_and_324_nl;
  wire [7:0] nl_pe_0_0_run_cmp_86_input_in_rsc_dat;
  assign input_reg_and_324_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_86_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_10_sva,
      pe_0_0_run_cmp_102_input_out_rsc_z, input_reg_and_324_nl);
  wire[0:0] psum_reg_and_351_nl;
  wire [15:0] nl_pe_0_0_run_cmp_86_psum_in_rsc_dat;
  assign psum_reg_and_351_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_86_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_11_sva,
      pe_0_0_run_cmp_87_psum_out_rsc_z, psum_reg_and_351_nl);
  wire [7:0] nl_pe_0_0_run_cmp_86_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_86_weight_rsc_dat = step_mux_174_itm_1;
  wire[0:0] input_reg_and_325_nl;
  wire [7:0] nl_pe_0_0_run_cmp_87_input_in_rsc_dat;
  assign input_reg_and_325_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_87_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_10_sva,
      pe_0_0_run_cmp_103_input_out_rsc_z, input_reg_and_325_nl);
  wire[0:0] psum_reg_and_352_nl;
  wire [15:0] nl_pe_0_0_run_cmp_87_psum_in_rsc_dat;
  assign psum_reg_and_352_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_87_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_11_sva, pe_0_0_run_cmp_88_psum_out_rsc_z,
      psum_reg_and_352_nl);
  wire [7:0] nl_pe_0_0_run_cmp_87_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_87_weight_rsc_dat = step_mux_158_itm_1;
  wire[0:0] input_reg_and_326_nl;
  wire [7:0] nl_pe_0_0_run_cmp_88_input_in_rsc_dat;
  assign input_reg_and_326_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_88_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_10_sva,
      pe_0_0_run_cmp_104_input_out_rsc_z, input_reg_and_326_nl);
  wire[0:0] psum_reg_and_353_nl;
  wire [15:0] nl_pe_0_0_run_cmp_88_psum_in_rsc_dat;
  assign psum_reg_and_353_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_88_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_11_sva, pe_0_0_run_cmp_89_psum_out_rsc_z,
      psum_reg_and_353_nl);
  wire [7:0] nl_pe_0_0_run_cmp_88_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_88_weight_rsc_dat = step_mux_142_itm_1;
  wire[0:0] input_reg_and_327_nl;
  wire [7:0] nl_pe_0_0_run_cmp_89_input_in_rsc_dat;
  assign input_reg_and_327_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_89_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_10_sva,
      pe_0_0_run_cmp_105_input_out_rsc_z, input_reg_and_327_nl);
  wire[0:0] psum_reg_and_354_nl;
  wire [15:0] nl_pe_0_0_run_cmp_89_psum_in_rsc_dat;
  assign psum_reg_and_354_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_89_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_11_sva, pe_0_0_run_cmp_90_psum_out_rsc_z,
      psum_reg_and_354_nl);
  wire [7:0] nl_pe_0_0_run_cmp_89_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_89_weight_rsc_dat = step_mux_126_itm_1;
  wire[0:0] input_reg_and_328_nl;
  wire [7:0] nl_pe_0_0_run_cmp_90_input_in_rsc_dat;
  assign input_reg_and_328_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_90_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_10_sva,
      pe_0_0_run_cmp_106_input_out_rsc_z, input_reg_and_328_nl);
  wire[0:0] psum_reg_and_355_nl;
  wire [15:0] nl_pe_0_0_run_cmp_90_psum_in_rsc_dat;
  assign psum_reg_and_355_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_90_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_11_sva, pe_0_0_run_cmp_91_psum_out_rsc_z,
      psum_reg_and_355_nl);
  wire [7:0] nl_pe_0_0_run_cmp_90_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_90_weight_rsc_dat = step_mux_110_itm_1;
  wire[0:0] input_reg_and_329_nl;
  wire [7:0] nl_pe_0_0_run_cmp_91_input_in_rsc_dat;
  assign input_reg_and_329_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_91_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_10_sva,
      pe_0_0_run_cmp_107_input_out_rsc_z, input_reg_and_329_nl);
  wire[0:0] psum_reg_and_356_nl;
  wire [15:0] nl_pe_0_0_run_cmp_91_psum_in_rsc_dat;
  assign psum_reg_and_356_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_91_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_11_sva, pe_0_0_run_cmp_92_psum_out_rsc_z,
      psum_reg_and_356_nl);
  wire [7:0] nl_pe_0_0_run_cmp_91_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_91_weight_rsc_dat = step_mux_94_itm_1;
  wire[0:0] input_reg_and_330_nl;
  wire [7:0] nl_pe_0_0_run_cmp_92_input_in_rsc_dat;
  assign input_reg_and_330_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_92_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_10_sva,
      pe_0_0_run_cmp_108_input_out_rsc_z, input_reg_and_330_nl);
  wire[0:0] psum_reg_and_357_nl;
  wire [15:0] nl_pe_0_0_run_cmp_92_psum_in_rsc_dat;
  assign psum_reg_and_357_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_92_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_11_sva, pe_0_0_run_cmp_93_psum_out_rsc_z,
      psum_reg_and_357_nl);
  wire [7:0] nl_pe_0_0_run_cmp_92_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_92_weight_rsc_dat = step_mux_78_itm_1;
  wire[0:0] input_reg_and_331_nl;
  wire [7:0] nl_pe_0_0_run_cmp_93_input_in_rsc_dat;
  assign input_reg_and_331_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_93_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_10_sva,
      pe_0_0_run_cmp_109_input_out_rsc_z, input_reg_and_331_nl);
  wire[0:0] psum_reg_and_358_nl;
  wire [15:0] nl_pe_0_0_run_cmp_93_psum_in_rsc_dat;
  assign psum_reg_and_358_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_93_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_11_sva, pe_0_0_run_cmp_94_psum_out_rsc_z,
      psum_reg_and_358_nl);
  wire [7:0] nl_pe_0_0_run_cmp_93_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_93_weight_rsc_dat = step_mux_62_itm_1;
  wire[0:0] input_reg_and_332_nl;
  wire [7:0] nl_pe_0_0_run_cmp_94_input_in_rsc_dat;
  assign input_reg_and_332_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_94_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_10_sva,
      pe_0_0_run_cmp_110_input_out_rsc_z, input_reg_and_332_nl);
  wire[0:0] psum_reg_and_359_nl;
  wire [15:0] nl_pe_0_0_run_cmp_94_psum_in_rsc_dat;
  assign psum_reg_and_359_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_94_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_11_sva, pe_0_0_run_cmp_95_psum_out_rsc_z,
      psum_reg_and_359_nl);
  wire [7:0] nl_pe_0_0_run_cmp_94_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_94_weight_rsc_dat = step_mux_46_itm_1;
  wire[0:0] input_reg_and_333_nl;
  wire [7:0] nl_pe_0_0_run_cmp_95_input_in_rsc_dat;
  assign input_reg_and_333_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_95_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_10_sva,
      pe_0_0_run_cmp_111_input_out_rsc_z, input_reg_and_333_nl);
  wire[0:0] psum_reg_and_360_nl;
  wire [15:0] nl_pe_0_0_run_cmp_95_psum_in_rsc_dat;
  assign psum_reg_and_360_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_95_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_11_sva, pe_0_0_run_cmp_96_psum_out_rsc_z,
      psum_reg_and_360_nl);
  wire [7:0] nl_pe_0_0_run_cmp_95_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_95_weight_rsc_dat = step_mux_30_itm_1;
  wire[0:0] input_reg_and_334_nl;
  wire [7:0] nl_pe_0_0_run_cmp_96_input_in_rsc_dat;
  assign input_reg_and_334_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_96_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_10_sva,
      pe_0_0_run_cmp_112_input_out_rsc_z, input_reg_and_334_nl);
  wire [7:0] nl_pe_0_0_run_cmp_96_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_96_weight_rsc_dat = step_mux_14_itm_1;
  wire[0:0] input_reg_and_335_nl;
  wire [7:0] nl_pe_0_0_run_cmp_97_input_in_rsc_dat;
  assign input_reg_and_335_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_97_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_9_sva,
      pe_0_0_run_cmp_113_input_out_rsc_z, input_reg_and_335_nl);
  wire[0:0] psum_reg_and_361_nl;
  wire [15:0] nl_pe_0_0_run_cmp_97_psum_in_rsc_dat;
  assign psum_reg_and_361_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_97_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_10_sva,
      pe_0_0_run_cmp_98_psum_out_rsc_z, psum_reg_and_361_nl);
  wire [7:0] nl_pe_0_0_run_cmp_97_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_97_weight_rsc_dat = step_mux_253_itm_1;
  wire[0:0] input_reg_and_336_nl;
  wire [7:0] nl_pe_0_0_run_cmp_98_input_in_rsc_dat;
  assign input_reg_and_336_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_98_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_9_sva,
      pe_0_0_run_cmp_114_input_out_rsc_z, input_reg_and_336_nl);
  wire[0:0] psum_reg_and_362_nl;
  wire [15:0] nl_pe_0_0_run_cmp_98_psum_in_rsc_dat;
  assign psum_reg_and_362_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_98_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_10_sva,
      pe_0_0_run_cmp_99_psum_out_rsc_z, psum_reg_and_362_nl);
  wire [7:0] nl_pe_0_0_run_cmp_98_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_98_weight_rsc_dat = step_mux_237_itm_1;
  wire[0:0] input_reg_and_337_nl;
  wire [7:0] nl_pe_0_0_run_cmp_99_input_in_rsc_dat;
  assign input_reg_and_337_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_99_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_9_sva,
      pe_0_0_run_cmp_115_input_out_rsc_z, input_reg_and_337_nl);
  wire[0:0] psum_reg_and_363_nl;
  wire [15:0] nl_pe_0_0_run_cmp_99_psum_in_rsc_dat;
  assign psum_reg_and_363_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_99_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_10_sva,
      pe_0_0_run_cmp_100_psum_out_rsc_z, psum_reg_and_363_nl);
  wire [7:0] nl_pe_0_0_run_cmp_99_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_99_weight_rsc_dat = step_mux_221_itm_1;
  wire[0:0] input_reg_and_338_nl;
  wire [7:0] nl_pe_0_0_run_cmp_100_input_in_rsc_dat;
  assign input_reg_and_338_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_100_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_9_sva,
      pe_0_0_run_cmp_116_input_out_rsc_z, input_reg_and_338_nl);
  wire[0:0] psum_reg_and_364_nl;
  wire [15:0] nl_pe_0_0_run_cmp_100_psum_in_rsc_dat;
  assign psum_reg_and_364_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_100_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_10_sva,
      pe_0_0_run_cmp_101_psum_out_rsc_z, psum_reg_and_364_nl);
  wire [7:0] nl_pe_0_0_run_cmp_100_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_100_weight_rsc_dat = step_mux_205_itm_1;
  wire[0:0] input_reg_and_339_nl;
  wire [7:0] nl_pe_0_0_run_cmp_101_input_in_rsc_dat;
  assign input_reg_and_339_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_101_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_9_sva,
      pe_0_0_run_cmp_117_input_out_rsc_z, input_reg_and_339_nl);
  wire[0:0] psum_reg_and_365_nl;
  wire [15:0] nl_pe_0_0_run_cmp_101_psum_in_rsc_dat;
  assign psum_reg_and_365_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_101_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_10_sva,
      pe_0_0_run_cmp_102_psum_out_rsc_z, psum_reg_and_365_nl);
  wire [7:0] nl_pe_0_0_run_cmp_101_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_101_weight_rsc_dat = step_mux_189_itm_1;
  wire[0:0] input_reg_and_340_nl;
  wire [7:0] nl_pe_0_0_run_cmp_102_input_in_rsc_dat;
  assign input_reg_and_340_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_102_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_9_sva,
      pe_0_0_run_cmp_118_input_out_rsc_z, input_reg_and_340_nl);
  wire[0:0] psum_reg_and_366_nl;
  wire [15:0] nl_pe_0_0_run_cmp_102_psum_in_rsc_dat;
  assign psum_reg_and_366_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_102_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_10_sva,
      pe_0_0_run_cmp_103_psum_out_rsc_z, psum_reg_and_366_nl);
  wire [7:0] nl_pe_0_0_run_cmp_102_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_102_weight_rsc_dat = step_mux_173_itm_1;
  wire[0:0] input_reg_and_341_nl;
  wire [7:0] nl_pe_0_0_run_cmp_103_input_in_rsc_dat;
  assign input_reg_and_341_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_103_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_9_sva,
      pe_0_0_run_cmp_119_input_out_rsc_z, input_reg_and_341_nl);
  wire[0:0] psum_reg_and_367_nl;
  wire [15:0] nl_pe_0_0_run_cmp_103_psum_in_rsc_dat;
  assign psum_reg_and_367_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_103_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_10_sva,
      pe_0_0_run_cmp_104_psum_out_rsc_z, psum_reg_and_367_nl);
  wire [7:0] nl_pe_0_0_run_cmp_103_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_103_weight_rsc_dat = step_mux_157_itm_1;
  wire[0:0] input_reg_and_342_nl;
  wire [7:0] nl_pe_0_0_run_cmp_104_input_in_rsc_dat;
  assign input_reg_and_342_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_104_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_9_sva,
      pe_0_0_run_cmp_120_input_out_rsc_z, input_reg_and_342_nl);
  wire[0:0] psum_reg_and_368_nl;
  wire [15:0] nl_pe_0_0_run_cmp_104_psum_in_rsc_dat;
  assign psum_reg_and_368_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_104_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_10_sva,
      pe_0_0_run_cmp_105_psum_out_rsc_z, psum_reg_and_368_nl);
  wire [7:0] nl_pe_0_0_run_cmp_104_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_104_weight_rsc_dat = step_mux_141_itm_1;
  wire[0:0] input_reg_and_343_nl;
  wire [7:0] nl_pe_0_0_run_cmp_105_input_in_rsc_dat;
  assign input_reg_and_343_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_105_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_9_sva,
      pe_0_0_run_cmp_121_input_out_rsc_z, input_reg_and_343_nl);
  wire[0:0] psum_reg_and_369_nl;
  wire [15:0] nl_pe_0_0_run_cmp_105_psum_in_rsc_dat;
  assign psum_reg_and_369_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_105_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_10_sva,
      pe_0_0_run_cmp_106_psum_out_rsc_z, psum_reg_and_369_nl);
  wire [7:0] nl_pe_0_0_run_cmp_105_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_105_weight_rsc_dat = step_mux_125_itm_1;
  wire[0:0] input_reg_and_344_nl;
  wire [7:0] nl_pe_0_0_run_cmp_106_input_in_rsc_dat;
  assign input_reg_and_344_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_106_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_9_sva,
      pe_0_0_run_cmp_122_input_out_rsc_z, input_reg_and_344_nl);
  wire[0:0] psum_reg_and_370_nl;
  wire [15:0] nl_pe_0_0_run_cmp_106_psum_in_rsc_dat;
  assign psum_reg_and_370_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_106_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_10_sva,
      pe_0_0_run_cmp_107_psum_out_rsc_z, psum_reg_and_370_nl);
  wire [7:0] nl_pe_0_0_run_cmp_106_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_106_weight_rsc_dat = step_mux_109_itm_1;
  wire[0:0] input_reg_and_345_nl;
  wire [7:0] nl_pe_0_0_run_cmp_107_input_in_rsc_dat;
  assign input_reg_and_345_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_107_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_9_sva,
      pe_0_0_run_cmp_123_input_out_rsc_z, input_reg_and_345_nl);
  wire[0:0] psum_reg_and_371_nl;
  wire [15:0] nl_pe_0_0_run_cmp_107_psum_in_rsc_dat;
  assign psum_reg_and_371_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_107_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_10_sva,
      pe_0_0_run_cmp_108_psum_out_rsc_z, psum_reg_and_371_nl);
  wire [7:0] nl_pe_0_0_run_cmp_107_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_107_weight_rsc_dat = step_mux_93_itm_1;
  wire[0:0] input_reg_and_346_nl;
  wire [7:0] nl_pe_0_0_run_cmp_108_input_in_rsc_dat;
  assign input_reg_and_346_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_108_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_9_sva,
      pe_0_0_run_cmp_124_input_out_rsc_z, input_reg_and_346_nl);
  wire[0:0] psum_reg_and_372_nl;
  wire [15:0] nl_pe_0_0_run_cmp_108_psum_in_rsc_dat;
  assign psum_reg_and_372_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_108_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_10_sva,
      pe_0_0_run_cmp_109_psum_out_rsc_z, psum_reg_and_372_nl);
  wire [7:0] nl_pe_0_0_run_cmp_108_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_108_weight_rsc_dat = step_mux_77_itm_1;
  wire[0:0] input_reg_and_347_nl;
  wire [7:0] nl_pe_0_0_run_cmp_109_input_in_rsc_dat;
  assign input_reg_and_347_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_109_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_9_sva,
      pe_0_0_run_cmp_125_input_out_rsc_z, input_reg_and_347_nl);
  wire[0:0] psum_reg_and_373_nl;
  wire [15:0] nl_pe_0_0_run_cmp_109_psum_in_rsc_dat;
  assign psum_reg_and_373_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_109_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_10_sva,
      pe_0_0_run_cmp_110_psum_out_rsc_z, psum_reg_and_373_nl);
  wire [7:0] nl_pe_0_0_run_cmp_109_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_109_weight_rsc_dat = step_mux_61_itm_1;
  wire[0:0] input_reg_and_348_nl;
  wire [7:0] nl_pe_0_0_run_cmp_110_input_in_rsc_dat;
  assign input_reg_and_348_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_110_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_9_sva,
      pe_0_0_run_cmp_126_input_out_rsc_z, input_reg_and_348_nl);
  wire[0:0] psum_reg_and_374_nl;
  wire [15:0] nl_pe_0_0_run_cmp_110_psum_in_rsc_dat;
  assign psum_reg_and_374_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_110_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_10_sva,
      pe_0_0_run_cmp_111_psum_out_rsc_z, psum_reg_and_374_nl);
  wire [7:0] nl_pe_0_0_run_cmp_110_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_110_weight_rsc_dat = step_mux_45_itm_1;
  wire[0:0] input_reg_and_349_nl;
  wire [7:0] nl_pe_0_0_run_cmp_111_input_in_rsc_dat;
  assign input_reg_and_349_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_111_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_9_sva,
      pe_0_0_run_cmp_127_input_out_rsc_z, input_reg_and_349_nl);
  wire[0:0] psum_reg_and_375_nl;
  wire [15:0] nl_pe_0_0_run_cmp_111_psum_in_rsc_dat;
  assign psum_reg_and_375_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_111_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_10_sva,
      pe_0_0_run_cmp_112_psum_out_rsc_z, psum_reg_and_375_nl);
  wire [7:0] nl_pe_0_0_run_cmp_111_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_111_weight_rsc_dat = step_mux_29_itm_1;
  wire[0:0] input_reg_and_350_nl;
  wire [7:0] nl_pe_0_0_run_cmp_112_input_in_rsc_dat;
  assign input_reg_and_350_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_112_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_9_sva,
      pe_0_0_run_cmp_128_input_out_rsc_z, input_reg_and_350_nl);
  wire [7:0] nl_pe_0_0_run_cmp_112_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_112_weight_rsc_dat = step_mux_13_itm_1;
  wire[0:0] input_reg_and_351_nl;
  wire [7:0] nl_pe_0_0_run_cmp_113_input_in_rsc_dat;
  assign input_reg_and_351_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_113_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_8_sva,
      pe_0_0_run_cmp_129_input_out_rsc_z, input_reg_and_351_nl);
  wire[0:0] psum_reg_and_376_nl;
  wire [15:0] nl_pe_0_0_run_cmp_113_psum_in_rsc_dat;
  assign psum_reg_and_376_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_113_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_9_sva,
      pe_0_0_run_cmp_114_psum_out_rsc_z, psum_reg_and_376_nl);
  wire [7:0] nl_pe_0_0_run_cmp_113_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_113_weight_rsc_dat = step_mux_252_itm_1;
  wire[0:0] input_reg_and_352_nl;
  wire [7:0] nl_pe_0_0_run_cmp_114_input_in_rsc_dat;
  assign input_reg_and_352_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_114_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_8_sva,
      pe_0_0_run_cmp_130_input_out_rsc_z, input_reg_and_352_nl);
  wire[0:0] psum_reg_and_377_nl;
  wire [15:0] nl_pe_0_0_run_cmp_114_psum_in_rsc_dat;
  assign psum_reg_and_377_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_114_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_9_sva,
      pe_0_0_run_cmp_115_psum_out_rsc_z, psum_reg_and_377_nl);
  wire [7:0] nl_pe_0_0_run_cmp_114_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_114_weight_rsc_dat = step_mux_236_itm_1;
  wire[0:0] input_reg_and_353_nl;
  wire [7:0] nl_pe_0_0_run_cmp_115_input_in_rsc_dat;
  assign input_reg_and_353_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_115_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_8_sva,
      pe_0_0_run_cmp_131_input_out_rsc_z, input_reg_and_353_nl);
  wire[0:0] psum_reg_and_378_nl;
  wire [15:0] nl_pe_0_0_run_cmp_115_psum_in_rsc_dat;
  assign psum_reg_and_378_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_115_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_9_sva,
      pe_0_0_run_cmp_116_psum_out_rsc_z, psum_reg_and_378_nl);
  wire [7:0] nl_pe_0_0_run_cmp_115_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_115_weight_rsc_dat = step_mux_220_itm_1;
  wire[0:0] input_reg_and_354_nl;
  wire [7:0] nl_pe_0_0_run_cmp_116_input_in_rsc_dat;
  assign input_reg_and_354_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_116_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_8_sva,
      pe_0_0_run_cmp_132_input_out_rsc_z, input_reg_and_354_nl);
  wire[0:0] psum_reg_and_379_nl;
  wire [15:0] nl_pe_0_0_run_cmp_116_psum_in_rsc_dat;
  assign psum_reg_and_379_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_116_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_9_sva,
      pe_0_0_run_cmp_117_psum_out_rsc_z, psum_reg_and_379_nl);
  wire [7:0] nl_pe_0_0_run_cmp_116_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_116_weight_rsc_dat = step_mux_204_itm_1;
  wire[0:0] input_reg_and_355_nl;
  wire [7:0] nl_pe_0_0_run_cmp_117_input_in_rsc_dat;
  assign input_reg_and_355_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_117_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_8_sva,
      pe_0_0_run_cmp_133_input_out_rsc_z, input_reg_and_355_nl);
  wire[0:0] psum_reg_and_380_nl;
  wire [15:0] nl_pe_0_0_run_cmp_117_psum_in_rsc_dat;
  assign psum_reg_and_380_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_117_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_9_sva,
      pe_0_0_run_cmp_118_psum_out_rsc_z, psum_reg_and_380_nl);
  wire [7:0] nl_pe_0_0_run_cmp_117_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_117_weight_rsc_dat = step_mux_188_itm_1;
  wire[0:0] input_reg_and_356_nl;
  wire [7:0] nl_pe_0_0_run_cmp_118_input_in_rsc_dat;
  assign input_reg_and_356_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_118_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_8_sva,
      pe_0_0_run_cmp_134_input_out_rsc_z, input_reg_and_356_nl);
  wire[0:0] psum_reg_and_381_nl;
  wire [15:0] nl_pe_0_0_run_cmp_118_psum_in_rsc_dat;
  assign psum_reg_and_381_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_118_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_9_sva,
      pe_0_0_run_cmp_119_psum_out_rsc_z, psum_reg_and_381_nl);
  wire [7:0] nl_pe_0_0_run_cmp_118_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_118_weight_rsc_dat = step_mux_172_itm_1;
  wire[0:0] input_reg_and_357_nl;
  wire [7:0] nl_pe_0_0_run_cmp_119_input_in_rsc_dat;
  assign input_reg_and_357_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_119_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_8_sva,
      pe_0_0_run_cmp_135_input_out_rsc_z, input_reg_and_357_nl);
  wire[0:0] psum_reg_and_382_nl;
  wire [15:0] nl_pe_0_0_run_cmp_119_psum_in_rsc_dat;
  assign psum_reg_and_382_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_119_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_9_sva, pe_0_0_run_cmp_120_psum_out_rsc_z,
      psum_reg_and_382_nl);
  wire [7:0] nl_pe_0_0_run_cmp_119_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_119_weight_rsc_dat = step_mux_156_itm_1;
  wire[0:0] input_reg_and_358_nl;
  wire [7:0] nl_pe_0_0_run_cmp_120_input_in_rsc_dat;
  assign input_reg_and_358_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_120_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_8_sva,
      pe_0_0_run_cmp_136_input_out_rsc_z, input_reg_and_358_nl);
  wire[0:0] psum_reg_and_383_nl;
  wire [15:0] nl_pe_0_0_run_cmp_120_psum_in_rsc_dat;
  assign psum_reg_and_383_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_120_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_9_sva, pe_0_0_run_cmp_121_psum_out_rsc_z,
      psum_reg_and_383_nl);
  wire [7:0] nl_pe_0_0_run_cmp_120_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_120_weight_rsc_dat = step_mux_140_itm_1;
  wire[0:0] input_reg_and_359_nl;
  wire [7:0] nl_pe_0_0_run_cmp_121_input_in_rsc_dat;
  assign input_reg_and_359_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_121_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_8_sva,
      pe_0_0_run_cmp_137_input_out_rsc_z, input_reg_and_359_nl);
  wire[0:0] psum_reg_and_384_nl;
  wire [15:0] nl_pe_0_0_run_cmp_121_psum_in_rsc_dat;
  assign psum_reg_and_384_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_121_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_9_sva, pe_0_0_run_cmp_122_psum_out_rsc_z,
      psum_reg_and_384_nl);
  wire [7:0] nl_pe_0_0_run_cmp_121_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_121_weight_rsc_dat = step_mux_124_itm_1;
  wire[0:0] input_reg_and_360_nl;
  wire [7:0] nl_pe_0_0_run_cmp_122_input_in_rsc_dat;
  assign input_reg_and_360_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_122_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_8_sva,
      pe_0_0_run_cmp_138_input_out_rsc_z, input_reg_and_360_nl);
  wire[0:0] psum_reg_and_385_nl;
  wire [15:0] nl_pe_0_0_run_cmp_122_psum_in_rsc_dat;
  assign psum_reg_and_385_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_122_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_9_sva, pe_0_0_run_cmp_123_psum_out_rsc_z,
      psum_reg_and_385_nl);
  wire [7:0] nl_pe_0_0_run_cmp_122_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_122_weight_rsc_dat = step_mux_108_itm_1;
  wire[0:0] input_reg_and_361_nl;
  wire [7:0] nl_pe_0_0_run_cmp_123_input_in_rsc_dat;
  assign input_reg_and_361_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_123_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_8_sva,
      pe_0_0_run_cmp_139_input_out_rsc_z, input_reg_and_361_nl);
  wire[0:0] psum_reg_and_386_nl;
  wire [15:0] nl_pe_0_0_run_cmp_123_psum_in_rsc_dat;
  assign psum_reg_and_386_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_123_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_9_sva, pe_0_0_run_cmp_124_psum_out_rsc_z,
      psum_reg_and_386_nl);
  wire [7:0] nl_pe_0_0_run_cmp_123_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_123_weight_rsc_dat = step_mux_92_itm_1;
  wire[0:0] input_reg_and_362_nl;
  wire [7:0] nl_pe_0_0_run_cmp_124_input_in_rsc_dat;
  assign input_reg_and_362_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_124_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_8_sva,
      pe_0_0_run_cmp_140_input_out_rsc_z, input_reg_and_362_nl);
  wire[0:0] psum_reg_and_387_nl;
  wire [15:0] nl_pe_0_0_run_cmp_124_psum_in_rsc_dat;
  assign psum_reg_and_387_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_124_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_9_sva, pe_0_0_run_cmp_125_psum_out_rsc_z,
      psum_reg_and_387_nl);
  wire [7:0] nl_pe_0_0_run_cmp_124_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_124_weight_rsc_dat = step_mux_76_itm_1;
  wire[0:0] input_reg_and_363_nl;
  wire [7:0] nl_pe_0_0_run_cmp_125_input_in_rsc_dat;
  assign input_reg_and_363_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_125_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_8_sva,
      pe_0_0_run_cmp_141_input_out_rsc_z, input_reg_and_363_nl);
  wire[0:0] psum_reg_and_388_nl;
  wire [15:0] nl_pe_0_0_run_cmp_125_psum_in_rsc_dat;
  assign psum_reg_and_388_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_125_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_9_sva, pe_0_0_run_cmp_126_psum_out_rsc_z,
      psum_reg_and_388_nl);
  wire [7:0] nl_pe_0_0_run_cmp_125_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_125_weight_rsc_dat = step_mux_60_itm_1;
  wire[0:0] input_reg_and_364_nl;
  wire [7:0] nl_pe_0_0_run_cmp_126_input_in_rsc_dat;
  assign input_reg_and_364_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_126_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_8_sva,
      pe_0_0_run_cmp_142_input_out_rsc_z, input_reg_and_364_nl);
  wire[0:0] psum_reg_and_389_nl;
  wire [15:0] nl_pe_0_0_run_cmp_126_psum_in_rsc_dat;
  assign psum_reg_and_389_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_126_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_9_sva, pe_0_0_run_cmp_127_psum_out_rsc_z,
      psum_reg_and_389_nl);
  wire [7:0] nl_pe_0_0_run_cmp_126_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_126_weight_rsc_dat = step_mux_44_itm_1;
  wire[0:0] input_reg_and_365_nl;
  wire [7:0] nl_pe_0_0_run_cmp_127_input_in_rsc_dat;
  assign input_reg_and_365_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_127_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_8_sva,
      pe_0_0_run_cmp_143_input_out_rsc_z, input_reg_and_365_nl);
  wire[0:0] psum_reg_and_390_nl;
  wire [15:0] nl_pe_0_0_run_cmp_127_psum_in_rsc_dat;
  assign psum_reg_and_390_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_127_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_9_sva, pe_0_0_run_cmp_128_psum_out_rsc_z,
      psum_reg_and_390_nl);
  wire [7:0] nl_pe_0_0_run_cmp_127_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_127_weight_rsc_dat = step_mux_28_itm_1;
  wire[0:0] input_reg_and_366_nl;
  wire [7:0] nl_pe_0_0_run_cmp_128_input_in_rsc_dat;
  assign input_reg_and_366_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_128_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_8_sva,
      pe_0_0_run_cmp_144_input_out_rsc_z, input_reg_and_366_nl);
  wire [7:0] nl_pe_0_0_run_cmp_128_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_128_weight_rsc_dat = step_mux_12_itm_1;
  wire[0:0] input_reg_and_367_nl;
  wire [7:0] nl_pe_0_0_run_cmp_129_input_in_rsc_dat;
  assign input_reg_and_367_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_129_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_7_sva,
      pe_0_0_run_cmp_145_input_out_rsc_z, input_reg_and_367_nl);
  wire[0:0] psum_reg_and_391_nl;
  wire [15:0] nl_pe_0_0_run_cmp_129_psum_in_rsc_dat;
  assign psum_reg_and_391_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_129_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_8_sva,
      pe_0_0_run_cmp_130_psum_out_rsc_z, psum_reg_and_391_nl);
  wire [7:0] nl_pe_0_0_run_cmp_129_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_129_weight_rsc_dat = step_mux_251_itm_1;
  wire[0:0] input_reg_and_368_nl;
  wire [7:0] nl_pe_0_0_run_cmp_130_input_in_rsc_dat;
  assign input_reg_and_368_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_130_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_7_sva,
      pe_0_0_run_cmp_146_input_out_rsc_z, input_reg_and_368_nl);
  wire[0:0] psum_reg_and_392_nl;
  wire [15:0] nl_pe_0_0_run_cmp_130_psum_in_rsc_dat;
  assign psum_reg_and_392_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_130_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_8_sva,
      pe_0_0_run_cmp_131_psum_out_rsc_z, psum_reg_and_392_nl);
  wire [7:0] nl_pe_0_0_run_cmp_130_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_130_weight_rsc_dat = step_mux_235_itm_1;
  wire[0:0] input_reg_and_369_nl;
  wire [7:0] nl_pe_0_0_run_cmp_131_input_in_rsc_dat;
  assign input_reg_and_369_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_131_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_7_sva,
      pe_0_0_run_cmp_147_input_out_rsc_z, input_reg_and_369_nl);
  wire[0:0] psum_reg_and_393_nl;
  wire [15:0] nl_pe_0_0_run_cmp_131_psum_in_rsc_dat;
  assign psum_reg_and_393_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_131_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_8_sva,
      pe_0_0_run_cmp_132_psum_out_rsc_z, psum_reg_and_393_nl);
  wire [7:0] nl_pe_0_0_run_cmp_131_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_131_weight_rsc_dat = step_mux_219_itm_1;
  wire[0:0] input_reg_and_370_nl;
  wire [7:0] nl_pe_0_0_run_cmp_132_input_in_rsc_dat;
  assign input_reg_and_370_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_132_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_7_sva,
      pe_0_0_run_cmp_148_input_out_rsc_z, input_reg_and_370_nl);
  wire[0:0] psum_reg_and_394_nl;
  wire [15:0] nl_pe_0_0_run_cmp_132_psum_in_rsc_dat;
  assign psum_reg_and_394_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_132_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_8_sva,
      pe_0_0_run_cmp_133_psum_out_rsc_z, psum_reg_and_394_nl);
  wire [7:0] nl_pe_0_0_run_cmp_132_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_132_weight_rsc_dat = step_mux_203_itm_1;
  wire[0:0] input_reg_and_371_nl;
  wire [7:0] nl_pe_0_0_run_cmp_133_input_in_rsc_dat;
  assign input_reg_and_371_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_133_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_7_sva,
      pe_0_0_run_cmp_149_input_out_rsc_z, input_reg_and_371_nl);
  wire[0:0] psum_reg_and_395_nl;
  wire [15:0] nl_pe_0_0_run_cmp_133_psum_in_rsc_dat;
  assign psum_reg_and_395_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_133_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_8_sva,
      pe_0_0_run_cmp_134_psum_out_rsc_z, psum_reg_and_395_nl);
  wire [7:0] nl_pe_0_0_run_cmp_133_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_133_weight_rsc_dat = step_mux_187_itm_1;
  wire[0:0] input_reg_and_372_nl;
  wire [7:0] nl_pe_0_0_run_cmp_134_input_in_rsc_dat;
  assign input_reg_and_372_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_134_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_7_sva,
      pe_0_0_run_cmp_150_input_out_rsc_z, input_reg_and_372_nl);
  wire[0:0] psum_reg_and_396_nl;
  wire [15:0] nl_pe_0_0_run_cmp_134_psum_in_rsc_dat;
  assign psum_reg_and_396_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_134_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_8_sva,
      pe_0_0_run_cmp_135_psum_out_rsc_z, psum_reg_and_396_nl);
  wire [7:0] nl_pe_0_0_run_cmp_134_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_134_weight_rsc_dat = step_mux_171_itm_1;
  wire[0:0] input_reg_and_373_nl;
  wire [7:0] nl_pe_0_0_run_cmp_135_input_in_rsc_dat;
  assign input_reg_and_373_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_135_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_7_sva,
      pe_0_0_run_cmp_151_input_out_rsc_z, input_reg_and_373_nl);
  wire[0:0] psum_reg_and_397_nl;
  wire [15:0] nl_pe_0_0_run_cmp_135_psum_in_rsc_dat;
  assign psum_reg_and_397_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_135_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_8_sva, pe_0_0_run_cmp_136_psum_out_rsc_z,
      psum_reg_and_397_nl);
  wire [7:0] nl_pe_0_0_run_cmp_135_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_135_weight_rsc_dat = step_mux_155_itm_1;
  wire[0:0] input_reg_and_374_nl;
  wire [7:0] nl_pe_0_0_run_cmp_136_input_in_rsc_dat;
  assign input_reg_and_374_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_136_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_7_sva,
      pe_0_0_run_cmp_152_input_out_rsc_z, input_reg_and_374_nl);
  wire[0:0] psum_reg_and_398_nl;
  wire [15:0] nl_pe_0_0_run_cmp_136_psum_in_rsc_dat;
  assign psum_reg_and_398_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_136_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_8_sva, pe_0_0_run_cmp_137_psum_out_rsc_z,
      psum_reg_and_398_nl);
  wire [7:0] nl_pe_0_0_run_cmp_136_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_136_weight_rsc_dat = step_mux_139_itm_1;
  wire[0:0] input_reg_and_375_nl;
  wire [7:0] nl_pe_0_0_run_cmp_137_input_in_rsc_dat;
  assign input_reg_and_375_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_137_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_7_sva,
      pe_0_0_run_cmp_153_input_out_rsc_z, input_reg_and_375_nl);
  wire[0:0] psum_reg_and_399_nl;
  wire [15:0] nl_pe_0_0_run_cmp_137_psum_in_rsc_dat;
  assign psum_reg_and_399_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_137_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_8_sva, pe_0_0_run_cmp_138_psum_out_rsc_z,
      psum_reg_and_399_nl);
  wire [7:0] nl_pe_0_0_run_cmp_137_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_137_weight_rsc_dat = step_mux_123_itm_1;
  wire[0:0] input_reg_and_376_nl;
  wire [7:0] nl_pe_0_0_run_cmp_138_input_in_rsc_dat;
  assign input_reg_and_376_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_138_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_7_sva,
      pe_0_0_run_cmp_154_input_out_rsc_z, input_reg_and_376_nl);
  wire[0:0] psum_reg_and_400_nl;
  wire [15:0] nl_pe_0_0_run_cmp_138_psum_in_rsc_dat;
  assign psum_reg_and_400_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_138_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_8_sva, pe_0_0_run_cmp_139_psum_out_rsc_z,
      psum_reg_and_400_nl);
  wire [7:0] nl_pe_0_0_run_cmp_138_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_138_weight_rsc_dat = step_mux_107_itm_1;
  wire[0:0] input_reg_and_377_nl;
  wire [7:0] nl_pe_0_0_run_cmp_139_input_in_rsc_dat;
  assign input_reg_and_377_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_139_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_7_sva,
      pe_0_0_run_cmp_155_input_out_rsc_z, input_reg_and_377_nl);
  wire[0:0] psum_reg_and_401_nl;
  wire [15:0] nl_pe_0_0_run_cmp_139_psum_in_rsc_dat;
  assign psum_reg_and_401_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_139_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_8_sva, pe_0_0_run_cmp_140_psum_out_rsc_z,
      psum_reg_and_401_nl);
  wire [7:0] nl_pe_0_0_run_cmp_139_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_139_weight_rsc_dat = step_mux_91_itm_1;
  wire[0:0] input_reg_and_378_nl;
  wire [7:0] nl_pe_0_0_run_cmp_140_input_in_rsc_dat;
  assign input_reg_and_378_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_140_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_7_sva,
      pe_0_0_run_cmp_156_input_out_rsc_z, input_reg_and_378_nl);
  wire[0:0] psum_reg_and_402_nl;
  wire [15:0] nl_pe_0_0_run_cmp_140_psum_in_rsc_dat;
  assign psum_reg_and_402_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_140_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_8_sva, pe_0_0_run_cmp_141_psum_out_rsc_z,
      psum_reg_and_402_nl);
  wire [7:0] nl_pe_0_0_run_cmp_140_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_140_weight_rsc_dat = step_mux_75_itm_1;
  wire[0:0] input_reg_and_379_nl;
  wire [7:0] nl_pe_0_0_run_cmp_141_input_in_rsc_dat;
  assign input_reg_and_379_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_141_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_7_sva,
      pe_0_0_run_cmp_157_input_out_rsc_z, input_reg_and_379_nl);
  wire[0:0] psum_reg_and_403_nl;
  wire [15:0] nl_pe_0_0_run_cmp_141_psum_in_rsc_dat;
  assign psum_reg_and_403_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_141_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_8_sva, pe_0_0_run_cmp_142_psum_out_rsc_z,
      psum_reg_and_403_nl);
  wire [7:0] nl_pe_0_0_run_cmp_141_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_141_weight_rsc_dat = step_mux_59_itm_1;
  wire[0:0] input_reg_and_380_nl;
  wire [7:0] nl_pe_0_0_run_cmp_142_input_in_rsc_dat;
  assign input_reg_and_380_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_142_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_7_sva,
      pe_0_0_run_cmp_158_input_out_rsc_z, input_reg_and_380_nl);
  wire[0:0] psum_reg_and_404_nl;
  wire [15:0] nl_pe_0_0_run_cmp_142_psum_in_rsc_dat;
  assign psum_reg_and_404_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_142_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_8_sva, pe_0_0_run_cmp_143_psum_out_rsc_z,
      psum_reg_and_404_nl);
  wire [7:0] nl_pe_0_0_run_cmp_142_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_142_weight_rsc_dat = step_mux_43_itm_1;
  wire[0:0] input_reg_and_381_nl;
  wire [7:0] nl_pe_0_0_run_cmp_143_input_in_rsc_dat;
  assign input_reg_and_381_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_143_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_7_sva,
      pe_0_0_run_cmp_159_input_out_rsc_z, input_reg_and_381_nl);
  wire[0:0] psum_reg_and_405_nl;
  wire [15:0] nl_pe_0_0_run_cmp_143_psum_in_rsc_dat;
  assign psum_reg_and_405_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_143_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_8_sva, pe_0_0_run_cmp_144_psum_out_rsc_z,
      psum_reg_and_405_nl);
  wire [7:0] nl_pe_0_0_run_cmp_143_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_143_weight_rsc_dat = step_mux_27_itm_1;
  wire[0:0] input_reg_and_382_nl;
  wire [7:0] nl_pe_0_0_run_cmp_144_input_in_rsc_dat;
  assign input_reg_and_382_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_144_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_7_sva,
      pe_0_0_run_cmp_160_input_out_rsc_z, input_reg_and_382_nl);
  wire [7:0] nl_pe_0_0_run_cmp_144_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_144_weight_rsc_dat = step_mux_11_itm_1;
  wire[0:0] input_reg_and_383_nl;
  wire [7:0] nl_pe_0_0_run_cmp_145_input_in_rsc_dat;
  assign input_reg_and_383_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_145_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_6_sva,
      pe_0_0_run_cmp_161_input_out_rsc_z, input_reg_and_383_nl);
  wire[0:0] psum_reg_and_406_nl;
  wire [15:0] nl_pe_0_0_run_cmp_145_psum_in_rsc_dat;
  assign psum_reg_and_406_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_145_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_7_sva,
      pe_0_0_run_cmp_146_psum_out_rsc_z, psum_reg_and_406_nl);
  wire [7:0] nl_pe_0_0_run_cmp_145_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_145_weight_rsc_dat = step_mux_250_itm_1;
  wire[0:0] input_reg_and_384_nl;
  wire [7:0] nl_pe_0_0_run_cmp_146_input_in_rsc_dat;
  assign input_reg_and_384_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_146_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_6_sva,
      pe_0_0_run_cmp_162_input_out_rsc_z, input_reg_and_384_nl);
  wire[0:0] psum_reg_and_407_nl;
  wire [15:0] nl_pe_0_0_run_cmp_146_psum_in_rsc_dat;
  assign psum_reg_and_407_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_146_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_7_sva,
      pe_0_0_run_cmp_147_psum_out_rsc_z, psum_reg_and_407_nl);
  wire [7:0] nl_pe_0_0_run_cmp_146_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_146_weight_rsc_dat = step_mux_234_itm_1;
  wire[0:0] input_reg_and_385_nl;
  wire [7:0] nl_pe_0_0_run_cmp_147_input_in_rsc_dat;
  assign input_reg_and_385_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_147_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_6_sva,
      pe_0_0_run_cmp_163_input_out_rsc_z, input_reg_and_385_nl);
  wire[0:0] psum_reg_and_408_nl;
  wire [15:0] nl_pe_0_0_run_cmp_147_psum_in_rsc_dat;
  assign psum_reg_and_408_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_147_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_7_sva,
      pe_0_0_run_cmp_148_psum_out_rsc_z, psum_reg_and_408_nl);
  wire [7:0] nl_pe_0_0_run_cmp_147_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_147_weight_rsc_dat = step_mux_218_itm_1;
  wire[0:0] input_reg_and_386_nl;
  wire [7:0] nl_pe_0_0_run_cmp_148_input_in_rsc_dat;
  assign input_reg_and_386_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_148_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_6_sva,
      pe_0_0_run_cmp_164_input_out_rsc_z, input_reg_and_386_nl);
  wire[0:0] psum_reg_and_409_nl;
  wire [15:0] nl_pe_0_0_run_cmp_148_psum_in_rsc_dat;
  assign psum_reg_and_409_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_148_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_7_sva,
      pe_0_0_run_cmp_149_psum_out_rsc_z, psum_reg_and_409_nl);
  wire [7:0] nl_pe_0_0_run_cmp_148_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_148_weight_rsc_dat = step_mux_202_itm_1;
  wire[0:0] input_reg_and_387_nl;
  wire [7:0] nl_pe_0_0_run_cmp_149_input_in_rsc_dat;
  assign input_reg_and_387_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_149_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_6_sva,
      pe_0_0_run_cmp_165_input_out_rsc_z, input_reg_and_387_nl);
  wire[0:0] psum_reg_and_410_nl;
  wire [15:0] nl_pe_0_0_run_cmp_149_psum_in_rsc_dat;
  assign psum_reg_and_410_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_149_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_7_sva,
      pe_0_0_run_cmp_150_psum_out_rsc_z, psum_reg_and_410_nl);
  wire [7:0] nl_pe_0_0_run_cmp_149_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_149_weight_rsc_dat = step_mux_186_itm_1;
  wire[0:0] input_reg_and_388_nl;
  wire [7:0] nl_pe_0_0_run_cmp_150_input_in_rsc_dat;
  assign input_reg_and_388_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_150_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_6_sva,
      pe_0_0_run_cmp_166_input_out_rsc_z, input_reg_and_388_nl);
  wire[0:0] psum_reg_and_411_nl;
  wire [15:0] nl_pe_0_0_run_cmp_150_psum_in_rsc_dat;
  assign psum_reg_and_411_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_150_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_7_sva,
      pe_0_0_run_cmp_151_psum_out_rsc_z, psum_reg_and_411_nl);
  wire [7:0] nl_pe_0_0_run_cmp_150_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_150_weight_rsc_dat = step_mux_170_itm_1;
  wire[0:0] input_reg_and_389_nl;
  wire [7:0] nl_pe_0_0_run_cmp_151_input_in_rsc_dat;
  assign input_reg_and_389_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_151_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_6_sva,
      pe_0_0_run_cmp_167_input_out_rsc_z, input_reg_and_389_nl);
  wire[0:0] psum_reg_and_412_nl;
  wire [15:0] nl_pe_0_0_run_cmp_151_psum_in_rsc_dat;
  assign psum_reg_and_412_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_151_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_7_sva, pe_0_0_run_cmp_152_psum_out_rsc_z,
      psum_reg_and_412_nl);
  wire [7:0] nl_pe_0_0_run_cmp_151_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_151_weight_rsc_dat = step_mux_154_itm_1;
  wire[0:0] input_reg_and_390_nl;
  wire [7:0] nl_pe_0_0_run_cmp_152_input_in_rsc_dat;
  assign input_reg_and_390_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_152_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_6_sva,
      pe_0_0_run_cmp_168_input_out_rsc_z, input_reg_and_390_nl);
  wire[0:0] psum_reg_and_413_nl;
  wire [15:0] nl_pe_0_0_run_cmp_152_psum_in_rsc_dat;
  assign psum_reg_and_413_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_152_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_7_sva, pe_0_0_run_cmp_153_psum_out_rsc_z,
      psum_reg_and_413_nl);
  wire [7:0] nl_pe_0_0_run_cmp_152_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_152_weight_rsc_dat = step_mux_138_itm_1;
  wire[0:0] input_reg_and_391_nl;
  wire [7:0] nl_pe_0_0_run_cmp_153_input_in_rsc_dat;
  assign input_reg_and_391_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_153_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_6_sva,
      pe_0_0_run_cmp_169_input_out_rsc_z, input_reg_and_391_nl);
  wire[0:0] psum_reg_and_414_nl;
  wire [15:0] nl_pe_0_0_run_cmp_153_psum_in_rsc_dat;
  assign psum_reg_and_414_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_153_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_7_sva, pe_0_0_run_cmp_154_psum_out_rsc_z,
      psum_reg_and_414_nl);
  wire [7:0] nl_pe_0_0_run_cmp_153_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_153_weight_rsc_dat = step_mux_122_itm_1;
  wire[0:0] input_reg_and_392_nl;
  wire [7:0] nl_pe_0_0_run_cmp_154_input_in_rsc_dat;
  assign input_reg_and_392_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_154_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_6_sva,
      pe_0_0_run_cmp_170_input_out_rsc_z, input_reg_and_392_nl);
  wire[0:0] psum_reg_and_415_nl;
  wire [15:0] nl_pe_0_0_run_cmp_154_psum_in_rsc_dat;
  assign psum_reg_and_415_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_154_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_7_sva, pe_0_0_run_cmp_155_psum_out_rsc_z,
      psum_reg_and_415_nl);
  wire [7:0] nl_pe_0_0_run_cmp_154_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_154_weight_rsc_dat = step_mux_106_itm_1;
  wire[0:0] input_reg_and_393_nl;
  wire [7:0] nl_pe_0_0_run_cmp_155_input_in_rsc_dat;
  assign input_reg_and_393_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_155_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_6_sva,
      pe_0_0_run_cmp_171_input_out_rsc_z, input_reg_and_393_nl);
  wire[0:0] psum_reg_and_416_nl;
  wire [15:0] nl_pe_0_0_run_cmp_155_psum_in_rsc_dat;
  assign psum_reg_and_416_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_155_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_7_sva, pe_0_0_run_cmp_156_psum_out_rsc_z,
      psum_reg_and_416_nl);
  wire [7:0] nl_pe_0_0_run_cmp_155_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_155_weight_rsc_dat = step_mux_90_itm_1;
  wire[0:0] input_reg_and_394_nl;
  wire [7:0] nl_pe_0_0_run_cmp_156_input_in_rsc_dat;
  assign input_reg_and_394_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_156_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_6_sva,
      pe_0_0_run_cmp_172_input_out_rsc_z, input_reg_and_394_nl);
  wire[0:0] psum_reg_and_417_nl;
  wire [15:0] nl_pe_0_0_run_cmp_156_psum_in_rsc_dat;
  assign psum_reg_and_417_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_156_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_7_sva, pe_0_0_run_cmp_157_psum_out_rsc_z,
      psum_reg_and_417_nl);
  wire [7:0] nl_pe_0_0_run_cmp_156_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_156_weight_rsc_dat = step_mux_74_itm_1;
  wire[0:0] input_reg_and_395_nl;
  wire [7:0] nl_pe_0_0_run_cmp_157_input_in_rsc_dat;
  assign input_reg_and_395_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_157_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_6_sva,
      pe_0_0_run_cmp_173_input_out_rsc_z, input_reg_and_395_nl);
  wire[0:0] psum_reg_and_418_nl;
  wire [15:0] nl_pe_0_0_run_cmp_157_psum_in_rsc_dat;
  assign psum_reg_and_418_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_157_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_7_sva, pe_0_0_run_cmp_158_psum_out_rsc_z,
      psum_reg_and_418_nl);
  wire [7:0] nl_pe_0_0_run_cmp_157_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_157_weight_rsc_dat = step_mux_58_itm_1;
  wire[0:0] input_reg_and_396_nl;
  wire [7:0] nl_pe_0_0_run_cmp_158_input_in_rsc_dat;
  assign input_reg_and_396_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_158_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_6_sva,
      pe_0_0_run_cmp_174_input_out_rsc_z, input_reg_and_396_nl);
  wire[0:0] psum_reg_and_419_nl;
  wire [15:0] nl_pe_0_0_run_cmp_158_psum_in_rsc_dat;
  assign psum_reg_and_419_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_158_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_7_sva, pe_0_0_run_cmp_159_psum_out_rsc_z,
      psum_reg_and_419_nl);
  wire [7:0] nl_pe_0_0_run_cmp_158_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_158_weight_rsc_dat = step_mux_42_itm_1;
  wire[0:0] input_reg_and_397_nl;
  wire [7:0] nl_pe_0_0_run_cmp_159_input_in_rsc_dat;
  assign input_reg_and_397_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_159_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_6_sva,
      pe_0_0_run_cmp_175_input_out_rsc_z, input_reg_and_397_nl);
  wire[0:0] psum_reg_and_420_nl;
  wire [15:0] nl_pe_0_0_run_cmp_159_psum_in_rsc_dat;
  assign psum_reg_and_420_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_159_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_7_sva, pe_0_0_run_cmp_160_psum_out_rsc_z,
      psum_reg_and_420_nl);
  wire [7:0] nl_pe_0_0_run_cmp_159_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_159_weight_rsc_dat = step_mux_26_itm_1;
  wire[0:0] input_reg_and_398_nl;
  wire [7:0] nl_pe_0_0_run_cmp_160_input_in_rsc_dat;
  assign input_reg_and_398_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_160_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_6_sva,
      pe_0_0_run_cmp_176_input_out_rsc_z, input_reg_and_398_nl);
  wire [7:0] nl_pe_0_0_run_cmp_160_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_160_weight_rsc_dat = step_mux_10_itm_1;
  wire[0:0] input_reg_and_399_nl;
  wire [7:0] nl_pe_0_0_run_cmp_161_input_in_rsc_dat;
  assign input_reg_and_399_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_161_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_5_sva,
      pe_0_0_run_cmp_177_input_out_rsc_z, input_reg_and_399_nl);
  wire[0:0] psum_reg_and_421_nl;
  wire [15:0] nl_pe_0_0_run_cmp_161_psum_in_rsc_dat;
  assign psum_reg_and_421_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_161_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_6_sva,
      pe_0_0_run_cmp_162_psum_out_rsc_z, psum_reg_and_421_nl);
  wire [7:0] nl_pe_0_0_run_cmp_161_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_161_weight_rsc_dat = step_mux_249_itm_1;
  wire[0:0] input_reg_and_400_nl;
  wire [7:0] nl_pe_0_0_run_cmp_162_input_in_rsc_dat;
  assign input_reg_and_400_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_162_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_5_sva,
      pe_0_0_run_cmp_178_input_out_rsc_z, input_reg_and_400_nl);
  wire[0:0] psum_reg_and_422_nl;
  wire [15:0] nl_pe_0_0_run_cmp_162_psum_in_rsc_dat;
  assign psum_reg_and_422_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_162_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_6_sva,
      pe_0_0_run_cmp_163_psum_out_rsc_z, psum_reg_and_422_nl);
  wire [7:0] nl_pe_0_0_run_cmp_162_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_162_weight_rsc_dat = step_mux_233_itm_1;
  wire[0:0] input_reg_and_401_nl;
  wire [7:0] nl_pe_0_0_run_cmp_163_input_in_rsc_dat;
  assign input_reg_and_401_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_163_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_5_sva,
      pe_0_0_run_cmp_179_input_out_rsc_z, input_reg_and_401_nl);
  wire[0:0] psum_reg_and_423_nl;
  wire [15:0] nl_pe_0_0_run_cmp_163_psum_in_rsc_dat;
  assign psum_reg_and_423_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_163_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_6_sva,
      pe_0_0_run_cmp_164_psum_out_rsc_z, psum_reg_and_423_nl);
  wire [7:0] nl_pe_0_0_run_cmp_163_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_163_weight_rsc_dat = step_mux_217_itm_1;
  wire[0:0] input_reg_and_402_nl;
  wire [7:0] nl_pe_0_0_run_cmp_164_input_in_rsc_dat;
  assign input_reg_and_402_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_164_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_5_sva,
      pe_0_0_run_cmp_180_input_out_rsc_z, input_reg_and_402_nl);
  wire[0:0] psum_reg_and_424_nl;
  wire [15:0] nl_pe_0_0_run_cmp_164_psum_in_rsc_dat;
  assign psum_reg_and_424_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_164_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_6_sva,
      pe_0_0_run_cmp_165_psum_out_rsc_z, psum_reg_and_424_nl);
  wire [7:0] nl_pe_0_0_run_cmp_164_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_164_weight_rsc_dat = step_mux_201_itm_1;
  wire[0:0] input_reg_and_403_nl;
  wire [7:0] nl_pe_0_0_run_cmp_165_input_in_rsc_dat;
  assign input_reg_and_403_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_165_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_5_sva,
      pe_0_0_run_cmp_181_input_out_rsc_z, input_reg_and_403_nl);
  wire[0:0] psum_reg_and_425_nl;
  wire [15:0] nl_pe_0_0_run_cmp_165_psum_in_rsc_dat;
  assign psum_reg_and_425_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_165_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_6_sva,
      pe_0_0_run_cmp_166_psum_out_rsc_z, psum_reg_and_425_nl);
  wire [7:0] nl_pe_0_0_run_cmp_165_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_165_weight_rsc_dat = step_mux_185_itm_1;
  wire[0:0] input_reg_and_404_nl;
  wire [7:0] nl_pe_0_0_run_cmp_166_input_in_rsc_dat;
  assign input_reg_and_404_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_166_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_5_sva,
      pe_0_0_run_cmp_182_input_out_rsc_z, input_reg_and_404_nl);
  wire[0:0] psum_reg_and_426_nl;
  wire [15:0] nl_pe_0_0_run_cmp_166_psum_in_rsc_dat;
  assign psum_reg_and_426_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_166_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_6_sva,
      pe_0_0_run_cmp_167_psum_out_rsc_z, psum_reg_and_426_nl);
  wire [7:0] nl_pe_0_0_run_cmp_166_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_166_weight_rsc_dat = step_mux_169_itm_1;
  wire[0:0] input_reg_and_405_nl;
  wire [7:0] nl_pe_0_0_run_cmp_167_input_in_rsc_dat;
  assign input_reg_and_405_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_167_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_5_sva,
      pe_0_0_run_cmp_183_input_out_rsc_z, input_reg_and_405_nl);
  wire[0:0] psum_reg_and_427_nl;
  wire [15:0] nl_pe_0_0_run_cmp_167_psum_in_rsc_dat;
  assign psum_reg_and_427_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_167_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_6_sva, pe_0_0_run_cmp_168_psum_out_rsc_z,
      psum_reg_and_427_nl);
  wire [7:0] nl_pe_0_0_run_cmp_167_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_167_weight_rsc_dat = step_mux_153_itm_1;
  wire[0:0] input_reg_and_406_nl;
  wire [7:0] nl_pe_0_0_run_cmp_168_input_in_rsc_dat;
  assign input_reg_and_406_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_168_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_5_sva,
      pe_0_0_run_cmp_184_input_out_rsc_z, input_reg_and_406_nl);
  wire[0:0] psum_reg_and_428_nl;
  wire [15:0] nl_pe_0_0_run_cmp_168_psum_in_rsc_dat;
  assign psum_reg_and_428_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_168_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_6_sva, pe_0_0_run_cmp_169_psum_out_rsc_z,
      psum_reg_and_428_nl);
  wire [7:0] nl_pe_0_0_run_cmp_168_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_168_weight_rsc_dat = step_mux_137_itm_1;
  wire[0:0] input_reg_and_407_nl;
  wire [7:0] nl_pe_0_0_run_cmp_169_input_in_rsc_dat;
  assign input_reg_and_407_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_169_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_5_sva,
      pe_0_0_run_cmp_185_input_out_rsc_z, input_reg_and_407_nl);
  wire[0:0] psum_reg_and_429_nl;
  wire [15:0] nl_pe_0_0_run_cmp_169_psum_in_rsc_dat;
  assign psum_reg_and_429_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_169_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_6_sva, pe_0_0_run_cmp_170_psum_out_rsc_z,
      psum_reg_and_429_nl);
  wire [7:0] nl_pe_0_0_run_cmp_169_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_169_weight_rsc_dat = step_mux_121_itm_1;
  wire[0:0] input_reg_and_408_nl;
  wire [7:0] nl_pe_0_0_run_cmp_170_input_in_rsc_dat;
  assign input_reg_and_408_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_170_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_5_sva,
      pe_0_0_run_cmp_186_input_out_rsc_z, input_reg_and_408_nl);
  wire[0:0] psum_reg_and_430_nl;
  wire [15:0] nl_pe_0_0_run_cmp_170_psum_in_rsc_dat;
  assign psum_reg_and_430_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_170_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_6_sva, pe_0_0_run_cmp_171_psum_out_rsc_z,
      psum_reg_and_430_nl);
  wire [7:0] nl_pe_0_0_run_cmp_170_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_170_weight_rsc_dat = step_mux_105_itm_1;
  wire[0:0] input_reg_and_409_nl;
  wire [7:0] nl_pe_0_0_run_cmp_171_input_in_rsc_dat;
  assign input_reg_and_409_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_171_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_5_sva,
      pe_0_0_run_cmp_187_input_out_rsc_z, input_reg_and_409_nl);
  wire[0:0] psum_reg_and_431_nl;
  wire [15:0] nl_pe_0_0_run_cmp_171_psum_in_rsc_dat;
  assign psum_reg_and_431_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_171_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_6_sva, pe_0_0_run_cmp_172_psum_out_rsc_z,
      psum_reg_and_431_nl);
  wire [7:0] nl_pe_0_0_run_cmp_171_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_171_weight_rsc_dat = step_mux_89_itm_1;
  wire[0:0] input_reg_and_410_nl;
  wire [7:0] nl_pe_0_0_run_cmp_172_input_in_rsc_dat;
  assign input_reg_and_410_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_172_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_5_sva,
      pe_0_0_run_cmp_188_input_out_rsc_z, input_reg_and_410_nl);
  wire[0:0] psum_reg_and_432_nl;
  wire [15:0] nl_pe_0_0_run_cmp_172_psum_in_rsc_dat;
  assign psum_reg_and_432_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_172_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_6_sva, pe_0_0_run_cmp_173_psum_out_rsc_z,
      psum_reg_and_432_nl);
  wire [7:0] nl_pe_0_0_run_cmp_172_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_172_weight_rsc_dat = step_mux_73_itm_1;
  wire[0:0] input_reg_and_411_nl;
  wire [7:0] nl_pe_0_0_run_cmp_173_input_in_rsc_dat;
  assign input_reg_and_411_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_173_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_5_sva,
      pe_0_0_run_cmp_189_input_out_rsc_z, input_reg_and_411_nl);
  wire[0:0] psum_reg_and_433_nl;
  wire [15:0] nl_pe_0_0_run_cmp_173_psum_in_rsc_dat;
  assign psum_reg_and_433_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_173_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_6_sva, pe_0_0_run_cmp_174_psum_out_rsc_z,
      psum_reg_and_433_nl);
  wire [7:0] nl_pe_0_0_run_cmp_173_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_173_weight_rsc_dat = step_mux_57_itm_1;
  wire[0:0] input_reg_and_412_nl;
  wire [7:0] nl_pe_0_0_run_cmp_174_input_in_rsc_dat;
  assign input_reg_and_412_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_174_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_5_sva,
      pe_0_0_run_cmp_190_input_out_rsc_z, input_reg_and_412_nl);
  wire[0:0] psum_reg_and_434_nl;
  wire [15:0] nl_pe_0_0_run_cmp_174_psum_in_rsc_dat;
  assign psum_reg_and_434_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_174_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_6_sva, pe_0_0_run_cmp_175_psum_out_rsc_z,
      psum_reg_and_434_nl);
  wire [7:0] nl_pe_0_0_run_cmp_174_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_174_weight_rsc_dat = step_mux_41_itm_1;
  wire[0:0] input_reg_and_413_nl;
  wire [7:0] nl_pe_0_0_run_cmp_175_input_in_rsc_dat;
  assign input_reg_and_413_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_175_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_5_sva,
      pe_0_0_run_cmp_191_input_out_rsc_z, input_reg_and_413_nl);
  wire[0:0] psum_reg_and_435_nl;
  wire [15:0] nl_pe_0_0_run_cmp_175_psum_in_rsc_dat;
  assign psum_reg_and_435_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_175_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_6_sva, pe_0_0_run_cmp_176_psum_out_rsc_z,
      psum_reg_and_435_nl);
  wire [7:0] nl_pe_0_0_run_cmp_175_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_175_weight_rsc_dat = step_mux_25_itm_1;
  wire[0:0] input_reg_and_414_nl;
  wire [7:0] nl_pe_0_0_run_cmp_176_input_in_rsc_dat;
  assign input_reg_and_414_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_176_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_5_sva,
      pe_0_0_run_cmp_192_input_out_rsc_z, input_reg_and_414_nl);
  wire [7:0] nl_pe_0_0_run_cmp_176_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_176_weight_rsc_dat = step_mux_9_itm_1;
  wire[0:0] input_reg_and_415_nl;
  wire [7:0] nl_pe_0_0_run_cmp_177_input_in_rsc_dat;
  assign input_reg_and_415_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_177_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_4_sva,
      pe_0_0_run_cmp_193_input_out_rsc_z, input_reg_and_415_nl);
  wire[0:0] psum_reg_and_436_nl;
  wire [15:0] nl_pe_0_0_run_cmp_177_psum_in_rsc_dat;
  assign psum_reg_and_436_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_177_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_5_sva,
      pe_0_0_run_cmp_178_psum_out_rsc_z, psum_reg_and_436_nl);
  wire [7:0] nl_pe_0_0_run_cmp_177_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_177_weight_rsc_dat = step_mux_248_itm_1;
  wire[0:0] input_reg_and_416_nl;
  wire [7:0] nl_pe_0_0_run_cmp_178_input_in_rsc_dat;
  assign input_reg_and_416_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_178_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_4_sva,
      pe_0_0_run_cmp_194_input_out_rsc_z, input_reg_and_416_nl);
  wire[0:0] psum_reg_and_437_nl;
  wire [15:0] nl_pe_0_0_run_cmp_178_psum_in_rsc_dat;
  assign psum_reg_and_437_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_178_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_5_sva,
      pe_0_0_run_cmp_179_psum_out_rsc_z, psum_reg_and_437_nl);
  wire [7:0] nl_pe_0_0_run_cmp_178_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_178_weight_rsc_dat = step_mux_232_itm_1;
  wire[0:0] input_reg_and_417_nl;
  wire [7:0] nl_pe_0_0_run_cmp_179_input_in_rsc_dat;
  assign input_reg_and_417_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_179_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_4_sva,
      pe_0_0_run_cmp_195_input_out_rsc_z, input_reg_and_417_nl);
  wire[0:0] psum_reg_and_438_nl;
  wire [15:0] nl_pe_0_0_run_cmp_179_psum_in_rsc_dat;
  assign psum_reg_and_438_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_179_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_5_sva,
      pe_0_0_run_cmp_180_psum_out_rsc_z, psum_reg_and_438_nl);
  wire [7:0] nl_pe_0_0_run_cmp_179_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_179_weight_rsc_dat = step_mux_216_itm_1;
  wire[0:0] input_reg_and_418_nl;
  wire [7:0] nl_pe_0_0_run_cmp_180_input_in_rsc_dat;
  assign input_reg_and_418_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_180_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_4_sva,
      pe_0_0_run_cmp_196_input_out_rsc_z, input_reg_and_418_nl);
  wire[0:0] psum_reg_and_439_nl;
  wire [15:0] nl_pe_0_0_run_cmp_180_psum_in_rsc_dat;
  assign psum_reg_and_439_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_180_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_5_sva,
      pe_0_0_run_cmp_181_psum_out_rsc_z, psum_reg_and_439_nl);
  wire [7:0] nl_pe_0_0_run_cmp_180_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_180_weight_rsc_dat = step_mux_200_itm_1;
  wire[0:0] input_reg_and_419_nl;
  wire [7:0] nl_pe_0_0_run_cmp_181_input_in_rsc_dat;
  assign input_reg_and_419_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_181_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_4_sva,
      pe_0_0_run_cmp_197_input_out_rsc_z, input_reg_and_419_nl);
  wire[0:0] psum_reg_and_440_nl;
  wire [15:0] nl_pe_0_0_run_cmp_181_psum_in_rsc_dat;
  assign psum_reg_and_440_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_181_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_5_sva,
      pe_0_0_run_cmp_182_psum_out_rsc_z, psum_reg_and_440_nl);
  wire [7:0] nl_pe_0_0_run_cmp_181_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_181_weight_rsc_dat = step_mux_184_itm_1;
  wire[0:0] input_reg_and_420_nl;
  wire [7:0] nl_pe_0_0_run_cmp_182_input_in_rsc_dat;
  assign input_reg_and_420_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_182_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_4_sva,
      pe_0_0_run_cmp_198_input_out_rsc_z, input_reg_and_420_nl);
  wire[0:0] psum_reg_and_441_nl;
  wire [15:0] nl_pe_0_0_run_cmp_182_psum_in_rsc_dat;
  assign psum_reg_and_441_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_182_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_5_sva,
      pe_0_0_run_cmp_183_psum_out_rsc_z, psum_reg_and_441_nl);
  wire [7:0] nl_pe_0_0_run_cmp_182_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_182_weight_rsc_dat = step_mux_168_itm_1;
  wire[0:0] input_reg_and_421_nl;
  wire [7:0] nl_pe_0_0_run_cmp_183_input_in_rsc_dat;
  assign input_reg_and_421_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_183_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_4_sva,
      pe_0_0_run_cmp_199_input_out_rsc_z, input_reg_and_421_nl);
  wire[0:0] psum_reg_and_442_nl;
  wire [15:0] nl_pe_0_0_run_cmp_183_psum_in_rsc_dat;
  assign psum_reg_and_442_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_183_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_5_sva, pe_0_0_run_cmp_184_psum_out_rsc_z,
      psum_reg_and_442_nl);
  wire [7:0] nl_pe_0_0_run_cmp_183_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_183_weight_rsc_dat = step_mux_152_itm_1;
  wire[0:0] input_reg_and_422_nl;
  wire [7:0] nl_pe_0_0_run_cmp_184_input_in_rsc_dat;
  assign input_reg_and_422_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_184_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_4_sva,
      pe_0_0_run_cmp_200_input_out_rsc_z, input_reg_and_422_nl);
  wire[0:0] psum_reg_and_443_nl;
  wire [15:0] nl_pe_0_0_run_cmp_184_psum_in_rsc_dat;
  assign psum_reg_and_443_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_184_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_5_sva, pe_0_0_run_cmp_185_psum_out_rsc_z,
      psum_reg_and_443_nl);
  wire [7:0] nl_pe_0_0_run_cmp_184_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_184_weight_rsc_dat = step_mux_136_itm_1;
  wire[0:0] input_reg_and_423_nl;
  wire [7:0] nl_pe_0_0_run_cmp_185_input_in_rsc_dat;
  assign input_reg_and_423_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_185_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_4_sva,
      pe_0_0_run_cmp_201_input_out_rsc_z, input_reg_and_423_nl);
  wire[0:0] psum_reg_and_444_nl;
  wire [15:0] nl_pe_0_0_run_cmp_185_psum_in_rsc_dat;
  assign psum_reg_and_444_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_185_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_5_sva, pe_0_0_run_cmp_186_psum_out_rsc_z,
      psum_reg_and_444_nl);
  wire [7:0] nl_pe_0_0_run_cmp_185_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_185_weight_rsc_dat = step_mux_120_itm_1;
  wire[0:0] input_reg_and_424_nl;
  wire [7:0] nl_pe_0_0_run_cmp_186_input_in_rsc_dat;
  assign input_reg_and_424_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_186_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_4_sva,
      pe_0_0_run_cmp_202_input_out_rsc_z, input_reg_and_424_nl);
  wire[0:0] psum_reg_and_445_nl;
  wire [15:0] nl_pe_0_0_run_cmp_186_psum_in_rsc_dat;
  assign psum_reg_and_445_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_186_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_5_sva, pe_0_0_run_cmp_187_psum_out_rsc_z,
      psum_reg_and_445_nl);
  wire [7:0] nl_pe_0_0_run_cmp_186_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_186_weight_rsc_dat = step_mux_104_itm_1;
  wire[0:0] input_reg_and_425_nl;
  wire [7:0] nl_pe_0_0_run_cmp_187_input_in_rsc_dat;
  assign input_reg_and_425_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_187_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_4_sva,
      pe_0_0_run_cmp_203_input_out_rsc_z, input_reg_and_425_nl);
  wire[0:0] psum_reg_and_446_nl;
  wire [15:0] nl_pe_0_0_run_cmp_187_psum_in_rsc_dat;
  assign psum_reg_and_446_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_187_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_5_sva, pe_0_0_run_cmp_188_psum_out_rsc_z,
      psum_reg_and_446_nl);
  wire [7:0] nl_pe_0_0_run_cmp_187_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_187_weight_rsc_dat = step_mux_88_itm_1;
  wire[0:0] input_reg_and_426_nl;
  wire [7:0] nl_pe_0_0_run_cmp_188_input_in_rsc_dat;
  assign input_reg_and_426_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_188_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_4_sva,
      pe_0_0_run_cmp_204_input_out_rsc_z, input_reg_and_426_nl);
  wire[0:0] psum_reg_and_447_nl;
  wire [15:0] nl_pe_0_0_run_cmp_188_psum_in_rsc_dat;
  assign psum_reg_and_447_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_188_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_5_sva, pe_0_0_run_cmp_189_psum_out_rsc_z,
      psum_reg_and_447_nl);
  wire [7:0] nl_pe_0_0_run_cmp_188_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_188_weight_rsc_dat = step_mux_72_itm_1;
  wire[0:0] input_reg_and_427_nl;
  wire [7:0] nl_pe_0_0_run_cmp_189_input_in_rsc_dat;
  assign input_reg_and_427_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_189_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_4_sva,
      pe_0_0_run_cmp_205_input_out_rsc_z, input_reg_and_427_nl);
  wire[0:0] psum_reg_and_448_nl;
  wire [15:0] nl_pe_0_0_run_cmp_189_psum_in_rsc_dat;
  assign psum_reg_and_448_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_189_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_5_sva, pe_0_0_run_cmp_190_psum_out_rsc_z,
      psum_reg_and_448_nl);
  wire [7:0] nl_pe_0_0_run_cmp_189_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_189_weight_rsc_dat = step_mux_56_itm_1;
  wire[0:0] input_reg_and_428_nl;
  wire [7:0] nl_pe_0_0_run_cmp_190_input_in_rsc_dat;
  assign input_reg_and_428_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_190_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_4_sva,
      pe_0_0_run_cmp_206_input_out_rsc_z, input_reg_and_428_nl);
  wire[0:0] psum_reg_and_449_nl;
  wire [15:0] nl_pe_0_0_run_cmp_190_psum_in_rsc_dat;
  assign psum_reg_and_449_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_190_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_5_sva, pe_0_0_run_cmp_191_psum_out_rsc_z,
      psum_reg_and_449_nl);
  wire [7:0] nl_pe_0_0_run_cmp_190_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_190_weight_rsc_dat = step_mux_40_itm_1;
  wire[0:0] input_reg_and_429_nl;
  wire [7:0] nl_pe_0_0_run_cmp_191_input_in_rsc_dat;
  assign input_reg_and_429_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_191_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_4_sva,
      pe_0_0_run_cmp_207_input_out_rsc_z, input_reg_and_429_nl);
  wire[0:0] psum_reg_and_450_nl;
  wire [15:0] nl_pe_0_0_run_cmp_191_psum_in_rsc_dat;
  assign psum_reg_and_450_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_191_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_5_sva, pe_0_0_run_cmp_192_psum_out_rsc_z,
      psum_reg_and_450_nl);
  wire [7:0] nl_pe_0_0_run_cmp_191_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_191_weight_rsc_dat = step_mux_24_itm_1;
  wire[0:0] input_reg_and_430_nl;
  wire [7:0] nl_pe_0_0_run_cmp_192_input_in_rsc_dat;
  assign input_reg_and_430_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_192_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_4_sva,
      pe_0_0_run_cmp_208_input_out_rsc_z, input_reg_and_430_nl);
  wire [7:0] nl_pe_0_0_run_cmp_192_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_192_weight_rsc_dat = step_mux_8_itm_1;
  wire[0:0] input_reg_and_431_nl;
  wire [7:0] nl_pe_0_0_run_cmp_193_input_in_rsc_dat;
  assign input_reg_and_431_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_193_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_3_sva,
      pe_0_0_run_cmp_209_input_out_rsc_z, input_reg_and_431_nl);
  wire[0:0] psum_reg_and_451_nl;
  wire [15:0] nl_pe_0_0_run_cmp_193_psum_in_rsc_dat;
  assign psum_reg_and_451_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_193_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_4_sva,
      pe_0_0_run_cmp_194_psum_out_rsc_z, psum_reg_and_451_nl);
  wire [7:0] nl_pe_0_0_run_cmp_193_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_193_weight_rsc_dat = step_mux_247_itm_1;
  wire[0:0] input_reg_and_432_nl;
  wire [7:0] nl_pe_0_0_run_cmp_194_input_in_rsc_dat;
  assign input_reg_and_432_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_194_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_3_sva,
      pe_0_0_run_cmp_210_input_out_rsc_z, input_reg_and_432_nl);
  wire[0:0] psum_reg_and_452_nl;
  wire [15:0] nl_pe_0_0_run_cmp_194_psum_in_rsc_dat;
  assign psum_reg_and_452_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_194_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_4_sva,
      pe_0_0_run_cmp_195_psum_out_rsc_z, psum_reg_and_452_nl);
  wire [7:0] nl_pe_0_0_run_cmp_194_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_194_weight_rsc_dat = step_mux_231_itm_1;
  wire[0:0] input_reg_and_433_nl;
  wire [7:0] nl_pe_0_0_run_cmp_195_input_in_rsc_dat;
  assign input_reg_and_433_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_195_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_3_sva,
      pe_0_0_run_cmp_211_input_out_rsc_z, input_reg_and_433_nl);
  wire[0:0] psum_reg_and_453_nl;
  wire [15:0] nl_pe_0_0_run_cmp_195_psum_in_rsc_dat;
  assign psum_reg_and_453_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_195_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_4_sva,
      pe_0_0_run_cmp_196_psum_out_rsc_z, psum_reg_and_453_nl);
  wire [7:0] nl_pe_0_0_run_cmp_195_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_195_weight_rsc_dat = step_mux_215_itm_1;
  wire[0:0] input_reg_and_434_nl;
  wire [7:0] nl_pe_0_0_run_cmp_196_input_in_rsc_dat;
  assign input_reg_and_434_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_196_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_3_sva,
      pe_0_0_run_cmp_212_input_out_rsc_z, input_reg_and_434_nl);
  wire[0:0] psum_reg_and_454_nl;
  wire [15:0] nl_pe_0_0_run_cmp_196_psum_in_rsc_dat;
  assign psum_reg_and_454_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_196_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_4_sva,
      pe_0_0_run_cmp_197_psum_out_rsc_z, psum_reg_and_454_nl);
  wire [7:0] nl_pe_0_0_run_cmp_196_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_196_weight_rsc_dat = step_mux_199_itm_1;
  wire[0:0] input_reg_and_435_nl;
  wire [7:0] nl_pe_0_0_run_cmp_197_input_in_rsc_dat;
  assign input_reg_and_435_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_197_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_3_sva,
      pe_0_0_run_cmp_213_input_out_rsc_z, input_reg_and_435_nl);
  wire[0:0] psum_reg_and_455_nl;
  wire [15:0] nl_pe_0_0_run_cmp_197_psum_in_rsc_dat;
  assign psum_reg_and_455_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_197_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_4_sva,
      pe_0_0_run_cmp_198_psum_out_rsc_z, psum_reg_and_455_nl);
  wire [7:0] nl_pe_0_0_run_cmp_197_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_197_weight_rsc_dat = step_mux_183_itm_1;
  wire[0:0] input_reg_and_436_nl;
  wire [7:0] nl_pe_0_0_run_cmp_198_input_in_rsc_dat;
  assign input_reg_and_436_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_198_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_3_sva,
      pe_0_0_run_cmp_214_input_out_rsc_z, input_reg_and_436_nl);
  wire[0:0] psum_reg_and_456_nl;
  wire [15:0] nl_pe_0_0_run_cmp_198_psum_in_rsc_dat;
  assign psum_reg_and_456_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_198_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_4_sva,
      pe_0_0_run_cmp_199_psum_out_rsc_z, psum_reg_and_456_nl);
  wire [7:0] nl_pe_0_0_run_cmp_198_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_198_weight_rsc_dat = step_mux_167_itm_1;
  wire[0:0] input_reg_and_437_nl;
  wire [7:0] nl_pe_0_0_run_cmp_199_input_in_rsc_dat;
  assign input_reg_and_437_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_199_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_3_sva,
      pe_0_0_run_cmp_215_input_out_rsc_z, input_reg_and_437_nl);
  wire[0:0] psum_reg_and_457_nl;
  wire [15:0] nl_pe_0_0_run_cmp_199_psum_in_rsc_dat;
  assign psum_reg_and_457_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_199_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_4_sva, pe_0_0_run_cmp_200_psum_out_rsc_z,
      psum_reg_and_457_nl);
  wire [7:0] nl_pe_0_0_run_cmp_199_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_199_weight_rsc_dat = step_mux_151_itm_1;
  wire[0:0] input_reg_and_438_nl;
  wire [7:0] nl_pe_0_0_run_cmp_200_input_in_rsc_dat;
  assign input_reg_and_438_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_200_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_3_sva,
      pe_0_0_run_cmp_216_input_out_rsc_z, input_reg_and_438_nl);
  wire[0:0] psum_reg_and_458_nl;
  wire [15:0] nl_pe_0_0_run_cmp_200_psum_in_rsc_dat;
  assign psum_reg_and_458_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_200_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_4_sva, pe_0_0_run_cmp_201_psum_out_rsc_z,
      psum_reg_and_458_nl);
  wire [7:0] nl_pe_0_0_run_cmp_200_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_200_weight_rsc_dat = step_mux_135_itm_1;
  wire[0:0] input_reg_and_439_nl;
  wire [7:0] nl_pe_0_0_run_cmp_201_input_in_rsc_dat;
  assign input_reg_and_439_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_201_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_3_sva,
      pe_0_0_run_cmp_217_input_out_rsc_z, input_reg_and_439_nl);
  wire[0:0] psum_reg_and_459_nl;
  wire [15:0] nl_pe_0_0_run_cmp_201_psum_in_rsc_dat;
  assign psum_reg_and_459_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_201_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_4_sva, pe_0_0_run_cmp_202_psum_out_rsc_z,
      psum_reg_and_459_nl);
  wire [7:0] nl_pe_0_0_run_cmp_201_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_201_weight_rsc_dat = step_mux_119_itm_1;
  wire[0:0] input_reg_and_440_nl;
  wire [7:0] nl_pe_0_0_run_cmp_202_input_in_rsc_dat;
  assign input_reg_and_440_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_202_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_3_sva,
      pe_0_0_run_cmp_218_input_out_rsc_z, input_reg_and_440_nl);
  wire[0:0] psum_reg_and_460_nl;
  wire [15:0] nl_pe_0_0_run_cmp_202_psum_in_rsc_dat;
  assign psum_reg_and_460_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_202_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_4_sva, pe_0_0_run_cmp_203_psum_out_rsc_z,
      psum_reg_and_460_nl);
  wire [7:0] nl_pe_0_0_run_cmp_202_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_202_weight_rsc_dat = step_mux_103_itm_1;
  wire[0:0] input_reg_and_441_nl;
  wire [7:0] nl_pe_0_0_run_cmp_203_input_in_rsc_dat;
  assign input_reg_and_441_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_203_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_3_sva,
      pe_0_0_run_cmp_219_input_out_rsc_z, input_reg_and_441_nl);
  wire[0:0] psum_reg_and_461_nl;
  wire [15:0] nl_pe_0_0_run_cmp_203_psum_in_rsc_dat;
  assign psum_reg_and_461_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_203_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_4_sva, pe_0_0_run_cmp_204_psum_out_rsc_z,
      psum_reg_and_461_nl);
  wire [7:0] nl_pe_0_0_run_cmp_203_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_203_weight_rsc_dat = step_mux_87_itm_1;
  wire[0:0] input_reg_and_442_nl;
  wire [7:0] nl_pe_0_0_run_cmp_204_input_in_rsc_dat;
  assign input_reg_and_442_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_204_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_3_sva,
      pe_0_0_run_cmp_220_input_out_rsc_z, input_reg_and_442_nl);
  wire[0:0] psum_reg_and_462_nl;
  wire [15:0] nl_pe_0_0_run_cmp_204_psum_in_rsc_dat;
  assign psum_reg_and_462_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_204_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_4_sva, pe_0_0_run_cmp_205_psum_out_rsc_z,
      psum_reg_and_462_nl);
  wire [7:0] nl_pe_0_0_run_cmp_204_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_204_weight_rsc_dat = step_mux_71_itm_1;
  wire[0:0] input_reg_and_443_nl;
  wire [7:0] nl_pe_0_0_run_cmp_205_input_in_rsc_dat;
  assign input_reg_and_443_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_205_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_3_sva,
      pe_0_0_run_cmp_221_input_out_rsc_z, input_reg_and_443_nl);
  wire[0:0] psum_reg_and_463_nl;
  wire [15:0] nl_pe_0_0_run_cmp_205_psum_in_rsc_dat;
  assign psum_reg_and_463_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_205_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_4_sva, pe_0_0_run_cmp_206_psum_out_rsc_z,
      psum_reg_and_463_nl);
  wire [7:0] nl_pe_0_0_run_cmp_205_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_205_weight_rsc_dat = step_mux_55_itm_1;
  wire[0:0] input_reg_and_444_nl;
  wire [7:0] nl_pe_0_0_run_cmp_206_input_in_rsc_dat;
  assign input_reg_and_444_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_206_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_3_sva,
      pe_0_0_run_cmp_222_input_out_rsc_z, input_reg_and_444_nl);
  wire[0:0] psum_reg_and_464_nl;
  wire [15:0] nl_pe_0_0_run_cmp_206_psum_in_rsc_dat;
  assign psum_reg_and_464_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_206_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_4_sva, pe_0_0_run_cmp_207_psum_out_rsc_z,
      psum_reg_and_464_nl);
  wire [7:0] nl_pe_0_0_run_cmp_206_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_206_weight_rsc_dat = step_mux_39_itm_1;
  wire[0:0] input_reg_and_445_nl;
  wire [7:0] nl_pe_0_0_run_cmp_207_input_in_rsc_dat;
  assign input_reg_and_445_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_207_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_3_sva,
      pe_0_0_run_cmp_223_input_out_rsc_z, input_reg_and_445_nl);
  wire[0:0] psum_reg_and_465_nl;
  wire [15:0] nl_pe_0_0_run_cmp_207_psum_in_rsc_dat;
  assign psum_reg_and_465_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_207_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_4_sva, pe_0_0_run_cmp_208_psum_out_rsc_z,
      psum_reg_and_465_nl);
  wire [7:0] nl_pe_0_0_run_cmp_207_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_207_weight_rsc_dat = step_mux_23_itm_1;
  wire[0:0] input_reg_and_446_nl;
  wire [7:0] nl_pe_0_0_run_cmp_208_input_in_rsc_dat;
  assign input_reg_and_446_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_208_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_3_sva,
      pe_0_0_run_cmp_224_input_out_rsc_z, input_reg_and_446_nl);
  wire [7:0] nl_pe_0_0_run_cmp_208_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_208_weight_rsc_dat = step_mux_7_itm_1;
  wire[0:0] input_reg_and_447_nl;
  wire [7:0] nl_pe_0_0_run_cmp_209_input_in_rsc_dat;
  assign input_reg_and_447_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_209_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_2_sva,
      pe_0_0_run_cmp_225_input_out_rsc_z, input_reg_and_447_nl);
  wire[0:0] psum_reg_and_466_nl;
  wire [15:0] nl_pe_0_0_run_cmp_209_psum_in_rsc_dat;
  assign psum_reg_and_466_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_209_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_3_sva,
      pe_0_0_run_cmp_210_psum_out_rsc_z, psum_reg_and_466_nl);
  wire [7:0] nl_pe_0_0_run_cmp_209_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_209_weight_rsc_dat = step_mux_246_itm_1;
  wire[0:0] input_reg_and_448_nl;
  wire [7:0] nl_pe_0_0_run_cmp_210_input_in_rsc_dat;
  assign input_reg_and_448_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_210_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_2_sva,
      pe_0_0_run_cmp_226_input_out_rsc_z, input_reg_and_448_nl);
  wire[0:0] psum_reg_and_467_nl;
  wire [15:0] nl_pe_0_0_run_cmp_210_psum_in_rsc_dat;
  assign psum_reg_and_467_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_210_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_3_sva,
      pe_0_0_run_cmp_211_psum_out_rsc_z, psum_reg_and_467_nl);
  wire [7:0] nl_pe_0_0_run_cmp_210_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_210_weight_rsc_dat = step_mux_230_itm_1;
  wire[0:0] input_reg_and_449_nl;
  wire [7:0] nl_pe_0_0_run_cmp_211_input_in_rsc_dat;
  assign input_reg_and_449_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_211_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_2_sva,
      pe_0_0_run_cmp_227_input_out_rsc_z, input_reg_and_449_nl);
  wire[0:0] psum_reg_and_468_nl;
  wire [15:0] nl_pe_0_0_run_cmp_211_psum_in_rsc_dat;
  assign psum_reg_and_468_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_211_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_3_sva,
      pe_0_0_run_cmp_212_psum_out_rsc_z, psum_reg_and_468_nl);
  wire [7:0] nl_pe_0_0_run_cmp_211_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_211_weight_rsc_dat = step_mux_214_itm_1;
  wire[0:0] input_reg_and_450_nl;
  wire [7:0] nl_pe_0_0_run_cmp_212_input_in_rsc_dat;
  assign input_reg_and_450_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_212_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_2_sva,
      pe_0_0_run_cmp_228_input_out_rsc_z, input_reg_and_450_nl);
  wire[0:0] psum_reg_and_469_nl;
  wire [15:0] nl_pe_0_0_run_cmp_212_psum_in_rsc_dat;
  assign psum_reg_and_469_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_212_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_3_sva,
      pe_0_0_run_cmp_213_psum_out_rsc_z, psum_reg_and_469_nl);
  wire [7:0] nl_pe_0_0_run_cmp_212_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_212_weight_rsc_dat = step_mux_198_itm_1;
  wire[0:0] input_reg_and_451_nl;
  wire [7:0] nl_pe_0_0_run_cmp_213_input_in_rsc_dat;
  assign input_reg_and_451_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_213_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_2_sva,
      pe_0_0_run_cmp_229_input_out_rsc_z, input_reg_and_451_nl);
  wire[0:0] psum_reg_and_470_nl;
  wire [15:0] nl_pe_0_0_run_cmp_213_psum_in_rsc_dat;
  assign psum_reg_and_470_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_213_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_3_sva,
      pe_0_0_run_cmp_214_psum_out_rsc_z, psum_reg_and_470_nl);
  wire [7:0] nl_pe_0_0_run_cmp_213_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_213_weight_rsc_dat = step_mux_182_itm_1;
  wire[0:0] input_reg_and_452_nl;
  wire [7:0] nl_pe_0_0_run_cmp_214_input_in_rsc_dat;
  assign input_reg_and_452_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_214_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_2_sva,
      pe_0_0_run_cmp_230_input_out_rsc_z, input_reg_and_452_nl);
  wire[0:0] psum_reg_and_471_nl;
  wire [15:0] nl_pe_0_0_run_cmp_214_psum_in_rsc_dat;
  assign psum_reg_and_471_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_214_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_3_sva,
      pe_0_0_run_cmp_215_psum_out_rsc_z, psum_reg_and_471_nl);
  wire [7:0] nl_pe_0_0_run_cmp_214_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_214_weight_rsc_dat = step_mux_166_itm_1;
  wire[0:0] input_reg_and_453_nl;
  wire [7:0] nl_pe_0_0_run_cmp_215_input_in_rsc_dat;
  assign input_reg_and_453_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_215_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_2_sva,
      pe_0_0_run_cmp_231_input_out_rsc_z, input_reg_and_453_nl);
  wire[0:0] psum_reg_and_472_nl;
  wire [15:0] nl_pe_0_0_run_cmp_215_psum_in_rsc_dat;
  assign psum_reg_and_472_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_215_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_3_sva, pe_0_0_run_cmp_216_psum_out_rsc_z,
      psum_reg_and_472_nl);
  wire [7:0] nl_pe_0_0_run_cmp_215_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_215_weight_rsc_dat = step_mux_150_itm_1;
  wire[0:0] input_reg_and_454_nl;
  wire [7:0] nl_pe_0_0_run_cmp_216_input_in_rsc_dat;
  assign input_reg_and_454_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_216_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_2_sva,
      pe_0_0_run_cmp_232_input_out_rsc_z, input_reg_and_454_nl);
  wire[0:0] psum_reg_and_473_nl;
  wire [15:0] nl_pe_0_0_run_cmp_216_psum_in_rsc_dat;
  assign psum_reg_and_473_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_216_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_3_sva, pe_0_0_run_cmp_217_psum_out_rsc_z,
      psum_reg_and_473_nl);
  wire [7:0] nl_pe_0_0_run_cmp_216_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_216_weight_rsc_dat = step_mux_134_itm_1;
  wire[0:0] input_reg_and_455_nl;
  wire [7:0] nl_pe_0_0_run_cmp_217_input_in_rsc_dat;
  assign input_reg_and_455_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_217_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_2_sva,
      pe_0_0_run_cmp_233_input_out_rsc_z, input_reg_and_455_nl);
  wire[0:0] psum_reg_and_474_nl;
  wire [15:0] nl_pe_0_0_run_cmp_217_psum_in_rsc_dat;
  assign psum_reg_and_474_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_217_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_3_sva, pe_0_0_run_cmp_218_psum_out_rsc_z,
      psum_reg_and_474_nl);
  wire [7:0] nl_pe_0_0_run_cmp_217_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_217_weight_rsc_dat = step_mux_118_itm_1;
  wire[0:0] input_reg_and_456_nl;
  wire [7:0] nl_pe_0_0_run_cmp_218_input_in_rsc_dat;
  assign input_reg_and_456_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_218_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_2_sva,
      pe_0_0_run_cmp_234_input_out_rsc_z, input_reg_and_456_nl);
  wire[0:0] psum_reg_and_475_nl;
  wire [15:0] nl_pe_0_0_run_cmp_218_psum_in_rsc_dat;
  assign psum_reg_and_475_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_218_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_3_sva, pe_0_0_run_cmp_219_psum_out_rsc_z,
      psum_reg_and_475_nl);
  wire [7:0] nl_pe_0_0_run_cmp_218_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_218_weight_rsc_dat = step_mux_102_itm_1;
  wire[0:0] input_reg_and_457_nl;
  wire [7:0] nl_pe_0_0_run_cmp_219_input_in_rsc_dat;
  assign input_reg_and_457_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_219_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_2_sva,
      pe_0_0_run_cmp_235_input_out_rsc_z, input_reg_and_457_nl);
  wire[0:0] psum_reg_and_476_nl;
  wire [15:0] nl_pe_0_0_run_cmp_219_psum_in_rsc_dat;
  assign psum_reg_and_476_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_219_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_3_sva, pe_0_0_run_cmp_220_psum_out_rsc_z,
      psum_reg_and_476_nl);
  wire [7:0] nl_pe_0_0_run_cmp_219_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_219_weight_rsc_dat = step_mux_86_itm_1;
  wire[0:0] input_reg_and_458_nl;
  wire [7:0] nl_pe_0_0_run_cmp_220_input_in_rsc_dat;
  assign input_reg_and_458_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_220_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_2_sva,
      pe_0_0_run_cmp_236_input_out_rsc_z, input_reg_and_458_nl);
  wire[0:0] psum_reg_and_477_nl;
  wire [15:0] nl_pe_0_0_run_cmp_220_psum_in_rsc_dat;
  assign psum_reg_and_477_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_220_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_3_sva, pe_0_0_run_cmp_221_psum_out_rsc_z,
      psum_reg_and_477_nl);
  wire [7:0] nl_pe_0_0_run_cmp_220_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_220_weight_rsc_dat = step_mux_70_itm_1;
  wire[0:0] input_reg_and_459_nl;
  wire [7:0] nl_pe_0_0_run_cmp_221_input_in_rsc_dat;
  assign input_reg_and_459_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_221_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_2_sva,
      pe_0_0_run_cmp_237_input_out_rsc_z, input_reg_and_459_nl);
  wire[0:0] psum_reg_and_478_nl;
  wire [15:0] nl_pe_0_0_run_cmp_221_psum_in_rsc_dat;
  assign psum_reg_and_478_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_221_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_3_sva, pe_0_0_run_cmp_222_psum_out_rsc_z,
      psum_reg_and_478_nl);
  wire [7:0] nl_pe_0_0_run_cmp_221_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_221_weight_rsc_dat = step_mux_54_itm_1;
  wire[0:0] input_reg_and_460_nl;
  wire [7:0] nl_pe_0_0_run_cmp_222_input_in_rsc_dat;
  assign input_reg_and_460_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_222_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_2_sva,
      pe_0_0_run_cmp_238_input_out_rsc_z, input_reg_and_460_nl);
  wire[0:0] psum_reg_and_479_nl;
  wire [15:0] nl_pe_0_0_run_cmp_222_psum_in_rsc_dat;
  assign psum_reg_and_479_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_222_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_3_sva, pe_0_0_run_cmp_223_psum_out_rsc_z,
      psum_reg_and_479_nl);
  wire [7:0] nl_pe_0_0_run_cmp_222_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_222_weight_rsc_dat = step_mux_38_itm_1;
  wire[0:0] input_reg_and_461_nl;
  wire [7:0] nl_pe_0_0_run_cmp_223_input_in_rsc_dat;
  assign input_reg_and_461_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_223_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_2_sva,
      pe_0_0_run_cmp_239_input_out_rsc_z, input_reg_and_461_nl);
  wire[0:0] psum_reg_and_480_nl;
  wire [15:0] nl_pe_0_0_run_cmp_223_psum_in_rsc_dat;
  assign psum_reg_and_480_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_223_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_3_sva, pe_0_0_run_cmp_224_psum_out_rsc_z,
      psum_reg_and_480_nl);
  wire [7:0] nl_pe_0_0_run_cmp_223_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_223_weight_rsc_dat = step_mux_22_itm_1;
  wire[0:0] input_reg_and_462_nl;
  wire [7:0] nl_pe_0_0_run_cmp_224_input_in_rsc_dat;
  assign input_reg_and_462_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_224_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_2_sva,
      pe_0_0_run_cmp_240_input_out_rsc_z, input_reg_and_462_nl);
  wire [7:0] nl_pe_0_0_run_cmp_224_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_224_weight_rsc_dat = step_mux_6_itm_1;
  wire[0:0] input_reg_and_463_nl;
  wire [7:0] nl_pe_0_0_run_cmp_225_input_in_rsc_dat;
  assign input_reg_and_463_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_225_input_in_rsc_dat = MUX_v_8_2_2(input_reg_16_1_sva,
      pe_0_0_run_cmp_241_input_out_rsc_z, input_reg_and_463_nl);
  wire[0:0] psum_reg_and_481_nl;
  wire [15:0] nl_pe_0_0_run_cmp_225_psum_in_rsc_dat;
  assign psum_reg_and_481_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_225_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_2_sva,
      pe_0_0_run_cmp_226_psum_out_rsc_z, psum_reg_and_481_nl);
  wire [7:0] nl_pe_0_0_run_cmp_225_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_225_weight_rsc_dat = step_mux_245_itm_1;
  wire[0:0] input_reg_and_464_nl;
  wire [7:0] nl_pe_0_0_run_cmp_226_input_in_rsc_dat;
  assign input_reg_and_464_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_226_input_in_rsc_dat = MUX_v_8_2_2(input_reg_15_1_sva,
      pe_0_0_run_cmp_242_input_out_rsc_z, input_reg_and_464_nl);
  wire[0:0] psum_reg_and_482_nl;
  wire [15:0] nl_pe_0_0_run_cmp_226_psum_in_rsc_dat;
  assign psum_reg_and_482_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_226_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_2_sva,
      pe_0_0_run_cmp_227_psum_out_rsc_z, psum_reg_and_482_nl);
  wire [7:0] nl_pe_0_0_run_cmp_226_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_226_weight_rsc_dat = step_mux_229_itm_1;
  wire[0:0] input_reg_and_465_nl;
  wire [7:0] nl_pe_0_0_run_cmp_227_input_in_rsc_dat;
  assign input_reg_and_465_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_227_input_in_rsc_dat = MUX_v_8_2_2(input_reg_14_1_sva,
      pe_0_0_run_cmp_243_input_out_rsc_z, input_reg_and_465_nl);
  wire[0:0] psum_reg_and_483_nl;
  wire [15:0] nl_pe_0_0_run_cmp_227_psum_in_rsc_dat;
  assign psum_reg_and_483_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_227_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_2_sva,
      pe_0_0_run_cmp_228_psum_out_rsc_z, psum_reg_and_483_nl);
  wire [7:0] nl_pe_0_0_run_cmp_227_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_227_weight_rsc_dat = step_mux_213_itm_1;
  wire[0:0] input_reg_and_466_nl;
  wire [7:0] nl_pe_0_0_run_cmp_228_input_in_rsc_dat;
  assign input_reg_and_466_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_228_input_in_rsc_dat = MUX_v_8_2_2(input_reg_13_1_sva,
      pe_0_0_run_cmp_244_input_out_rsc_z, input_reg_and_466_nl);
  wire[0:0] psum_reg_and_484_nl;
  wire [15:0] nl_pe_0_0_run_cmp_228_psum_in_rsc_dat;
  assign psum_reg_and_484_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_228_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_2_sva,
      pe_0_0_run_cmp_229_psum_out_rsc_z, psum_reg_and_484_nl);
  wire [7:0] nl_pe_0_0_run_cmp_228_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_228_weight_rsc_dat = step_mux_197_itm_1;
  wire[0:0] input_reg_and_467_nl;
  wire [7:0] nl_pe_0_0_run_cmp_229_input_in_rsc_dat;
  assign input_reg_and_467_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_229_input_in_rsc_dat = MUX_v_8_2_2(input_reg_12_1_sva,
      pe_0_0_run_cmp_245_input_out_rsc_z, input_reg_and_467_nl);
  wire[0:0] psum_reg_and_485_nl;
  wire [15:0] nl_pe_0_0_run_cmp_229_psum_in_rsc_dat;
  assign psum_reg_and_485_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_229_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_2_sva,
      pe_0_0_run_cmp_230_psum_out_rsc_z, psum_reg_and_485_nl);
  wire [7:0] nl_pe_0_0_run_cmp_229_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_229_weight_rsc_dat = step_mux_181_itm_1;
  wire[0:0] input_reg_and_468_nl;
  wire [7:0] nl_pe_0_0_run_cmp_230_input_in_rsc_dat;
  assign input_reg_and_468_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_230_input_in_rsc_dat = MUX_v_8_2_2(input_reg_11_1_sva,
      pe_0_0_run_cmp_246_input_out_rsc_z, input_reg_and_468_nl);
  wire[0:0] psum_reg_and_486_nl;
  wire [15:0] nl_pe_0_0_run_cmp_230_psum_in_rsc_dat;
  assign psum_reg_and_486_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_230_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_2_sva,
      pe_0_0_run_cmp_231_psum_out_rsc_z, psum_reg_and_486_nl);
  wire [7:0] nl_pe_0_0_run_cmp_230_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_230_weight_rsc_dat = step_mux_165_itm_1;
  wire[0:0] input_reg_and_469_nl;
  wire [7:0] nl_pe_0_0_run_cmp_231_input_in_rsc_dat;
  assign input_reg_and_469_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_231_input_in_rsc_dat = MUX_v_8_2_2(input_reg_10_1_sva,
      pe_0_0_run_cmp_247_input_out_rsc_z, input_reg_and_469_nl);
  wire[0:0] psum_reg_and_487_nl;
  wire [15:0] nl_pe_0_0_run_cmp_231_psum_in_rsc_dat;
  assign psum_reg_and_487_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_231_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_2_sva, pe_0_0_run_cmp_232_psum_out_rsc_z,
      psum_reg_and_487_nl);
  wire [7:0] nl_pe_0_0_run_cmp_231_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_231_weight_rsc_dat = step_mux_149_itm_1;
  wire[0:0] input_reg_and_470_nl;
  wire [7:0] nl_pe_0_0_run_cmp_232_input_in_rsc_dat;
  assign input_reg_and_470_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_232_input_in_rsc_dat = MUX_v_8_2_2(input_reg_9_1_sva,
      pe_0_0_run_cmp_248_input_out_rsc_z, input_reg_and_470_nl);
  wire[0:0] psum_reg_and_488_nl;
  wire [15:0] nl_pe_0_0_run_cmp_232_psum_in_rsc_dat;
  assign psum_reg_and_488_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_232_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_2_sva, pe_0_0_run_cmp_233_psum_out_rsc_z,
      psum_reg_and_488_nl);
  wire [7:0] nl_pe_0_0_run_cmp_232_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_232_weight_rsc_dat = step_mux_133_itm_1;
  wire[0:0] input_reg_and_471_nl;
  wire [7:0] nl_pe_0_0_run_cmp_233_input_in_rsc_dat;
  assign input_reg_and_471_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_233_input_in_rsc_dat = MUX_v_8_2_2(input_reg_8_1_sva,
      pe_0_0_run_cmp_249_input_out_rsc_z, input_reg_and_471_nl);
  wire[0:0] psum_reg_and_489_nl;
  wire [15:0] nl_pe_0_0_run_cmp_233_psum_in_rsc_dat;
  assign psum_reg_and_489_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_233_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_2_sva, pe_0_0_run_cmp_234_psum_out_rsc_z,
      psum_reg_and_489_nl);
  wire [7:0] nl_pe_0_0_run_cmp_233_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_233_weight_rsc_dat = step_mux_117_itm_1;
  wire[0:0] input_reg_and_472_nl;
  wire [7:0] nl_pe_0_0_run_cmp_234_input_in_rsc_dat;
  assign input_reg_and_472_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_234_input_in_rsc_dat = MUX_v_8_2_2(input_reg_7_1_sva,
      pe_0_0_run_cmp_250_input_out_rsc_z, input_reg_and_472_nl);
  wire[0:0] psum_reg_and_490_nl;
  wire [15:0] nl_pe_0_0_run_cmp_234_psum_in_rsc_dat;
  assign psum_reg_and_490_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_234_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_2_sva, pe_0_0_run_cmp_235_psum_out_rsc_z,
      psum_reg_and_490_nl);
  wire [7:0] nl_pe_0_0_run_cmp_234_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_234_weight_rsc_dat = step_mux_101_itm_1;
  wire[0:0] input_reg_and_473_nl;
  wire [7:0] nl_pe_0_0_run_cmp_235_input_in_rsc_dat;
  assign input_reg_and_473_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_235_input_in_rsc_dat = MUX_v_8_2_2(input_reg_6_1_sva,
      pe_0_0_run_cmp_251_input_out_rsc_z, input_reg_and_473_nl);
  wire[0:0] psum_reg_and_491_nl;
  wire [15:0] nl_pe_0_0_run_cmp_235_psum_in_rsc_dat;
  assign psum_reg_and_491_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_235_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_2_sva, pe_0_0_run_cmp_236_psum_out_rsc_z,
      psum_reg_and_491_nl);
  wire [7:0] nl_pe_0_0_run_cmp_235_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_235_weight_rsc_dat = step_mux_85_itm_1;
  wire[0:0] input_reg_and_474_nl;
  wire [7:0] nl_pe_0_0_run_cmp_236_input_in_rsc_dat;
  assign input_reg_and_474_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_236_input_in_rsc_dat = MUX_v_8_2_2(input_reg_5_1_sva,
      pe_0_0_run_cmp_252_input_out_rsc_z, input_reg_and_474_nl);
  wire[0:0] psum_reg_and_492_nl;
  wire [15:0] nl_pe_0_0_run_cmp_236_psum_in_rsc_dat;
  assign psum_reg_and_492_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_236_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_2_sva, pe_0_0_run_cmp_237_psum_out_rsc_z,
      psum_reg_and_492_nl);
  wire [7:0] nl_pe_0_0_run_cmp_236_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_236_weight_rsc_dat = step_mux_69_itm_1;
  wire[0:0] input_reg_and_475_nl;
  wire [7:0] nl_pe_0_0_run_cmp_237_input_in_rsc_dat;
  assign input_reg_and_475_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_237_input_in_rsc_dat = MUX_v_8_2_2(input_reg_4_1_sva,
      pe_0_0_run_cmp_253_input_out_rsc_z, input_reg_and_475_nl);
  wire[0:0] psum_reg_and_493_nl;
  wire [15:0] nl_pe_0_0_run_cmp_237_psum_in_rsc_dat;
  assign psum_reg_and_493_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_237_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_2_sva, pe_0_0_run_cmp_238_psum_out_rsc_z,
      psum_reg_and_493_nl);
  wire [7:0] nl_pe_0_0_run_cmp_237_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_237_weight_rsc_dat = step_mux_53_itm_1;
  wire[0:0] input_reg_and_476_nl;
  wire [7:0] nl_pe_0_0_run_cmp_238_input_in_rsc_dat;
  assign input_reg_and_476_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_238_input_in_rsc_dat = MUX_v_8_2_2(input_reg_3_1_sva,
      pe_0_0_run_cmp_254_input_out_rsc_z, input_reg_and_476_nl);
  wire[0:0] psum_reg_and_494_nl;
  wire [15:0] nl_pe_0_0_run_cmp_238_psum_in_rsc_dat;
  assign psum_reg_and_494_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_238_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_2_sva, pe_0_0_run_cmp_239_psum_out_rsc_z,
      psum_reg_and_494_nl);
  wire [7:0] nl_pe_0_0_run_cmp_238_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_238_weight_rsc_dat = step_mux_37_itm_1;
  wire[0:0] input_reg_and_477_nl;
  wire [7:0] nl_pe_0_0_run_cmp_239_input_in_rsc_dat;
  assign input_reg_and_477_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_239_input_in_rsc_dat = MUX_v_8_2_2(input_reg_2_1_sva,
      pe_0_0_run_cmp_255_input_out_rsc_z, input_reg_and_477_nl);
  wire[0:0] psum_reg_and_495_nl;
  wire [15:0] nl_pe_0_0_run_cmp_239_psum_in_rsc_dat;
  assign psum_reg_and_495_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_239_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_2_sva, pe_0_0_run_cmp_240_psum_out_rsc_z,
      psum_reg_and_495_nl);
  wire [7:0] nl_pe_0_0_run_cmp_239_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_239_weight_rsc_dat = step_mux_21_itm_1;
  wire[0:0] input_reg_and_478_nl;
  wire [7:0] nl_pe_0_0_run_cmp_240_input_in_rsc_dat;
  assign input_reg_and_478_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_240_input_in_rsc_dat = MUX_v_8_2_2(input_reg_1_1_sva,
      pe_0_0_run_cmp_input_out_rsc_z, input_reg_and_478_nl);
  wire [7:0] nl_pe_0_0_run_cmp_240_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_240_weight_rsc_dat = step_mux_5_itm_1;
  wire[0:0] psum_reg_and_496_nl;
  wire [15:0] nl_pe_0_0_run_cmp_241_psum_in_rsc_dat;
  assign psum_reg_and_496_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_241_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_15_1_sva,
      pe_0_0_run_cmp_242_psum_out_rsc_z, psum_reg_and_496_nl);
  wire [7:0] nl_pe_0_0_run_cmp_241_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_241_weight_rsc_dat = step_mux_244_itm_1;
  wire[0:0] psum_reg_and_497_nl;
  wire [15:0] nl_pe_0_0_run_cmp_242_psum_in_rsc_dat;
  assign psum_reg_and_497_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_242_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_14_1_sva,
      pe_0_0_run_cmp_243_psum_out_rsc_z, psum_reg_and_497_nl);
  wire [7:0] nl_pe_0_0_run_cmp_242_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_242_weight_rsc_dat = step_mux_228_itm_1;
  wire[0:0] psum_reg_and_498_nl;
  wire [15:0] nl_pe_0_0_run_cmp_243_psum_in_rsc_dat;
  assign psum_reg_and_498_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_243_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_13_1_sva,
      pe_0_0_run_cmp_244_psum_out_rsc_z, psum_reg_and_498_nl);
  wire [7:0] nl_pe_0_0_run_cmp_243_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_243_weight_rsc_dat = step_mux_212_itm_1;
  wire[0:0] psum_reg_and_499_nl;
  wire [15:0] nl_pe_0_0_run_cmp_244_psum_in_rsc_dat;
  assign psum_reg_and_499_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_244_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_12_1_sva,
      pe_0_0_run_cmp_245_psum_out_rsc_z, psum_reg_and_499_nl);
  wire [7:0] nl_pe_0_0_run_cmp_244_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_244_weight_rsc_dat = step_mux_196_itm_1;
  wire[0:0] psum_reg_and_500_nl;
  wire [15:0] nl_pe_0_0_run_cmp_245_psum_in_rsc_dat;
  assign psum_reg_and_500_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_245_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_11_1_sva,
      pe_0_0_run_cmp_246_psum_out_rsc_z, psum_reg_and_500_nl);
  wire [7:0] nl_pe_0_0_run_cmp_245_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_245_weight_rsc_dat = step_mux_180_itm_1;
  wire[0:0] psum_reg_and_501_nl;
  wire [15:0] nl_pe_0_0_run_cmp_246_psum_in_rsc_dat;
  assign psum_reg_and_501_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_246_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_10_1_sva,
      pe_0_0_run_cmp_247_psum_out_rsc_z, psum_reg_and_501_nl);
  wire [7:0] nl_pe_0_0_run_cmp_246_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_246_weight_rsc_dat = step_mux_164_itm_1;
  wire[0:0] psum_reg_and_502_nl;
  wire [15:0] nl_pe_0_0_run_cmp_247_psum_in_rsc_dat;
  assign psum_reg_and_502_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_247_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_9_1_sva, pe_0_0_run_cmp_248_psum_out_rsc_z,
      psum_reg_and_502_nl);
  wire [7:0] nl_pe_0_0_run_cmp_247_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_247_weight_rsc_dat = step_mux_148_itm_1;
  wire[0:0] psum_reg_and_503_nl;
  wire [15:0] nl_pe_0_0_run_cmp_248_psum_in_rsc_dat;
  assign psum_reg_and_503_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_248_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_8_1_sva, pe_0_0_run_cmp_249_psum_out_rsc_z,
      psum_reg_and_503_nl);
  wire [7:0] nl_pe_0_0_run_cmp_248_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_248_weight_rsc_dat = step_mux_132_itm_1;
  wire[0:0] psum_reg_and_504_nl;
  wire [15:0] nl_pe_0_0_run_cmp_249_psum_in_rsc_dat;
  assign psum_reg_and_504_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_249_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_7_1_sva, pe_0_0_run_cmp_250_psum_out_rsc_z,
      psum_reg_and_504_nl);
  wire [7:0] nl_pe_0_0_run_cmp_249_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_249_weight_rsc_dat = step_mux_116_itm_1;
  wire[0:0] psum_reg_and_505_nl;
  wire [15:0] nl_pe_0_0_run_cmp_250_psum_in_rsc_dat;
  assign psum_reg_and_505_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_250_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_6_1_sva, pe_0_0_run_cmp_251_psum_out_rsc_z,
      psum_reg_and_505_nl);
  wire [7:0] nl_pe_0_0_run_cmp_250_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_250_weight_rsc_dat = step_mux_100_itm_1;
  wire[0:0] psum_reg_and_506_nl;
  wire [15:0] nl_pe_0_0_run_cmp_251_psum_in_rsc_dat;
  assign psum_reg_and_506_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_251_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_5_1_sva, pe_0_0_run_cmp_252_psum_out_rsc_z,
      psum_reg_and_506_nl);
  wire [7:0] nl_pe_0_0_run_cmp_251_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_251_weight_rsc_dat = step_mux_84_itm_1;
  wire[0:0] psum_reg_and_507_nl;
  wire [15:0] nl_pe_0_0_run_cmp_252_psum_in_rsc_dat;
  assign psum_reg_and_507_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_252_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_4_1_sva, pe_0_0_run_cmp_253_psum_out_rsc_z,
      psum_reg_and_507_nl);
  wire [7:0] nl_pe_0_0_run_cmp_252_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_252_weight_rsc_dat = step_mux_68_itm_1;
  wire[0:0] psum_reg_and_508_nl;
  wire [15:0] nl_pe_0_0_run_cmp_253_psum_in_rsc_dat;
  assign psum_reg_and_508_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_253_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_3_1_sva, pe_0_0_run_cmp_254_psum_out_rsc_z,
      psum_reg_and_508_nl);
  wire [7:0] nl_pe_0_0_run_cmp_253_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_253_weight_rsc_dat = step_mux_52_itm_1;
  wire[0:0] psum_reg_and_509_nl;
  wire [15:0] nl_pe_0_0_run_cmp_254_psum_in_rsc_dat;
  assign psum_reg_and_509_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_254_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_2_1_sva, pe_0_0_run_cmp_255_psum_out_rsc_z,
      psum_reg_and_509_nl);
  wire [7:0] nl_pe_0_0_run_cmp_254_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_254_weight_rsc_dat = step_mux_36_itm_1;
  wire[0:0] psum_reg_and_510_nl;
  wire [15:0] nl_pe_0_0_run_cmp_255_psum_in_rsc_dat;
  assign psum_reg_and_510_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_pe_0_0_run_cmp_255_psum_in_rsc_dat = MUX_v_16_2_2(psum_reg_1_1_sva, pe_0_0_run_cmp_psum_out_rsc_z,
      psum_reg_and_510_nl);
  wire [7:0] nl_pe_0_0_run_cmp_255_weight_rsc_dat;
  assign nl_pe_0_0_run_cmp_255_weight_rsc_dat = step_mux_20_itm_1;
  wire[0:0] step_if_2_aelse_1_not_16_nl;
  wire [15:0] nl_accum_fifo_0_run_cmp_input_rsc_dat;
  assign step_if_2_aelse_1_not_16_nl = ~ step_and_10_psp;
  assign nl_accum_fifo_0_run_cmp_input_rsc_dat = MUX_v_16_2_2(16'b0000000000000000,
      accumulation_buffer_rsc_0_0_i_q_d_mxwt, (step_if_2_aelse_1_not_16_nl));
  wire[0:0] psum_reg_and_511_nl;
  wire [15:0] nl_accum_fifo_0_run_cmp_1_input_rsc_dat;
  assign psum_reg_and_511_nl = and_dcpl_10 & (fsm_output[1]);
  assign nl_accum_fifo_0_run_cmp_1_input_rsc_dat = MUX_v_16_2_2(psum_reg_16_16_sva,
      pe_0_0_run_cmp_1_psum_out_rsc_z, psum_reg_and_511_nl);
  wire [7:0] nl_input_fifo_0_run_cmp_input_rsc_dat;
  assign nl_input_fifo_0_run_cmp_input_rsc_dat = step_in_col_value_lpi_1_dfm_mx0[7:0];
  wire [255:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat
      = {output_rsci_idat_255_240 , output_rsci_idat_239_224 , output_rsci_idat_223_208
      , output_rsci_idat_207_192 , output_rsci_idat_191_176 , output_rsci_idat_175_160
      , output_rsci_idat_159_144 , output_rsci_idat_143_128 , output_rsci_idat_127_112
      , output_rsci_idat_111_96 , output_rsci_idat_95_80 , output_rsci_idat_79_64
      , output_rsci_idat_63_48 , output_rsci_idat_47_32 , output_rsci_idat_31_16
      , output_rsci_idat_15_0};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_radr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_radr_d_run
      = {2'b0, step_step_lpi_1_dfm_1[5:0]};
  wire [7:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run
      = {2'b0, step_if_3_for_1_operator_16_false_acc_cse_sva_3};
  Fifo_ODTYPE_16  accum_fifo_15_rsci (
      .input_rsc_dat(nl_accum_fifo_15_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_15_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_16  output_fifo_0_rsci (
      .input_rsc_dat(nl_output_fifo_0_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_0_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_15  accum_fifo_14_rsci (
      .input_rsc_dat(nl_accum_fifo_14_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_15  output_fifo_1_rsci (
      .input_rsc_dat(nl_output_fifo_1_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_14  accum_fifo_13_rsci (
      .input_rsc_dat(nl_accum_fifo_13_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_14  output_fifo_2_rsci (
      .input_rsc_dat(nl_output_fifo_2_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_13  accum_fifo_12_rsci (
      .input_rsc_dat(nl_accum_fifo_12_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_13  output_fifo_3_rsci (
      .input_rsc_dat(nl_output_fifo_3_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_12  accum_fifo_11_rsci (
      .input_rsc_dat(nl_accum_fifo_11_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_12  output_fifo_4_rsci (
      .input_rsc_dat(nl_output_fifo_4_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_11  accum_fifo_10_rsci (
      .input_rsc_dat(nl_accum_fifo_10_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_11  output_fifo_5_rsci (
      .input_rsc_dat(nl_output_fifo_5_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_10  accum_fifo_9_rsci (
      .input_rsc_dat(nl_accum_fifo_9_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_10  output_fifo_6_rsci (
      .input_rsc_dat(nl_output_fifo_6_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_9  accum_fifo_8_rsci (
      .input_rsc_dat(nl_accum_fifo_8_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_9  output_fifo_7_rsci (
      .input_rsc_dat(nl_output_fifo_7_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_8  accum_fifo_7_rsci (
      .input_rsc_dat(nl_accum_fifo_7_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_8  output_fifo_8_rsci (
      .input_rsc_dat(nl_output_fifo_8_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_7  accum_fifo_6_rsci (
      .input_rsc_dat(nl_accum_fifo_6_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_7  output_fifo_9_rsci (
      .input_rsc_dat(nl_output_fifo_9_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_6  accum_fifo_5_rsci (
      .input_rsc_dat(nl_accum_fifo_5_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_6  output_fifo_10_rsci (
      .input_rsc_dat(nl_output_fifo_10_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_5  accum_fifo_4_rsci (
      .input_rsc_dat(nl_accum_fifo_4_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_5  output_fifo_11_rsci (
      .input_rsc_dat(nl_output_fifo_11_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_4  accum_fifo_3_rsci (
      .input_rsc_dat(nl_accum_fifo_3_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_4  output_fifo_12_rsci (
      .input_rsc_dat(nl_output_fifo_12_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_3  accum_fifo_2_rsci (
      .input_rsc_dat(nl_accum_fifo_2_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_3  output_fifo_13_rsci (
      .input_rsc_dat(nl_output_fifo_13_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_2  accum_fifo_1_rsci (
      .input_rsc_dat(nl_accum_fifo_1_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_2  output_fifo_14_rsci (
      .input_rsc_dat(nl_output_fifo_14_rsci_input_rsc_dat[15:0]),
      .output_rsc_z(output_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_IDTYPE_16  input_fifo_15_rsci (
      .input_rsc_dat(nl_input_fifo_15_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_15_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_15  input_fifo_14_rsci (
      .input_rsc_dat(nl_input_fifo_14_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_14_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_14  input_fifo_13_rsci (
      .input_rsc_dat(nl_input_fifo_13_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_13_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_13  input_fifo_12_rsci (
      .input_rsc_dat(nl_input_fifo_12_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_12_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_12  input_fifo_11_rsci (
      .input_rsc_dat(nl_input_fifo_11_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_11_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_11  input_fifo_10_rsci (
      .input_rsc_dat(nl_input_fifo_10_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_10_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_10  input_fifo_9_rsci (
      .input_rsc_dat(nl_input_fifo_9_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_9_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_9  input_fifo_8_rsci (
      .input_rsc_dat(nl_input_fifo_8_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_8_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_8  input_fifo_7_rsci (
      .input_rsc_dat(nl_input_fifo_7_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_7_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_7  input_fifo_6_rsci (
      .input_rsc_dat(nl_input_fifo_6_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_6_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_6  input_fifo_5_rsci (
      .input_rsc_dat(nl_input_fifo_5_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_5_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_5  input_fifo_4_rsci (
      .input_rsc_dat(nl_input_fifo_4_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_4_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_4  input_fifo_3_rsci (
      .input_rsc_dat(nl_input_fifo_3_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_3_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_3  input_fifo_2_rsci (
      .input_rsc_dat(nl_input_fifo_2_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_2_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_IDTYPE_2  input_fifo_1_rsci (
      .input_rsc_dat(nl_input_fifo_1_rsci_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_1_rsci_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp (
      .input_in_rsc_dat(input_fifo_0_run_cmp_output_rsc_z),
      .psum_in_rsc_dat(accum_fifo_0_run_cmp_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_1 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_1_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_1_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_1_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_1_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_1_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_2 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_2_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_2_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_2_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_2_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_2_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_3 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_3_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_3_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_3_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_3_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_3_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_4 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_4_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_4_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_4_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_4_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_4_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_5 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_5_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_5_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_5_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_5_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_5_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_6 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_6_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_6_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_6_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_6_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_6_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_7 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_7_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_7_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_7_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_7_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_7_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_8 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_8_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_8_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_8_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_8_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_8_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_9 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_9_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_9_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_9_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_9_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_9_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_10 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_10_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_10_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_10_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_10_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_10_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_11 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_11_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_11_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_11_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_11_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_11_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_12 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_12_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_12_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_12_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_12_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_12_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_13 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_13_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_13_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_13_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_13_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_13_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_14 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_14_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_14_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_14_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_14_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_14_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_15 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_15_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_15_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_15_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_15_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_15_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_16 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_16_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_15_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_16_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_16_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_16_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_17 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_17_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_17_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_17_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_17_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_17_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_18 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_18_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_18_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_18_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_18_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_18_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_19 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_19_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_19_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_19_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_19_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_19_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_20 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_20_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_20_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_20_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_20_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_20_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_21 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_21_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_21_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_21_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_21_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_21_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_22 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_22_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_22_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_22_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_22_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_22_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_23 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_23_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_23_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_23_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_23_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_23_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_24 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_24_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_24_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_24_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_24_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_24_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_25 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_25_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_25_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_25_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_25_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_25_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_26 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_26_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_26_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_26_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_26_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_26_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_27 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_27_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_27_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_27_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_27_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_27_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_28 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_28_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_28_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_28_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_28_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_28_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_29 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_29_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_29_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_29_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_29_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_29_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_30 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_30_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_30_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_30_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_30_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_30_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_31 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_31_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_31_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_31_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_31_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_31_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_32 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_32_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_14_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_32_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_32_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_32_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_33 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_33_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_33_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_33_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_33_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_33_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_34 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_34_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_34_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_34_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_34_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_34_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_35 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_35_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_35_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_35_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_35_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_35_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_36 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_36_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_36_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_36_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_36_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_36_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_37 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_37_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_37_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_37_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_37_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_37_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_38 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_38_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_38_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_38_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_38_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_38_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_39 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_39_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_39_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_39_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_39_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_39_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_40 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_40_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_40_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_40_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_40_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_40_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_41 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_41_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_41_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_41_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_41_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_41_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_42 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_42_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_42_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_42_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_42_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_42_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_43 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_43_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_43_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_43_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_43_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_43_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_44 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_44_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_44_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_44_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_44_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_44_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_45 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_45_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_45_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_45_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_45_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_45_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_46 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_46_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_46_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_46_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_46_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_46_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_47 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_47_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_47_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_47_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_47_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_47_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_48 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_48_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_13_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_48_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_48_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_48_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_49 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_49_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_49_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_49_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_49_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_49_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_50 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_50_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_50_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_50_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_50_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_50_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_51 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_51_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_51_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_51_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_51_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_51_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_52 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_52_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_52_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_52_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_52_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_52_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_53 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_53_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_53_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_53_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_53_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_53_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_54 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_54_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_54_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_54_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_54_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_54_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_55 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_55_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_55_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_55_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_55_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_55_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_56 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_56_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_56_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_56_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_56_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_56_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_57 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_57_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_57_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_57_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_57_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_57_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_58 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_58_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_58_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_58_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_58_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_58_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_59 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_59_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_59_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_59_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_59_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_59_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_60 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_60_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_60_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_60_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_60_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_60_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_61 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_61_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_61_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_61_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_61_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_61_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_62 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_62_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_62_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_62_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_62_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_62_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_63 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_63_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_63_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_63_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_63_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_63_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_64 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_64_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_12_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_64_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_64_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_64_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_65 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_65_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_65_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_65_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_65_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_65_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_66 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_66_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_66_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_66_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_66_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_66_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_67 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_67_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_67_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_67_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_67_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_67_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_68 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_68_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_68_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_68_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_68_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_68_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_69 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_69_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_69_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_69_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_69_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_69_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_70 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_70_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_70_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_70_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_70_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_70_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_71 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_71_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_71_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_71_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_71_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_71_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_72 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_72_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_72_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_72_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_72_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_72_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_73 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_73_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_73_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_73_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_73_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_73_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_74 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_74_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_74_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_74_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_74_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_74_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_75 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_75_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_75_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_75_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_75_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_75_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_76 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_76_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_76_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_76_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_76_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_76_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_77 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_77_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_77_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_77_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_77_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_77_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_78 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_78_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_78_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_78_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_78_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_78_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_79 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_79_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_79_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_79_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_79_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_79_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_80 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_80_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_11_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_80_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_80_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_80_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_81 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_81_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_81_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_81_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_81_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_81_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_82 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_82_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_82_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_82_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_82_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_82_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_83 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_83_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_83_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_83_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_83_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_83_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_84 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_84_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_84_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_84_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_84_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_84_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_85 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_85_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_85_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_85_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_85_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_85_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_86 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_86_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_86_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_86_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_86_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_86_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_87 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_87_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_87_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_87_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_87_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_87_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_88 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_88_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_88_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_88_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_88_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_88_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_89 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_89_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_89_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_89_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_89_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_89_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_90 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_90_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_90_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_90_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_90_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_90_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_91 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_91_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_91_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_91_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_91_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_91_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_92 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_92_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_92_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_92_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_92_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_92_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_93 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_93_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_93_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_93_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_93_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_93_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_94 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_94_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_94_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_94_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_94_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_94_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_95 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_95_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_95_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_95_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_95_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_95_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_96 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_96_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_10_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_96_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_96_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_96_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_97 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_97_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_97_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_97_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_97_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_97_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_98 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_98_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_98_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_98_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_98_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_98_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_99 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_99_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_99_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_99_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_99_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_99_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_100 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_100_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_100_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_100_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_100_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_100_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_101 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_101_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_101_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_101_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_101_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_101_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_102 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_102_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_102_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_102_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_102_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_102_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_103 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_103_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_103_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_103_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_103_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_103_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_104 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_104_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_104_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_104_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_104_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_104_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_105 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_105_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_105_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_105_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_105_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_105_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_106 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_106_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_106_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_106_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_106_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_106_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_107 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_107_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_107_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_107_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_107_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_107_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_108 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_108_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_108_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_108_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_108_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_108_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_109 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_109_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_109_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_109_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_109_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_109_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_110 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_110_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_110_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_110_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_110_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_110_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_111 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_111_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_111_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_111_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_111_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_111_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_112 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_112_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_9_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_112_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_112_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_112_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_113 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_113_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_113_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_113_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_113_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_113_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_114 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_114_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_114_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_114_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_114_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_114_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_115 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_115_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_115_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_115_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_115_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_115_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_116 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_116_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_116_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_116_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_116_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_116_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_117 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_117_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_117_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_117_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_117_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_117_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_118 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_118_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_118_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_118_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_118_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_118_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_119 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_119_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_119_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_119_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_119_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_119_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_120 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_120_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_120_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_120_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_120_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_120_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_121 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_121_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_121_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_121_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_121_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_121_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_122 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_122_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_122_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_122_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_122_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_122_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_123 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_123_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_123_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_123_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_123_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_123_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_124 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_124_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_124_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_124_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_124_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_124_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_125 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_125_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_125_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_125_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_125_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_125_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_126 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_126_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_126_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_126_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_126_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_126_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_127 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_127_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_127_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_127_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_127_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_127_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_128 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_128_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_8_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_128_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_128_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_128_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_129 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_129_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_129_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_129_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_129_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_129_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_130 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_130_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_130_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_130_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_130_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_130_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_131 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_131_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_131_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_131_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_131_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_131_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_132 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_132_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_132_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_132_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_132_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_132_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_133 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_133_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_133_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_133_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_133_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_133_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_134 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_134_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_134_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_134_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_134_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_134_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_135 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_135_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_135_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_135_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_135_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_135_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_136 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_136_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_136_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_136_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_136_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_136_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_137 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_137_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_137_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_137_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_137_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_137_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_138 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_138_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_138_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_138_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_138_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_138_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_139 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_139_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_139_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_139_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_139_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_139_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_140 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_140_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_140_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_140_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_140_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_140_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_141 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_141_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_141_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_141_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_141_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_141_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_142 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_142_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_142_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_142_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_142_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_142_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_143 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_143_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_143_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_143_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_143_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_143_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_144 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_144_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_7_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_144_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_144_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_144_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_145 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_145_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_145_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_145_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_145_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_145_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_146 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_146_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_146_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_146_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_146_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_146_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_147 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_147_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_147_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_147_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_147_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_147_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_148 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_148_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_148_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_148_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_148_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_148_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_149 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_149_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_149_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_149_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_149_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_149_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_150 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_150_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_150_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_150_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_150_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_150_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_151 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_151_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_151_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_151_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_151_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_151_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_152 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_152_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_152_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_152_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_152_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_152_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_153 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_153_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_153_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_153_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_153_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_153_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_154 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_154_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_154_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_154_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_154_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_154_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_155 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_155_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_155_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_155_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_155_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_155_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_156 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_156_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_156_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_156_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_156_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_156_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_157 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_157_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_157_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_157_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_157_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_157_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_158 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_158_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_158_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_158_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_158_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_158_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_159 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_159_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_159_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_159_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_159_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_159_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_160 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_160_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_6_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_160_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_160_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_160_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_161 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_161_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_161_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_161_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_161_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_161_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_162 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_162_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_162_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_162_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_162_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_162_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_163 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_163_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_163_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_163_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_163_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_163_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_164 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_164_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_164_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_164_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_164_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_164_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_165 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_165_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_165_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_165_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_165_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_165_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_166 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_166_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_166_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_166_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_166_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_166_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_167 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_167_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_167_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_167_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_167_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_167_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_168 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_168_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_168_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_168_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_168_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_168_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_169 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_169_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_169_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_169_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_169_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_169_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_170 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_170_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_170_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_170_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_170_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_170_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_171 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_171_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_171_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_171_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_171_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_171_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_172 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_172_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_172_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_172_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_172_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_172_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_173 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_173_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_173_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_173_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_173_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_173_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_174 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_174_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_174_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_174_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_174_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_174_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_175 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_175_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_175_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_175_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_175_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_175_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_176 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_176_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_5_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_176_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_176_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_176_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_177 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_177_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_177_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_177_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_177_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_177_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_178 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_178_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_178_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_178_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_178_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_178_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_179 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_179_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_179_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_179_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_179_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_179_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_180 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_180_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_180_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_180_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_180_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_180_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_181 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_181_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_181_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_181_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_181_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_181_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_182 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_182_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_182_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_182_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_182_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_182_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_183 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_183_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_183_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_183_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_183_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_183_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_184 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_184_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_184_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_184_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_184_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_184_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_185 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_185_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_185_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_185_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_185_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_185_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_186 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_186_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_186_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_186_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_186_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_186_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_187 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_187_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_187_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_187_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_187_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_187_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_188 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_188_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_188_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_188_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_188_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_188_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_189 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_189_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_189_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_189_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_189_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_189_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_190 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_190_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_190_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_190_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_190_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_190_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_191 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_191_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_191_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_191_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_191_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_191_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_192 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_192_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_4_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_192_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_192_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_192_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_193 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_193_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_193_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_193_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_193_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_193_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_194 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_194_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_194_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_194_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_194_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_194_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_195 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_195_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_195_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_195_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_195_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_195_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_196 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_196_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_196_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_196_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_196_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_196_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_197 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_197_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_197_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_197_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_197_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_197_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_198 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_198_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_198_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_198_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_198_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_198_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_199 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_199_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_199_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_199_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_199_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_199_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_200 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_200_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_200_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_200_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_200_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_200_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_201 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_201_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_201_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_201_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_201_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_201_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_202 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_202_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_202_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_202_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_202_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_202_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_203 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_203_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_203_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_203_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_203_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_203_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_204 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_204_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_204_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_204_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_204_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_204_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_205 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_205_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_205_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_205_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_205_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_205_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_206 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_206_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_206_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_206_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_206_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_206_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_207 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_207_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_207_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_207_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_207_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_207_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_208 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_208_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_3_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_208_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_208_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_208_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_209 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_209_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_209_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_209_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_209_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_209_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_210 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_210_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_210_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_210_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_210_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_210_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_211 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_211_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_211_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_211_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_211_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_211_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_212 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_212_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_212_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_212_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_212_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_212_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_213 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_213_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_213_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_213_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_213_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_213_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_214 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_214_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_214_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_214_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_214_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_214_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_215 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_215_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_215_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_215_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_215_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_215_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_216 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_216_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_216_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_216_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_216_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_216_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_217 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_217_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_217_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_217_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_217_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_217_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_218 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_218_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_218_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_218_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_218_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_218_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_219 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_219_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_219_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_219_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_219_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_219_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_220 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_220_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_220_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_220_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_220_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_220_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_221 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_221_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_221_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_221_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_221_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_221_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_222 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_222_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_222_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_222_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_222_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_222_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_223 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_223_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_223_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_223_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_223_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_223_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_224 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_224_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_2_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_224_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_224_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_224_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_225 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_225_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_225_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_225_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_225_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_225_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_226 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_226_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_226_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_226_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_226_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_226_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_227 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_227_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_227_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_227_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_227_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_227_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_228 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_228_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_228_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_228_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_228_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_228_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_229 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_229_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_229_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_229_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_229_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_229_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_230 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_230_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_230_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_230_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_230_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_230_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_231 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_231_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_231_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_231_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_231_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_231_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_232 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_232_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_232_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_232_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_232_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_232_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_233 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_233_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_233_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_233_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_233_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_233_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_234 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_234_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_234_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_234_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_234_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_234_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_235 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_235_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_235_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_235_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_235_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_235_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_236 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_236_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_236_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_236_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_236_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_236_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_237 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_237_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_237_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_237_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_237_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_237_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_238 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_238_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_238_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_238_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_238_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_238_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_239 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_239_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_239_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_239_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_239_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_239_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_240 (
      .input_in_rsc_dat(nl_pe_0_0_run_cmp_240_input_in_rsc_dat[7:0]),
      .psum_in_rsc_dat(accum_fifo_1_rsci_output_rsc_z),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_240_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_240_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_240_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_241 (
      .input_in_rsc_dat(input_fifo_15_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_241_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_241_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_241_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_241_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_242 (
      .input_in_rsc_dat(input_fifo_14_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_242_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_242_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_242_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_242_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_243 (
      .input_in_rsc_dat(input_fifo_13_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_243_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_243_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_243_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_243_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_244 (
      .input_in_rsc_dat(input_fifo_12_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_244_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_244_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_244_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_244_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_245 (
      .input_in_rsc_dat(input_fifo_11_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_245_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_245_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_245_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_245_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_246 (
      .input_in_rsc_dat(input_fifo_10_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_246_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_246_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_246_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_246_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_247 (
      .input_in_rsc_dat(input_fifo_9_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_247_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_247_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_247_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_247_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_248 (
      .input_in_rsc_dat(input_fifo_8_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_248_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_248_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_248_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_248_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_249 (
      .input_in_rsc_dat(input_fifo_7_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_249_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_249_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_249_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_249_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_250 (
      .input_in_rsc_dat(input_fifo_6_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_250_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_250_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_250_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_250_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_251 (
      .input_in_rsc_dat(input_fifo_5_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_251_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_251_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_251_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_251_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_252 (
      .input_in_rsc_dat(input_fifo_4_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_252_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_252_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_252_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_252_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_253 (
      .input_in_rsc_dat(input_fifo_3_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_253_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_253_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_253_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_253_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_254 (
      .input_in_rsc_dat(input_fifo_2_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_254_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_254_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_254_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_254_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  ProcessingElement_IDTYPE_ODTYPE  pe_0_0_run_cmp_255 (
      .input_in_rsc_dat(input_fifo_1_rsci_output_rsc_z),
      .psum_in_rsc_dat(nl_pe_0_0_run_cmp_255_psum_in_rsc_dat[15:0]),
      .weight_rsc_dat(nl_pe_0_0_run_cmp_255_weight_rsc_dat[7:0]),
      .input_out_rsc_z(pe_0_0_run_cmp_255_input_out_rsc_z),
      .psum_out_rsc_z(pe_0_0_run_cmp_255_psum_out_rsc_z),
      .clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .arst_n(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_ODTYPE_1  accum_fifo_0_run_cmp (
      .input_rsc_dat(nl_accum_fifo_0_run_cmp_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_0_run_cmp_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  Fifo_ODTYPE_1  accum_fifo_0_run_cmp_1 (
      .input_rsc_dat(nl_accum_fifo_0_run_cmp_1_input_rsc_dat[15:0]),
      .output_rsc_z(accum_fifo_0_run_cmp_1_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_1)
    );
  Fifo_IDTYPE_1  input_fifo_0_run_cmp (
      .input_rsc_dat(nl_input_fifo_0_run_cmp_input_rsc_dat[7:0]),
      .output_rsc_z(input_fifo_0_run_cmp_output_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ccs_ccore_arst(arst_n),
      .ccs_ccore_start_rsc_dat(and_dcpl_4)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_input_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .run_wen(run_wen),
      .input_rsci_oswt(reg_input_rsci_irdy_run_psct_cse),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .input_rsci_idat_mxwt(input_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_weight_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weight_rsc_dat(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .run_wen(run_wen),
      .weight_rsci_oswt(reg_weight_rsci_irdy_run_psct_cse),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .weight_rsci_idat_mxwt(weight_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .run_wen(run_wen),
      .output_rsci_oswt(reg_output_rsci_ivld_run_psct_cse),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .output_rsci_idat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_output_rsci_inst_output_rsci_idat[255:0])
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_loopIndicesIn_rsci_oswt_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_loopIndicesIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(reg_loopIndicesIn_rsci_oswt_cse),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_0_i_radr_d(accumulation_buffer_rsc_0_0_i_radr_d_reg),
      .accumulation_buffer_rsc_0_0_i_wadr_d(accumulation_buffer_rsc_0_0_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_0_i_q_d(accumulation_buffer_rsc_0_0_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_0_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_0_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_0_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_0_i_1_inst_accumulation_buffer_rsc_0_0_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_0_i_q_d_mxwt(accumulation_buffer_rsc_0_0_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_0_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_0_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_0_i_we_d_pff(accumulation_buffer_rsc_0_0_i_we_d_iff),
      .accumulation_buffer_rsc_0_0_i_re_d_pff(accumulation_buffer_rsc_0_0_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_1_i_radr_d(accumulation_buffer_rsc_0_1_i_radr_d_reg),
      .accumulation_buffer_rsc_0_1_i_wadr_d(accumulation_buffer_rsc_0_1_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_1_i_q_d(accumulation_buffer_rsc_0_1_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_1_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_1_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_1_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_1_i_1_inst_accumulation_buffer_rsc_0_1_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_1_i_q_d_mxwt(accumulation_buffer_rsc_0_1_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_1_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_1_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_1_i_we_d_pff(accumulation_buffer_rsc_0_1_i_we_d_iff),
      .accumulation_buffer_rsc_0_1_i_re_d_pff(accumulation_buffer_rsc_0_1_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_2_i_radr_d(accumulation_buffer_rsc_0_2_i_radr_d_reg),
      .accumulation_buffer_rsc_0_2_i_wadr_d(accumulation_buffer_rsc_0_2_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_2_i_q_d(accumulation_buffer_rsc_0_2_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_2_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_2_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_2_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_2_i_1_inst_accumulation_buffer_rsc_0_2_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_2_i_q_d_mxwt(accumulation_buffer_rsc_0_2_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_2_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_2_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_2_i_we_d_pff(accumulation_buffer_rsc_0_2_i_we_d_iff),
      .accumulation_buffer_rsc_0_2_i_re_d_pff(accumulation_buffer_rsc_0_2_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_3_i_radr_d(accumulation_buffer_rsc_0_3_i_radr_d_reg),
      .accumulation_buffer_rsc_0_3_i_wadr_d(accumulation_buffer_rsc_0_3_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_3_i_q_d(accumulation_buffer_rsc_0_3_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_3_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_3_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_3_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_3_i_1_inst_accumulation_buffer_rsc_0_3_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_3_i_q_d_mxwt(accumulation_buffer_rsc_0_3_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_3_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_3_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_3_i_we_d_pff(accumulation_buffer_rsc_0_3_i_we_d_iff),
      .accumulation_buffer_rsc_0_3_i_re_d_pff(accumulation_buffer_rsc_0_3_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_4_i_radr_d(accumulation_buffer_rsc_0_4_i_radr_d_reg),
      .accumulation_buffer_rsc_0_4_i_wadr_d(accumulation_buffer_rsc_0_4_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_4_i_q_d(accumulation_buffer_rsc_0_4_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_4_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_4_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_4_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_4_i_1_inst_accumulation_buffer_rsc_0_4_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_4_i_q_d_mxwt(accumulation_buffer_rsc_0_4_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_4_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_4_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_4_i_we_d_pff(accumulation_buffer_rsc_0_4_i_we_d_iff),
      .accumulation_buffer_rsc_0_4_i_re_d_pff(accumulation_buffer_rsc_0_4_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_5_i_radr_d(accumulation_buffer_rsc_0_5_i_radr_d_reg),
      .accumulation_buffer_rsc_0_5_i_wadr_d(accumulation_buffer_rsc_0_5_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_5_i_q_d(accumulation_buffer_rsc_0_5_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_5_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_5_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_5_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_5_i_1_inst_accumulation_buffer_rsc_0_5_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_5_i_q_d_mxwt(accumulation_buffer_rsc_0_5_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_5_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_5_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_5_i_we_d_pff(accumulation_buffer_rsc_0_5_i_we_d_iff),
      .accumulation_buffer_rsc_0_5_i_re_d_pff(accumulation_buffer_rsc_0_5_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_6_i_radr_d(accumulation_buffer_rsc_0_6_i_radr_d_reg),
      .accumulation_buffer_rsc_0_6_i_wadr_d(accumulation_buffer_rsc_0_6_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_6_i_q_d(accumulation_buffer_rsc_0_6_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_6_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_6_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_6_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_6_i_1_inst_accumulation_buffer_rsc_0_6_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_6_i_q_d_mxwt(accumulation_buffer_rsc_0_6_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_6_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_6_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_6_i_we_d_pff(accumulation_buffer_rsc_0_6_i_we_d_iff),
      .accumulation_buffer_rsc_0_6_i_re_d_pff(accumulation_buffer_rsc_0_6_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_7_i_radr_d(accumulation_buffer_rsc_0_7_i_radr_d_reg),
      .accumulation_buffer_rsc_0_7_i_wadr_d(accumulation_buffer_rsc_0_7_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_7_i_q_d(accumulation_buffer_rsc_0_7_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_7_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_7_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_7_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_7_i_1_inst_accumulation_buffer_rsc_0_7_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_7_i_q_d_mxwt(accumulation_buffer_rsc_0_7_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_7_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_7_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_7_i_we_d_pff(accumulation_buffer_rsc_0_7_i_we_d_iff),
      .accumulation_buffer_rsc_0_7_i_re_d_pff(accumulation_buffer_rsc_0_7_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_8_i_radr_d(accumulation_buffer_rsc_0_8_i_radr_d_reg),
      .accumulation_buffer_rsc_0_8_i_wadr_d(accumulation_buffer_rsc_0_8_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_8_i_q_d(accumulation_buffer_rsc_0_8_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_8_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_8_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_8_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_8_i_1_inst_accumulation_buffer_rsc_0_8_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_8_i_q_d_mxwt(accumulation_buffer_rsc_0_8_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_8_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_8_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_8_i_we_d_pff(accumulation_buffer_rsc_0_8_i_we_d_iff),
      .accumulation_buffer_rsc_0_8_i_re_d_pff(accumulation_buffer_rsc_0_8_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_9_i_radr_d(accumulation_buffer_rsc_0_9_i_radr_d_reg),
      .accumulation_buffer_rsc_0_9_i_wadr_d(accumulation_buffer_rsc_0_9_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_9_i_q_d(accumulation_buffer_rsc_0_9_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_9_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_9_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_9_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_9_i_1_inst_accumulation_buffer_rsc_0_9_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_9_i_q_d_mxwt(accumulation_buffer_rsc_0_9_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_9_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_9_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_9_i_we_d_pff(accumulation_buffer_rsc_0_9_i_we_d_iff),
      .accumulation_buffer_rsc_0_9_i_re_d_pff(accumulation_buffer_rsc_0_9_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_10_i_radr_d(accumulation_buffer_rsc_0_10_i_radr_d_reg),
      .accumulation_buffer_rsc_0_10_i_wadr_d(accumulation_buffer_rsc_0_10_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_10_i_q_d(accumulation_buffer_rsc_0_10_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_10_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_10_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_10_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_10_i_1_inst_accumulation_buffer_rsc_0_10_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_10_i_q_d_mxwt(accumulation_buffer_rsc_0_10_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_10_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_10_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_10_i_we_d_pff(accumulation_buffer_rsc_0_10_i_we_d_iff),
      .accumulation_buffer_rsc_0_10_i_re_d_pff(accumulation_buffer_rsc_0_10_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_11_i_radr_d(accumulation_buffer_rsc_0_11_i_radr_d_reg),
      .accumulation_buffer_rsc_0_11_i_wadr_d(accumulation_buffer_rsc_0_11_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_11_i_q_d(accumulation_buffer_rsc_0_11_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_11_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_11_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_11_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_11_i_1_inst_accumulation_buffer_rsc_0_11_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_11_i_q_d_mxwt(accumulation_buffer_rsc_0_11_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_11_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_11_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_11_i_we_d_pff(accumulation_buffer_rsc_0_11_i_we_d_iff),
      .accumulation_buffer_rsc_0_11_i_re_d_pff(accumulation_buffer_rsc_0_11_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_12_i_radr_d(accumulation_buffer_rsc_0_12_i_radr_d_reg),
      .accumulation_buffer_rsc_0_12_i_wadr_d(accumulation_buffer_rsc_0_12_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_12_i_q_d(accumulation_buffer_rsc_0_12_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_12_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_12_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_12_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_12_i_1_inst_accumulation_buffer_rsc_0_12_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_12_i_q_d_mxwt(accumulation_buffer_rsc_0_12_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_12_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_12_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_12_i_we_d_pff(accumulation_buffer_rsc_0_12_i_we_d_iff),
      .accumulation_buffer_rsc_0_12_i_re_d_pff(accumulation_buffer_rsc_0_12_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_13_i_radr_d(accumulation_buffer_rsc_0_13_i_radr_d_reg),
      .accumulation_buffer_rsc_0_13_i_wadr_d(accumulation_buffer_rsc_0_13_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_13_i_q_d(accumulation_buffer_rsc_0_13_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_13_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_13_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_13_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_13_i_1_inst_accumulation_buffer_rsc_0_13_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_13_i_q_d_mxwt(accumulation_buffer_rsc_0_13_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_13_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_13_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_13_i_we_d_pff(accumulation_buffer_rsc_0_13_i_we_d_iff),
      .accumulation_buffer_rsc_0_13_i_re_d_pff(accumulation_buffer_rsc_0_13_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_14_i_radr_d(accumulation_buffer_rsc_0_14_i_radr_d_reg),
      .accumulation_buffer_rsc_0_14_i_wadr_d(accumulation_buffer_rsc_0_14_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_14_i_q_d(accumulation_buffer_rsc_0_14_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_14_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_14_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_14_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_14_i_1_inst_accumulation_buffer_rsc_0_14_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_14_i_q_d_mxwt(accumulation_buffer_rsc_0_14_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_14_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_14_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_14_i_we_d_pff(accumulation_buffer_rsc_0_14_i_we_d_iff),
      .accumulation_buffer_rsc_0_14_i_re_d_pff(accumulation_buffer_rsc_0_14_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1
      SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulation_buffer_rsc_0_15_i_radr_d(accumulation_buffer_rsc_0_15_i_radr_d_reg),
      .accumulation_buffer_rsc_0_15_i_wadr_d(accumulation_buffer_rsc_0_15_i_wadr_d_reg),
      .accumulation_buffer_rsc_0_15_i_q_d(accumulation_buffer_rsc_0_15_i_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .accumulation_buffer_rsc_0_15_i_oswt(reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .accumulation_buffer_rsc_0_15_i_radr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_radr_d_run[7:0]),
      .accumulation_buffer_rsc_0_15_i_wadr_d_run(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_accumulation_buffer_rsc_0_15_i_1_inst_accumulation_buffer_rsc_0_15_i_wadr_d_run[7:0]),
      .accumulation_buffer_rsc_0_15_i_q_d_mxwt(accumulation_buffer_rsc_0_15_i_q_d_mxwt),
      .accumulation_buffer_rsc_0_15_i_oswt_pff(and_1019_rmff),
      .accumulation_buffer_rsc_0_15_i_iswt0_1_pff(and_12_rmff),
      .accumulation_buffer_rsc_0_15_i_we_d_pff(accumulation_buffer_rsc_0_15_i_we_d_iff),
      .accumulation_buffer_rsc_0_15_i_re_d_pff(accumulation_buffer_rsc_0_15_i_re_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_wait_dp_inst
      (
      .ensig_cgo_iro(and_23_rmff),
      .ensig_cgo_iro_1(and_27_rmff),
      .run_wen(run_wen),
      .ensig_cgo(reg_ensig_cgo_303_cse),
      .accum_fifo_15_rsci_ccs_ccore_en(accum_fifo_15_rsci_ccs_ccore_en),
      .ensig_cgo_1(reg_ensig_cgo_302_cse),
      .output_fifo_0_rsci_ccs_ccore_en(output_fifo_0_rsci_ccs_ccore_en)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .input_rsci_wen_comp(input_rsci_wen_comp),
      .weight_rsci_wen_comp(weight_rsci_wen_comp),
      .output_rsci_wen_comp(output_rsci_wen_comp),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign output_and_cse = run_wen & (~((~ main_stage_0_4) | reg_step_not_mdf_sva_3_cse
      | operator_16_false_slc_operator_16_false_acc_16_itm_3 | (~ step_if_3_if_step_if_3_if_and_1_itm_3)));
  assign and_23_rmff = (and_dcpl_4 | and_dcpl_1) & (fsm_output[1]);
  assign and_27_rmff = (and_dcpl_10 | and_dcpl_1) & (fsm_output[1]);
  assign and_12_rmff = and_dcpl_10 & (~ operator_16_false_slc_operator_16_false_acc_16_itm_3);
  assign and_1019_rmff = and_dcpl_13 & (~ step_if_2_if_step_if_2_if_nor_1_tmp) &
      (fsm_output[1]);
  assign step_and_241_cse = run_wen & (~ (fsm_output[0]));
  assign psum_reg_and_cse = run_wen & ((~ main_stage_0_3) | step_not_mdf_sva_st_2);
  assign step_if_3_if_and_cse = run_wen & and_dcpl_1 & (~ operator_16_false_slc_operator_16_false_acc_16_itm_2);
  assign step_and_499_cse = run_wen & and_dcpl_4;
  assign and_1562_cse = run_wen & operator_32_false_acc_itm_31;
  assign or_1168_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b1000)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_290_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_62));
  assign mux_11_nl = MUX_s_1_2_2((or_1168_nl), (nor_290_nl), step_and_128_psp);
  assign weight_reg_and_cse = run_wen & (or_dcpl_8 | or_dcpl_4 | (step_step_lpi_1[0]))
      & (~((mux_11_nl) | or_dcpl_74));
  assign mux_12_nl = MUX_s_1_2_2(not_tmp_36, or_tmp_3, step_and_psp);
  assign weight_reg_and_1_cse = run_wen & or_dcpl_13 & (~((~ (mux_12_nl)) | or_dcpl_74));
  assign step_if_for_and_20_cse = step_and_241_cse & or_dcpl_7 & (~((~(main_stage_0_2
      & operator_16_false_slc_operator_16_false_acc_12_svs_st_1)) | step_not_mdf_sva_st_1));
  assign or_1167_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b1001)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_289_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_61));
  assign mux_42_nl = MUX_s_1_2_2((or_1167_nl), (nor_289_nl), step_and_144_psp);
  assign weight_reg_and_32_cse = run_wen & (or_dcpl_8 | or_dcpl_14) & (~((mux_42_nl)
      | or_dcpl_74));
  assign or_1166_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b0001)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_288_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_71));
  assign mux_43_nl = MUX_s_1_2_2((or_1166_nl), (nor_288_nl), step_and_16_psp);
  assign weight_reg_and_33_cse = run_wen & (or_dcpl_17 | or_dcpl_14) & (~((mux_43_nl)
      | or_dcpl_74));
  assign or_1165_nl = step_not_mdf_sva_st_1 | (~ (step_step_lpi_1_dfm_1_3_0[3]))
      | (step_step_lpi_1_dfm_1_3_0[2]) | (step_step_lpi_1_dfm_1_3_0[0]) | or_dcpl_48;
  assign nor_287_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_60));
  assign mux_74_nl = MUX_s_1_2_2((or_1165_nl), (nor_287_nl), step_and_160_psp);
  assign weight_reg_and_64_cse = run_wen & (or_dcpl_8 | or_dcpl_20) & (~((mux_74_nl)
      | or_dcpl_74));
  assign or_1164_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0[3]) | (step_step_lpi_1_dfm_1_3_0[2])
      | (step_step_lpi_1_dfm_1_3_0[0]) | or_dcpl_48;
  assign nor_286_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_70));
  assign mux_75_nl = MUX_s_1_2_2((or_1164_nl), (nor_286_nl), step_and_32_psp);
  assign weight_reg_and_65_cse = run_wen & (or_dcpl_17 | or_dcpl_20) & (~((mux_75_nl)
      | or_dcpl_74));
  assign or_1163_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0[3:2]!=2'b10)
      | or_dcpl_49;
  assign nor_285_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_59));
  assign mux_106_nl = MUX_s_1_2_2((or_1163_nl), (nor_285_nl), step_and_176_psp);
  assign weight_reg_and_96_cse = run_wen & (or_dcpl_8 | or_dcpl_23) & (~((mux_106_nl)
      | or_dcpl_74));
  assign or_1162_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0[3:2]!=2'b00)
      | or_dcpl_49;
  assign nor_284_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_69));
  assign mux_107_nl = MUX_s_1_2_2((or_1162_nl), (nor_284_nl), step_and_48_psp);
  assign weight_reg_and_97_cse = run_wen & (or_dcpl_17 | or_dcpl_23) & (~((mux_107_nl)
      | or_dcpl_74));
  assign or_1161_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b1100)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_283_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_57));
  assign mux_138_nl = MUX_s_1_2_2((or_1161_nl), (nor_283_nl), step_and_192_psp);
  assign weight_reg_and_128_cse = run_wen & (or_dcpl_8 | or_dcpl_27) & (~((mux_138_nl)
      | or_dcpl_74));
  assign or_1160_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b0100)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_282_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_67));
  assign mux_139_nl = MUX_s_1_2_2((or_1160_nl), (nor_282_nl), step_and_64_psp);
  assign weight_reg_and_129_cse = run_wen & (or_dcpl_17 | or_dcpl_27) & (~((mux_139_nl)
      | or_dcpl_74));
  assign or_1159_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b1101)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_281_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_55));
  assign mux_170_nl = MUX_s_1_2_2((or_1159_nl), (nor_281_nl), step_and_208_psp);
  assign weight_reg_and_160_cse = run_wen & (or_dcpl_8 | or_dcpl_30) & (~((mux_170_nl)
      | or_dcpl_74));
  assign or_1158_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b0101)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign nor_280_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_66));
  assign mux_171_nl = MUX_s_1_2_2((or_1158_nl), (nor_280_nl), step_and_80_psp);
  assign weight_reg_and_161_cse = run_wen & (or_dcpl_17 | or_dcpl_30) & (~((mux_171_nl)
      | or_dcpl_74));
  assign or_1157_nl = step_not_mdf_sva_st_1 | (~ (step_step_lpi_1_dfm_1_3_0[3]))
      | (~ (step_step_lpi_1_dfm_1_3_0[2])) | (step_step_lpi_1_dfm_1_3_0[0]) | or_dcpl_48;
  assign nor_279_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_52));
  assign mux_202_nl = MUX_s_1_2_2((or_1157_nl), (nor_279_nl), step_and_224_psp);
  assign weight_reg_and_192_cse = run_wen & (or_dcpl_8 | or_dcpl_34) & (~((mux_202_nl)
      | or_dcpl_74));
  assign mux_203_nl = MUX_s_1_2_2(not_tmp_251, or_tmp_39, step_and_96_psp);
  assign weight_reg_and_193_cse = run_wen & or_dcpl_36 & (~((~ (mux_203_nl)) | or_dcpl_74));
  assign or_1156_nl = step_not_mdf_sva_st_1 | or_dcpl_50;
  assign nor_278_nl = ~(step_not_mdf_sva_st_1 | ((step_step_lpi_1_dfm_1_3_0==4'b1111)
      & operator_16_false_slc_operator_16_false_acc_12_svs_st_1));
  assign mux_234_nl = MUX_s_1_2_2((or_1156_nl), (nor_278_nl), step_and_240_psp);
  assign weight_reg_and_224_cse = run_wen & (or_dcpl_8 | or_dcpl_37) & (~((mux_234_nl)
      | or_dcpl_74));
  assign or_1155_nl = step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0[3]) | (~((step_step_lpi_1_dfm_1_3_0[2:0]==3'b111)
      & operator_16_false_slc_operator_16_false_acc_12_svs_st_1));
  assign nor_277_nl = ~(step_not_mdf_sva_st_1 | (~ or_dcpl_64));
  assign mux_235_nl = MUX_s_1_2_2((or_1155_nl), (nor_277_nl), step_and_112_psp);
  assign weight_reg_and_225_cse = run_wen & (or_dcpl_17 | or_dcpl_37) & (~((mux_235_nl)
      | or_dcpl_74));
  assign step_if_3_if_and_1_cse = run_wen & and_dcpl_4 & (~ operator_16_false_slc_operator_16_false_acc_16_itm_1);
  assign step_and_757_cse = step_and_241_cse & (~ operator_32_false_acc_itm_31) &
      (~ or_dcpl_74);
  assign nl_operator_32_false_acc_1_nl = conv_u2u_32_33(~ step_mul_itm) + conv_u2u_16_33(step_step_lpi_1_dfm_1);
  assign operator_32_false_acc_1_nl = nl_operator_32_false_acc_1_nl[32:0];
  assign nl_operator_32_false_acc_nl = (readslicef_33_32_1((operator_32_false_acc_1_nl)))
      + 32'b01111111111111111111111111110001;
  assign operator_32_false_acc_nl = nl_operator_32_false_acc_nl[31:0];
  assign operator_32_false_acc_itm_31 = readslicef_32_1_31((operator_32_false_acc_nl));
  assign nl_operator_16_false_acc_nl = conv_u2u_12_13(step_step_lpi_1_dfm_1[15:4])
      + 13'b1111111111111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[12:0];
  assign operator_16_false_acc_itm_12_1 = readslicef_13_1_12((operator_16_false_acc_nl));
  assign loopIndicesIn_crt_lpi_1_dfm_mx0 = MUX_v_48_2_2(loopIndicesIn_crt_lpi_1_dfm,
      loopIndicesIn_rsci_idat_mxwt, exitL_exit_step_sva);
  assign paramsIn_crt_lpi_1_dfm_127_80_mx0 = MUX_v_48_2_2(paramsIn_crt_lpi_1_dfm_127_80,
      (paramsIn_rsci_idat_mxwt[79:32]), exitL_exit_step_sva);
  assign paramsIn_crt_lpi_1_dfm_63_32_mx0 = MUX_v_32_2_2(paramsIn_crt_lpi_1_dfm_63_32,
      (paramsIn_rsci_idat_mxwt[31:0]), exitL_exit_step_sva);
  assign step_if_for_and_stg_2_0_sva_mx1w0 = step_if_for_and_stg_1_0_sva_1 & (~ (step_step_lpi_1_dfm_1_3_0[2]));
  assign step_if_for_and_stg_2_0_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_0_sva,
      step_if_for_and_stg_2_0_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_1_sva_mx1w0 = step_if_for_and_stg_1_1_sva_1 & (~ (step_step_lpi_1_dfm_1_3_0[2]));
  assign step_if_for_and_stg_2_1_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_1_sva,
      step_if_for_and_stg_2_1_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_2_sva_mx1w0 = step_if_for_and_stg_1_2_sva_1 & (~ (step_step_lpi_1_dfm_1_3_0[2]));
  assign step_if_for_and_stg_2_2_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_2_sva,
      step_if_for_and_stg_2_2_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_3_sva_mx1w0 = step_if_for_and_stg_1_3_sva_1 & (~ (step_step_lpi_1_dfm_1_3_0[2]));
  assign step_if_for_and_stg_2_3_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_3_sva,
      step_if_for_and_stg_2_3_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_4_sva_mx1w0 = step_if_for_and_stg_1_0_sva_1 & (step_step_lpi_1_dfm_1_3_0[2]);
  assign step_if_for_and_stg_2_4_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_4_sva,
      step_if_for_and_stg_2_4_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_5_sva_mx1w0 = step_if_for_and_stg_1_1_sva_1 & (step_step_lpi_1_dfm_1_3_0[2]);
  assign step_if_for_and_stg_2_5_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_5_sva,
      step_if_for_and_stg_2_5_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_6_sva_mx1w0 = step_if_for_and_stg_1_2_sva_1 & (step_step_lpi_1_dfm_1_3_0[2]);
  assign step_if_for_and_stg_2_6_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_6_sva,
      step_if_for_and_stg_2_6_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_if_for_and_stg_2_7_sva_mx1w0 = step_if_for_and_stg_1_3_sva_1 & (step_step_lpi_1_dfm_1_3_0[2]);
  assign step_if_for_and_stg_2_7_sva_mx1 = MUX_s_1_2_2(step_if_for_and_stg_2_7_sva,
      step_if_for_and_stg_2_7_sva_mx1w0, operator_16_false_slc_operator_16_false_acc_12_svs_st_1);
  assign step_and_96_psp_1 = step_if_for_and_stg_2_6_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
      & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
  assign step_and_psp_1 = step_if_for_and_stg_2_0_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
      & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
  assign step_if_2_if_step_if_2_if_nor_1_tmp = ~((loopIndicesIn_crt_lpi_1_dfm_mx0!=48'b000000000000000000000000000000000000000000000000));
  assign nl_step_if_1_acc_nl = ({17'b10000000000000000 , step_step_lpi_1_dfm_1})
      + conv_u2u_32_33(~ step_mul_itm) + 33'b000000000000000000000000000000001;
  assign step_if_1_acc_nl = nl_step_if_1_acc_nl[32:0];
  assign step_if_1_acc_itm_32_1 = readslicef_33_1_32((step_if_1_acc_nl));
  assign nl_operator_16_false_acc_nl_1 = conv_u2s_16_17(step_step_lpi_1_dfm_1) +
      17'b11111111111100001;
  assign operator_16_false_acc_nl_1 = nl_operator_16_false_acc_nl_1[16:0];
  assign operator_16_false_acc_itm_16_1 = readslicef_17_1_16((operator_16_false_acc_nl_1));
  assign step_in_col_value_lpi_1_dfm_mx0 = MUX_v_128_2_2(step_in_col_value_lpi_1,
      input_rsci_idat_mxwt, step_if_1_acc_cse_32);
  assign step_not_12_nl = ~ exitL_exit_step_sva;
  assign step_step_lpi_1_dfm_1 = MUX_v_16_2_2(16'b0000000000000000, step_step_lpi_1,
      (step_not_12_nl));
  assign nl_operator_16_false_2_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_lpi_1_dfm_127_80_mx0[31:16])
      + 17'b11111111111111111;
  assign operator_16_false_2_acc_psp_sva_1 = nl_operator_16_false_2_acc_psp_sva_1[16:0];
  assign nl_operator_16_false_1_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_lpi_1_dfm_127_80_mx0[15:0])
      + 17'b11111111111111111;
  assign operator_16_false_1_acc_psp_sva_1 = nl_operator_16_false_1_acc_psp_sva_1[16:0];
  assign step_if_for_and_stg_1_0_sva_1 = ~((step_step_lpi_1_dfm_1_3_0[1:0]!=2'b00));
  assign step_if_for_and_stg_1_1_sva_1 = (step_step_lpi_1_dfm_1_3_0[1:0]==2'b01);
  assign step_if_for_and_stg_1_2_sva_1 = (step_step_lpi_1_dfm_1_3_0[1:0]==2'b10);
  assign step_if_for_and_stg_1_3_sva_1 = (step_step_lpi_1_dfm_1_3_0[1:0]==2'b11);
  assign nl_operator_16_false_3_acc_psp_sva_1 = conv_u2s_16_17(paramsIn_crt_lpi_1_dfm_127_80_mx0[47:32])
      + 17'b11111111111111111;
  assign operator_16_false_3_acc_psp_sva_1 = nl_operator_16_false_3_acc_psp_sva_1[16:0];
  assign step_mul_itm = conv_u2u_32_32((paramsIn_crt_lpi_1_dfm_63_32_mx0[31:16])
      * (paramsIn_crt_lpi_1_dfm_63_32_mx0[15:0]));
  assign and_dcpl_1 = main_stage_0_3 & (~ step_not_mdf_sva_st_2);
  assign and_dcpl_4 = main_stage_0_2 & (~ step_not_mdf_sva_st_1);
  assign or_dcpl_4 = (step_step_lpi_1[2:1]!=2'b00);
  assign or_dcpl_7 = ~(operator_32_false_acc_itm_31 & operator_16_false_acc_itm_12_1);
  assign or_dcpl_8 = or_dcpl_7 | exitL_exit_step_sva | (~ (step_step_lpi_1[3]));
  assign or_dcpl_13 = (~((~((step_step_lpi_1[3:0]!=4'b0000))) | exitL_exit_step_sva))
      | or_dcpl_7;
  assign or_dcpl_14 = or_dcpl_4 | (~ (step_step_lpi_1[0]));
  assign or_dcpl_17 = or_dcpl_7 | exitL_exit_step_sva | (step_step_lpi_1[3]);
  assign or_dcpl_19 = (step_step_lpi_1[2:1]!=2'b01);
  assign or_dcpl_20 = or_dcpl_19 | (step_step_lpi_1[0]);
  assign or_dcpl_23 = or_dcpl_19 | (~ (step_step_lpi_1[0]));
  assign or_dcpl_26 = (step_step_lpi_1[2:1]!=2'b10);
  assign or_dcpl_27 = or_dcpl_26 | (step_step_lpi_1[0]);
  assign or_dcpl_30 = or_dcpl_26 | (~ (step_step_lpi_1[0]));
  assign or_dcpl_33 = ~((step_step_lpi_1[2:1]==2'b11));
  assign or_dcpl_34 = or_dcpl_33 | (step_step_lpi_1[0]);
  assign or_dcpl_36 = or_dcpl_17 | or_dcpl_34;
  assign or_dcpl_37 = or_dcpl_33 | (~ (step_step_lpi_1[0]));
  assign and_dcpl_10 = main_stage_0_4 & (~ reg_step_not_mdf_sva_3_cse);
  assign and_dcpl_13 = operator_32_false_acc_itm_31 & step_if_1_acc_itm_32_1;
  assign or_dcpl_47 = ~((step_step_lpi_1_dfm_1_3_0[3:2]==2'b11));
  assign or_dcpl_48 = ~(operator_16_false_slc_operator_16_false_acc_12_svs_st_1 &
      (step_step_lpi_1_dfm_1_3_0[1]));
  assign or_dcpl_49 = or_dcpl_48 | (~ (step_step_lpi_1_dfm_1_3_0[0]));
  assign or_dcpl_50 = or_dcpl_49 | or_dcpl_47;
  assign or_dcpl_51 = or_dcpl_48 | (step_step_lpi_1_dfm_1_3_0[0]);
  assign or_dcpl_52 = or_dcpl_51 | or_dcpl_47;
  assign or_dcpl_53 = (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1)
      | (step_step_lpi_1_dfm_1_3_0[1]);
  assign or_dcpl_54 = or_dcpl_53 | (~ (step_step_lpi_1_dfm_1_3_0[0]));
  assign or_dcpl_55 = or_dcpl_54 | or_dcpl_47;
  assign or_dcpl_56 = or_dcpl_53 | (step_step_lpi_1_dfm_1_3_0[0]);
  assign or_dcpl_57 = or_dcpl_56 | or_dcpl_47;
  assign or_dcpl_58 = (step_step_lpi_1_dfm_1_3_0[3:2]!=2'b10);
  assign or_dcpl_59 = or_dcpl_49 | or_dcpl_58;
  assign or_dcpl_60 = or_dcpl_51 | or_dcpl_58;
  assign or_dcpl_61 = or_dcpl_54 | or_dcpl_58;
  assign or_dcpl_62 = or_dcpl_56 | or_dcpl_58;
  assign or_dcpl_63 = (step_step_lpi_1_dfm_1_3_0[3:2]!=2'b01);
  assign or_dcpl_64 = or_dcpl_49 | or_dcpl_63;
  assign or_dcpl_65 = or_dcpl_51 | or_dcpl_63;
  assign or_dcpl_66 = or_dcpl_54 | or_dcpl_63;
  assign or_dcpl_67 = or_dcpl_56 | or_dcpl_63;
  assign or_dcpl_68 = (step_step_lpi_1_dfm_1_3_0[3:2]!=2'b00);
  assign or_dcpl_69 = or_dcpl_49 | or_dcpl_68;
  assign or_dcpl_70 = or_dcpl_51 | or_dcpl_68;
  assign or_dcpl_71 = or_dcpl_54 | or_dcpl_68;
  assign or_dcpl_72 = or_dcpl_56 | or_dcpl_68;
  assign and_dcpl_18 = and_dcpl_4 & (~ operator_32_false_acc_itm_31);
  assign or_dcpl_74 = (~ main_stage_0_2) | step_not_mdf_sva_st_1;
  assign or_tmp_3 = step_not_mdf_sva_st_1 | (~ or_dcpl_72);
  assign not_tmp_36 = ~(step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0!=4'b0000)
      | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1));
  assign or_tmp_39 = step_not_mdf_sva_st_1 | (~ or_dcpl_65);
  assign not_tmp_251 = ~(step_not_mdf_sva_st_1 | (step_step_lpi_1_dfm_1_3_0[3]) |
      (~ (step_step_lpi_1_dfm_1_3_0[2])) | (step_step_lpi_1_dfm_1_3_0[0]) | or_dcpl_48);
  assign or_tmp_47 = operator_32_false_acc_itm_31 & (fsm_output[1]);
  assign accumulation_buffer_rsc_0_0_i_radr_d = accumulation_buffer_rsc_0_0_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_wadr_d = accumulation_buffer_rsc_0_0_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_0_i_d_d = output_fifo_0_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_0_i_we_d_pff = accumulation_buffer_rsc_0_0_i_we_d_iff;
  assign accumulation_buffer_rsc_0_0_i_re_d_pff = accumulation_buffer_rsc_0_0_i_re_d_iff;
  assign accumulation_buffer_rsc_0_1_i_radr_d = accumulation_buffer_rsc_0_1_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_wadr_d = accumulation_buffer_rsc_0_1_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_1_i_d_d = output_fifo_1_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_1_i_we_d_pff = accumulation_buffer_rsc_0_1_i_we_d_iff;
  assign accumulation_buffer_rsc_0_1_i_re_d_pff = accumulation_buffer_rsc_0_1_i_re_d_iff;
  assign accumulation_buffer_rsc_0_2_i_radr_d = accumulation_buffer_rsc_0_2_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_wadr_d = accumulation_buffer_rsc_0_2_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_2_i_d_d = output_fifo_2_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_2_i_we_d_pff = accumulation_buffer_rsc_0_2_i_we_d_iff;
  assign accumulation_buffer_rsc_0_2_i_re_d_pff = accumulation_buffer_rsc_0_2_i_re_d_iff;
  assign accumulation_buffer_rsc_0_3_i_radr_d = accumulation_buffer_rsc_0_3_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_wadr_d = accumulation_buffer_rsc_0_3_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_3_i_d_d = output_fifo_3_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_3_i_we_d_pff = accumulation_buffer_rsc_0_3_i_we_d_iff;
  assign accumulation_buffer_rsc_0_3_i_re_d_pff = accumulation_buffer_rsc_0_3_i_re_d_iff;
  assign accumulation_buffer_rsc_0_4_i_radr_d = accumulation_buffer_rsc_0_4_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_wadr_d = accumulation_buffer_rsc_0_4_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_4_i_d_d = output_fifo_4_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_4_i_we_d_pff = accumulation_buffer_rsc_0_4_i_we_d_iff;
  assign accumulation_buffer_rsc_0_4_i_re_d_pff = accumulation_buffer_rsc_0_4_i_re_d_iff;
  assign accumulation_buffer_rsc_0_5_i_radr_d = accumulation_buffer_rsc_0_5_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_wadr_d = accumulation_buffer_rsc_0_5_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_5_i_d_d = output_fifo_5_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_5_i_we_d_pff = accumulation_buffer_rsc_0_5_i_we_d_iff;
  assign accumulation_buffer_rsc_0_5_i_re_d_pff = accumulation_buffer_rsc_0_5_i_re_d_iff;
  assign accumulation_buffer_rsc_0_6_i_radr_d = accumulation_buffer_rsc_0_6_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_wadr_d = accumulation_buffer_rsc_0_6_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_6_i_d_d = output_fifo_6_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_6_i_we_d_pff = accumulation_buffer_rsc_0_6_i_we_d_iff;
  assign accumulation_buffer_rsc_0_6_i_re_d_pff = accumulation_buffer_rsc_0_6_i_re_d_iff;
  assign accumulation_buffer_rsc_0_7_i_radr_d = accumulation_buffer_rsc_0_7_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_wadr_d = accumulation_buffer_rsc_0_7_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_7_i_d_d = output_fifo_7_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_7_i_we_d_pff = accumulation_buffer_rsc_0_7_i_we_d_iff;
  assign accumulation_buffer_rsc_0_7_i_re_d_pff = accumulation_buffer_rsc_0_7_i_re_d_iff;
  assign accumulation_buffer_rsc_0_8_i_radr_d = accumulation_buffer_rsc_0_8_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_wadr_d = accumulation_buffer_rsc_0_8_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_8_i_d_d = output_fifo_8_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_8_i_we_d_pff = accumulation_buffer_rsc_0_8_i_we_d_iff;
  assign accumulation_buffer_rsc_0_8_i_re_d_pff = accumulation_buffer_rsc_0_8_i_re_d_iff;
  assign accumulation_buffer_rsc_0_9_i_radr_d = accumulation_buffer_rsc_0_9_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_wadr_d = accumulation_buffer_rsc_0_9_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_9_i_d_d = output_fifo_9_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_9_i_we_d_pff = accumulation_buffer_rsc_0_9_i_we_d_iff;
  assign accumulation_buffer_rsc_0_9_i_re_d_pff = accumulation_buffer_rsc_0_9_i_re_d_iff;
  assign accumulation_buffer_rsc_0_10_i_radr_d = accumulation_buffer_rsc_0_10_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_wadr_d = accumulation_buffer_rsc_0_10_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_10_i_d_d = output_fifo_10_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_10_i_we_d_pff = accumulation_buffer_rsc_0_10_i_we_d_iff;
  assign accumulation_buffer_rsc_0_10_i_re_d_pff = accumulation_buffer_rsc_0_10_i_re_d_iff;
  assign accumulation_buffer_rsc_0_11_i_radr_d = accumulation_buffer_rsc_0_11_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_wadr_d = accumulation_buffer_rsc_0_11_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_11_i_d_d = output_fifo_11_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_11_i_we_d_pff = accumulation_buffer_rsc_0_11_i_we_d_iff;
  assign accumulation_buffer_rsc_0_11_i_re_d_pff = accumulation_buffer_rsc_0_11_i_re_d_iff;
  assign accumulation_buffer_rsc_0_12_i_radr_d = accumulation_buffer_rsc_0_12_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_wadr_d = accumulation_buffer_rsc_0_12_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_12_i_d_d = output_fifo_12_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_12_i_we_d_pff = accumulation_buffer_rsc_0_12_i_we_d_iff;
  assign accumulation_buffer_rsc_0_12_i_re_d_pff = accumulation_buffer_rsc_0_12_i_re_d_iff;
  assign accumulation_buffer_rsc_0_13_i_radr_d = accumulation_buffer_rsc_0_13_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_wadr_d = accumulation_buffer_rsc_0_13_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_13_i_d_d = output_fifo_13_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_13_i_we_d_pff = accumulation_buffer_rsc_0_13_i_we_d_iff;
  assign accumulation_buffer_rsc_0_13_i_re_d_pff = accumulation_buffer_rsc_0_13_i_re_d_iff;
  assign accumulation_buffer_rsc_0_14_i_radr_d = accumulation_buffer_rsc_0_14_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_wadr_d = accumulation_buffer_rsc_0_14_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_14_i_d_d = output_fifo_14_rsci_output_rsc_z;
  assign accumulation_buffer_rsc_0_14_i_we_d_pff = accumulation_buffer_rsc_0_14_i_we_d_iff;
  assign accumulation_buffer_rsc_0_14_i_re_d_pff = accumulation_buffer_rsc_0_14_i_re_d_iff;
  assign accumulation_buffer_rsc_0_15_i_radr_d = accumulation_buffer_rsc_0_15_i_radr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_wadr_d = accumulation_buffer_rsc_0_15_i_wadr_d_reg;
  assign accumulation_buffer_rsc_0_15_i_d_d = accum_fifo_0_run_cmp_1_output_rsc_z;
  assign accumulation_buffer_rsc_0_15_i_we_d_pff = accumulation_buffer_rsc_0_15_i_we_d_iff;
  assign accumulation_buffer_rsc_0_15_i_re_d_pff = accumulation_buffer_rsc_0_15_i_re_d_iff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_loopIndicesIn_rsci_oswt_cse <= 1'b0;
      reg_ensig_cgo_303_cse <= 1'b0;
      reg_ensig_cgo_302_cse <= 1'b0;
      reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse
          <= 1'b0;
      reg_output_rsci_ivld_run_psct_cse <= 1'b0;
      reg_weight_rsci_irdy_run_psct_cse <= 1'b0;
      reg_input_rsci_irdy_run_psct_cse <= 1'b0;
      step_not_mdf_sva_st_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_loopIndicesIn_rsci_oswt_cse <= ~ or_tmp_47;
      reg_ensig_cgo_303_cse <= and_23_rmff;
      reg_ensig_cgo_302_cse <= and_27_rmff;
      reg_accumulation_buffer_rsc_0_15_i_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse
          <= and_1019_rmff;
      reg_output_rsci_ivld_run_psct_cse <= and_dcpl_10 & (~ operator_16_false_slc_operator_16_false_acc_16_itm_3)
          & step_if_3_if_step_if_3_if_and_1_itm_3;
      reg_weight_rsci_irdy_run_psct_cse <= operator_32_false_acc_itm_31 & operator_16_false_acc_itm_12_1
          & (fsm_output[1]);
      reg_input_rsci_irdy_run_psct_cse <= and_dcpl_13 & (fsm_output[1]);
      step_not_mdf_sva_st_1 <= ~ operator_32_false_acc_itm_31;
      main_stage_0_2 <= fsm_output[1];
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_rsci_idat_15_0 <= 16'b0000000000000000;
      output_rsci_idat_31_16 <= 16'b0000000000000000;
      output_rsci_idat_47_32 <= 16'b0000000000000000;
      output_rsci_idat_63_48 <= 16'b0000000000000000;
      output_rsci_idat_79_64 <= 16'b0000000000000000;
      output_rsci_idat_95_80 <= 16'b0000000000000000;
      output_rsci_idat_111_96 <= 16'b0000000000000000;
      output_rsci_idat_127_112 <= 16'b0000000000000000;
      output_rsci_idat_143_128 <= 16'b0000000000000000;
      output_rsci_idat_159_144 <= 16'b0000000000000000;
      output_rsci_idat_175_160 <= 16'b0000000000000000;
      output_rsci_idat_191_176 <= 16'b0000000000000000;
      output_rsci_idat_207_192 <= 16'b0000000000000000;
      output_rsci_idat_223_208 <= 16'b0000000000000000;
      output_rsci_idat_239_224 <= 16'b0000000000000000;
      output_rsci_idat_255_240 <= 16'b0000000000000000;
    end
    else if ( output_and_cse ) begin
      output_rsci_idat_15_0 <= output_fifo_0_rsci_output_rsc_z;
      output_rsci_idat_31_16 <= output_fifo_1_rsci_output_rsc_z;
      output_rsci_idat_47_32 <= output_fifo_2_rsci_output_rsc_z;
      output_rsci_idat_63_48 <= output_fifo_3_rsci_output_rsc_z;
      output_rsci_idat_79_64 <= output_fifo_4_rsci_output_rsc_z;
      output_rsci_idat_95_80 <= output_fifo_5_rsci_output_rsc_z;
      output_rsci_idat_111_96 <= output_fifo_6_rsci_output_rsc_z;
      output_rsci_idat_127_112 <= output_fifo_7_rsci_output_rsc_z;
      output_rsci_idat_143_128 <= output_fifo_8_rsci_output_rsc_z;
      output_rsci_idat_159_144 <= output_fifo_9_rsci_output_rsc_z;
      output_rsci_idat_175_160 <= output_fifo_10_rsci_output_rsc_z;
      output_rsci_idat_191_176 <= output_fifo_11_rsci_output_rsc_z;
      output_rsci_idat_207_192 <= output_fifo_12_rsci_output_rsc_z;
      output_rsci_idat_223_208 <= output_fifo_13_rsci_output_rsc_z;
      output_rsci_idat_239_224 <= output_fifo_14_rsci_output_rsc_z;
      output_rsci_idat_255_240 <= accum_fifo_0_run_cmp_1_output_rsc_z;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exit_step_sva <= 1'b1;
    end
    else if ( step_and_241_cse ) begin
      exitL_exit_step_sva <= ~ operator_32_false_acc_itm_31;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psum_reg_16_16_sva <= 16'b0000000000000000;
      psum_reg_16_15_sva <= 16'b0000000000000000;
      psum_reg_16_14_sva <= 16'b0000000000000000;
      psum_reg_16_13_sva <= 16'b0000000000000000;
      psum_reg_16_12_sva <= 16'b0000000000000000;
      psum_reg_16_11_sva <= 16'b0000000000000000;
      psum_reg_16_10_sva <= 16'b0000000000000000;
      psum_reg_16_9_sva <= 16'b0000000000000000;
      psum_reg_16_8_sva <= 16'b0000000000000000;
      psum_reg_16_7_sva <= 16'b0000000000000000;
      psum_reg_16_6_sva <= 16'b0000000000000000;
      psum_reg_16_5_sva <= 16'b0000000000000000;
      psum_reg_16_4_sva <= 16'b0000000000000000;
      psum_reg_16_3_sva <= 16'b0000000000000000;
      psum_reg_16_2_sva <= 16'b0000000000000000;
      psum_reg_16_1_sva <= 16'b0000000000000000;
      psum_reg_15_16_sva <= 16'b0000000000000000;
      psum_reg_15_15_sva <= 16'b0000000000000000;
      psum_reg_15_14_sva <= 16'b0000000000000000;
      psum_reg_15_13_sva <= 16'b0000000000000000;
      psum_reg_15_12_sva <= 16'b0000000000000000;
      psum_reg_15_11_sva <= 16'b0000000000000000;
      psum_reg_15_10_sva <= 16'b0000000000000000;
      psum_reg_15_9_sva <= 16'b0000000000000000;
      psum_reg_15_8_sva <= 16'b0000000000000000;
      psum_reg_15_7_sva <= 16'b0000000000000000;
      psum_reg_15_6_sva <= 16'b0000000000000000;
      psum_reg_15_5_sva <= 16'b0000000000000000;
      psum_reg_15_4_sva <= 16'b0000000000000000;
      psum_reg_15_3_sva <= 16'b0000000000000000;
      psum_reg_15_2_sva <= 16'b0000000000000000;
      psum_reg_15_1_sva <= 16'b0000000000000000;
      psum_reg_14_16_sva <= 16'b0000000000000000;
      psum_reg_14_15_sva <= 16'b0000000000000000;
      psum_reg_14_14_sva <= 16'b0000000000000000;
      psum_reg_14_13_sva <= 16'b0000000000000000;
      psum_reg_14_12_sva <= 16'b0000000000000000;
      psum_reg_14_11_sva <= 16'b0000000000000000;
      psum_reg_14_10_sva <= 16'b0000000000000000;
      psum_reg_14_9_sva <= 16'b0000000000000000;
      psum_reg_14_8_sva <= 16'b0000000000000000;
      psum_reg_14_7_sva <= 16'b0000000000000000;
      psum_reg_14_6_sva <= 16'b0000000000000000;
      psum_reg_14_5_sva <= 16'b0000000000000000;
      psum_reg_14_4_sva <= 16'b0000000000000000;
      psum_reg_14_3_sva <= 16'b0000000000000000;
      psum_reg_14_2_sva <= 16'b0000000000000000;
      psum_reg_14_1_sva <= 16'b0000000000000000;
      psum_reg_13_16_sva <= 16'b0000000000000000;
      psum_reg_13_15_sva <= 16'b0000000000000000;
      psum_reg_13_14_sva <= 16'b0000000000000000;
      psum_reg_13_13_sva <= 16'b0000000000000000;
      psum_reg_13_12_sva <= 16'b0000000000000000;
      psum_reg_13_11_sva <= 16'b0000000000000000;
      psum_reg_13_10_sva <= 16'b0000000000000000;
      psum_reg_13_9_sva <= 16'b0000000000000000;
      psum_reg_13_8_sva <= 16'b0000000000000000;
      psum_reg_13_7_sva <= 16'b0000000000000000;
      psum_reg_13_6_sva <= 16'b0000000000000000;
      psum_reg_13_5_sva <= 16'b0000000000000000;
      psum_reg_13_4_sva <= 16'b0000000000000000;
      psum_reg_13_3_sva <= 16'b0000000000000000;
      psum_reg_13_2_sva <= 16'b0000000000000000;
      psum_reg_13_1_sva <= 16'b0000000000000000;
      psum_reg_12_16_sva <= 16'b0000000000000000;
      psum_reg_12_15_sva <= 16'b0000000000000000;
      psum_reg_12_14_sva <= 16'b0000000000000000;
      psum_reg_12_13_sva <= 16'b0000000000000000;
      psum_reg_12_12_sva <= 16'b0000000000000000;
      psum_reg_12_11_sva <= 16'b0000000000000000;
      psum_reg_12_10_sva <= 16'b0000000000000000;
      psum_reg_12_9_sva <= 16'b0000000000000000;
      psum_reg_12_8_sva <= 16'b0000000000000000;
      psum_reg_12_7_sva <= 16'b0000000000000000;
      psum_reg_12_6_sva <= 16'b0000000000000000;
      psum_reg_12_5_sva <= 16'b0000000000000000;
      psum_reg_12_4_sva <= 16'b0000000000000000;
      psum_reg_12_3_sva <= 16'b0000000000000000;
      psum_reg_12_2_sva <= 16'b0000000000000000;
      psum_reg_12_1_sva <= 16'b0000000000000000;
      psum_reg_11_16_sva <= 16'b0000000000000000;
      psum_reg_11_15_sva <= 16'b0000000000000000;
      psum_reg_11_14_sva <= 16'b0000000000000000;
      psum_reg_11_13_sva <= 16'b0000000000000000;
      psum_reg_11_12_sva <= 16'b0000000000000000;
      psum_reg_11_11_sva <= 16'b0000000000000000;
      psum_reg_11_10_sva <= 16'b0000000000000000;
      psum_reg_11_9_sva <= 16'b0000000000000000;
      psum_reg_11_8_sva <= 16'b0000000000000000;
      psum_reg_11_7_sva <= 16'b0000000000000000;
      psum_reg_11_6_sva <= 16'b0000000000000000;
      psum_reg_11_5_sva <= 16'b0000000000000000;
      psum_reg_11_4_sva <= 16'b0000000000000000;
      psum_reg_11_3_sva <= 16'b0000000000000000;
      psum_reg_11_2_sva <= 16'b0000000000000000;
      psum_reg_11_1_sva <= 16'b0000000000000000;
      psum_reg_10_16_sva <= 16'b0000000000000000;
      psum_reg_10_15_sva <= 16'b0000000000000000;
      psum_reg_10_14_sva <= 16'b0000000000000000;
      psum_reg_10_13_sva <= 16'b0000000000000000;
      psum_reg_10_12_sva <= 16'b0000000000000000;
      psum_reg_10_11_sva <= 16'b0000000000000000;
      psum_reg_10_10_sva <= 16'b0000000000000000;
      psum_reg_10_9_sva <= 16'b0000000000000000;
      psum_reg_10_8_sva <= 16'b0000000000000000;
      psum_reg_10_7_sva <= 16'b0000000000000000;
      psum_reg_10_6_sva <= 16'b0000000000000000;
      psum_reg_10_5_sva <= 16'b0000000000000000;
      psum_reg_10_4_sva <= 16'b0000000000000000;
      psum_reg_10_3_sva <= 16'b0000000000000000;
      psum_reg_10_2_sva <= 16'b0000000000000000;
      psum_reg_10_1_sva <= 16'b0000000000000000;
      psum_reg_9_16_sva <= 16'b0000000000000000;
      psum_reg_9_15_sva <= 16'b0000000000000000;
      psum_reg_9_14_sva <= 16'b0000000000000000;
      psum_reg_9_13_sva <= 16'b0000000000000000;
      psum_reg_9_12_sva <= 16'b0000000000000000;
      psum_reg_9_11_sva <= 16'b0000000000000000;
      psum_reg_9_10_sva <= 16'b0000000000000000;
      psum_reg_9_9_sva <= 16'b0000000000000000;
      psum_reg_9_8_sva <= 16'b0000000000000000;
      psum_reg_9_7_sva <= 16'b0000000000000000;
      psum_reg_9_6_sva <= 16'b0000000000000000;
      psum_reg_9_5_sva <= 16'b0000000000000000;
      psum_reg_9_4_sva <= 16'b0000000000000000;
      psum_reg_9_3_sva <= 16'b0000000000000000;
      psum_reg_9_2_sva <= 16'b0000000000000000;
      psum_reg_9_1_sva <= 16'b0000000000000000;
      psum_reg_8_16_sva <= 16'b0000000000000000;
      psum_reg_8_15_sva <= 16'b0000000000000000;
      psum_reg_8_14_sva <= 16'b0000000000000000;
      psum_reg_8_13_sva <= 16'b0000000000000000;
      psum_reg_8_12_sva <= 16'b0000000000000000;
      psum_reg_8_11_sva <= 16'b0000000000000000;
      psum_reg_8_10_sva <= 16'b0000000000000000;
      psum_reg_8_9_sva <= 16'b0000000000000000;
      psum_reg_8_8_sva <= 16'b0000000000000000;
      psum_reg_8_7_sva <= 16'b0000000000000000;
      psum_reg_8_6_sva <= 16'b0000000000000000;
      psum_reg_8_5_sva <= 16'b0000000000000000;
      psum_reg_8_4_sva <= 16'b0000000000000000;
      psum_reg_8_3_sva <= 16'b0000000000000000;
      psum_reg_8_2_sva <= 16'b0000000000000000;
      psum_reg_8_1_sva <= 16'b0000000000000000;
      psum_reg_7_16_sva <= 16'b0000000000000000;
      psum_reg_7_15_sva <= 16'b0000000000000000;
      psum_reg_7_14_sva <= 16'b0000000000000000;
      psum_reg_7_13_sva <= 16'b0000000000000000;
      psum_reg_7_12_sva <= 16'b0000000000000000;
      psum_reg_7_11_sva <= 16'b0000000000000000;
      psum_reg_7_10_sva <= 16'b0000000000000000;
      psum_reg_7_9_sva <= 16'b0000000000000000;
      psum_reg_7_8_sva <= 16'b0000000000000000;
      psum_reg_7_7_sva <= 16'b0000000000000000;
      psum_reg_7_6_sva <= 16'b0000000000000000;
      psum_reg_7_5_sva <= 16'b0000000000000000;
      psum_reg_7_4_sva <= 16'b0000000000000000;
      psum_reg_7_3_sva <= 16'b0000000000000000;
      psum_reg_7_2_sva <= 16'b0000000000000000;
      psum_reg_7_1_sva <= 16'b0000000000000000;
      psum_reg_6_16_sva <= 16'b0000000000000000;
      psum_reg_6_15_sva <= 16'b0000000000000000;
      psum_reg_6_14_sva <= 16'b0000000000000000;
      psum_reg_6_13_sva <= 16'b0000000000000000;
      psum_reg_6_12_sva <= 16'b0000000000000000;
      psum_reg_6_11_sva <= 16'b0000000000000000;
      psum_reg_6_10_sva <= 16'b0000000000000000;
      psum_reg_6_9_sva <= 16'b0000000000000000;
      psum_reg_6_8_sva <= 16'b0000000000000000;
      psum_reg_6_7_sva <= 16'b0000000000000000;
      psum_reg_6_6_sva <= 16'b0000000000000000;
      psum_reg_6_5_sva <= 16'b0000000000000000;
      psum_reg_6_4_sva <= 16'b0000000000000000;
      psum_reg_6_3_sva <= 16'b0000000000000000;
      psum_reg_6_2_sva <= 16'b0000000000000000;
      psum_reg_6_1_sva <= 16'b0000000000000000;
      psum_reg_5_16_sva <= 16'b0000000000000000;
      psum_reg_5_15_sva <= 16'b0000000000000000;
      psum_reg_5_14_sva <= 16'b0000000000000000;
      psum_reg_5_13_sva <= 16'b0000000000000000;
      psum_reg_5_12_sva <= 16'b0000000000000000;
      psum_reg_5_11_sva <= 16'b0000000000000000;
      psum_reg_5_10_sva <= 16'b0000000000000000;
      psum_reg_5_9_sva <= 16'b0000000000000000;
      psum_reg_5_8_sva <= 16'b0000000000000000;
      psum_reg_5_7_sva <= 16'b0000000000000000;
      psum_reg_5_6_sva <= 16'b0000000000000000;
      psum_reg_5_5_sva <= 16'b0000000000000000;
      psum_reg_5_4_sva <= 16'b0000000000000000;
      psum_reg_5_3_sva <= 16'b0000000000000000;
      psum_reg_5_2_sva <= 16'b0000000000000000;
      psum_reg_5_1_sva <= 16'b0000000000000000;
      psum_reg_4_16_sva <= 16'b0000000000000000;
      psum_reg_4_15_sva <= 16'b0000000000000000;
      psum_reg_4_14_sva <= 16'b0000000000000000;
      psum_reg_4_13_sva <= 16'b0000000000000000;
      psum_reg_4_12_sva <= 16'b0000000000000000;
      psum_reg_4_11_sva <= 16'b0000000000000000;
      psum_reg_4_10_sva <= 16'b0000000000000000;
      psum_reg_4_9_sva <= 16'b0000000000000000;
      psum_reg_4_8_sva <= 16'b0000000000000000;
      psum_reg_4_7_sva <= 16'b0000000000000000;
      psum_reg_4_6_sva <= 16'b0000000000000000;
      psum_reg_4_5_sva <= 16'b0000000000000000;
      psum_reg_4_4_sva <= 16'b0000000000000000;
      psum_reg_4_3_sva <= 16'b0000000000000000;
      psum_reg_4_2_sva <= 16'b0000000000000000;
      psum_reg_4_1_sva <= 16'b0000000000000000;
      psum_reg_3_16_sva <= 16'b0000000000000000;
      psum_reg_3_15_sva <= 16'b0000000000000000;
      psum_reg_3_14_sva <= 16'b0000000000000000;
      psum_reg_3_13_sva <= 16'b0000000000000000;
      psum_reg_3_12_sva <= 16'b0000000000000000;
      psum_reg_3_11_sva <= 16'b0000000000000000;
      psum_reg_3_10_sva <= 16'b0000000000000000;
      psum_reg_3_9_sva <= 16'b0000000000000000;
      psum_reg_3_8_sva <= 16'b0000000000000000;
      psum_reg_3_7_sva <= 16'b0000000000000000;
      psum_reg_3_6_sva <= 16'b0000000000000000;
      psum_reg_3_5_sva <= 16'b0000000000000000;
      psum_reg_3_4_sva <= 16'b0000000000000000;
      psum_reg_3_3_sva <= 16'b0000000000000000;
      psum_reg_3_2_sva <= 16'b0000000000000000;
      psum_reg_3_1_sva <= 16'b0000000000000000;
      psum_reg_2_16_sva <= 16'b0000000000000000;
      psum_reg_2_15_sva <= 16'b0000000000000000;
      psum_reg_2_14_sva <= 16'b0000000000000000;
      psum_reg_2_13_sva <= 16'b0000000000000000;
      psum_reg_2_12_sva <= 16'b0000000000000000;
      psum_reg_2_11_sva <= 16'b0000000000000000;
      psum_reg_2_10_sva <= 16'b0000000000000000;
      psum_reg_2_9_sva <= 16'b0000000000000000;
      psum_reg_2_8_sva <= 16'b0000000000000000;
      psum_reg_2_7_sva <= 16'b0000000000000000;
      psum_reg_2_6_sva <= 16'b0000000000000000;
      psum_reg_2_5_sva <= 16'b0000000000000000;
      psum_reg_2_4_sva <= 16'b0000000000000000;
      psum_reg_2_3_sva <= 16'b0000000000000000;
      psum_reg_2_2_sva <= 16'b0000000000000000;
      psum_reg_2_1_sva <= 16'b0000000000000000;
      psum_reg_1_16_sva <= 16'b0000000000000000;
      psum_reg_1_15_sva <= 16'b0000000000000000;
      psum_reg_1_14_sva <= 16'b0000000000000000;
      psum_reg_1_13_sva <= 16'b0000000000000000;
      psum_reg_1_12_sva <= 16'b0000000000000000;
      psum_reg_1_11_sva <= 16'b0000000000000000;
      psum_reg_1_10_sva <= 16'b0000000000000000;
      psum_reg_1_9_sva <= 16'b0000000000000000;
      psum_reg_1_8_sva <= 16'b0000000000000000;
      psum_reg_1_7_sva <= 16'b0000000000000000;
      psum_reg_1_6_sva <= 16'b0000000000000000;
      psum_reg_1_5_sva <= 16'b0000000000000000;
      psum_reg_1_4_sva <= 16'b0000000000000000;
      psum_reg_1_3_sva <= 16'b0000000000000000;
      psum_reg_1_2_sva <= 16'b0000000000000000;
      psum_reg_1_1_sva <= 16'b0000000000000000;
      input_reg_16_15_sva <= 8'b00000000;
      input_reg_16_14_sva <= 8'b00000000;
      input_reg_16_13_sva <= 8'b00000000;
      input_reg_16_12_sva <= 8'b00000000;
      input_reg_16_11_sva <= 8'b00000000;
      input_reg_16_10_sva <= 8'b00000000;
      input_reg_16_9_sva <= 8'b00000000;
      input_reg_16_8_sva <= 8'b00000000;
      input_reg_16_7_sva <= 8'b00000000;
      input_reg_16_6_sva <= 8'b00000000;
      input_reg_16_5_sva <= 8'b00000000;
      input_reg_16_4_sva <= 8'b00000000;
      input_reg_16_3_sva <= 8'b00000000;
      input_reg_16_2_sva <= 8'b00000000;
      input_reg_16_1_sva <= 8'b00000000;
      input_reg_15_15_sva <= 8'b00000000;
      input_reg_15_14_sva <= 8'b00000000;
      input_reg_15_13_sva <= 8'b00000000;
      input_reg_15_12_sva <= 8'b00000000;
      input_reg_15_11_sva <= 8'b00000000;
      input_reg_15_10_sva <= 8'b00000000;
      input_reg_15_9_sva <= 8'b00000000;
      input_reg_15_8_sva <= 8'b00000000;
      input_reg_15_7_sva <= 8'b00000000;
      input_reg_15_6_sva <= 8'b00000000;
      input_reg_15_5_sva <= 8'b00000000;
      input_reg_15_4_sva <= 8'b00000000;
      input_reg_15_3_sva <= 8'b00000000;
      input_reg_15_2_sva <= 8'b00000000;
      input_reg_15_1_sva <= 8'b00000000;
      input_reg_14_15_sva <= 8'b00000000;
      input_reg_14_14_sva <= 8'b00000000;
      input_reg_14_13_sva <= 8'b00000000;
      input_reg_14_12_sva <= 8'b00000000;
      input_reg_14_11_sva <= 8'b00000000;
      input_reg_14_10_sva <= 8'b00000000;
      input_reg_14_9_sva <= 8'b00000000;
      input_reg_14_8_sva <= 8'b00000000;
      input_reg_14_7_sva <= 8'b00000000;
      input_reg_14_6_sva <= 8'b00000000;
      input_reg_14_5_sva <= 8'b00000000;
      input_reg_14_4_sva <= 8'b00000000;
      input_reg_14_3_sva <= 8'b00000000;
      input_reg_14_2_sva <= 8'b00000000;
      input_reg_14_1_sva <= 8'b00000000;
      input_reg_13_15_sva <= 8'b00000000;
      input_reg_13_14_sva <= 8'b00000000;
      input_reg_13_13_sva <= 8'b00000000;
      input_reg_13_12_sva <= 8'b00000000;
      input_reg_13_11_sva <= 8'b00000000;
      input_reg_13_10_sva <= 8'b00000000;
      input_reg_13_9_sva <= 8'b00000000;
      input_reg_13_8_sva <= 8'b00000000;
      input_reg_13_7_sva <= 8'b00000000;
      input_reg_13_6_sva <= 8'b00000000;
      input_reg_13_5_sva <= 8'b00000000;
      input_reg_13_4_sva <= 8'b00000000;
      input_reg_13_3_sva <= 8'b00000000;
      input_reg_13_2_sva <= 8'b00000000;
      input_reg_13_1_sva <= 8'b00000000;
      input_reg_12_15_sva <= 8'b00000000;
      input_reg_12_14_sva <= 8'b00000000;
      input_reg_12_13_sva <= 8'b00000000;
      input_reg_12_12_sva <= 8'b00000000;
      input_reg_12_11_sva <= 8'b00000000;
      input_reg_12_10_sva <= 8'b00000000;
      input_reg_12_9_sva <= 8'b00000000;
      input_reg_12_8_sva <= 8'b00000000;
      input_reg_12_7_sva <= 8'b00000000;
      input_reg_12_6_sva <= 8'b00000000;
      input_reg_12_5_sva <= 8'b00000000;
      input_reg_12_4_sva <= 8'b00000000;
      input_reg_12_3_sva <= 8'b00000000;
      input_reg_12_2_sva <= 8'b00000000;
      input_reg_12_1_sva <= 8'b00000000;
      input_reg_11_15_sva <= 8'b00000000;
      input_reg_11_14_sva <= 8'b00000000;
      input_reg_11_13_sva <= 8'b00000000;
      input_reg_11_12_sva <= 8'b00000000;
      input_reg_11_11_sva <= 8'b00000000;
      input_reg_11_10_sva <= 8'b00000000;
      input_reg_11_9_sva <= 8'b00000000;
      input_reg_11_8_sva <= 8'b00000000;
      input_reg_11_7_sva <= 8'b00000000;
      input_reg_11_6_sva <= 8'b00000000;
      input_reg_11_5_sva <= 8'b00000000;
      input_reg_11_4_sva <= 8'b00000000;
      input_reg_11_3_sva <= 8'b00000000;
      input_reg_11_2_sva <= 8'b00000000;
      input_reg_11_1_sva <= 8'b00000000;
      input_reg_10_15_sva <= 8'b00000000;
      input_reg_10_14_sva <= 8'b00000000;
      input_reg_10_13_sva <= 8'b00000000;
      input_reg_10_12_sva <= 8'b00000000;
      input_reg_10_11_sva <= 8'b00000000;
      input_reg_10_10_sva <= 8'b00000000;
      input_reg_10_9_sva <= 8'b00000000;
      input_reg_10_8_sva <= 8'b00000000;
      input_reg_10_7_sva <= 8'b00000000;
      input_reg_10_6_sva <= 8'b00000000;
      input_reg_10_5_sva <= 8'b00000000;
      input_reg_10_4_sva <= 8'b00000000;
      input_reg_10_3_sva <= 8'b00000000;
      input_reg_10_2_sva <= 8'b00000000;
      input_reg_10_1_sva <= 8'b00000000;
      input_reg_9_15_sva <= 8'b00000000;
      input_reg_9_14_sva <= 8'b00000000;
      input_reg_9_13_sva <= 8'b00000000;
      input_reg_9_12_sva <= 8'b00000000;
      input_reg_9_11_sva <= 8'b00000000;
      input_reg_9_10_sva <= 8'b00000000;
      input_reg_9_9_sva <= 8'b00000000;
      input_reg_9_8_sva <= 8'b00000000;
      input_reg_9_7_sva <= 8'b00000000;
      input_reg_9_6_sva <= 8'b00000000;
      input_reg_9_5_sva <= 8'b00000000;
      input_reg_9_4_sva <= 8'b00000000;
      input_reg_9_3_sva <= 8'b00000000;
      input_reg_9_2_sva <= 8'b00000000;
      input_reg_9_1_sva <= 8'b00000000;
      input_reg_8_15_sva <= 8'b00000000;
      input_reg_8_14_sva <= 8'b00000000;
      input_reg_8_13_sva <= 8'b00000000;
      input_reg_8_12_sva <= 8'b00000000;
      input_reg_8_11_sva <= 8'b00000000;
      input_reg_8_10_sva <= 8'b00000000;
      input_reg_8_9_sva <= 8'b00000000;
      input_reg_8_8_sva <= 8'b00000000;
      input_reg_8_7_sva <= 8'b00000000;
      input_reg_8_6_sva <= 8'b00000000;
      input_reg_8_5_sva <= 8'b00000000;
      input_reg_8_4_sva <= 8'b00000000;
      input_reg_8_3_sva <= 8'b00000000;
      input_reg_8_2_sva <= 8'b00000000;
      input_reg_8_1_sva <= 8'b00000000;
      input_reg_7_15_sva <= 8'b00000000;
      input_reg_7_14_sva <= 8'b00000000;
      input_reg_7_13_sva <= 8'b00000000;
      input_reg_7_12_sva <= 8'b00000000;
      input_reg_7_11_sva <= 8'b00000000;
      input_reg_7_10_sva <= 8'b00000000;
      input_reg_7_9_sva <= 8'b00000000;
      input_reg_7_8_sva <= 8'b00000000;
      input_reg_7_7_sva <= 8'b00000000;
      input_reg_7_6_sva <= 8'b00000000;
      input_reg_7_5_sva <= 8'b00000000;
      input_reg_7_4_sva <= 8'b00000000;
      input_reg_7_3_sva <= 8'b00000000;
      input_reg_7_2_sva <= 8'b00000000;
      input_reg_7_1_sva <= 8'b00000000;
      input_reg_6_15_sva <= 8'b00000000;
      input_reg_6_14_sva <= 8'b00000000;
      input_reg_6_13_sva <= 8'b00000000;
      input_reg_6_12_sva <= 8'b00000000;
      input_reg_6_11_sva <= 8'b00000000;
      input_reg_6_10_sva <= 8'b00000000;
      input_reg_6_9_sva <= 8'b00000000;
      input_reg_6_8_sva <= 8'b00000000;
      input_reg_6_7_sva <= 8'b00000000;
      input_reg_6_6_sva <= 8'b00000000;
      input_reg_6_5_sva <= 8'b00000000;
      input_reg_6_4_sva <= 8'b00000000;
      input_reg_6_3_sva <= 8'b00000000;
      input_reg_6_2_sva <= 8'b00000000;
      input_reg_6_1_sva <= 8'b00000000;
      input_reg_5_15_sva <= 8'b00000000;
      input_reg_5_14_sva <= 8'b00000000;
      input_reg_5_13_sva <= 8'b00000000;
      input_reg_5_12_sva <= 8'b00000000;
      input_reg_5_11_sva <= 8'b00000000;
      input_reg_5_10_sva <= 8'b00000000;
      input_reg_5_9_sva <= 8'b00000000;
      input_reg_5_8_sva <= 8'b00000000;
      input_reg_5_7_sva <= 8'b00000000;
      input_reg_5_6_sva <= 8'b00000000;
      input_reg_5_5_sva <= 8'b00000000;
      input_reg_5_4_sva <= 8'b00000000;
      input_reg_5_3_sva <= 8'b00000000;
      input_reg_5_2_sva <= 8'b00000000;
      input_reg_5_1_sva <= 8'b00000000;
      input_reg_4_15_sva <= 8'b00000000;
      input_reg_4_14_sva <= 8'b00000000;
      input_reg_4_13_sva <= 8'b00000000;
      input_reg_4_12_sva <= 8'b00000000;
      input_reg_4_11_sva <= 8'b00000000;
      input_reg_4_10_sva <= 8'b00000000;
      input_reg_4_9_sva <= 8'b00000000;
      input_reg_4_8_sva <= 8'b00000000;
      input_reg_4_7_sva <= 8'b00000000;
      input_reg_4_6_sva <= 8'b00000000;
      input_reg_4_5_sva <= 8'b00000000;
      input_reg_4_4_sva <= 8'b00000000;
      input_reg_4_3_sva <= 8'b00000000;
      input_reg_4_2_sva <= 8'b00000000;
      input_reg_4_1_sva <= 8'b00000000;
      input_reg_3_15_sva <= 8'b00000000;
      input_reg_3_14_sva <= 8'b00000000;
      input_reg_3_13_sva <= 8'b00000000;
      input_reg_3_12_sva <= 8'b00000000;
      input_reg_3_11_sva <= 8'b00000000;
      input_reg_3_10_sva <= 8'b00000000;
      input_reg_3_9_sva <= 8'b00000000;
      input_reg_3_8_sva <= 8'b00000000;
      input_reg_3_7_sva <= 8'b00000000;
      input_reg_3_6_sva <= 8'b00000000;
      input_reg_3_5_sva <= 8'b00000000;
      input_reg_3_4_sva <= 8'b00000000;
      input_reg_3_3_sva <= 8'b00000000;
      input_reg_3_2_sva <= 8'b00000000;
      input_reg_3_1_sva <= 8'b00000000;
      input_reg_2_15_sva <= 8'b00000000;
      input_reg_2_14_sva <= 8'b00000000;
      input_reg_2_13_sva <= 8'b00000000;
      input_reg_2_12_sva <= 8'b00000000;
      input_reg_2_11_sva <= 8'b00000000;
      input_reg_2_10_sva <= 8'b00000000;
      input_reg_2_9_sva <= 8'b00000000;
      input_reg_2_8_sva <= 8'b00000000;
      input_reg_2_7_sva <= 8'b00000000;
      input_reg_2_6_sva <= 8'b00000000;
      input_reg_2_5_sva <= 8'b00000000;
      input_reg_2_4_sva <= 8'b00000000;
      input_reg_2_3_sva <= 8'b00000000;
      input_reg_2_2_sva <= 8'b00000000;
      input_reg_2_1_sva <= 8'b00000000;
      input_reg_1_15_sva <= 8'b00000000;
      input_reg_1_14_sva <= 8'b00000000;
      input_reg_1_13_sva <= 8'b00000000;
      input_reg_1_12_sva <= 8'b00000000;
      input_reg_1_11_sva <= 8'b00000000;
      input_reg_1_10_sva <= 8'b00000000;
      input_reg_1_9_sva <= 8'b00000000;
      input_reg_1_8_sva <= 8'b00000000;
      input_reg_1_7_sva <= 8'b00000000;
      input_reg_1_6_sva <= 8'b00000000;
      input_reg_1_5_sva <= 8'b00000000;
      input_reg_1_4_sva <= 8'b00000000;
      input_reg_1_3_sva <= 8'b00000000;
      input_reg_1_2_sva <= 8'b00000000;
      input_reg_1_1_sva <= 8'b00000000;
    end
    else if ( psum_reg_and_cse ) begin
      psum_reg_16_16_sva <= MUX_v_16_2_2(psum_reg_16_16_sva, pe_0_0_run_cmp_1_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_15_sva <= MUX_v_16_2_2(psum_reg_16_15_sva, pe_0_0_run_cmp_17_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_14_sva <= MUX_v_16_2_2(psum_reg_16_14_sva, pe_0_0_run_cmp_33_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_13_sva <= MUX_v_16_2_2(psum_reg_16_13_sva, pe_0_0_run_cmp_49_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_12_sva <= MUX_v_16_2_2(psum_reg_16_12_sva, pe_0_0_run_cmp_65_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_11_sva <= MUX_v_16_2_2(psum_reg_16_11_sva, pe_0_0_run_cmp_81_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_10_sva <= MUX_v_16_2_2(psum_reg_16_10_sva, pe_0_0_run_cmp_97_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_9_sva <= MUX_v_16_2_2(psum_reg_16_9_sva, pe_0_0_run_cmp_113_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_8_sva <= MUX_v_16_2_2(psum_reg_16_8_sva, pe_0_0_run_cmp_129_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_7_sva <= MUX_v_16_2_2(psum_reg_16_7_sva, pe_0_0_run_cmp_145_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_6_sva <= MUX_v_16_2_2(psum_reg_16_6_sva, pe_0_0_run_cmp_161_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_5_sva <= MUX_v_16_2_2(psum_reg_16_5_sva, pe_0_0_run_cmp_177_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_4_sva <= MUX_v_16_2_2(psum_reg_16_4_sva, pe_0_0_run_cmp_193_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_3_sva <= MUX_v_16_2_2(psum_reg_16_3_sva, pe_0_0_run_cmp_209_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_2_sva <= MUX_v_16_2_2(psum_reg_16_2_sva, pe_0_0_run_cmp_225_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_16_1_sva <= MUX_v_16_2_2(psum_reg_16_1_sva, pe_0_0_run_cmp_241_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_16_sva <= MUX_v_16_2_2(psum_reg_15_16_sva, pe_0_0_run_cmp_2_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_15_sva <= MUX_v_16_2_2(psum_reg_15_15_sva, pe_0_0_run_cmp_18_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_14_sva <= MUX_v_16_2_2(psum_reg_15_14_sva, pe_0_0_run_cmp_34_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_13_sva <= MUX_v_16_2_2(psum_reg_15_13_sva, pe_0_0_run_cmp_50_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_12_sva <= MUX_v_16_2_2(psum_reg_15_12_sva, pe_0_0_run_cmp_66_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_11_sva <= MUX_v_16_2_2(psum_reg_15_11_sva, pe_0_0_run_cmp_82_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_10_sva <= MUX_v_16_2_2(psum_reg_15_10_sva, pe_0_0_run_cmp_98_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_9_sva <= MUX_v_16_2_2(psum_reg_15_9_sva, pe_0_0_run_cmp_114_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_8_sva <= MUX_v_16_2_2(psum_reg_15_8_sva, pe_0_0_run_cmp_130_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_7_sva <= MUX_v_16_2_2(psum_reg_15_7_sva, pe_0_0_run_cmp_146_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_6_sva <= MUX_v_16_2_2(psum_reg_15_6_sva, pe_0_0_run_cmp_162_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_5_sva <= MUX_v_16_2_2(psum_reg_15_5_sva, pe_0_0_run_cmp_178_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_4_sva <= MUX_v_16_2_2(psum_reg_15_4_sva, pe_0_0_run_cmp_194_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_3_sva <= MUX_v_16_2_2(psum_reg_15_3_sva, pe_0_0_run_cmp_210_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_2_sva <= MUX_v_16_2_2(psum_reg_15_2_sva, pe_0_0_run_cmp_226_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_15_1_sva <= MUX_v_16_2_2(psum_reg_15_1_sva, pe_0_0_run_cmp_242_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_16_sva <= MUX_v_16_2_2(psum_reg_14_16_sva, pe_0_0_run_cmp_3_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_15_sva <= MUX_v_16_2_2(psum_reg_14_15_sva, pe_0_0_run_cmp_19_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_14_sva <= MUX_v_16_2_2(psum_reg_14_14_sva, pe_0_0_run_cmp_35_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_13_sva <= MUX_v_16_2_2(psum_reg_14_13_sva, pe_0_0_run_cmp_51_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_12_sva <= MUX_v_16_2_2(psum_reg_14_12_sva, pe_0_0_run_cmp_67_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_11_sva <= MUX_v_16_2_2(psum_reg_14_11_sva, pe_0_0_run_cmp_83_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_10_sva <= MUX_v_16_2_2(psum_reg_14_10_sva, pe_0_0_run_cmp_99_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_9_sva <= MUX_v_16_2_2(psum_reg_14_9_sva, pe_0_0_run_cmp_115_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_8_sva <= MUX_v_16_2_2(psum_reg_14_8_sva, pe_0_0_run_cmp_131_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_7_sva <= MUX_v_16_2_2(psum_reg_14_7_sva, pe_0_0_run_cmp_147_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_6_sva <= MUX_v_16_2_2(psum_reg_14_6_sva, pe_0_0_run_cmp_163_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_5_sva <= MUX_v_16_2_2(psum_reg_14_5_sva, pe_0_0_run_cmp_179_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_4_sva <= MUX_v_16_2_2(psum_reg_14_4_sva, pe_0_0_run_cmp_195_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_3_sva <= MUX_v_16_2_2(psum_reg_14_3_sva, pe_0_0_run_cmp_211_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_2_sva <= MUX_v_16_2_2(psum_reg_14_2_sva, pe_0_0_run_cmp_227_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_14_1_sva <= MUX_v_16_2_2(psum_reg_14_1_sva, pe_0_0_run_cmp_243_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_16_sva <= MUX_v_16_2_2(psum_reg_13_16_sva, pe_0_0_run_cmp_4_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_15_sva <= MUX_v_16_2_2(psum_reg_13_15_sva, pe_0_0_run_cmp_20_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_14_sva <= MUX_v_16_2_2(psum_reg_13_14_sva, pe_0_0_run_cmp_36_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_13_sva <= MUX_v_16_2_2(psum_reg_13_13_sva, pe_0_0_run_cmp_52_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_12_sva <= MUX_v_16_2_2(psum_reg_13_12_sva, pe_0_0_run_cmp_68_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_11_sva <= MUX_v_16_2_2(psum_reg_13_11_sva, pe_0_0_run_cmp_84_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_10_sva <= MUX_v_16_2_2(psum_reg_13_10_sva, pe_0_0_run_cmp_100_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_9_sva <= MUX_v_16_2_2(psum_reg_13_9_sva, pe_0_0_run_cmp_116_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_8_sva <= MUX_v_16_2_2(psum_reg_13_8_sva, pe_0_0_run_cmp_132_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_7_sva <= MUX_v_16_2_2(psum_reg_13_7_sva, pe_0_0_run_cmp_148_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_6_sva <= MUX_v_16_2_2(psum_reg_13_6_sva, pe_0_0_run_cmp_164_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_5_sva <= MUX_v_16_2_2(psum_reg_13_5_sva, pe_0_0_run_cmp_180_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_4_sva <= MUX_v_16_2_2(psum_reg_13_4_sva, pe_0_0_run_cmp_196_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_3_sva <= MUX_v_16_2_2(psum_reg_13_3_sva, pe_0_0_run_cmp_212_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_2_sva <= MUX_v_16_2_2(psum_reg_13_2_sva, pe_0_0_run_cmp_228_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_13_1_sva <= MUX_v_16_2_2(psum_reg_13_1_sva, pe_0_0_run_cmp_244_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_16_sva <= MUX_v_16_2_2(psum_reg_12_16_sva, pe_0_0_run_cmp_5_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_15_sva <= MUX_v_16_2_2(psum_reg_12_15_sva, pe_0_0_run_cmp_21_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_14_sva <= MUX_v_16_2_2(psum_reg_12_14_sva, pe_0_0_run_cmp_37_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_13_sva <= MUX_v_16_2_2(psum_reg_12_13_sva, pe_0_0_run_cmp_53_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_12_sva <= MUX_v_16_2_2(psum_reg_12_12_sva, pe_0_0_run_cmp_69_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_11_sva <= MUX_v_16_2_2(psum_reg_12_11_sva, pe_0_0_run_cmp_85_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_10_sva <= MUX_v_16_2_2(psum_reg_12_10_sva, pe_0_0_run_cmp_101_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_9_sva <= MUX_v_16_2_2(psum_reg_12_9_sva, pe_0_0_run_cmp_117_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_8_sva <= MUX_v_16_2_2(psum_reg_12_8_sva, pe_0_0_run_cmp_133_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_7_sva <= MUX_v_16_2_2(psum_reg_12_7_sva, pe_0_0_run_cmp_149_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_6_sva <= MUX_v_16_2_2(psum_reg_12_6_sva, pe_0_0_run_cmp_165_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_5_sva <= MUX_v_16_2_2(psum_reg_12_5_sva, pe_0_0_run_cmp_181_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_4_sva <= MUX_v_16_2_2(psum_reg_12_4_sva, pe_0_0_run_cmp_197_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_3_sva <= MUX_v_16_2_2(psum_reg_12_3_sva, pe_0_0_run_cmp_213_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_2_sva <= MUX_v_16_2_2(psum_reg_12_2_sva, pe_0_0_run_cmp_229_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_12_1_sva <= MUX_v_16_2_2(psum_reg_12_1_sva, pe_0_0_run_cmp_245_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_16_sva <= MUX_v_16_2_2(psum_reg_11_16_sva, pe_0_0_run_cmp_6_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_15_sva <= MUX_v_16_2_2(psum_reg_11_15_sva, pe_0_0_run_cmp_22_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_14_sva <= MUX_v_16_2_2(psum_reg_11_14_sva, pe_0_0_run_cmp_38_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_13_sva <= MUX_v_16_2_2(psum_reg_11_13_sva, pe_0_0_run_cmp_54_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_12_sva <= MUX_v_16_2_2(psum_reg_11_12_sva, pe_0_0_run_cmp_70_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_11_sva <= MUX_v_16_2_2(psum_reg_11_11_sva, pe_0_0_run_cmp_86_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_10_sva <= MUX_v_16_2_2(psum_reg_11_10_sva, pe_0_0_run_cmp_102_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_9_sva <= MUX_v_16_2_2(psum_reg_11_9_sva, pe_0_0_run_cmp_118_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_8_sva <= MUX_v_16_2_2(psum_reg_11_8_sva, pe_0_0_run_cmp_134_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_7_sva <= MUX_v_16_2_2(psum_reg_11_7_sva, pe_0_0_run_cmp_150_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_6_sva <= MUX_v_16_2_2(psum_reg_11_6_sva, pe_0_0_run_cmp_166_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_5_sva <= MUX_v_16_2_2(psum_reg_11_5_sva, pe_0_0_run_cmp_182_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_4_sva <= MUX_v_16_2_2(psum_reg_11_4_sva, pe_0_0_run_cmp_198_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_3_sva <= MUX_v_16_2_2(psum_reg_11_3_sva, pe_0_0_run_cmp_214_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_2_sva <= MUX_v_16_2_2(psum_reg_11_2_sva, pe_0_0_run_cmp_230_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_11_1_sva <= MUX_v_16_2_2(psum_reg_11_1_sva, pe_0_0_run_cmp_246_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_16_sva <= MUX_v_16_2_2(psum_reg_10_16_sva, pe_0_0_run_cmp_7_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_15_sva <= MUX_v_16_2_2(psum_reg_10_15_sva, pe_0_0_run_cmp_23_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_14_sva <= MUX_v_16_2_2(psum_reg_10_14_sva, pe_0_0_run_cmp_39_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_13_sva <= MUX_v_16_2_2(psum_reg_10_13_sva, pe_0_0_run_cmp_55_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_12_sva <= MUX_v_16_2_2(psum_reg_10_12_sva, pe_0_0_run_cmp_71_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_11_sva <= MUX_v_16_2_2(psum_reg_10_11_sva, pe_0_0_run_cmp_87_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_10_sva <= MUX_v_16_2_2(psum_reg_10_10_sva, pe_0_0_run_cmp_103_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_9_sva <= MUX_v_16_2_2(psum_reg_10_9_sva, pe_0_0_run_cmp_119_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_8_sva <= MUX_v_16_2_2(psum_reg_10_8_sva, pe_0_0_run_cmp_135_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_7_sva <= MUX_v_16_2_2(psum_reg_10_7_sva, pe_0_0_run_cmp_151_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_6_sva <= MUX_v_16_2_2(psum_reg_10_6_sva, pe_0_0_run_cmp_167_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_5_sva <= MUX_v_16_2_2(psum_reg_10_5_sva, pe_0_0_run_cmp_183_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_4_sva <= MUX_v_16_2_2(psum_reg_10_4_sva, pe_0_0_run_cmp_199_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_3_sva <= MUX_v_16_2_2(psum_reg_10_3_sva, pe_0_0_run_cmp_215_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_2_sva <= MUX_v_16_2_2(psum_reg_10_2_sva, pe_0_0_run_cmp_231_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_10_1_sva <= MUX_v_16_2_2(psum_reg_10_1_sva, pe_0_0_run_cmp_247_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_16_sva <= MUX_v_16_2_2(psum_reg_9_16_sva, pe_0_0_run_cmp_8_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_15_sva <= MUX_v_16_2_2(psum_reg_9_15_sva, pe_0_0_run_cmp_24_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_14_sva <= MUX_v_16_2_2(psum_reg_9_14_sva, pe_0_0_run_cmp_40_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_13_sva <= MUX_v_16_2_2(psum_reg_9_13_sva, pe_0_0_run_cmp_56_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_12_sva <= MUX_v_16_2_2(psum_reg_9_12_sva, pe_0_0_run_cmp_72_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_11_sva <= MUX_v_16_2_2(psum_reg_9_11_sva, pe_0_0_run_cmp_88_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_10_sva <= MUX_v_16_2_2(psum_reg_9_10_sva, pe_0_0_run_cmp_104_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_9_sva <= MUX_v_16_2_2(psum_reg_9_9_sva, pe_0_0_run_cmp_120_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_8_sva <= MUX_v_16_2_2(psum_reg_9_8_sva, pe_0_0_run_cmp_136_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_7_sva <= MUX_v_16_2_2(psum_reg_9_7_sva, pe_0_0_run_cmp_152_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_6_sva <= MUX_v_16_2_2(psum_reg_9_6_sva, pe_0_0_run_cmp_168_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_5_sva <= MUX_v_16_2_2(psum_reg_9_5_sva, pe_0_0_run_cmp_184_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_4_sva <= MUX_v_16_2_2(psum_reg_9_4_sva, pe_0_0_run_cmp_200_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_3_sva <= MUX_v_16_2_2(psum_reg_9_3_sva, pe_0_0_run_cmp_216_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_2_sva <= MUX_v_16_2_2(psum_reg_9_2_sva, pe_0_0_run_cmp_232_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_9_1_sva <= MUX_v_16_2_2(psum_reg_9_1_sva, pe_0_0_run_cmp_248_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_16_sva <= MUX_v_16_2_2(psum_reg_8_16_sva, pe_0_0_run_cmp_9_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_15_sva <= MUX_v_16_2_2(psum_reg_8_15_sva, pe_0_0_run_cmp_25_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_14_sva <= MUX_v_16_2_2(psum_reg_8_14_sva, pe_0_0_run_cmp_41_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_13_sva <= MUX_v_16_2_2(psum_reg_8_13_sva, pe_0_0_run_cmp_57_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_12_sva <= MUX_v_16_2_2(psum_reg_8_12_sva, pe_0_0_run_cmp_73_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_11_sva <= MUX_v_16_2_2(psum_reg_8_11_sva, pe_0_0_run_cmp_89_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_10_sva <= MUX_v_16_2_2(psum_reg_8_10_sva, pe_0_0_run_cmp_105_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_9_sva <= MUX_v_16_2_2(psum_reg_8_9_sva, pe_0_0_run_cmp_121_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_8_sva <= MUX_v_16_2_2(psum_reg_8_8_sva, pe_0_0_run_cmp_137_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_7_sva <= MUX_v_16_2_2(psum_reg_8_7_sva, pe_0_0_run_cmp_153_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_6_sva <= MUX_v_16_2_2(psum_reg_8_6_sva, pe_0_0_run_cmp_169_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_5_sva <= MUX_v_16_2_2(psum_reg_8_5_sva, pe_0_0_run_cmp_185_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_4_sva <= MUX_v_16_2_2(psum_reg_8_4_sva, pe_0_0_run_cmp_201_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_3_sva <= MUX_v_16_2_2(psum_reg_8_3_sva, pe_0_0_run_cmp_217_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_2_sva <= MUX_v_16_2_2(psum_reg_8_2_sva, pe_0_0_run_cmp_233_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_8_1_sva <= MUX_v_16_2_2(psum_reg_8_1_sva, pe_0_0_run_cmp_249_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_16_sva <= MUX_v_16_2_2(psum_reg_7_16_sva, pe_0_0_run_cmp_10_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_15_sva <= MUX_v_16_2_2(psum_reg_7_15_sva, pe_0_0_run_cmp_26_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_14_sva <= MUX_v_16_2_2(psum_reg_7_14_sva, pe_0_0_run_cmp_42_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_13_sva <= MUX_v_16_2_2(psum_reg_7_13_sva, pe_0_0_run_cmp_58_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_12_sva <= MUX_v_16_2_2(psum_reg_7_12_sva, pe_0_0_run_cmp_74_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_11_sva <= MUX_v_16_2_2(psum_reg_7_11_sva, pe_0_0_run_cmp_90_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_10_sva <= MUX_v_16_2_2(psum_reg_7_10_sva, pe_0_0_run_cmp_106_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_9_sva <= MUX_v_16_2_2(psum_reg_7_9_sva, pe_0_0_run_cmp_122_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_8_sva <= MUX_v_16_2_2(psum_reg_7_8_sva, pe_0_0_run_cmp_138_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_7_sva <= MUX_v_16_2_2(psum_reg_7_7_sva, pe_0_0_run_cmp_154_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_6_sva <= MUX_v_16_2_2(psum_reg_7_6_sva, pe_0_0_run_cmp_170_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_5_sva <= MUX_v_16_2_2(psum_reg_7_5_sva, pe_0_0_run_cmp_186_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_4_sva <= MUX_v_16_2_2(psum_reg_7_4_sva, pe_0_0_run_cmp_202_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_3_sva <= MUX_v_16_2_2(psum_reg_7_3_sva, pe_0_0_run_cmp_218_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_2_sva <= MUX_v_16_2_2(psum_reg_7_2_sva, pe_0_0_run_cmp_234_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_7_1_sva <= MUX_v_16_2_2(psum_reg_7_1_sva, pe_0_0_run_cmp_250_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_16_sva <= MUX_v_16_2_2(psum_reg_6_16_sva, pe_0_0_run_cmp_11_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_15_sva <= MUX_v_16_2_2(psum_reg_6_15_sva, pe_0_0_run_cmp_27_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_14_sva <= MUX_v_16_2_2(psum_reg_6_14_sva, pe_0_0_run_cmp_43_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_13_sva <= MUX_v_16_2_2(psum_reg_6_13_sva, pe_0_0_run_cmp_59_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_12_sva <= MUX_v_16_2_2(psum_reg_6_12_sva, pe_0_0_run_cmp_75_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_11_sva <= MUX_v_16_2_2(psum_reg_6_11_sva, pe_0_0_run_cmp_91_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_10_sva <= MUX_v_16_2_2(psum_reg_6_10_sva, pe_0_0_run_cmp_107_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_9_sva <= MUX_v_16_2_2(psum_reg_6_9_sva, pe_0_0_run_cmp_123_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_8_sva <= MUX_v_16_2_2(psum_reg_6_8_sva, pe_0_0_run_cmp_139_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_7_sva <= MUX_v_16_2_2(psum_reg_6_7_sva, pe_0_0_run_cmp_155_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_6_sva <= MUX_v_16_2_2(psum_reg_6_6_sva, pe_0_0_run_cmp_171_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_5_sva <= MUX_v_16_2_2(psum_reg_6_5_sva, pe_0_0_run_cmp_187_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_4_sva <= MUX_v_16_2_2(psum_reg_6_4_sva, pe_0_0_run_cmp_203_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_3_sva <= MUX_v_16_2_2(psum_reg_6_3_sva, pe_0_0_run_cmp_219_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_2_sva <= MUX_v_16_2_2(psum_reg_6_2_sva, pe_0_0_run_cmp_235_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_6_1_sva <= MUX_v_16_2_2(psum_reg_6_1_sva, pe_0_0_run_cmp_251_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_16_sva <= MUX_v_16_2_2(psum_reg_5_16_sva, pe_0_0_run_cmp_12_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_15_sva <= MUX_v_16_2_2(psum_reg_5_15_sva, pe_0_0_run_cmp_28_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_14_sva <= MUX_v_16_2_2(psum_reg_5_14_sva, pe_0_0_run_cmp_44_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_13_sva <= MUX_v_16_2_2(psum_reg_5_13_sva, pe_0_0_run_cmp_60_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_12_sva <= MUX_v_16_2_2(psum_reg_5_12_sva, pe_0_0_run_cmp_76_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_11_sva <= MUX_v_16_2_2(psum_reg_5_11_sva, pe_0_0_run_cmp_92_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_10_sva <= MUX_v_16_2_2(psum_reg_5_10_sva, pe_0_0_run_cmp_108_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_9_sva <= MUX_v_16_2_2(psum_reg_5_9_sva, pe_0_0_run_cmp_124_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_8_sva <= MUX_v_16_2_2(psum_reg_5_8_sva, pe_0_0_run_cmp_140_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_7_sva <= MUX_v_16_2_2(psum_reg_5_7_sva, pe_0_0_run_cmp_156_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_6_sva <= MUX_v_16_2_2(psum_reg_5_6_sva, pe_0_0_run_cmp_172_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_5_sva <= MUX_v_16_2_2(psum_reg_5_5_sva, pe_0_0_run_cmp_188_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_4_sva <= MUX_v_16_2_2(psum_reg_5_4_sva, pe_0_0_run_cmp_204_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_3_sva <= MUX_v_16_2_2(psum_reg_5_3_sva, pe_0_0_run_cmp_220_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_2_sva <= MUX_v_16_2_2(psum_reg_5_2_sva, pe_0_0_run_cmp_236_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_5_1_sva <= MUX_v_16_2_2(psum_reg_5_1_sva, pe_0_0_run_cmp_252_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_16_sva <= MUX_v_16_2_2(psum_reg_4_16_sva, pe_0_0_run_cmp_13_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_15_sva <= MUX_v_16_2_2(psum_reg_4_15_sva, pe_0_0_run_cmp_29_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_14_sva <= MUX_v_16_2_2(psum_reg_4_14_sva, pe_0_0_run_cmp_45_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_13_sva <= MUX_v_16_2_2(psum_reg_4_13_sva, pe_0_0_run_cmp_61_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_12_sva <= MUX_v_16_2_2(psum_reg_4_12_sva, pe_0_0_run_cmp_77_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_11_sva <= MUX_v_16_2_2(psum_reg_4_11_sva, pe_0_0_run_cmp_93_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_10_sva <= MUX_v_16_2_2(psum_reg_4_10_sva, pe_0_0_run_cmp_109_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_9_sva <= MUX_v_16_2_2(psum_reg_4_9_sva, pe_0_0_run_cmp_125_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_8_sva <= MUX_v_16_2_2(psum_reg_4_8_sva, pe_0_0_run_cmp_141_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_7_sva <= MUX_v_16_2_2(psum_reg_4_7_sva, pe_0_0_run_cmp_157_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_6_sva <= MUX_v_16_2_2(psum_reg_4_6_sva, pe_0_0_run_cmp_173_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_5_sva <= MUX_v_16_2_2(psum_reg_4_5_sva, pe_0_0_run_cmp_189_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_4_sva <= MUX_v_16_2_2(psum_reg_4_4_sva, pe_0_0_run_cmp_205_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_3_sva <= MUX_v_16_2_2(psum_reg_4_3_sva, pe_0_0_run_cmp_221_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_2_sva <= MUX_v_16_2_2(psum_reg_4_2_sva, pe_0_0_run_cmp_237_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_4_1_sva <= MUX_v_16_2_2(psum_reg_4_1_sva, pe_0_0_run_cmp_253_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_16_sva <= MUX_v_16_2_2(psum_reg_3_16_sva, pe_0_0_run_cmp_14_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_15_sva <= MUX_v_16_2_2(psum_reg_3_15_sva, pe_0_0_run_cmp_30_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_14_sva <= MUX_v_16_2_2(psum_reg_3_14_sva, pe_0_0_run_cmp_46_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_13_sva <= MUX_v_16_2_2(psum_reg_3_13_sva, pe_0_0_run_cmp_62_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_12_sva <= MUX_v_16_2_2(psum_reg_3_12_sva, pe_0_0_run_cmp_78_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_11_sva <= MUX_v_16_2_2(psum_reg_3_11_sva, pe_0_0_run_cmp_94_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_10_sva <= MUX_v_16_2_2(psum_reg_3_10_sva, pe_0_0_run_cmp_110_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_9_sva <= MUX_v_16_2_2(psum_reg_3_9_sva, pe_0_0_run_cmp_126_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_8_sva <= MUX_v_16_2_2(psum_reg_3_8_sva, pe_0_0_run_cmp_142_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_7_sva <= MUX_v_16_2_2(psum_reg_3_7_sva, pe_0_0_run_cmp_158_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_6_sva <= MUX_v_16_2_2(psum_reg_3_6_sva, pe_0_0_run_cmp_174_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_5_sva <= MUX_v_16_2_2(psum_reg_3_5_sva, pe_0_0_run_cmp_190_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_4_sva <= MUX_v_16_2_2(psum_reg_3_4_sva, pe_0_0_run_cmp_206_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_3_sva <= MUX_v_16_2_2(psum_reg_3_3_sva, pe_0_0_run_cmp_222_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_2_sva <= MUX_v_16_2_2(psum_reg_3_2_sva, pe_0_0_run_cmp_238_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_3_1_sva <= MUX_v_16_2_2(psum_reg_3_1_sva, pe_0_0_run_cmp_254_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_16_sva <= MUX_v_16_2_2(psum_reg_2_16_sva, pe_0_0_run_cmp_15_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_15_sva <= MUX_v_16_2_2(psum_reg_2_15_sva, pe_0_0_run_cmp_31_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_14_sva <= MUX_v_16_2_2(psum_reg_2_14_sva, pe_0_0_run_cmp_47_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_13_sva <= MUX_v_16_2_2(psum_reg_2_13_sva, pe_0_0_run_cmp_63_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_12_sva <= MUX_v_16_2_2(psum_reg_2_12_sva, pe_0_0_run_cmp_79_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_11_sva <= MUX_v_16_2_2(psum_reg_2_11_sva, pe_0_0_run_cmp_95_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_10_sva <= MUX_v_16_2_2(psum_reg_2_10_sva, pe_0_0_run_cmp_111_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_9_sva <= MUX_v_16_2_2(psum_reg_2_9_sva, pe_0_0_run_cmp_127_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_8_sva <= MUX_v_16_2_2(psum_reg_2_8_sva, pe_0_0_run_cmp_143_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_7_sva <= MUX_v_16_2_2(psum_reg_2_7_sva, pe_0_0_run_cmp_159_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_6_sva <= MUX_v_16_2_2(psum_reg_2_6_sva, pe_0_0_run_cmp_175_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_5_sva <= MUX_v_16_2_2(psum_reg_2_5_sva, pe_0_0_run_cmp_191_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_4_sva <= MUX_v_16_2_2(psum_reg_2_4_sva, pe_0_0_run_cmp_207_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_3_sva <= MUX_v_16_2_2(psum_reg_2_3_sva, pe_0_0_run_cmp_223_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_2_sva <= MUX_v_16_2_2(psum_reg_2_2_sva, pe_0_0_run_cmp_239_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_2_1_sva <= MUX_v_16_2_2(psum_reg_2_1_sva, pe_0_0_run_cmp_255_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_16_sva <= MUX_v_16_2_2(psum_reg_1_16_sva, pe_0_0_run_cmp_16_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_15_sva <= MUX_v_16_2_2(psum_reg_1_15_sva, pe_0_0_run_cmp_32_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_14_sva <= MUX_v_16_2_2(psum_reg_1_14_sva, pe_0_0_run_cmp_48_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_13_sva <= MUX_v_16_2_2(psum_reg_1_13_sva, pe_0_0_run_cmp_64_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_12_sva <= MUX_v_16_2_2(psum_reg_1_12_sva, pe_0_0_run_cmp_80_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_11_sva <= MUX_v_16_2_2(psum_reg_1_11_sva, pe_0_0_run_cmp_96_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_10_sva <= MUX_v_16_2_2(psum_reg_1_10_sva, pe_0_0_run_cmp_112_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_9_sva <= MUX_v_16_2_2(psum_reg_1_9_sva, pe_0_0_run_cmp_128_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_8_sva <= MUX_v_16_2_2(psum_reg_1_8_sva, pe_0_0_run_cmp_144_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_7_sva <= MUX_v_16_2_2(psum_reg_1_7_sva, pe_0_0_run_cmp_160_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_6_sva <= MUX_v_16_2_2(psum_reg_1_6_sva, pe_0_0_run_cmp_176_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_5_sva <= MUX_v_16_2_2(psum_reg_1_5_sva, pe_0_0_run_cmp_192_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_4_sva <= MUX_v_16_2_2(psum_reg_1_4_sva, pe_0_0_run_cmp_208_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_3_sva <= MUX_v_16_2_2(psum_reg_1_3_sva, pe_0_0_run_cmp_224_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_2_sva <= MUX_v_16_2_2(psum_reg_1_2_sva, pe_0_0_run_cmp_240_psum_out_rsc_z,
          and_dcpl_10);
      psum_reg_1_1_sva <= MUX_v_16_2_2(psum_reg_1_1_sva, pe_0_0_run_cmp_psum_out_rsc_z,
          and_dcpl_10);
      input_reg_16_15_sva <= MUX_v_8_2_2(input_reg_16_15_sva, pe_0_0_run_cmp_17_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_14_sva <= MUX_v_8_2_2(input_reg_16_14_sva, pe_0_0_run_cmp_33_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_13_sva <= MUX_v_8_2_2(input_reg_16_13_sva, pe_0_0_run_cmp_49_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_12_sva <= MUX_v_8_2_2(input_reg_16_12_sva, pe_0_0_run_cmp_65_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_11_sva <= MUX_v_8_2_2(input_reg_16_11_sva, pe_0_0_run_cmp_81_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_10_sva <= MUX_v_8_2_2(input_reg_16_10_sva, pe_0_0_run_cmp_97_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_9_sva <= MUX_v_8_2_2(input_reg_16_9_sva, pe_0_0_run_cmp_113_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_8_sva <= MUX_v_8_2_2(input_reg_16_8_sva, pe_0_0_run_cmp_129_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_7_sva <= MUX_v_8_2_2(input_reg_16_7_sva, pe_0_0_run_cmp_145_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_6_sva <= MUX_v_8_2_2(input_reg_16_6_sva, pe_0_0_run_cmp_161_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_5_sva <= MUX_v_8_2_2(input_reg_16_5_sva, pe_0_0_run_cmp_177_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_4_sva <= MUX_v_8_2_2(input_reg_16_4_sva, pe_0_0_run_cmp_193_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_3_sva <= MUX_v_8_2_2(input_reg_16_3_sva, pe_0_0_run_cmp_209_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_2_sva <= MUX_v_8_2_2(input_reg_16_2_sva, pe_0_0_run_cmp_225_input_out_rsc_z,
          and_dcpl_10);
      input_reg_16_1_sva <= MUX_v_8_2_2(input_reg_16_1_sva, pe_0_0_run_cmp_241_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_15_sva <= MUX_v_8_2_2(input_reg_15_15_sva, pe_0_0_run_cmp_18_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_14_sva <= MUX_v_8_2_2(input_reg_15_14_sva, pe_0_0_run_cmp_34_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_13_sva <= MUX_v_8_2_2(input_reg_15_13_sva, pe_0_0_run_cmp_50_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_12_sva <= MUX_v_8_2_2(input_reg_15_12_sva, pe_0_0_run_cmp_66_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_11_sva <= MUX_v_8_2_2(input_reg_15_11_sva, pe_0_0_run_cmp_82_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_10_sva <= MUX_v_8_2_2(input_reg_15_10_sva, pe_0_0_run_cmp_98_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_9_sva <= MUX_v_8_2_2(input_reg_15_9_sva, pe_0_0_run_cmp_114_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_8_sva <= MUX_v_8_2_2(input_reg_15_8_sva, pe_0_0_run_cmp_130_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_7_sva <= MUX_v_8_2_2(input_reg_15_7_sva, pe_0_0_run_cmp_146_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_6_sva <= MUX_v_8_2_2(input_reg_15_6_sva, pe_0_0_run_cmp_162_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_5_sva <= MUX_v_8_2_2(input_reg_15_5_sva, pe_0_0_run_cmp_178_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_4_sva <= MUX_v_8_2_2(input_reg_15_4_sva, pe_0_0_run_cmp_194_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_3_sva <= MUX_v_8_2_2(input_reg_15_3_sva, pe_0_0_run_cmp_210_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_2_sva <= MUX_v_8_2_2(input_reg_15_2_sva, pe_0_0_run_cmp_226_input_out_rsc_z,
          and_dcpl_10);
      input_reg_15_1_sva <= MUX_v_8_2_2(input_reg_15_1_sva, pe_0_0_run_cmp_242_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_15_sva <= MUX_v_8_2_2(input_reg_14_15_sva, pe_0_0_run_cmp_19_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_14_sva <= MUX_v_8_2_2(input_reg_14_14_sva, pe_0_0_run_cmp_35_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_13_sva <= MUX_v_8_2_2(input_reg_14_13_sva, pe_0_0_run_cmp_51_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_12_sva <= MUX_v_8_2_2(input_reg_14_12_sva, pe_0_0_run_cmp_67_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_11_sva <= MUX_v_8_2_2(input_reg_14_11_sva, pe_0_0_run_cmp_83_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_10_sva <= MUX_v_8_2_2(input_reg_14_10_sva, pe_0_0_run_cmp_99_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_9_sva <= MUX_v_8_2_2(input_reg_14_9_sva, pe_0_0_run_cmp_115_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_8_sva <= MUX_v_8_2_2(input_reg_14_8_sva, pe_0_0_run_cmp_131_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_7_sva <= MUX_v_8_2_2(input_reg_14_7_sva, pe_0_0_run_cmp_147_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_6_sva <= MUX_v_8_2_2(input_reg_14_6_sva, pe_0_0_run_cmp_163_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_5_sva <= MUX_v_8_2_2(input_reg_14_5_sva, pe_0_0_run_cmp_179_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_4_sva <= MUX_v_8_2_2(input_reg_14_4_sva, pe_0_0_run_cmp_195_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_3_sva <= MUX_v_8_2_2(input_reg_14_3_sva, pe_0_0_run_cmp_211_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_2_sva <= MUX_v_8_2_2(input_reg_14_2_sva, pe_0_0_run_cmp_227_input_out_rsc_z,
          and_dcpl_10);
      input_reg_14_1_sva <= MUX_v_8_2_2(input_reg_14_1_sva, pe_0_0_run_cmp_243_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_15_sva <= MUX_v_8_2_2(input_reg_13_15_sva, pe_0_0_run_cmp_20_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_14_sva <= MUX_v_8_2_2(input_reg_13_14_sva, pe_0_0_run_cmp_36_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_13_sva <= MUX_v_8_2_2(input_reg_13_13_sva, pe_0_0_run_cmp_52_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_12_sva <= MUX_v_8_2_2(input_reg_13_12_sva, pe_0_0_run_cmp_68_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_11_sva <= MUX_v_8_2_2(input_reg_13_11_sva, pe_0_0_run_cmp_84_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_10_sva <= MUX_v_8_2_2(input_reg_13_10_sva, pe_0_0_run_cmp_100_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_9_sva <= MUX_v_8_2_2(input_reg_13_9_sva, pe_0_0_run_cmp_116_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_8_sva <= MUX_v_8_2_2(input_reg_13_8_sva, pe_0_0_run_cmp_132_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_7_sva <= MUX_v_8_2_2(input_reg_13_7_sva, pe_0_0_run_cmp_148_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_6_sva <= MUX_v_8_2_2(input_reg_13_6_sva, pe_0_0_run_cmp_164_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_5_sva <= MUX_v_8_2_2(input_reg_13_5_sva, pe_0_0_run_cmp_180_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_4_sva <= MUX_v_8_2_2(input_reg_13_4_sva, pe_0_0_run_cmp_196_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_3_sva <= MUX_v_8_2_2(input_reg_13_3_sva, pe_0_0_run_cmp_212_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_2_sva <= MUX_v_8_2_2(input_reg_13_2_sva, pe_0_0_run_cmp_228_input_out_rsc_z,
          and_dcpl_10);
      input_reg_13_1_sva <= MUX_v_8_2_2(input_reg_13_1_sva, pe_0_0_run_cmp_244_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_15_sva <= MUX_v_8_2_2(input_reg_12_15_sva, pe_0_0_run_cmp_21_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_14_sva <= MUX_v_8_2_2(input_reg_12_14_sva, pe_0_0_run_cmp_37_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_13_sva <= MUX_v_8_2_2(input_reg_12_13_sva, pe_0_0_run_cmp_53_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_12_sva <= MUX_v_8_2_2(input_reg_12_12_sva, pe_0_0_run_cmp_69_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_11_sva <= MUX_v_8_2_2(input_reg_12_11_sva, pe_0_0_run_cmp_85_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_10_sva <= MUX_v_8_2_2(input_reg_12_10_sva, pe_0_0_run_cmp_101_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_9_sva <= MUX_v_8_2_2(input_reg_12_9_sva, pe_0_0_run_cmp_117_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_8_sva <= MUX_v_8_2_2(input_reg_12_8_sva, pe_0_0_run_cmp_133_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_7_sva <= MUX_v_8_2_2(input_reg_12_7_sva, pe_0_0_run_cmp_149_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_6_sva <= MUX_v_8_2_2(input_reg_12_6_sva, pe_0_0_run_cmp_165_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_5_sva <= MUX_v_8_2_2(input_reg_12_5_sva, pe_0_0_run_cmp_181_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_4_sva <= MUX_v_8_2_2(input_reg_12_4_sva, pe_0_0_run_cmp_197_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_3_sva <= MUX_v_8_2_2(input_reg_12_3_sva, pe_0_0_run_cmp_213_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_2_sva <= MUX_v_8_2_2(input_reg_12_2_sva, pe_0_0_run_cmp_229_input_out_rsc_z,
          and_dcpl_10);
      input_reg_12_1_sva <= MUX_v_8_2_2(input_reg_12_1_sva, pe_0_0_run_cmp_245_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_15_sva <= MUX_v_8_2_2(input_reg_11_15_sva, pe_0_0_run_cmp_22_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_14_sva <= MUX_v_8_2_2(input_reg_11_14_sva, pe_0_0_run_cmp_38_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_13_sva <= MUX_v_8_2_2(input_reg_11_13_sva, pe_0_0_run_cmp_54_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_12_sva <= MUX_v_8_2_2(input_reg_11_12_sva, pe_0_0_run_cmp_70_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_11_sva <= MUX_v_8_2_2(input_reg_11_11_sva, pe_0_0_run_cmp_86_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_10_sva <= MUX_v_8_2_2(input_reg_11_10_sva, pe_0_0_run_cmp_102_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_9_sva <= MUX_v_8_2_2(input_reg_11_9_sva, pe_0_0_run_cmp_118_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_8_sva <= MUX_v_8_2_2(input_reg_11_8_sva, pe_0_0_run_cmp_134_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_7_sva <= MUX_v_8_2_2(input_reg_11_7_sva, pe_0_0_run_cmp_150_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_6_sva <= MUX_v_8_2_2(input_reg_11_6_sva, pe_0_0_run_cmp_166_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_5_sva <= MUX_v_8_2_2(input_reg_11_5_sva, pe_0_0_run_cmp_182_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_4_sva <= MUX_v_8_2_2(input_reg_11_4_sva, pe_0_0_run_cmp_198_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_3_sva <= MUX_v_8_2_2(input_reg_11_3_sva, pe_0_0_run_cmp_214_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_2_sva <= MUX_v_8_2_2(input_reg_11_2_sva, pe_0_0_run_cmp_230_input_out_rsc_z,
          and_dcpl_10);
      input_reg_11_1_sva <= MUX_v_8_2_2(input_reg_11_1_sva, pe_0_0_run_cmp_246_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_15_sva <= MUX_v_8_2_2(input_reg_10_15_sva, pe_0_0_run_cmp_23_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_14_sva <= MUX_v_8_2_2(input_reg_10_14_sva, pe_0_0_run_cmp_39_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_13_sva <= MUX_v_8_2_2(input_reg_10_13_sva, pe_0_0_run_cmp_55_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_12_sva <= MUX_v_8_2_2(input_reg_10_12_sva, pe_0_0_run_cmp_71_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_11_sva <= MUX_v_8_2_2(input_reg_10_11_sva, pe_0_0_run_cmp_87_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_10_sva <= MUX_v_8_2_2(input_reg_10_10_sva, pe_0_0_run_cmp_103_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_9_sva <= MUX_v_8_2_2(input_reg_10_9_sva, pe_0_0_run_cmp_119_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_8_sva <= MUX_v_8_2_2(input_reg_10_8_sva, pe_0_0_run_cmp_135_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_7_sva <= MUX_v_8_2_2(input_reg_10_7_sva, pe_0_0_run_cmp_151_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_6_sva <= MUX_v_8_2_2(input_reg_10_6_sva, pe_0_0_run_cmp_167_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_5_sva <= MUX_v_8_2_2(input_reg_10_5_sva, pe_0_0_run_cmp_183_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_4_sva <= MUX_v_8_2_2(input_reg_10_4_sva, pe_0_0_run_cmp_199_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_3_sva <= MUX_v_8_2_2(input_reg_10_3_sva, pe_0_0_run_cmp_215_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_2_sva <= MUX_v_8_2_2(input_reg_10_2_sva, pe_0_0_run_cmp_231_input_out_rsc_z,
          and_dcpl_10);
      input_reg_10_1_sva <= MUX_v_8_2_2(input_reg_10_1_sva, pe_0_0_run_cmp_247_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_15_sva <= MUX_v_8_2_2(input_reg_9_15_sva, pe_0_0_run_cmp_24_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_14_sva <= MUX_v_8_2_2(input_reg_9_14_sva, pe_0_0_run_cmp_40_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_13_sva <= MUX_v_8_2_2(input_reg_9_13_sva, pe_0_0_run_cmp_56_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_12_sva <= MUX_v_8_2_2(input_reg_9_12_sva, pe_0_0_run_cmp_72_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_11_sva <= MUX_v_8_2_2(input_reg_9_11_sva, pe_0_0_run_cmp_88_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_10_sva <= MUX_v_8_2_2(input_reg_9_10_sva, pe_0_0_run_cmp_104_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_9_sva <= MUX_v_8_2_2(input_reg_9_9_sva, pe_0_0_run_cmp_120_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_8_sva <= MUX_v_8_2_2(input_reg_9_8_sva, pe_0_0_run_cmp_136_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_7_sva <= MUX_v_8_2_2(input_reg_9_7_sva, pe_0_0_run_cmp_152_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_6_sva <= MUX_v_8_2_2(input_reg_9_6_sva, pe_0_0_run_cmp_168_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_5_sva <= MUX_v_8_2_2(input_reg_9_5_sva, pe_0_0_run_cmp_184_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_4_sva <= MUX_v_8_2_2(input_reg_9_4_sva, pe_0_0_run_cmp_200_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_3_sva <= MUX_v_8_2_2(input_reg_9_3_sva, pe_0_0_run_cmp_216_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_2_sva <= MUX_v_8_2_2(input_reg_9_2_sva, pe_0_0_run_cmp_232_input_out_rsc_z,
          and_dcpl_10);
      input_reg_9_1_sva <= MUX_v_8_2_2(input_reg_9_1_sva, pe_0_0_run_cmp_248_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_15_sva <= MUX_v_8_2_2(input_reg_8_15_sva, pe_0_0_run_cmp_25_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_14_sva <= MUX_v_8_2_2(input_reg_8_14_sva, pe_0_0_run_cmp_41_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_13_sva <= MUX_v_8_2_2(input_reg_8_13_sva, pe_0_0_run_cmp_57_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_12_sva <= MUX_v_8_2_2(input_reg_8_12_sva, pe_0_0_run_cmp_73_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_11_sva <= MUX_v_8_2_2(input_reg_8_11_sva, pe_0_0_run_cmp_89_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_10_sva <= MUX_v_8_2_2(input_reg_8_10_sva, pe_0_0_run_cmp_105_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_9_sva <= MUX_v_8_2_2(input_reg_8_9_sva, pe_0_0_run_cmp_121_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_8_sva <= MUX_v_8_2_2(input_reg_8_8_sva, pe_0_0_run_cmp_137_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_7_sva <= MUX_v_8_2_2(input_reg_8_7_sva, pe_0_0_run_cmp_153_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_6_sva <= MUX_v_8_2_2(input_reg_8_6_sva, pe_0_0_run_cmp_169_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_5_sva <= MUX_v_8_2_2(input_reg_8_5_sva, pe_0_0_run_cmp_185_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_4_sva <= MUX_v_8_2_2(input_reg_8_4_sva, pe_0_0_run_cmp_201_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_3_sva <= MUX_v_8_2_2(input_reg_8_3_sva, pe_0_0_run_cmp_217_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_2_sva <= MUX_v_8_2_2(input_reg_8_2_sva, pe_0_0_run_cmp_233_input_out_rsc_z,
          and_dcpl_10);
      input_reg_8_1_sva <= MUX_v_8_2_2(input_reg_8_1_sva, pe_0_0_run_cmp_249_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_15_sva <= MUX_v_8_2_2(input_reg_7_15_sva, pe_0_0_run_cmp_26_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_14_sva <= MUX_v_8_2_2(input_reg_7_14_sva, pe_0_0_run_cmp_42_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_13_sva <= MUX_v_8_2_2(input_reg_7_13_sva, pe_0_0_run_cmp_58_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_12_sva <= MUX_v_8_2_2(input_reg_7_12_sva, pe_0_0_run_cmp_74_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_11_sva <= MUX_v_8_2_2(input_reg_7_11_sva, pe_0_0_run_cmp_90_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_10_sva <= MUX_v_8_2_2(input_reg_7_10_sva, pe_0_0_run_cmp_106_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_9_sva <= MUX_v_8_2_2(input_reg_7_9_sva, pe_0_0_run_cmp_122_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_8_sva <= MUX_v_8_2_2(input_reg_7_8_sva, pe_0_0_run_cmp_138_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_7_sva <= MUX_v_8_2_2(input_reg_7_7_sva, pe_0_0_run_cmp_154_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_6_sva <= MUX_v_8_2_2(input_reg_7_6_sva, pe_0_0_run_cmp_170_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_5_sva <= MUX_v_8_2_2(input_reg_7_5_sva, pe_0_0_run_cmp_186_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_4_sva <= MUX_v_8_2_2(input_reg_7_4_sva, pe_0_0_run_cmp_202_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_3_sva <= MUX_v_8_2_2(input_reg_7_3_sva, pe_0_0_run_cmp_218_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_2_sva <= MUX_v_8_2_2(input_reg_7_2_sva, pe_0_0_run_cmp_234_input_out_rsc_z,
          and_dcpl_10);
      input_reg_7_1_sva <= MUX_v_8_2_2(input_reg_7_1_sva, pe_0_0_run_cmp_250_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_15_sva <= MUX_v_8_2_2(input_reg_6_15_sva, pe_0_0_run_cmp_27_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_14_sva <= MUX_v_8_2_2(input_reg_6_14_sva, pe_0_0_run_cmp_43_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_13_sva <= MUX_v_8_2_2(input_reg_6_13_sva, pe_0_0_run_cmp_59_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_12_sva <= MUX_v_8_2_2(input_reg_6_12_sva, pe_0_0_run_cmp_75_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_11_sva <= MUX_v_8_2_2(input_reg_6_11_sva, pe_0_0_run_cmp_91_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_10_sva <= MUX_v_8_2_2(input_reg_6_10_sva, pe_0_0_run_cmp_107_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_9_sva <= MUX_v_8_2_2(input_reg_6_9_sva, pe_0_0_run_cmp_123_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_8_sva <= MUX_v_8_2_2(input_reg_6_8_sva, pe_0_0_run_cmp_139_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_7_sva <= MUX_v_8_2_2(input_reg_6_7_sva, pe_0_0_run_cmp_155_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_6_sva <= MUX_v_8_2_2(input_reg_6_6_sva, pe_0_0_run_cmp_171_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_5_sva <= MUX_v_8_2_2(input_reg_6_5_sva, pe_0_0_run_cmp_187_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_4_sva <= MUX_v_8_2_2(input_reg_6_4_sva, pe_0_0_run_cmp_203_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_3_sva <= MUX_v_8_2_2(input_reg_6_3_sva, pe_0_0_run_cmp_219_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_2_sva <= MUX_v_8_2_2(input_reg_6_2_sva, pe_0_0_run_cmp_235_input_out_rsc_z,
          and_dcpl_10);
      input_reg_6_1_sva <= MUX_v_8_2_2(input_reg_6_1_sva, pe_0_0_run_cmp_251_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_15_sva <= MUX_v_8_2_2(input_reg_5_15_sva, pe_0_0_run_cmp_28_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_14_sva <= MUX_v_8_2_2(input_reg_5_14_sva, pe_0_0_run_cmp_44_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_13_sva <= MUX_v_8_2_2(input_reg_5_13_sva, pe_0_0_run_cmp_60_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_12_sva <= MUX_v_8_2_2(input_reg_5_12_sva, pe_0_0_run_cmp_76_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_11_sva <= MUX_v_8_2_2(input_reg_5_11_sva, pe_0_0_run_cmp_92_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_10_sva <= MUX_v_8_2_2(input_reg_5_10_sva, pe_0_0_run_cmp_108_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_9_sva <= MUX_v_8_2_2(input_reg_5_9_sva, pe_0_0_run_cmp_124_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_8_sva <= MUX_v_8_2_2(input_reg_5_8_sva, pe_0_0_run_cmp_140_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_7_sva <= MUX_v_8_2_2(input_reg_5_7_sva, pe_0_0_run_cmp_156_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_6_sva <= MUX_v_8_2_2(input_reg_5_6_sva, pe_0_0_run_cmp_172_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_5_sva <= MUX_v_8_2_2(input_reg_5_5_sva, pe_0_0_run_cmp_188_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_4_sva <= MUX_v_8_2_2(input_reg_5_4_sva, pe_0_0_run_cmp_204_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_3_sva <= MUX_v_8_2_2(input_reg_5_3_sva, pe_0_0_run_cmp_220_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_2_sva <= MUX_v_8_2_2(input_reg_5_2_sva, pe_0_0_run_cmp_236_input_out_rsc_z,
          and_dcpl_10);
      input_reg_5_1_sva <= MUX_v_8_2_2(input_reg_5_1_sva, pe_0_0_run_cmp_252_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_15_sva <= MUX_v_8_2_2(input_reg_4_15_sva, pe_0_0_run_cmp_29_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_14_sva <= MUX_v_8_2_2(input_reg_4_14_sva, pe_0_0_run_cmp_45_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_13_sva <= MUX_v_8_2_2(input_reg_4_13_sva, pe_0_0_run_cmp_61_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_12_sva <= MUX_v_8_2_2(input_reg_4_12_sva, pe_0_0_run_cmp_77_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_11_sva <= MUX_v_8_2_2(input_reg_4_11_sva, pe_0_0_run_cmp_93_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_10_sva <= MUX_v_8_2_2(input_reg_4_10_sva, pe_0_0_run_cmp_109_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_9_sva <= MUX_v_8_2_2(input_reg_4_9_sva, pe_0_0_run_cmp_125_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_8_sva <= MUX_v_8_2_2(input_reg_4_8_sva, pe_0_0_run_cmp_141_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_7_sva <= MUX_v_8_2_2(input_reg_4_7_sva, pe_0_0_run_cmp_157_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_6_sva <= MUX_v_8_2_2(input_reg_4_6_sva, pe_0_0_run_cmp_173_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_5_sva <= MUX_v_8_2_2(input_reg_4_5_sva, pe_0_0_run_cmp_189_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_4_sva <= MUX_v_8_2_2(input_reg_4_4_sva, pe_0_0_run_cmp_205_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_3_sva <= MUX_v_8_2_2(input_reg_4_3_sva, pe_0_0_run_cmp_221_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_2_sva <= MUX_v_8_2_2(input_reg_4_2_sva, pe_0_0_run_cmp_237_input_out_rsc_z,
          and_dcpl_10);
      input_reg_4_1_sva <= MUX_v_8_2_2(input_reg_4_1_sva, pe_0_0_run_cmp_253_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_15_sva <= MUX_v_8_2_2(input_reg_3_15_sva, pe_0_0_run_cmp_30_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_14_sva <= MUX_v_8_2_2(input_reg_3_14_sva, pe_0_0_run_cmp_46_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_13_sva <= MUX_v_8_2_2(input_reg_3_13_sva, pe_0_0_run_cmp_62_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_12_sva <= MUX_v_8_2_2(input_reg_3_12_sva, pe_0_0_run_cmp_78_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_11_sva <= MUX_v_8_2_2(input_reg_3_11_sva, pe_0_0_run_cmp_94_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_10_sva <= MUX_v_8_2_2(input_reg_3_10_sva, pe_0_0_run_cmp_110_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_9_sva <= MUX_v_8_2_2(input_reg_3_9_sva, pe_0_0_run_cmp_126_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_8_sva <= MUX_v_8_2_2(input_reg_3_8_sva, pe_0_0_run_cmp_142_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_7_sva <= MUX_v_8_2_2(input_reg_3_7_sva, pe_0_0_run_cmp_158_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_6_sva <= MUX_v_8_2_2(input_reg_3_6_sva, pe_0_0_run_cmp_174_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_5_sva <= MUX_v_8_2_2(input_reg_3_5_sva, pe_0_0_run_cmp_190_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_4_sva <= MUX_v_8_2_2(input_reg_3_4_sva, pe_0_0_run_cmp_206_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_3_sva <= MUX_v_8_2_2(input_reg_3_3_sva, pe_0_0_run_cmp_222_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_2_sva <= MUX_v_8_2_2(input_reg_3_2_sva, pe_0_0_run_cmp_238_input_out_rsc_z,
          and_dcpl_10);
      input_reg_3_1_sva <= MUX_v_8_2_2(input_reg_3_1_sva, pe_0_0_run_cmp_254_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_15_sva <= MUX_v_8_2_2(input_reg_2_15_sva, pe_0_0_run_cmp_31_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_14_sva <= MUX_v_8_2_2(input_reg_2_14_sva, pe_0_0_run_cmp_47_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_13_sva <= MUX_v_8_2_2(input_reg_2_13_sva, pe_0_0_run_cmp_63_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_12_sva <= MUX_v_8_2_2(input_reg_2_12_sva, pe_0_0_run_cmp_79_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_11_sva <= MUX_v_8_2_2(input_reg_2_11_sva, pe_0_0_run_cmp_95_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_10_sva <= MUX_v_8_2_2(input_reg_2_10_sva, pe_0_0_run_cmp_111_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_9_sva <= MUX_v_8_2_2(input_reg_2_9_sva, pe_0_0_run_cmp_127_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_8_sva <= MUX_v_8_2_2(input_reg_2_8_sva, pe_0_0_run_cmp_143_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_7_sva <= MUX_v_8_2_2(input_reg_2_7_sva, pe_0_0_run_cmp_159_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_6_sva <= MUX_v_8_2_2(input_reg_2_6_sva, pe_0_0_run_cmp_175_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_5_sva <= MUX_v_8_2_2(input_reg_2_5_sva, pe_0_0_run_cmp_191_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_4_sva <= MUX_v_8_2_2(input_reg_2_4_sva, pe_0_0_run_cmp_207_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_3_sva <= MUX_v_8_2_2(input_reg_2_3_sva, pe_0_0_run_cmp_223_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_2_sva <= MUX_v_8_2_2(input_reg_2_2_sva, pe_0_0_run_cmp_239_input_out_rsc_z,
          and_dcpl_10);
      input_reg_2_1_sva <= MUX_v_8_2_2(input_reg_2_1_sva, pe_0_0_run_cmp_255_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_15_sva <= MUX_v_8_2_2(input_reg_1_15_sva, pe_0_0_run_cmp_32_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_14_sva <= MUX_v_8_2_2(input_reg_1_14_sva, pe_0_0_run_cmp_48_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_13_sva <= MUX_v_8_2_2(input_reg_1_13_sva, pe_0_0_run_cmp_64_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_12_sva <= MUX_v_8_2_2(input_reg_1_12_sva, pe_0_0_run_cmp_80_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_11_sva <= MUX_v_8_2_2(input_reg_1_11_sva, pe_0_0_run_cmp_96_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_10_sva <= MUX_v_8_2_2(input_reg_1_10_sva, pe_0_0_run_cmp_112_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_9_sva <= MUX_v_8_2_2(input_reg_1_9_sva, pe_0_0_run_cmp_128_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_8_sva <= MUX_v_8_2_2(input_reg_1_8_sva, pe_0_0_run_cmp_144_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_7_sva <= MUX_v_8_2_2(input_reg_1_7_sva, pe_0_0_run_cmp_160_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_6_sva <= MUX_v_8_2_2(input_reg_1_6_sva, pe_0_0_run_cmp_176_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_5_sva <= MUX_v_8_2_2(input_reg_1_5_sva, pe_0_0_run_cmp_192_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_4_sva <= MUX_v_8_2_2(input_reg_1_4_sva, pe_0_0_run_cmp_208_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_3_sva <= MUX_v_8_2_2(input_reg_1_3_sva, pe_0_0_run_cmp_224_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_2_sva <= MUX_v_8_2_2(input_reg_1_2_sva, pe_0_0_run_cmp_240_input_out_rsc_z,
          and_dcpl_10);
      input_reg_1_1_sva <= MUX_v_8_2_2(input_reg_1_1_sva, pe_0_0_run_cmp_input_out_rsc_z,
          and_dcpl_10);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_if_3_if_step_if_3_if_and_1_itm_3 <= 1'b0;
      step_if_3_for_1_operator_16_false_acc_cse_sva_3 <= 6'b000000;
    end
    else if ( step_if_3_if_and_cse ) begin
      step_if_3_if_step_if_3_if_and_1_itm_3 <= step_if_3_if_step_if_3_if_and_1_itm_2;
      step_if_3_for_1_operator_16_false_acc_cse_sva_3 <= step_if_3_for_1_operator_16_false_acc_cse_sva_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_slc_operator_16_false_acc_16_itm_3 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_1 ) begin
      operator_16_false_slc_operator_16_false_acc_16_itm_3 <= operator_16_false_slc_operator_16_false_acc_16_itm_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_step_not_mdf_sva_3_cse <= 1'b0;
    end
    else if ( run_wen & main_stage_0_3 ) begin
      reg_step_not_mdf_sva_3_cse <= step_not_mdf_sva_st_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_mux_259_itm_1 <= 8'b00000000;
      step_mux_243_itm_1 <= 8'b00000000;
      step_mux_227_itm_1 <= 8'b00000000;
      step_mux_211_itm_1 <= 8'b00000000;
      step_mux_195_itm_1 <= 8'b00000000;
      step_mux_179_itm_1 <= 8'b00000000;
      step_mux_163_itm_1 <= 8'b00000000;
      step_mux_147_itm_1 <= 8'b00000000;
      step_mux_131_itm_1 <= 8'b00000000;
      step_mux_115_itm_1 <= 8'b00000000;
      step_mux_99_itm_1 <= 8'b00000000;
      step_mux_83_itm_1 <= 8'b00000000;
      step_mux_67_itm_1 <= 8'b00000000;
      step_mux_51_itm_1 <= 8'b00000000;
      step_mux_35_itm_1 <= 8'b00000000;
      step_mux_19_itm_1 <= 8'b00000000;
      step_mux_258_itm_1 <= 8'b00000000;
      step_mux_242_itm_1 <= 8'b00000000;
      step_mux_226_itm_1 <= 8'b00000000;
      step_mux_210_itm_1 <= 8'b00000000;
      step_mux_194_itm_1 <= 8'b00000000;
      step_mux_178_itm_1 <= 8'b00000000;
      step_mux_162_itm_1 <= 8'b00000000;
      step_mux_146_itm_1 <= 8'b00000000;
      step_mux_130_itm_1 <= 8'b00000000;
      step_mux_114_itm_1 <= 8'b00000000;
      step_mux_98_itm_1 <= 8'b00000000;
      step_mux_82_itm_1 <= 8'b00000000;
      step_mux_66_itm_1 <= 8'b00000000;
      step_mux_50_itm_1 <= 8'b00000000;
      step_mux_34_itm_1 <= 8'b00000000;
      step_mux_18_itm_1 <= 8'b00000000;
      step_mux_257_itm_1 <= 8'b00000000;
      step_mux_241_itm_1 <= 8'b00000000;
      step_mux_225_itm_1 <= 8'b00000000;
      step_mux_209_itm_1 <= 8'b00000000;
      step_mux_193_itm_1 <= 8'b00000000;
      step_mux_177_itm_1 <= 8'b00000000;
      step_mux_161_itm_1 <= 8'b00000000;
      step_mux_145_itm_1 <= 8'b00000000;
      step_mux_129_itm_1 <= 8'b00000000;
      step_mux_113_itm_1 <= 8'b00000000;
      step_mux_97_itm_1 <= 8'b00000000;
      step_mux_81_itm_1 <= 8'b00000000;
      step_mux_65_itm_1 <= 8'b00000000;
      step_mux_49_itm_1 <= 8'b00000000;
      step_mux_33_itm_1 <= 8'b00000000;
      step_mux_17_itm_1 <= 8'b00000000;
      step_mux_256_itm_1 <= 8'b00000000;
      step_mux_240_itm_1 <= 8'b00000000;
      step_mux_224_itm_1 <= 8'b00000000;
      step_mux_208_itm_1 <= 8'b00000000;
      step_mux_192_itm_1 <= 8'b00000000;
      step_mux_176_itm_1 <= 8'b00000000;
      step_mux_160_itm_1 <= 8'b00000000;
      step_mux_144_itm_1 <= 8'b00000000;
      step_mux_128_itm_1 <= 8'b00000000;
      step_mux_112_itm_1 <= 8'b00000000;
      step_mux_96_itm_1 <= 8'b00000000;
      step_mux_80_itm_1 <= 8'b00000000;
      step_mux_64_itm_1 <= 8'b00000000;
      step_mux_48_itm_1 <= 8'b00000000;
      step_mux_32_itm_1 <= 8'b00000000;
      step_mux_16_itm_1 <= 8'b00000000;
      step_mux_255_itm_1 <= 8'b00000000;
      step_mux_239_itm_1 <= 8'b00000000;
      step_mux_223_itm_1 <= 8'b00000000;
      step_mux_207_itm_1 <= 8'b00000000;
      step_mux_191_itm_1 <= 8'b00000000;
      step_mux_175_itm_1 <= 8'b00000000;
      step_mux_159_itm_1 <= 8'b00000000;
      step_mux_143_itm_1 <= 8'b00000000;
      step_mux_127_itm_1 <= 8'b00000000;
      step_mux_111_itm_1 <= 8'b00000000;
      step_mux_95_itm_1 <= 8'b00000000;
      step_mux_79_itm_1 <= 8'b00000000;
      step_mux_63_itm_1 <= 8'b00000000;
      step_mux_47_itm_1 <= 8'b00000000;
      step_mux_31_itm_1 <= 8'b00000000;
      step_mux_15_itm_1 <= 8'b00000000;
      step_mux_254_itm_1 <= 8'b00000000;
      step_mux_238_itm_1 <= 8'b00000000;
      step_mux_222_itm_1 <= 8'b00000000;
      step_mux_206_itm_1 <= 8'b00000000;
      step_mux_190_itm_1 <= 8'b00000000;
      step_mux_174_itm_1 <= 8'b00000000;
      step_mux_158_itm_1 <= 8'b00000000;
      step_mux_142_itm_1 <= 8'b00000000;
      step_mux_126_itm_1 <= 8'b00000000;
      step_mux_110_itm_1 <= 8'b00000000;
      step_mux_94_itm_1 <= 8'b00000000;
      step_mux_78_itm_1 <= 8'b00000000;
      step_mux_62_itm_1 <= 8'b00000000;
      step_mux_46_itm_1 <= 8'b00000000;
      step_mux_30_itm_1 <= 8'b00000000;
      step_mux_14_itm_1 <= 8'b00000000;
      step_mux_253_itm_1 <= 8'b00000000;
      step_mux_237_itm_1 <= 8'b00000000;
      step_mux_221_itm_1 <= 8'b00000000;
      step_mux_205_itm_1 <= 8'b00000000;
      step_mux_189_itm_1 <= 8'b00000000;
      step_mux_173_itm_1 <= 8'b00000000;
      step_mux_157_itm_1 <= 8'b00000000;
      step_mux_141_itm_1 <= 8'b00000000;
      step_mux_125_itm_1 <= 8'b00000000;
      step_mux_109_itm_1 <= 8'b00000000;
      step_mux_93_itm_1 <= 8'b00000000;
      step_mux_77_itm_1 <= 8'b00000000;
      step_mux_61_itm_1 <= 8'b00000000;
      step_mux_45_itm_1 <= 8'b00000000;
      step_mux_29_itm_1 <= 8'b00000000;
      step_mux_13_itm_1 <= 8'b00000000;
      step_mux_252_itm_1 <= 8'b00000000;
      step_mux_236_itm_1 <= 8'b00000000;
      step_mux_220_itm_1 <= 8'b00000000;
      step_mux_204_itm_1 <= 8'b00000000;
      step_mux_188_itm_1 <= 8'b00000000;
      step_mux_172_itm_1 <= 8'b00000000;
      step_mux_156_itm_1 <= 8'b00000000;
      step_mux_140_itm_1 <= 8'b00000000;
      step_mux_124_itm_1 <= 8'b00000000;
      step_mux_108_itm_1 <= 8'b00000000;
      step_mux_92_itm_1 <= 8'b00000000;
      step_mux_76_itm_1 <= 8'b00000000;
      step_mux_60_itm_1 <= 8'b00000000;
      step_mux_44_itm_1 <= 8'b00000000;
      step_mux_28_itm_1 <= 8'b00000000;
      step_mux_12_itm_1 <= 8'b00000000;
      step_mux_251_itm_1 <= 8'b00000000;
      step_mux_235_itm_1 <= 8'b00000000;
      step_mux_219_itm_1 <= 8'b00000000;
      step_mux_203_itm_1 <= 8'b00000000;
      step_mux_187_itm_1 <= 8'b00000000;
      step_mux_171_itm_1 <= 8'b00000000;
      step_mux_155_itm_1 <= 8'b00000000;
      step_mux_139_itm_1 <= 8'b00000000;
      step_mux_123_itm_1 <= 8'b00000000;
      step_mux_107_itm_1 <= 8'b00000000;
      step_mux_91_itm_1 <= 8'b00000000;
      step_mux_75_itm_1 <= 8'b00000000;
      step_mux_59_itm_1 <= 8'b00000000;
      step_mux_43_itm_1 <= 8'b00000000;
      step_mux_27_itm_1 <= 8'b00000000;
      step_mux_11_itm_1 <= 8'b00000000;
      step_mux_250_itm_1 <= 8'b00000000;
      step_mux_234_itm_1 <= 8'b00000000;
      step_mux_218_itm_1 <= 8'b00000000;
      step_mux_202_itm_1 <= 8'b00000000;
      step_mux_186_itm_1 <= 8'b00000000;
      step_mux_170_itm_1 <= 8'b00000000;
      step_mux_154_itm_1 <= 8'b00000000;
      step_mux_138_itm_1 <= 8'b00000000;
      step_mux_122_itm_1 <= 8'b00000000;
      step_mux_106_itm_1 <= 8'b00000000;
      step_mux_90_itm_1 <= 8'b00000000;
      step_mux_74_itm_1 <= 8'b00000000;
      step_mux_58_itm_1 <= 8'b00000000;
      step_mux_42_itm_1 <= 8'b00000000;
      step_mux_26_itm_1 <= 8'b00000000;
      step_mux_10_itm_1 <= 8'b00000000;
      step_mux_249_itm_1 <= 8'b00000000;
      step_mux_233_itm_1 <= 8'b00000000;
      step_mux_217_itm_1 <= 8'b00000000;
      step_mux_201_itm_1 <= 8'b00000000;
      step_mux_185_itm_1 <= 8'b00000000;
      step_mux_169_itm_1 <= 8'b00000000;
      step_mux_153_itm_1 <= 8'b00000000;
      step_mux_137_itm_1 <= 8'b00000000;
      step_mux_121_itm_1 <= 8'b00000000;
      step_mux_105_itm_1 <= 8'b00000000;
      step_mux_89_itm_1 <= 8'b00000000;
      step_mux_73_itm_1 <= 8'b00000000;
      step_mux_57_itm_1 <= 8'b00000000;
      step_mux_41_itm_1 <= 8'b00000000;
      step_mux_25_itm_1 <= 8'b00000000;
      step_mux_9_itm_1 <= 8'b00000000;
      step_mux_248_itm_1 <= 8'b00000000;
      step_mux_232_itm_1 <= 8'b00000000;
      step_mux_216_itm_1 <= 8'b00000000;
      step_mux_200_itm_1 <= 8'b00000000;
      step_mux_184_itm_1 <= 8'b00000000;
      step_mux_168_itm_1 <= 8'b00000000;
      step_mux_152_itm_1 <= 8'b00000000;
      step_mux_136_itm_1 <= 8'b00000000;
      step_mux_120_itm_1 <= 8'b00000000;
      step_mux_104_itm_1 <= 8'b00000000;
      step_mux_88_itm_1 <= 8'b00000000;
      step_mux_72_itm_1 <= 8'b00000000;
      step_mux_56_itm_1 <= 8'b00000000;
      step_mux_40_itm_1 <= 8'b00000000;
      step_mux_24_itm_1 <= 8'b00000000;
      step_mux_8_itm_1 <= 8'b00000000;
      step_mux_247_itm_1 <= 8'b00000000;
      step_mux_231_itm_1 <= 8'b00000000;
      step_mux_215_itm_1 <= 8'b00000000;
      step_mux_199_itm_1 <= 8'b00000000;
      step_mux_183_itm_1 <= 8'b00000000;
      step_mux_167_itm_1 <= 8'b00000000;
      step_mux_151_itm_1 <= 8'b00000000;
      step_mux_135_itm_1 <= 8'b00000000;
      step_mux_119_itm_1 <= 8'b00000000;
      step_mux_103_itm_1 <= 8'b00000000;
      step_mux_87_itm_1 <= 8'b00000000;
      step_mux_71_itm_1 <= 8'b00000000;
      step_mux_55_itm_1 <= 8'b00000000;
      step_mux_39_itm_1 <= 8'b00000000;
      step_mux_23_itm_1 <= 8'b00000000;
      step_mux_7_itm_1 <= 8'b00000000;
      step_mux_246_itm_1 <= 8'b00000000;
      step_mux_230_itm_1 <= 8'b00000000;
      step_mux_214_itm_1 <= 8'b00000000;
      step_mux_198_itm_1 <= 8'b00000000;
      step_mux_182_itm_1 <= 8'b00000000;
      step_mux_166_itm_1 <= 8'b00000000;
      step_mux_150_itm_1 <= 8'b00000000;
      step_mux_134_itm_1 <= 8'b00000000;
      step_mux_118_itm_1 <= 8'b00000000;
      step_mux_102_itm_1 <= 8'b00000000;
      step_mux_86_itm_1 <= 8'b00000000;
      step_mux_70_itm_1 <= 8'b00000000;
      step_mux_54_itm_1 <= 8'b00000000;
      step_mux_38_itm_1 <= 8'b00000000;
      step_mux_22_itm_1 <= 8'b00000000;
      step_mux_6_itm_1 <= 8'b00000000;
      step_mux_245_itm_1 <= 8'b00000000;
      step_mux_229_itm_1 <= 8'b00000000;
      step_mux_213_itm_1 <= 8'b00000000;
      step_mux_197_itm_1 <= 8'b00000000;
      step_mux_181_itm_1 <= 8'b00000000;
      step_mux_165_itm_1 <= 8'b00000000;
      step_mux_149_itm_1 <= 8'b00000000;
      step_mux_133_itm_1 <= 8'b00000000;
      step_mux_117_itm_1 <= 8'b00000000;
      step_mux_101_itm_1 <= 8'b00000000;
      step_mux_85_itm_1 <= 8'b00000000;
      step_mux_69_itm_1 <= 8'b00000000;
      step_mux_53_itm_1 <= 8'b00000000;
      step_mux_37_itm_1 <= 8'b00000000;
      step_mux_21_itm_1 <= 8'b00000000;
      step_mux_5_itm_1 <= 8'b00000000;
      step_mux_244_itm_1 <= 8'b00000000;
      step_mux_228_itm_1 <= 8'b00000000;
      step_mux_212_itm_1 <= 8'b00000000;
      step_mux_196_itm_1 <= 8'b00000000;
      step_mux_180_itm_1 <= 8'b00000000;
      step_mux_164_itm_1 <= 8'b00000000;
      step_mux_148_itm_1 <= 8'b00000000;
      step_mux_132_itm_1 <= 8'b00000000;
      step_mux_116_itm_1 <= 8'b00000000;
      step_mux_100_itm_1 <= 8'b00000000;
      step_mux_84_itm_1 <= 8'b00000000;
      step_mux_68_itm_1 <= 8'b00000000;
      step_mux_52_itm_1 <= 8'b00000000;
      step_mux_36_itm_1 <= 8'b00000000;
      step_mux_20_itm_1 <= 8'b00000000;
      step_mux_4_itm_1 <= 8'b00000000;
      operator_16_false_slc_operator_16_false_acc_16_itm_2 <= 1'b0;
    end
    else if ( step_and_499_cse ) begin
      step_mux_259_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_15_15_sva,
          or_dcpl_50);
      step_mux_243_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_14_15_sva,
          or_dcpl_52);
      step_mux_227_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_13_15_sva,
          or_dcpl_55);
      step_mux_211_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_12_15_sva,
          or_dcpl_57);
      step_mux_195_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_11_15_sva,
          or_dcpl_59);
      step_mux_179_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_10_15_sva,
          or_dcpl_60);
      step_mux_163_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_9_15_sva,
          or_dcpl_61);
      step_mux_147_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_8_15_sva,
          or_dcpl_62);
      step_mux_131_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_7_15_sva,
          or_dcpl_64);
      step_mux_115_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_6_15_sva,
          or_dcpl_65);
      step_mux_99_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_5_15_sva,
          or_dcpl_66);
      step_mux_83_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_4_15_sva,
          or_dcpl_67);
      step_mux_67_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_3_15_sva,
          or_dcpl_69);
      step_mux_51_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_2_15_sva,
          or_dcpl_70);
      step_mux_35_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_1_15_sva,
          or_dcpl_71);
      step_mux_19_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[127:120]), weight_reg_0_15_sva,
          or_dcpl_72);
      step_mux_258_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_15_14_sva,
          or_dcpl_50);
      step_mux_242_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_14_14_sva,
          or_dcpl_52);
      step_mux_226_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_13_14_sva,
          or_dcpl_55);
      step_mux_210_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_12_14_sva,
          or_dcpl_57);
      step_mux_194_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_11_14_sva,
          or_dcpl_59);
      step_mux_178_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_10_14_sva,
          or_dcpl_60);
      step_mux_162_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_9_14_sva,
          or_dcpl_61);
      step_mux_146_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_8_14_sva,
          or_dcpl_62);
      step_mux_130_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_7_14_sva,
          or_dcpl_64);
      step_mux_114_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_6_14_sva,
          or_dcpl_65);
      step_mux_98_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_5_14_sva,
          or_dcpl_66);
      step_mux_82_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_4_14_sva,
          or_dcpl_67);
      step_mux_66_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_3_14_sva,
          or_dcpl_69);
      step_mux_50_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_2_14_sva,
          or_dcpl_70);
      step_mux_34_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_1_14_sva,
          or_dcpl_71);
      step_mux_18_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[119:112]), weight_reg_0_14_sva,
          or_dcpl_72);
      step_mux_257_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_15_13_sva,
          or_dcpl_50);
      step_mux_241_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_14_13_sva,
          or_dcpl_52);
      step_mux_225_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_13_13_sva,
          or_dcpl_55);
      step_mux_209_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_12_13_sva,
          or_dcpl_57);
      step_mux_193_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_11_13_sva,
          or_dcpl_59);
      step_mux_177_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_10_13_sva,
          or_dcpl_60);
      step_mux_161_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_9_13_sva,
          or_dcpl_61);
      step_mux_145_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_8_13_sva,
          or_dcpl_62);
      step_mux_129_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_7_13_sva,
          or_dcpl_64);
      step_mux_113_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_6_13_sva,
          or_dcpl_65);
      step_mux_97_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_5_13_sva,
          or_dcpl_66);
      step_mux_81_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_4_13_sva,
          or_dcpl_67);
      step_mux_65_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_3_13_sva,
          or_dcpl_69);
      step_mux_49_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_2_13_sva,
          or_dcpl_70);
      step_mux_33_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_1_13_sva,
          or_dcpl_71);
      step_mux_17_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[111:104]), weight_reg_0_13_sva,
          or_dcpl_72);
      step_mux_256_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_15_12_sva,
          or_dcpl_50);
      step_mux_240_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_14_12_sva,
          or_dcpl_52);
      step_mux_224_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_13_12_sva,
          or_dcpl_55);
      step_mux_208_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_12_12_sva,
          or_dcpl_57);
      step_mux_192_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_11_12_sva,
          or_dcpl_59);
      step_mux_176_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_10_12_sva,
          or_dcpl_60);
      step_mux_160_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_9_12_sva,
          or_dcpl_61);
      step_mux_144_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_8_12_sva,
          or_dcpl_62);
      step_mux_128_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_7_12_sva,
          or_dcpl_64);
      step_mux_112_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_6_12_sva,
          or_dcpl_65);
      step_mux_96_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_5_12_sva,
          or_dcpl_66);
      step_mux_80_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_4_12_sva,
          or_dcpl_67);
      step_mux_64_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_3_12_sva,
          or_dcpl_69);
      step_mux_48_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_2_12_sva,
          or_dcpl_70);
      step_mux_32_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_1_12_sva,
          or_dcpl_71);
      step_mux_16_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[103:96]), weight_reg_0_12_sva,
          or_dcpl_72);
      step_mux_255_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_15_11_sva,
          or_dcpl_50);
      step_mux_239_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_14_11_sva,
          or_dcpl_52);
      step_mux_223_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_13_11_sva,
          or_dcpl_55);
      step_mux_207_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_12_11_sva,
          or_dcpl_57);
      step_mux_191_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_11_11_sva,
          or_dcpl_59);
      step_mux_175_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_10_11_sva,
          or_dcpl_60);
      step_mux_159_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_9_11_sva,
          or_dcpl_61);
      step_mux_143_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_8_11_sva,
          or_dcpl_62);
      step_mux_127_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_7_11_sva,
          or_dcpl_64);
      step_mux_111_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_6_11_sva,
          or_dcpl_65);
      step_mux_95_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_5_11_sva,
          or_dcpl_66);
      step_mux_79_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_4_11_sva,
          or_dcpl_67);
      step_mux_63_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_3_11_sva,
          or_dcpl_69);
      step_mux_47_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_2_11_sva,
          or_dcpl_70);
      step_mux_31_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_1_11_sva,
          or_dcpl_71);
      step_mux_15_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[95:88]), weight_reg_0_11_sva,
          or_dcpl_72);
      step_mux_254_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_15_10_sva,
          or_dcpl_50);
      step_mux_238_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_14_10_sva,
          or_dcpl_52);
      step_mux_222_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_13_10_sva,
          or_dcpl_55);
      step_mux_206_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_12_10_sva,
          or_dcpl_57);
      step_mux_190_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_11_10_sva,
          or_dcpl_59);
      step_mux_174_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_10_10_sva,
          or_dcpl_60);
      step_mux_158_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_9_10_sva,
          or_dcpl_61);
      step_mux_142_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_8_10_sva,
          or_dcpl_62);
      step_mux_126_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_7_10_sva,
          or_dcpl_64);
      step_mux_110_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_6_10_sva,
          or_dcpl_65);
      step_mux_94_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_5_10_sva,
          or_dcpl_66);
      step_mux_78_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_4_10_sva,
          or_dcpl_67);
      step_mux_62_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_3_10_sva,
          or_dcpl_69);
      step_mux_46_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_2_10_sva,
          or_dcpl_70);
      step_mux_30_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_1_10_sva,
          or_dcpl_71);
      step_mux_14_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[87:80]), weight_reg_0_10_sva,
          or_dcpl_72);
      step_mux_253_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_15_9_sva,
          or_dcpl_50);
      step_mux_237_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_14_9_sva,
          or_dcpl_52);
      step_mux_221_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_13_9_sva,
          or_dcpl_55);
      step_mux_205_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_12_9_sva,
          or_dcpl_57);
      step_mux_189_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_11_9_sva,
          or_dcpl_59);
      step_mux_173_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_10_9_sva,
          or_dcpl_60);
      step_mux_157_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_9_9_sva,
          or_dcpl_61);
      step_mux_141_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_8_9_sva,
          or_dcpl_62);
      step_mux_125_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_7_9_sva,
          or_dcpl_64);
      step_mux_109_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_6_9_sva,
          or_dcpl_65);
      step_mux_93_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_5_9_sva,
          or_dcpl_66);
      step_mux_77_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_4_9_sva,
          or_dcpl_67);
      step_mux_61_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_3_9_sva,
          or_dcpl_69);
      step_mux_45_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_2_9_sva,
          or_dcpl_70);
      step_mux_29_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_1_9_sva,
          or_dcpl_71);
      step_mux_13_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[79:72]), weight_reg_0_9_sva,
          or_dcpl_72);
      step_mux_252_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_15_8_sva,
          or_dcpl_50);
      step_mux_236_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_14_8_sva,
          or_dcpl_52);
      step_mux_220_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_13_8_sva,
          or_dcpl_55);
      step_mux_204_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_12_8_sva,
          or_dcpl_57);
      step_mux_188_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_11_8_sva,
          or_dcpl_59);
      step_mux_172_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_10_8_sva,
          or_dcpl_60);
      step_mux_156_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_9_8_sva,
          or_dcpl_61);
      step_mux_140_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_8_8_sva,
          or_dcpl_62);
      step_mux_124_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_7_8_sva,
          or_dcpl_64);
      step_mux_108_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_6_8_sva,
          or_dcpl_65);
      step_mux_92_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_5_8_sva,
          or_dcpl_66);
      step_mux_76_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_4_8_sva,
          or_dcpl_67);
      step_mux_60_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_3_8_sva,
          or_dcpl_69);
      step_mux_44_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_2_8_sva,
          or_dcpl_70);
      step_mux_28_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_1_8_sva,
          or_dcpl_71);
      step_mux_12_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[71:64]), weight_reg_0_8_sva,
          or_dcpl_72);
      step_mux_251_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_15_7_sva,
          or_dcpl_50);
      step_mux_235_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_14_7_sva,
          or_dcpl_52);
      step_mux_219_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_13_7_sva,
          or_dcpl_55);
      step_mux_203_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_12_7_sva,
          or_dcpl_57);
      step_mux_187_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_11_7_sva,
          or_dcpl_59);
      step_mux_171_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_10_7_sva,
          or_dcpl_60);
      step_mux_155_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_9_7_sva,
          or_dcpl_61);
      step_mux_139_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_8_7_sva,
          or_dcpl_62);
      step_mux_123_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_7_7_sva,
          or_dcpl_64);
      step_mux_107_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_6_7_sva,
          or_dcpl_65);
      step_mux_91_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_5_7_sva,
          or_dcpl_66);
      step_mux_75_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_4_7_sva,
          or_dcpl_67);
      step_mux_59_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_3_7_sva,
          or_dcpl_69);
      step_mux_43_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_2_7_sva,
          or_dcpl_70);
      step_mux_27_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_1_7_sva,
          or_dcpl_71);
      step_mux_11_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[63:56]), weight_reg_0_7_sva,
          or_dcpl_72);
      step_mux_250_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_15_6_sva,
          or_dcpl_50);
      step_mux_234_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_14_6_sva,
          or_dcpl_52);
      step_mux_218_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_13_6_sva,
          or_dcpl_55);
      step_mux_202_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_12_6_sva,
          or_dcpl_57);
      step_mux_186_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_11_6_sva,
          or_dcpl_59);
      step_mux_170_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_10_6_sva,
          or_dcpl_60);
      step_mux_154_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_9_6_sva,
          or_dcpl_61);
      step_mux_138_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_8_6_sva,
          or_dcpl_62);
      step_mux_122_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_7_6_sva,
          or_dcpl_64);
      step_mux_106_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_6_6_sva,
          or_dcpl_65);
      step_mux_90_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_5_6_sva,
          or_dcpl_66);
      step_mux_74_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_4_6_sva,
          or_dcpl_67);
      step_mux_58_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_3_6_sva,
          or_dcpl_69);
      step_mux_42_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_2_6_sva,
          or_dcpl_70);
      step_mux_26_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_1_6_sva,
          or_dcpl_71);
      step_mux_10_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[55:48]), weight_reg_0_6_sva,
          or_dcpl_72);
      step_mux_249_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_15_5_sva,
          or_dcpl_50);
      step_mux_233_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_14_5_sva,
          or_dcpl_52);
      step_mux_217_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_13_5_sva,
          or_dcpl_55);
      step_mux_201_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_12_5_sva,
          or_dcpl_57);
      step_mux_185_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_11_5_sva,
          or_dcpl_59);
      step_mux_169_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_10_5_sva,
          or_dcpl_60);
      step_mux_153_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_9_5_sva,
          or_dcpl_61);
      step_mux_137_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_8_5_sva,
          or_dcpl_62);
      step_mux_121_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_7_5_sva,
          or_dcpl_64);
      step_mux_105_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_6_5_sva,
          or_dcpl_65);
      step_mux_89_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_5_5_sva,
          or_dcpl_66);
      step_mux_73_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_4_5_sva,
          or_dcpl_67);
      step_mux_57_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_3_5_sva,
          or_dcpl_69);
      step_mux_41_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_2_5_sva,
          or_dcpl_70);
      step_mux_25_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_1_5_sva,
          or_dcpl_71);
      step_mux_9_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[47:40]), weight_reg_0_5_sva,
          or_dcpl_72);
      step_mux_248_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_15_4_sva,
          or_dcpl_50);
      step_mux_232_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_14_4_sva,
          or_dcpl_52);
      step_mux_216_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_13_4_sva,
          or_dcpl_55);
      step_mux_200_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_12_4_sva,
          or_dcpl_57);
      step_mux_184_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_11_4_sva,
          or_dcpl_59);
      step_mux_168_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_10_4_sva,
          or_dcpl_60);
      step_mux_152_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_9_4_sva,
          or_dcpl_61);
      step_mux_136_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_8_4_sva,
          or_dcpl_62);
      step_mux_120_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_7_4_sva,
          or_dcpl_64);
      step_mux_104_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_6_4_sva,
          or_dcpl_65);
      step_mux_88_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_5_4_sva,
          or_dcpl_66);
      step_mux_72_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_4_4_sva,
          or_dcpl_67);
      step_mux_56_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_3_4_sva,
          or_dcpl_69);
      step_mux_40_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_2_4_sva,
          or_dcpl_70);
      step_mux_24_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_1_4_sva,
          or_dcpl_71);
      step_mux_8_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[39:32]), weight_reg_0_4_sva,
          or_dcpl_72);
      step_mux_247_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_15_3_sva,
          or_dcpl_50);
      step_mux_231_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_14_3_sva,
          or_dcpl_52);
      step_mux_215_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_13_3_sva,
          or_dcpl_55);
      step_mux_199_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_12_3_sva,
          or_dcpl_57);
      step_mux_183_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_11_3_sva,
          or_dcpl_59);
      step_mux_167_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_10_3_sva,
          or_dcpl_60);
      step_mux_151_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_9_3_sva,
          or_dcpl_61);
      step_mux_135_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_8_3_sva,
          or_dcpl_62);
      step_mux_119_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_7_3_sva,
          or_dcpl_64);
      step_mux_103_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_6_3_sva,
          or_dcpl_65);
      step_mux_87_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_5_3_sva,
          or_dcpl_66);
      step_mux_71_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_4_3_sva,
          or_dcpl_67);
      step_mux_55_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_3_3_sva,
          or_dcpl_69);
      step_mux_39_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_2_3_sva,
          or_dcpl_70);
      step_mux_23_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_1_3_sva,
          or_dcpl_71);
      step_mux_7_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[31:24]), weight_reg_0_3_sva,
          or_dcpl_72);
      step_mux_246_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_15_2_sva,
          or_dcpl_50);
      step_mux_230_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_14_2_sva,
          or_dcpl_52);
      step_mux_214_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_13_2_sva,
          or_dcpl_55);
      step_mux_198_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_12_2_sva,
          or_dcpl_57);
      step_mux_182_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_11_2_sva,
          or_dcpl_59);
      step_mux_166_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_10_2_sva,
          or_dcpl_60);
      step_mux_150_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_9_2_sva,
          or_dcpl_61);
      step_mux_134_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_8_2_sva,
          or_dcpl_62);
      step_mux_118_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_7_2_sva,
          or_dcpl_64);
      step_mux_102_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_6_2_sva,
          or_dcpl_65);
      step_mux_86_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_5_2_sva,
          or_dcpl_66);
      step_mux_70_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_4_2_sva,
          or_dcpl_67);
      step_mux_54_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_3_2_sva,
          or_dcpl_69);
      step_mux_38_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_2_2_sva,
          or_dcpl_70);
      step_mux_22_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_1_2_sva,
          or_dcpl_71);
      step_mux_6_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[23:16]), weight_reg_0_2_sva,
          or_dcpl_72);
      step_mux_245_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_15_1_sva,
          or_dcpl_50);
      step_mux_229_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_14_1_sva,
          or_dcpl_52);
      step_mux_213_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_13_1_sva,
          or_dcpl_55);
      step_mux_197_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_12_1_sva,
          or_dcpl_57);
      step_mux_181_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_11_1_sva,
          or_dcpl_59);
      step_mux_165_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_10_1_sva,
          or_dcpl_60);
      step_mux_149_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_9_1_sva,
          or_dcpl_61);
      step_mux_133_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_8_1_sva,
          or_dcpl_62);
      step_mux_117_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_7_1_sva,
          or_dcpl_64);
      step_mux_101_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_6_1_sva,
          or_dcpl_65);
      step_mux_85_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_5_1_sva,
          or_dcpl_66);
      step_mux_69_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_4_1_sva,
          or_dcpl_67);
      step_mux_53_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_3_1_sva,
          or_dcpl_69);
      step_mux_37_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_2_1_sva,
          or_dcpl_70);
      step_mux_21_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_1_1_sva,
          or_dcpl_71);
      step_mux_5_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[15:8]), weight_reg_0_1_sva,
          or_dcpl_72);
      step_mux_244_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_15_0_sva,
          or_dcpl_50);
      step_mux_228_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_14_0_sva,
          or_dcpl_52);
      step_mux_212_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_13_0_sva,
          or_dcpl_55);
      step_mux_196_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_12_0_sva,
          or_dcpl_57);
      step_mux_180_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_11_0_sva,
          or_dcpl_59);
      step_mux_164_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_10_0_sva,
          or_dcpl_60);
      step_mux_148_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_9_0_sva,
          or_dcpl_61);
      step_mux_132_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_8_0_sva,
          or_dcpl_62);
      step_mux_116_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_7_0_sva,
          or_dcpl_64);
      step_mux_100_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_6_0_sva,
          or_dcpl_65);
      step_mux_84_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_5_0_sva,
          or_dcpl_66);
      step_mux_68_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_4_0_sva,
          or_dcpl_67);
      step_mux_52_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_3_0_sva,
          or_dcpl_69);
      step_mux_36_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_2_0_sva,
          or_dcpl_70);
      step_mux_20_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_1_0_sva,
          or_dcpl_71);
      step_mux_4_itm_1 <= MUX_v_8_2_2((weight_rsci_idat_mxwt[7:0]), weight_reg_0_0_sva,
          or_dcpl_72);
      operator_16_false_slc_operator_16_false_acc_16_itm_2 <= operator_16_false_slc_operator_16_false_acc_16_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_not_mdf_sva_st_2 <= 1'b0;
    end
    else if ( run_wen & main_stage_0_2 ) begin
      step_not_mdf_sva_st_2 <= step_not_mdf_sva_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_in_col_value_lpi_1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(operator_32_false_acc_itm_31 & step_if_1_acc_itm_32_1))
        ) begin
      step_in_col_value_lpi_1 <= MUX_v_128_2_2(input_rsci_idat_mxwt, step_in_col_value_lpi_1,
          or_73_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_16_false_slc_operator_16_false_acc_12_svs_st_1 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_47 | and_dcpl_18) ) begin
      operator_16_false_slc_operator_16_false_acc_12_svs_st_1 <= MUX_s_1_2_2(operator_16_false_acc_itm_12_1,
          step_and_psp_1, and_dcpl_18);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_crt_lpi_1_dfm <= 48'b000000000000000000000000000000000000000000000000;
      paramsIn_crt_lpi_1_dfm_63_32 <= 32'b00000000000000000000000000000000;
      step_step_lpi_1 <= 16'b0000000000000000;
      step_step_lpi_1_dfm_1_3_0 <= 4'b0000;
      operator_16_false_slc_operator_16_false_acc_16_itm_1 <= 1'b0;
    end
    else if ( and_1562_cse ) begin
      loopIndicesIn_crt_lpi_1_dfm <= loopIndicesIn_crt_lpi_1_dfm_mx0;
      paramsIn_crt_lpi_1_dfm_63_32 <= paramsIn_crt_lpi_1_dfm_63_32_mx0;
      step_step_lpi_1 <= nl_step_step_lpi_1[15:0];
      step_step_lpi_1_dfm_1_3_0 <= step_step_lpi_1_dfm_1[3:0];
      operator_16_false_slc_operator_16_false_acc_16_itm_1 <= operator_16_false_acc_itm_16_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_lpi_1_dfm_127_80 <= 48'b000000000000000000000000000000000000000000000000;
    end
    else if ( operator_32_false_acc_itm_31 & run_wen & exitL_exit_step_sva ) begin
      paramsIn_crt_lpi_1_dfm_127_80 <= paramsIn_crt_lpi_1_dfm_127_80_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_8_15_sva <= 8'b00000000;
      weight_reg_8_14_sva <= 8'b00000000;
      weight_reg_8_13_sva <= 8'b00000000;
      weight_reg_8_12_sva <= 8'b00000000;
      weight_reg_8_11_sva <= 8'b00000000;
      weight_reg_8_10_sva <= 8'b00000000;
      weight_reg_8_9_sva <= 8'b00000000;
      weight_reg_8_8_sva <= 8'b00000000;
      weight_reg_8_7_sva <= 8'b00000000;
      weight_reg_8_6_sva <= 8'b00000000;
      weight_reg_8_5_sva <= 8'b00000000;
      weight_reg_8_4_sva <= 8'b00000000;
      weight_reg_8_3_sva <= 8'b00000000;
      weight_reg_8_2_sva <= 8'b00000000;
      weight_reg_8_1_sva <= 8'b00000000;
      weight_reg_8_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_cse ) begin
      weight_reg_8_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_8_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_8_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_8_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_8_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_8_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_8_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_8_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_8_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_8_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_8_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_8_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_8_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_8_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_8_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_8_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_0_15_sva <= 8'b00000000;
      weight_reg_0_14_sva <= 8'b00000000;
      weight_reg_0_13_sva <= 8'b00000000;
      weight_reg_0_12_sva <= 8'b00000000;
      weight_reg_0_11_sva <= 8'b00000000;
      weight_reg_0_9_sva <= 8'b00000000;
      weight_reg_0_8_sva <= 8'b00000000;
      weight_reg_0_7_sva <= 8'b00000000;
      weight_reg_0_6_sva <= 8'b00000000;
      weight_reg_0_5_sva <= 8'b00000000;
      weight_reg_0_4_sva <= 8'b00000000;
      weight_reg_0_3_sva <= 8'b00000000;
      weight_reg_0_2_sva <= 8'b00000000;
      weight_reg_0_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_1_cse ) begin
      weight_reg_0_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_0_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_0_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_0_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_0_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_0_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_0_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_0_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_0_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_0_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_0_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_0_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_0_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_0_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_0_10_sva <= 8'b00000000;
    end
    else if ( run_wen & or_dcpl_13 & (~((~ (mux_22_nl)) | or_dcpl_74)) ) begin
      weight_reg_0_10_sva <= weight_rsci_idat_mxwt[87:80];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_0_1_sva <= 8'b00000000;
    end
    else if ( run_wen & or_dcpl_13 & (~((~((~((step_step_lpi_1_dfm_1_3_0[1:0]!=2'b00)
        | or_dcpl_68)) | step_not_mdf_sva_st_1)) | or_dcpl_74 | (~ operator_16_false_slc_operator_16_false_acc_12_svs_st_1)))
        ) begin
      weight_reg_0_1_sva <= weight_rsci_idat_mxwt[15:8];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_if_for_and_stg_2_0_sva <= 1'b0;
      step_if_for_and_stg_2_1_sva <= 1'b0;
      step_if_for_and_stg_2_2_sva <= 1'b0;
      step_if_for_and_stg_2_3_sva <= 1'b0;
      step_if_for_and_stg_2_4_sva <= 1'b0;
      step_if_for_and_stg_2_5_sva <= 1'b0;
      step_if_for_and_stg_2_6_sva <= 1'b0;
      step_if_for_and_stg_2_7_sva <= 1'b0;
    end
    else if ( step_if_for_and_20_cse ) begin
      step_if_for_and_stg_2_0_sva <= step_if_for_and_stg_2_0_sva_mx1w0;
      step_if_for_and_stg_2_1_sva <= step_if_for_and_stg_2_1_sva_mx1w0;
      step_if_for_and_stg_2_2_sva <= step_if_for_and_stg_2_2_sva_mx1w0;
      step_if_for_and_stg_2_3_sva <= step_if_for_and_stg_2_3_sva_mx1w0;
      step_if_for_and_stg_2_4_sva <= step_if_for_and_stg_2_4_sva_mx1w0;
      step_if_for_and_stg_2_5_sva <= step_if_for_and_stg_2_5_sva_mx1w0;
      step_if_for_and_stg_2_6_sva <= step_if_for_and_stg_2_6_sva_mx1w0;
      step_if_for_and_stg_2_7_sva <= step_if_for_and_stg_2_7_sva_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_9_15_sva <= 8'b00000000;
      weight_reg_9_14_sva <= 8'b00000000;
      weight_reg_9_13_sva <= 8'b00000000;
      weight_reg_9_12_sva <= 8'b00000000;
      weight_reg_9_11_sva <= 8'b00000000;
      weight_reg_9_10_sva <= 8'b00000000;
      weight_reg_9_9_sva <= 8'b00000000;
      weight_reg_9_8_sva <= 8'b00000000;
      weight_reg_9_7_sva <= 8'b00000000;
      weight_reg_9_6_sva <= 8'b00000000;
      weight_reg_9_5_sva <= 8'b00000000;
      weight_reg_9_4_sva <= 8'b00000000;
      weight_reg_9_3_sva <= 8'b00000000;
      weight_reg_9_2_sva <= 8'b00000000;
      weight_reg_9_1_sva <= 8'b00000000;
      weight_reg_9_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_32_cse ) begin
      weight_reg_9_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_9_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_9_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_9_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_9_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_9_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_9_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_9_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_9_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_9_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_9_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_9_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_9_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_9_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_9_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_9_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_1_15_sva <= 8'b00000000;
      weight_reg_1_14_sva <= 8'b00000000;
      weight_reg_1_13_sva <= 8'b00000000;
      weight_reg_1_12_sva <= 8'b00000000;
      weight_reg_1_11_sva <= 8'b00000000;
      weight_reg_1_10_sva <= 8'b00000000;
      weight_reg_1_9_sva <= 8'b00000000;
      weight_reg_1_8_sva <= 8'b00000000;
      weight_reg_1_7_sva <= 8'b00000000;
      weight_reg_1_6_sva <= 8'b00000000;
      weight_reg_1_5_sva <= 8'b00000000;
      weight_reg_1_4_sva <= 8'b00000000;
      weight_reg_1_3_sva <= 8'b00000000;
      weight_reg_1_2_sva <= 8'b00000000;
      weight_reg_1_1_sva <= 8'b00000000;
      weight_reg_1_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_33_cse ) begin
      weight_reg_1_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_1_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_1_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_1_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_1_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_1_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_1_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_1_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_1_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_1_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_1_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_1_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_1_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_1_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_1_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_1_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_10_15_sva <= 8'b00000000;
      weight_reg_10_14_sva <= 8'b00000000;
      weight_reg_10_13_sva <= 8'b00000000;
      weight_reg_10_12_sva <= 8'b00000000;
      weight_reg_10_11_sva <= 8'b00000000;
      weight_reg_10_10_sva <= 8'b00000000;
      weight_reg_10_9_sva <= 8'b00000000;
      weight_reg_10_8_sva <= 8'b00000000;
      weight_reg_10_7_sva <= 8'b00000000;
      weight_reg_10_6_sva <= 8'b00000000;
      weight_reg_10_5_sva <= 8'b00000000;
      weight_reg_10_4_sva <= 8'b00000000;
      weight_reg_10_3_sva <= 8'b00000000;
      weight_reg_10_2_sva <= 8'b00000000;
      weight_reg_10_1_sva <= 8'b00000000;
      weight_reg_10_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_64_cse ) begin
      weight_reg_10_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_10_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_10_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_10_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_10_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_10_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_10_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_10_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_10_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_10_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_10_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_10_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_10_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_10_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_10_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_10_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_2_15_sva <= 8'b00000000;
      weight_reg_2_14_sva <= 8'b00000000;
      weight_reg_2_13_sva <= 8'b00000000;
      weight_reg_2_12_sva <= 8'b00000000;
      weight_reg_2_11_sva <= 8'b00000000;
      weight_reg_2_10_sva <= 8'b00000000;
      weight_reg_2_9_sva <= 8'b00000000;
      weight_reg_2_8_sva <= 8'b00000000;
      weight_reg_2_7_sva <= 8'b00000000;
      weight_reg_2_6_sva <= 8'b00000000;
      weight_reg_2_5_sva <= 8'b00000000;
      weight_reg_2_4_sva <= 8'b00000000;
      weight_reg_2_3_sva <= 8'b00000000;
      weight_reg_2_2_sva <= 8'b00000000;
      weight_reg_2_1_sva <= 8'b00000000;
      weight_reg_2_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_65_cse ) begin
      weight_reg_2_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_2_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_2_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_2_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_2_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_2_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_2_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_2_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_2_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_2_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_2_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_2_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_2_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_2_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_2_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_2_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_11_15_sva <= 8'b00000000;
      weight_reg_11_14_sva <= 8'b00000000;
      weight_reg_11_13_sva <= 8'b00000000;
      weight_reg_11_12_sva <= 8'b00000000;
      weight_reg_11_11_sva <= 8'b00000000;
      weight_reg_11_10_sva <= 8'b00000000;
      weight_reg_11_9_sva <= 8'b00000000;
      weight_reg_11_8_sva <= 8'b00000000;
      weight_reg_11_7_sva <= 8'b00000000;
      weight_reg_11_6_sva <= 8'b00000000;
      weight_reg_11_5_sva <= 8'b00000000;
      weight_reg_11_4_sva <= 8'b00000000;
      weight_reg_11_3_sva <= 8'b00000000;
      weight_reg_11_2_sva <= 8'b00000000;
      weight_reg_11_1_sva <= 8'b00000000;
      weight_reg_11_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_96_cse ) begin
      weight_reg_11_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_11_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_11_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_11_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_11_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_11_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_11_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_11_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_11_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_11_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_11_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_11_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_11_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_11_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_11_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_11_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_3_15_sva <= 8'b00000000;
      weight_reg_3_14_sva <= 8'b00000000;
      weight_reg_3_13_sva <= 8'b00000000;
      weight_reg_3_12_sva <= 8'b00000000;
      weight_reg_3_11_sva <= 8'b00000000;
      weight_reg_3_10_sva <= 8'b00000000;
      weight_reg_3_9_sva <= 8'b00000000;
      weight_reg_3_8_sva <= 8'b00000000;
      weight_reg_3_7_sva <= 8'b00000000;
      weight_reg_3_6_sva <= 8'b00000000;
      weight_reg_3_5_sva <= 8'b00000000;
      weight_reg_3_4_sva <= 8'b00000000;
      weight_reg_3_3_sva <= 8'b00000000;
      weight_reg_3_2_sva <= 8'b00000000;
      weight_reg_3_1_sva <= 8'b00000000;
      weight_reg_3_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_97_cse ) begin
      weight_reg_3_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_3_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_3_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_3_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_3_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_3_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_3_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_3_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_3_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_3_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_3_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_3_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_3_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_3_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_3_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_3_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_12_15_sva <= 8'b00000000;
      weight_reg_12_14_sva <= 8'b00000000;
      weight_reg_12_13_sva <= 8'b00000000;
      weight_reg_12_12_sva <= 8'b00000000;
      weight_reg_12_11_sva <= 8'b00000000;
      weight_reg_12_10_sva <= 8'b00000000;
      weight_reg_12_9_sva <= 8'b00000000;
      weight_reg_12_8_sva <= 8'b00000000;
      weight_reg_12_7_sva <= 8'b00000000;
      weight_reg_12_6_sva <= 8'b00000000;
      weight_reg_12_5_sva <= 8'b00000000;
      weight_reg_12_4_sva <= 8'b00000000;
      weight_reg_12_3_sva <= 8'b00000000;
      weight_reg_12_2_sva <= 8'b00000000;
      weight_reg_12_1_sva <= 8'b00000000;
      weight_reg_12_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_128_cse ) begin
      weight_reg_12_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_12_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_12_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_12_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_12_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_12_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_12_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_12_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_12_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_12_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_12_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_12_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_12_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_12_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_12_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_12_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_4_15_sva <= 8'b00000000;
      weight_reg_4_14_sva <= 8'b00000000;
      weight_reg_4_13_sva <= 8'b00000000;
      weight_reg_4_12_sva <= 8'b00000000;
      weight_reg_4_11_sva <= 8'b00000000;
      weight_reg_4_10_sva <= 8'b00000000;
      weight_reg_4_9_sva <= 8'b00000000;
      weight_reg_4_8_sva <= 8'b00000000;
      weight_reg_4_7_sva <= 8'b00000000;
      weight_reg_4_6_sva <= 8'b00000000;
      weight_reg_4_5_sva <= 8'b00000000;
      weight_reg_4_4_sva <= 8'b00000000;
      weight_reg_4_3_sva <= 8'b00000000;
      weight_reg_4_2_sva <= 8'b00000000;
      weight_reg_4_1_sva <= 8'b00000000;
      weight_reg_4_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_129_cse ) begin
      weight_reg_4_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_4_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_4_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_4_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_4_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_4_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_4_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_4_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_4_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_4_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_4_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_4_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_4_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_4_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_4_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_4_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_13_15_sva <= 8'b00000000;
      weight_reg_13_14_sva <= 8'b00000000;
      weight_reg_13_13_sva <= 8'b00000000;
      weight_reg_13_12_sva <= 8'b00000000;
      weight_reg_13_11_sva <= 8'b00000000;
      weight_reg_13_10_sva <= 8'b00000000;
      weight_reg_13_9_sva <= 8'b00000000;
      weight_reg_13_8_sva <= 8'b00000000;
      weight_reg_13_7_sva <= 8'b00000000;
      weight_reg_13_6_sva <= 8'b00000000;
      weight_reg_13_5_sva <= 8'b00000000;
      weight_reg_13_4_sva <= 8'b00000000;
      weight_reg_13_3_sva <= 8'b00000000;
      weight_reg_13_2_sva <= 8'b00000000;
      weight_reg_13_1_sva <= 8'b00000000;
      weight_reg_13_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_160_cse ) begin
      weight_reg_13_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_13_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_13_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_13_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_13_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_13_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_13_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_13_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_13_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_13_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_13_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_13_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_13_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_13_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_13_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_13_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_5_15_sva <= 8'b00000000;
      weight_reg_5_14_sva <= 8'b00000000;
      weight_reg_5_13_sva <= 8'b00000000;
      weight_reg_5_12_sva <= 8'b00000000;
      weight_reg_5_11_sva <= 8'b00000000;
      weight_reg_5_10_sva <= 8'b00000000;
      weight_reg_5_9_sva <= 8'b00000000;
      weight_reg_5_8_sva <= 8'b00000000;
      weight_reg_5_7_sva <= 8'b00000000;
      weight_reg_5_6_sva <= 8'b00000000;
      weight_reg_5_5_sva <= 8'b00000000;
      weight_reg_5_4_sva <= 8'b00000000;
      weight_reg_5_3_sva <= 8'b00000000;
      weight_reg_5_2_sva <= 8'b00000000;
      weight_reg_5_1_sva <= 8'b00000000;
      weight_reg_5_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_161_cse ) begin
      weight_reg_5_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_5_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_5_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_5_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_5_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_5_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_5_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_5_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_5_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_5_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_5_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_5_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_5_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_5_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_5_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_5_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_14_15_sva <= 8'b00000000;
      weight_reg_14_14_sva <= 8'b00000000;
      weight_reg_14_13_sva <= 8'b00000000;
      weight_reg_14_12_sva <= 8'b00000000;
      weight_reg_14_11_sva <= 8'b00000000;
      weight_reg_14_10_sva <= 8'b00000000;
      weight_reg_14_9_sva <= 8'b00000000;
      weight_reg_14_8_sva <= 8'b00000000;
      weight_reg_14_7_sva <= 8'b00000000;
      weight_reg_14_6_sva <= 8'b00000000;
      weight_reg_14_5_sva <= 8'b00000000;
      weight_reg_14_4_sva <= 8'b00000000;
      weight_reg_14_3_sva <= 8'b00000000;
      weight_reg_14_2_sva <= 8'b00000000;
      weight_reg_14_1_sva <= 8'b00000000;
      weight_reg_14_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_192_cse ) begin
      weight_reg_14_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_14_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_14_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_14_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_14_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_14_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_14_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_14_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_14_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_14_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_14_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_14_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_14_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_14_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_14_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_14_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_6_15_sva <= 8'b00000000;
      weight_reg_6_14_sva <= 8'b00000000;
      weight_reg_6_13_sva <= 8'b00000000;
      weight_reg_6_12_sva <= 8'b00000000;
      weight_reg_6_11_sva <= 8'b00000000;
      weight_reg_6_10_sva <= 8'b00000000;
      weight_reg_6_9_sva <= 8'b00000000;
      weight_reg_6_8_sva <= 8'b00000000;
      weight_reg_6_7_sva <= 8'b00000000;
      weight_reg_6_6_sva <= 8'b00000000;
      weight_reg_6_5_sva <= 8'b00000000;
      weight_reg_6_3_sva <= 8'b00000000;
      weight_reg_6_2_sva <= 8'b00000000;
      weight_reg_6_1_sva <= 8'b00000000;
      weight_reg_6_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_193_cse ) begin
      weight_reg_6_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_6_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_6_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_6_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_6_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_6_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_6_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_6_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_6_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_6_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_6_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_6_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_6_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_6_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_6_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_6_4_sva <= 8'b00000000;
    end
    else if ( run_wen & or_dcpl_36 & (~((~ (mux_225_nl)) | or_dcpl_74)) ) begin
      weight_reg_6_4_sva <= weight_rsci_idat_mxwt[39:32];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_15_15_sva <= 8'b00000000;
      weight_reg_15_14_sva <= 8'b00000000;
      weight_reg_15_13_sva <= 8'b00000000;
      weight_reg_15_12_sva <= 8'b00000000;
      weight_reg_15_11_sva <= 8'b00000000;
      weight_reg_15_10_sva <= 8'b00000000;
      weight_reg_15_9_sva <= 8'b00000000;
      weight_reg_15_8_sva <= 8'b00000000;
      weight_reg_15_7_sva <= 8'b00000000;
      weight_reg_15_6_sva <= 8'b00000000;
      weight_reg_15_5_sva <= 8'b00000000;
      weight_reg_15_4_sva <= 8'b00000000;
      weight_reg_15_3_sva <= 8'b00000000;
      weight_reg_15_2_sva <= 8'b00000000;
      weight_reg_15_1_sva <= 8'b00000000;
      weight_reg_15_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_224_cse ) begin
      weight_reg_15_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_15_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_15_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_15_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_15_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_15_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_15_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_15_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_15_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_15_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_15_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_15_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_15_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_15_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_15_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_15_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weight_reg_7_15_sva <= 8'b00000000;
      weight_reg_7_14_sva <= 8'b00000000;
      weight_reg_7_13_sva <= 8'b00000000;
      weight_reg_7_12_sva <= 8'b00000000;
      weight_reg_7_11_sva <= 8'b00000000;
      weight_reg_7_10_sva <= 8'b00000000;
      weight_reg_7_9_sva <= 8'b00000000;
      weight_reg_7_8_sva <= 8'b00000000;
      weight_reg_7_7_sva <= 8'b00000000;
      weight_reg_7_6_sva <= 8'b00000000;
      weight_reg_7_5_sva <= 8'b00000000;
      weight_reg_7_4_sva <= 8'b00000000;
      weight_reg_7_3_sva <= 8'b00000000;
      weight_reg_7_2_sva <= 8'b00000000;
      weight_reg_7_1_sva <= 8'b00000000;
      weight_reg_7_0_sva <= 8'b00000000;
    end
    else if ( weight_reg_and_225_cse ) begin
      weight_reg_7_15_sva <= weight_rsci_idat_mxwt[127:120];
      weight_reg_7_14_sva <= weight_rsci_idat_mxwt[119:112];
      weight_reg_7_13_sva <= weight_rsci_idat_mxwt[111:104];
      weight_reg_7_12_sva <= weight_rsci_idat_mxwt[103:96];
      weight_reg_7_11_sva <= weight_rsci_idat_mxwt[95:88];
      weight_reg_7_10_sva <= weight_rsci_idat_mxwt[87:80];
      weight_reg_7_9_sva <= weight_rsci_idat_mxwt[79:72];
      weight_reg_7_8_sva <= weight_rsci_idat_mxwt[71:64];
      weight_reg_7_7_sva <= weight_rsci_idat_mxwt[63:56];
      weight_reg_7_6_sva <= weight_rsci_idat_mxwt[55:48];
      weight_reg_7_5_sva <= weight_rsci_idat_mxwt[47:40];
      weight_reg_7_4_sva <= weight_rsci_idat_mxwt[39:32];
      weight_reg_7_3_sva <= weight_rsci_idat_mxwt[31:24];
      weight_reg_7_2_sva <= weight_rsci_idat_mxwt[23:16];
      weight_reg_7_1_sva <= weight_rsci_idat_mxwt[15:8];
      weight_reg_7_0_sva <= weight_rsci_idat_mxwt[7:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_if_3_if_step_if_3_if_and_1_itm_2 <= 1'b0;
      step_if_3_for_1_operator_16_false_acc_cse_sva_2 <= 6'b000000;
    end
    else if ( step_if_3_if_and_1_cse ) begin
      step_if_3_if_step_if_3_if_and_1_itm_2 <= step_and_100_psp;
      step_if_3_for_1_operator_16_false_acc_cse_sva_2 <= step_if_3_for_1_operator_16_false_acc_cse_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_and_240_psp <= 1'b0;
      step_and_224_psp <= 1'b0;
      step_and_208_psp <= 1'b0;
      step_and_192_psp <= 1'b0;
      step_and_176_psp <= 1'b0;
      step_and_160_psp <= 1'b0;
      step_and_144_psp <= 1'b0;
      step_and_128_psp <= 1'b0;
      step_and_112_psp <= 1'b0;
      step_and_96_psp <= 1'b0;
      step_and_80_psp <= 1'b0;
      step_and_64_psp <= 1'b0;
      step_and_48_psp <= 1'b0;
      step_and_32_psp <= 1'b0;
      step_and_16_psp <= 1'b0;
      step_and_psp <= 1'b0;
    end
    else if ( step_and_757_cse ) begin
      step_and_240_psp <= step_if_for_and_stg_2_7_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_224_psp <= step_if_for_and_stg_2_6_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_208_psp <= step_if_for_and_stg_2_5_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_192_psp <= step_if_for_and_stg_2_4_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_176_psp <= step_if_for_and_stg_2_3_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_160_psp <= step_if_for_and_stg_2_2_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_144_psp <= step_if_for_and_stg_2_1_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_128_psp <= step_if_for_and_stg_2_0_sva_mx1 & (step_step_lpi_1_dfm_1_3_0[3])
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_112_psp <= step_if_for_and_stg_2_7_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_96_psp <= step_and_96_psp_1;
      step_and_80_psp <= step_if_for_and_stg_2_5_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_64_psp <= step_if_for_and_stg_2_4_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_48_psp <= step_if_for_and_stg_2_3_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_32_psp <= step_if_for_and_stg_2_2_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_16_psp <= step_if_for_and_stg_2_1_sva_mx1 & (~ (step_step_lpi_1_dfm_1_3_0[3]))
          & operator_16_false_slc_operator_16_false_acc_12_svs_st_1;
      step_and_psp <= step_and_psp_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_and_100_psp <= 1'b0;
    end
    else if ( step_and_241_cse & (~(operator_32_false_acc_itm_31 & operator_16_false_acc_itm_16_1))
        & (and_dcpl_18 | operator_32_false_acc_itm_31) ) begin
      step_and_100_psp <= MUX_s_1_2_2(step_and_96_psp_1, (step_if_3_if_step_if_3_if_and_1_nl),
          operator_32_false_acc_itm_31);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_and_10_psp <= 1'b0;
    end
    else if ( step_and_241_cse & ((~ operator_32_false_acc_itm_31) | step_if_1_acc_itm_32_1)
        ) begin
      step_and_10_psp <= MUX1HOT_s_1_3_2(step_and_psp_1, step_if_2_if_step_if_2_if_nor_1_tmp,
          step_and_10_psp, {and_dcpl_18 , operator_32_false_acc_itm_31 , (and_19_nl)});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_if_1_acc_cse_32 <= 1'b0;
    end
    else if ( run_wen & (~((~ operator_32_false_acc_itm_31) | (fsm_output[0]))) )
        begin
      step_if_1_acc_cse_32 <= step_if_1_acc_itm_32_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      step_if_3_for_1_operator_16_false_acc_cse_sva_1 <= 6'b000000;
    end
    else if ( run_wen & operator_32_false_acc_itm_31 & (~ operator_16_false_acc_itm_16_1)
        ) begin
      step_if_3_for_1_operator_16_false_acc_cse_sva_1 <= nl_step_if_3_for_1_operator_16_false_acc_cse_sva_1[5:0];
    end
  end
  assign or_73_nl = step_not_mdf_sva_st_1 | (~ step_if_1_acc_cse_32);
  assign nl_step_step_lpi_1  = step_step_lpi_1_dfm_1 + 16'b0000000000000001;
  assign mux_22_nl = MUX_s_1_2_2(not_tmp_36, or_tmp_3, step_and_10_psp);
  assign mux_225_nl = MUX_s_1_2_2(not_tmp_251, or_tmp_39, step_and_100_psp);
  assign step_if_3_if_step_if_3_if_and_1_nl = (~(((loopIndicesIn_crt_lpi_1_dfm_mx0[47:32])
      != (operator_16_false_3_acc_psp_sva_1[15:0])) | (operator_16_false_3_acc_psp_sva_1[16])))
      & (~(((loopIndicesIn_crt_lpi_1_dfm_mx0[31:16]) != (operator_16_false_2_acc_psp_sva_1[15:0]))
      | (operator_16_false_2_acc_psp_sva_1[16]))) & (~(((loopIndicesIn_crt_lpi_1_dfm_mx0[15:0])
      != (operator_16_false_1_acc_psp_sva_1[15:0])) | (operator_16_false_1_acc_psp_sva_1[16])));
  assign and_19_nl = or_dcpl_74 & (~ operator_32_false_acc_itm_31);
  assign nl_step_if_3_for_1_operator_16_false_acc_cse_sva_1  = (step_step_lpi_1_dfm_1[5:0])
      + 6'b100001;

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [47:0] MUX_v_48_2_2;
    input [47:0] input_0;
    input [47:0] input_1;
    input [0:0] sel;
    reg [47:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_48_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_32_1_31;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_32_1_31 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [16:0] conv_u2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2s_16_17 =  {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_16_33 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_33 = {{17{1'b0}}, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct (
  clk, arst_n, input_rsc_dat_value, input_rsc_vld, input_rsc_rdy, weight_rsc_dat_value,
      weight_rsc_vld, weight_rsc_rdy, output_rsc_dat_value, output_rsc_vld, output_rsc_rdy,
      paramsIn_rsc_dat_STRIDE, paramsIn_rsc_dat_FY, paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1,
      paramsIn_rsc_dat_OC1, paramsIn_rsc_dat_OX0, paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1,
      paramsIn_rsc_dat_OY1, paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat_fy_idx,
      loopIndicesIn_rsc_dat_fx_idx, loopIndicesIn_rsc_dat_ic1_idx, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat_value;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat_value;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat_value;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] loopIndicesIn_rsc_dat_fy_idx;
  input [15:0] loopIndicesIn_rsc_dat_fx_idx;
  input [15:0] loopIndicesIn_rsc_dat_ic1_idx;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;


  // Interconnect Declarations
  wire [7:0] accumulation_buffer_rsc_0_0_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_0_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_0_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_0_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_1_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_1_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_1_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_1_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_2_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_2_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_2_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_2_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_3_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_3_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_3_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_3_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_4_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_4_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_4_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_4_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_5_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_5_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_5_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_5_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_6_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_6_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_6_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_6_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_7_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_7_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_7_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_7_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_8_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_8_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_8_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_8_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_9_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_9_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_9_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_9_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_10_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_10_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_10_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_10_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_11_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_11_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_11_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_11_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_12_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_12_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_12_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_12_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_13_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_13_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_13_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_13_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_14_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_14_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_14_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_14_i_q_d;
  wire [7:0] accumulation_buffer_rsc_0_15_i_radr_d;
  wire [7:0] accumulation_buffer_rsc_0_15_i_wadr_d;
  wire [15:0] accumulation_buffer_rsc_0_15_i_d_d;
  wire [15:0] accumulation_buffer_rsc_0_15_i_q_d;
  wire accumulation_buffer_rsc_0_0_we;
  wire [15:0] accumulation_buffer_rsc_0_0_d;
  wire [7:0] accumulation_buffer_rsc_0_0_wadr;
  wire [15:0] accumulation_buffer_rsc_0_0_q;
  wire accumulation_buffer_rsc_0_0_re;
  wire [7:0] accumulation_buffer_rsc_0_0_radr;
  wire accumulation_buffer_rsc_0_1_we;
  wire [15:0] accumulation_buffer_rsc_0_1_d;
  wire [7:0] accumulation_buffer_rsc_0_1_wadr;
  wire [15:0] accumulation_buffer_rsc_0_1_q;
  wire accumulation_buffer_rsc_0_1_re;
  wire [7:0] accumulation_buffer_rsc_0_1_radr;
  wire accumulation_buffer_rsc_0_2_we;
  wire [15:0] accumulation_buffer_rsc_0_2_d;
  wire [7:0] accumulation_buffer_rsc_0_2_wadr;
  wire [15:0] accumulation_buffer_rsc_0_2_q;
  wire accumulation_buffer_rsc_0_2_re;
  wire [7:0] accumulation_buffer_rsc_0_2_radr;
  wire accumulation_buffer_rsc_0_3_we;
  wire [15:0] accumulation_buffer_rsc_0_3_d;
  wire [7:0] accumulation_buffer_rsc_0_3_wadr;
  wire [15:0] accumulation_buffer_rsc_0_3_q;
  wire accumulation_buffer_rsc_0_3_re;
  wire [7:0] accumulation_buffer_rsc_0_3_radr;
  wire accumulation_buffer_rsc_0_4_we;
  wire [15:0] accumulation_buffer_rsc_0_4_d;
  wire [7:0] accumulation_buffer_rsc_0_4_wadr;
  wire [15:0] accumulation_buffer_rsc_0_4_q;
  wire accumulation_buffer_rsc_0_4_re;
  wire [7:0] accumulation_buffer_rsc_0_4_radr;
  wire accumulation_buffer_rsc_0_5_we;
  wire [15:0] accumulation_buffer_rsc_0_5_d;
  wire [7:0] accumulation_buffer_rsc_0_5_wadr;
  wire [15:0] accumulation_buffer_rsc_0_5_q;
  wire accumulation_buffer_rsc_0_5_re;
  wire [7:0] accumulation_buffer_rsc_0_5_radr;
  wire accumulation_buffer_rsc_0_6_we;
  wire [15:0] accumulation_buffer_rsc_0_6_d;
  wire [7:0] accumulation_buffer_rsc_0_6_wadr;
  wire [15:0] accumulation_buffer_rsc_0_6_q;
  wire accumulation_buffer_rsc_0_6_re;
  wire [7:0] accumulation_buffer_rsc_0_6_radr;
  wire accumulation_buffer_rsc_0_7_we;
  wire [15:0] accumulation_buffer_rsc_0_7_d;
  wire [7:0] accumulation_buffer_rsc_0_7_wadr;
  wire [15:0] accumulation_buffer_rsc_0_7_q;
  wire accumulation_buffer_rsc_0_7_re;
  wire [7:0] accumulation_buffer_rsc_0_7_radr;
  wire accumulation_buffer_rsc_0_8_we;
  wire [15:0] accumulation_buffer_rsc_0_8_d;
  wire [7:0] accumulation_buffer_rsc_0_8_wadr;
  wire [15:0] accumulation_buffer_rsc_0_8_q;
  wire accumulation_buffer_rsc_0_8_re;
  wire [7:0] accumulation_buffer_rsc_0_8_radr;
  wire accumulation_buffer_rsc_0_9_we;
  wire [15:0] accumulation_buffer_rsc_0_9_d;
  wire [7:0] accumulation_buffer_rsc_0_9_wadr;
  wire [15:0] accumulation_buffer_rsc_0_9_q;
  wire accumulation_buffer_rsc_0_9_re;
  wire [7:0] accumulation_buffer_rsc_0_9_radr;
  wire accumulation_buffer_rsc_0_10_we;
  wire [15:0] accumulation_buffer_rsc_0_10_d;
  wire [7:0] accumulation_buffer_rsc_0_10_wadr;
  wire [15:0] accumulation_buffer_rsc_0_10_q;
  wire accumulation_buffer_rsc_0_10_re;
  wire [7:0] accumulation_buffer_rsc_0_10_radr;
  wire accumulation_buffer_rsc_0_11_we;
  wire [15:0] accumulation_buffer_rsc_0_11_d;
  wire [7:0] accumulation_buffer_rsc_0_11_wadr;
  wire [15:0] accumulation_buffer_rsc_0_11_q;
  wire accumulation_buffer_rsc_0_11_re;
  wire [7:0] accumulation_buffer_rsc_0_11_radr;
  wire accumulation_buffer_rsc_0_12_we;
  wire [15:0] accumulation_buffer_rsc_0_12_d;
  wire [7:0] accumulation_buffer_rsc_0_12_wadr;
  wire [15:0] accumulation_buffer_rsc_0_12_q;
  wire accumulation_buffer_rsc_0_12_re;
  wire [7:0] accumulation_buffer_rsc_0_12_radr;
  wire accumulation_buffer_rsc_0_13_we;
  wire [15:0] accumulation_buffer_rsc_0_13_d;
  wire [7:0] accumulation_buffer_rsc_0_13_wadr;
  wire [15:0] accumulation_buffer_rsc_0_13_q;
  wire accumulation_buffer_rsc_0_13_re;
  wire [7:0] accumulation_buffer_rsc_0_13_radr;
  wire accumulation_buffer_rsc_0_14_we;
  wire [15:0] accumulation_buffer_rsc_0_14_d;
  wire [7:0] accumulation_buffer_rsc_0_14_wadr;
  wire [15:0] accumulation_buffer_rsc_0_14_q;
  wire accumulation_buffer_rsc_0_14_re;
  wire [7:0] accumulation_buffer_rsc_0_14_radr;
  wire accumulation_buffer_rsc_0_15_we;
  wire [15:0] accumulation_buffer_rsc_0_15_d;
  wire [7:0] accumulation_buffer_rsc_0_15_wadr;
  wire [15:0] accumulation_buffer_rsc_0_15_q;
  wire accumulation_buffer_rsc_0_15_re;
  wire [7:0] accumulation_buffer_rsc_0_15_radr;
  wire [255:0] output_rsc_dat;
  wire accumulation_buffer_rsc_0_0_i_we_d_iff;
  wire accumulation_buffer_rsc_0_0_i_re_d_iff;
  wire accumulation_buffer_rsc_0_1_i_we_d_iff;
  wire accumulation_buffer_rsc_0_1_i_re_d_iff;
  wire accumulation_buffer_rsc_0_2_i_we_d_iff;
  wire accumulation_buffer_rsc_0_2_i_re_d_iff;
  wire accumulation_buffer_rsc_0_3_i_we_d_iff;
  wire accumulation_buffer_rsc_0_3_i_re_d_iff;
  wire accumulation_buffer_rsc_0_4_i_we_d_iff;
  wire accumulation_buffer_rsc_0_4_i_re_d_iff;
  wire accumulation_buffer_rsc_0_5_i_we_d_iff;
  wire accumulation_buffer_rsc_0_5_i_re_d_iff;
  wire accumulation_buffer_rsc_0_6_i_we_d_iff;
  wire accumulation_buffer_rsc_0_6_i_re_d_iff;
  wire accumulation_buffer_rsc_0_7_i_we_d_iff;
  wire accumulation_buffer_rsc_0_7_i_re_d_iff;
  wire accumulation_buffer_rsc_0_8_i_we_d_iff;
  wire accumulation_buffer_rsc_0_8_i_re_d_iff;
  wire accumulation_buffer_rsc_0_9_i_we_d_iff;
  wire accumulation_buffer_rsc_0_9_i_re_d_iff;
  wire accumulation_buffer_rsc_0_10_i_we_d_iff;
  wire accumulation_buffer_rsc_0_10_i_re_d_iff;
  wire accumulation_buffer_rsc_0_11_i_we_d_iff;
  wire accumulation_buffer_rsc_0_11_i_re_d_iff;
  wire accumulation_buffer_rsc_0_12_i_we_d_iff;
  wire accumulation_buffer_rsc_0_12_i_re_d_iff;
  wire accumulation_buffer_rsc_0_13_i_we_d_iff;
  wire accumulation_buffer_rsc_0_13_i_re_d_iff;
  wire accumulation_buffer_rsc_0_14_i_we_d_iff;
  wire accumulation_buffer_rsc_0_14_i_re_d_iff;
  wire accumulation_buffer_rsc_0_15_i_we_d_iff;
  wire accumulation_buffer_rsc_0_15_i_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat
      = {paramsIn_rsc_dat_STRIDE , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1
      , paramsIn_rsc_dat_OC1 , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1
      , paramsIn_rsc_dat_OY1};
  wire [47:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat
      = {loopIndicesIn_rsc_dat_fy_idx , loopIndicesIn_rsc_dat_fx_idx , loopIndicesIn_rsc_dat_ic1_idx};
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_0_comp (
      .radr(accumulation_buffer_rsc_0_0_radr),
      .wadr(accumulation_buffer_rsc_0_0_wadr),
      .d(accumulation_buffer_rsc_0_0_d),
      .we(accumulation_buffer_rsc_0_0_we),
      .re(accumulation_buffer_rsc_0_0_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_0_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_1_comp (
      .radr(accumulation_buffer_rsc_0_1_radr),
      .wadr(accumulation_buffer_rsc_0_1_wadr),
      .d(accumulation_buffer_rsc_0_1_d),
      .we(accumulation_buffer_rsc_0_1_we),
      .re(accumulation_buffer_rsc_0_1_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_1_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_2_comp (
      .radr(accumulation_buffer_rsc_0_2_radr),
      .wadr(accumulation_buffer_rsc_0_2_wadr),
      .d(accumulation_buffer_rsc_0_2_d),
      .we(accumulation_buffer_rsc_0_2_we),
      .re(accumulation_buffer_rsc_0_2_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_2_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_3_comp (
      .radr(accumulation_buffer_rsc_0_3_radr),
      .wadr(accumulation_buffer_rsc_0_3_wadr),
      .d(accumulation_buffer_rsc_0_3_d),
      .we(accumulation_buffer_rsc_0_3_we),
      .re(accumulation_buffer_rsc_0_3_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_3_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_4_comp (
      .radr(accumulation_buffer_rsc_0_4_radr),
      .wadr(accumulation_buffer_rsc_0_4_wadr),
      .d(accumulation_buffer_rsc_0_4_d),
      .we(accumulation_buffer_rsc_0_4_we),
      .re(accumulation_buffer_rsc_0_4_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_4_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_5_comp (
      .radr(accumulation_buffer_rsc_0_5_radr),
      .wadr(accumulation_buffer_rsc_0_5_wadr),
      .d(accumulation_buffer_rsc_0_5_d),
      .we(accumulation_buffer_rsc_0_5_we),
      .re(accumulation_buffer_rsc_0_5_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_5_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_6_comp (
      .radr(accumulation_buffer_rsc_0_6_radr),
      .wadr(accumulation_buffer_rsc_0_6_wadr),
      .d(accumulation_buffer_rsc_0_6_d),
      .we(accumulation_buffer_rsc_0_6_we),
      .re(accumulation_buffer_rsc_0_6_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_6_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_7_comp (
      .radr(accumulation_buffer_rsc_0_7_radr),
      .wadr(accumulation_buffer_rsc_0_7_wadr),
      .d(accumulation_buffer_rsc_0_7_d),
      .we(accumulation_buffer_rsc_0_7_we),
      .re(accumulation_buffer_rsc_0_7_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_7_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_8_comp (
      .radr(accumulation_buffer_rsc_0_8_radr),
      .wadr(accumulation_buffer_rsc_0_8_wadr),
      .d(accumulation_buffer_rsc_0_8_d),
      .we(accumulation_buffer_rsc_0_8_we),
      .re(accumulation_buffer_rsc_0_8_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_8_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_9_comp (
      .radr(accumulation_buffer_rsc_0_9_radr),
      .wadr(accumulation_buffer_rsc_0_9_wadr),
      .d(accumulation_buffer_rsc_0_9_d),
      .we(accumulation_buffer_rsc_0_9_we),
      .re(accumulation_buffer_rsc_0_9_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_9_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_10_comp (
      .radr(accumulation_buffer_rsc_0_10_radr),
      .wadr(accumulation_buffer_rsc_0_10_wadr),
      .d(accumulation_buffer_rsc_0_10_d),
      .we(accumulation_buffer_rsc_0_10_we),
      .re(accumulation_buffer_rsc_0_10_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_10_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_11_comp (
      .radr(accumulation_buffer_rsc_0_11_radr),
      .wadr(accumulation_buffer_rsc_0_11_wadr),
      .d(accumulation_buffer_rsc_0_11_d),
      .we(accumulation_buffer_rsc_0_11_we),
      .re(accumulation_buffer_rsc_0_11_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_11_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_12_comp (
      .radr(accumulation_buffer_rsc_0_12_radr),
      .wadr(accumulation_buffer_rsc_0_12_wadr),
      .d(accumulation_buffer_rsc_0_12_d),
      .we(accumulation_buffer_rsc_0_12_we),
      .re(accumulation_buffer_rsc_0_12_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_12_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_13_comp (
      .radr(accumulation_buffer_rsc_0_13_radr),
      .wadr(accumulation_buffer_rsc_0_13_wadr),
      .d(accumulation_buffer_rsc_0_13_d),
      .we(accumulation_buffer_rsc_0_13_we),
      .re(accumulation_buffer_rsc_0_13_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_13_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_14_comp (
      .radr(accumulation_buffer_rsc_0_14_radr),
      .wadr(accumulation_buffer_rsc_0_14_wadr),
      .d(accumulation_buffer_rsc_0_14_d),
      .we(accumulation_buffer_rsc_0_14_we),
      .re(accumulation_buffer_rsc_0_14_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_14_q)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd8),
  .depth(32'sd256)) accumulation_buffer_rsc_0_15_comp (
      .radr(accumulation_buffer_rsc_0_15_radr),
      .wadr(accumulation_buffer_rsc_0_15_wadr),
      .d(accumulation_buffer_rsc_0_15_d),
      .we(accumulation_buffer_rsc_0_15_we),
      .re(accumulation_buffer_rsc_0_15_re),
      .clk(clk),
      .q(accumulation_buffer_rsc_0_15_q)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_149_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_0_i (
      .we(accumulation_buffer_rsc_0_0_we),
      .d(accumulation_buffer_rsc_0_0_d),
      .wadr(accumulation_buffer_rsc_0_0_wadr),
      .q(accumulation_buffer_rsc_0_0_q),
      .re(accumulation_buffer_rsc_0_0_re),
      .radr(accumulation_buffer_rsc_0_0_radr),
      .radr_d(accumulation_buffer_rsc_0_0_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_0_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_0_i_d_d),
      .we_d(accumulation_buffer_rsc_0_0_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_0_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_0_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_0_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_0_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_150_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_1_i (
      .we(accumulation_buffer_rsc_0_1_we),
      .d(accumulation_buffer_rsc_0_1_d),
      .wadr(accumulation_buffer_rsc_0_1_wadr),
      .q(accumulation_buffer_rsc_0_1_q),
      .re(accumulation_buffer_rsc_0_1_re),
      .radr(accumulation_buffer_rsc_0_1_radr),
      .radr_d(accumulation_buffer_rsc_0_1_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_1_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_1_i_d_d),
      .we_d(accumulation_buffer_rsc_0_1_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_1_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_1_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_1_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_1_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_151_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_2_i (
      .we(accumulation_buffer_rsc_0_2_we),
      .d(accumulation_buffer_rsc_0_2_d),
      .wadr(accumulation_buffer_rsc_0_2_wadr),
      .q(accumulation_buffer_rsc_0_2_q),
      .re(accumulation_buffer_rsc_0_2_re),
      .radr(accumulation_buffer_rsc_0_2_radr),
      .radr_d(accumulation_buffer_rsc_0_2_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_2_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_2_i_d_d),
      .we_d(accumulation_buffer_rsc_0_2_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_2_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_2_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_2_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_2_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_152_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_3_i (
      .we(accumulation_buffer_rsc_0_3_we),
      .d(accumulation_buffer_rsc_0_3_d),
      .wadr(accumulation_buffer_rsc_0_3_wadr),
      .q(accumulation_buffer_rsc_0_3_q),
      .re(accumulation_buffer_rsc_0_3_re),
      .radr(accumulation_buffer_rsc_0_3_radr),
      .radr_d(accumulation_buffer_rsc_0_3_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_3_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_3_i_d_d),
      .we_d(accumulation_buffer_rsc_0_3_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_3_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_3_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_3_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_3_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_153_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_4_i (
      .we(accumulation_buffer_rsc_0_4_we),
      .d(accumulation_buffer_rsc_0_4_d),
      .wadr(accumulation_buffer_rsc_0_4_wadr),
      .q(accumulation_buffer_rsc_0_4_q),
      .re(accumulation_buffer_rsc_0_4_re),
      .radr(accumulation_buffer_rsc_0_4_radr),
      .radr_d(accumulation_buffer_rsc_0_4_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_4_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_4_i_d_d),
      .we_d(accumulation_buffer_rsc_0_4_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_4_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_4_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_4_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_4_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_154_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_5_i (
      .we(accumulation_buffer_rsc_0_5_we),
      .d(accumulation_buffer_rsc_0_5_d),
      .wadr(accumulation_buffer_rsc_0_5_wadr),
      .q(accumulation_buffer_rsc_0_5_q),
      .re(accumulation_buffer_rsc_0_5_re),
      .radr(accumulation_buffer_rsc_0_5_radr),
      .radr_d(accumulation_buffer_rsc_0_5_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_5_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_5_i_d_d),
      .we_d(accumulation_buffer_rsc_0_5_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_5_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_5_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_5_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_5_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_155_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_6_i (
      .we(accumulation_buffer_rsc_0_6_we),
      .d(accumulation_buffer_rsc_0_6_d),
      .wadr(accumulation_buffer_rsc_0_6_wadr),
      .q(accumulation_buffer_rsc_0_6_q),
      .re(accumulation_buffer_rsc_0_6_re),
      .radr(accumulation_buffer_rsc_0_6_radr),
      .radr_d(accumulation_buffer_rsc_0_6_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_6_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_6_i_d_d),
      .we_d(accumulation_buffer_rsc_0_6_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_6_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_6_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_6_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_6_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_156_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_7_i (
      .we(accumulation_buffer_rsc_0_7_we),
      .d(accumulation_buffer_rsc_0_7_d),
      .wadr(accumulation_buffer_rsc_0_7_wadr),
      .q(accumulation_buffer_rsc_0_7_q),
      .re(accumulation_buffer_rsc_0_7_re),
      .radr(accumulation_buffer_rsc_0_7_radr),
      .radr_d(accumulation_buffer_rsc_0_7_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_7_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_7_i_d_d),
      .we_d(accumulation_buffer_rsc_0_7_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_7_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_7_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_7_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_7_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_157_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_8_i (
      .we(accumulation_buffer_rsc_0_8_we),
      .d(accumulation_buffer_rsc_0_8_d),
      .wadr(accumulation_buffer_rsc_0_8_wadr),
      .q(accumulation_buffer_rsc_0_8_q),
      .re(accumulation_buffer_rsc_0_8_re),
      .radr(accumulation_buffer_rsc_0_8_radr),
      .radr_d(accumulation_buffer_rsc_0_8_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_8_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_8_i_d_d),
      .we_d(accumulation_buffer_rsc_0_8_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_8_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_8_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_8_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_8_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_158_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_9_i (
      .we(accumulation_buffer_rsc_0_9_we),
      .d(accumulation_buffer_rsc_0_9_d),
      .wadr(accumulation_buffer_rsc_0_9_wadr),
      .q(accumulation_buffer_rsc_0_9_q),
      .re(accumulation_buffer_rsc_0_9_re),
      .radr(accumulation_buffer_rsc_0_9_radr),
      .radr_d(accumulation_buffer_rsc_0_9_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_9_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_9_i_d_d),
      .we_d(accumulation_buffer_rsc_0_9_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_9_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_9_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_9_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_9_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_159_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_10_i (
      .we(accumulation_buffer_rsc_0_10_we),
      .d(accumulation_buffer_rsc_0_10_d),
      .wadr(accumulation_buffer_rsc_0_10_wadr),
      .q(accumulation_buffer_rsc_0_10_q),
      .re(accumulation_buffer_rsc_0_10_re),
      .radr(accumulation_buffer_rsc_0_10_radr),
      .radr_d(accumulation_buffer_rsc_0_10_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_10_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_10_i_d_d),
      .we_d(accumulation_buffer_rsc_0_10_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_10_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_10_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_10_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_10_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_160_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_11_i (
      .we(accumulation_buffer_rsc_0_11_we),
      .d(accumulation_buffer_rsc_0_11_d),
      .wadr(accumulation_buffer_rsc_0_11_wadr),
      .q(accumulation_buffer_rsc_0_11_q),
      .re(accumulation_buffer_rsc_0_11_re),
      .radr(accumulation_buffer_rsc_0_11_radr),
      .radr_d(accumulation_buffer_rsc_0_11_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_11_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_11_i_d_d),
      .we_d(accumulation_buffer_rsc_0_11_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_11_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_11_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_11_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_11_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_161_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_12_i (
      .we(accumulation_buffer_rsc_0_12_we),
      .d(accumulation_buffer_rsc_0_12_d),
      .wadr(accumulation_buffer_rsc_0_12_wadr),
      .q(accumulation_buffer_rsc_0_12_q),
      .re(accumulation_buffer_rsc_0_12_re),
      .radr(accumulation_buffer_rsc_0_12_radr),
      .radr_d(accumulation_buffer_rsc_0_12_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_12_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_12_i_d_d),
      .we_d(accumulation_buffer_rsc_0_12_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_12_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_12_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_12_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_12_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_162_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_13_i (
      .we(accumulation_buffer_rsc_0_13_we),
      .d(accumulation_buffer_rsc_0_13_d),
      .wadr(accumulation_buffer_rsc_0_13_wadr),
      .q(accumulation_buffer_rsc_0_13_q),
      .re(accumulation_buffer_rsc_0_13_re),
      .radr(accumulation_buffer_rsc_0_13_radr),
      .radr_d(accumulation_buffer_rsc_0_13_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_13_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_13_i_d_d),
      .we_d(accumulation_buffer_rsc_0_13_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_13_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_13_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_13_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_13_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_163_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_14_i (
      .we(accumulation_buffer_rsc_0_14_we),
      .d(accumulation_buffer_rsc_0_14_d),
      .wadr(accumulation_buffer_rsc_0_14_wadr),
      .q(accumulation_buffer_rsc_0_14_q),
      .re(accumulation_buffer_rsc_0_14_re),
      .radr(accumulation_buffer_rsc_0_14_radr),
      .radr_d(accumulation_buffer_rsc_0_14_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_14_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_14_i_d_d),
      .we_d(accumulation_buffer_rsc_0_14_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_14_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_14_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_14_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_14_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_164_16_8_256_256_16_5_gen
      accumulation_buffer_rsc_0_15_i (
      .we(accumulation_buffer_rsc_0_15_we),
      .d(accumulation_buffer_rsc_0_15_d),
      .wadr(accumulation_buffer_rsc_0_15_wadr),
      .q(accumulation_buffer_rsc_0_15_q),
      .re(accumulation_buffer_rsc_0_15_re),
      .radr(accumulation_buffer_rsc_0_15_radr),
      .radr_d(accumulation_buffer_rsc_0_15_i_radr_d),
      .wadr_d(accumulation_buffer_rsc_0_15_i_wadr_d),
      .d_d(accumulation_buffer_rsc_0_15_i_d_d),
      .we_d(accumulation_buffer_rsc_0_15_i_we_d_iff),
      .re_d(accumulation_buffer_rsc_0_15_i_re_d_iff),
      .q_d(accumulation_buffer_rsc_0_15_i_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(accumulation_buffer_rsc_0_15_i_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(accumulation_buffer_rsc_0_15_i_we_d_iff)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat_value),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .weight_rsc_dat(weight_rsc_dat_value),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .output_rsc_dat(output_rsc_dat),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .loopIndicesIn_rsc_dat(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_run_inst_loopIndicesIn_rsc_dat[47:0]),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .accumulation_buffer_rsc_0_0_i_radr_d(accumulation_buffer_rsc_0_0_i_radr_d),
      .accumulation_buffer_rsc_0_0_i_wadr_d(accumulation_buffer_rsc_0_0_i_wadr_d),
      .accumulation_buffer_rsc_0_0_i_d_d(accumulation_buffer_rsc_0_0_i_d_d),
      .accumulation_buffer_rsc_0_0_i_q_d(accumulation_buffer_rsc_0_0_i_q_d),
      .accumulation_buffer_rsc_0_1_i_radr_d(accumulation_buffer_rsc_0_1_i_radr_d),
      .accumulation_buffer_rsc_0_1_i_wadr_d(accumulation_buffer_rsc_0_1_i_wadr_d),
      .accumulation_buffer_rsc_0_1_i_d_d(accumulation_buffer_rsc_0_1_i_d_d),
      .accumulation_buffer_rsc_0_1_i_q_d(accumulation_buffer_rsc_0_1_i_q_d),
      .accumulation_buffer_rsc_0_2_i_radr_d(accumulation_buffer_rsc_0_2_i_radr_d),
      .accumulation_buffer_rsc_0_2_i_wadr_d(accumulation_buffer_rsc_0_2_i_wadr_d),
      .accumulation_buffer_rsc_0_2_i_d_d(accumulation_buffer_rsc_0_2_i_d_d),
      .accumulation_buffer_rsc_0_2_i_q_d(accumulation_buffer_rsc_0_2_i_q_d),
      .accumulation_buffer_rsc_0_3_i_radr_d(accumulation_buffer_rsc_0_3_i_radr_d),
      .accumulation_buffer_rsc_0_3_i_wadr_d(accumulation_buffer_rsc_0_3_i_wadr_d),
      .accumulation_buffer_rsc_0_3_i_d_d(accumulation_buffer_rsc_0_3_i_d_d),
      .accumulation_buffer_rsc_0_3_i_q_d(accumulation_buffer_rsc_0_3_i_q_d),
      .accumulation_buffer_rsc_0_4_i_radr_d(accumulation_buffer_rsc_0_4_i_radr_d),
      .accumulation_buffer_rsc_0_4_i_wadr_d(accumulation_buffer_rsc_0_4_i_wadr_d),
      .accumulation_buffer_rsc_0_4_i_d_d(accumulation_buffer_rsc_0_4_i_d_d),
      .accumulation_buffer_rsc_0_4_i_q_d(accumulation_buffer_rsc_0_4_i_q_d),
      .accumulation_buffer_rsc_0_5_i_radr_d(accumulation_buffer_rsc_0_5_i_radr_d),
      .accumulation_buffer_rsc_0_5_i_wadr_d(accumulation_buffer_rsc_0_5_i_wadr_d),
      .accumulation_buffer_rsc_0_5_i_d_d(accumulation_buffer_rsc_0_5_i_d_d),
      .accumulation_buffer_rsc_0_5_i_q_d(accumulation_buffer_rsc_0_5_i_q_d),
      .accumulation_buffer_rsc_0_6_i_radr_d(accumulation_buffer_rsc_0_6_i_radr_d),
      .accumulation_buffer_rsc_0_6_i_wadr_d(accumulation_buffer_rsc_0_6_i_wadr_d),
      .accumulation_buffer_rsc_0_6_i_d_d(accumulation_buffer_rsc_0_6_i_d_d),
      .accumulation_buffer_rsc_0_6_i_q_d(accumulation_buffer_rsc_0_6_i_q_d),
      .accumulation_buffer_rsc_0_7_i_radr_d(accumulation_buffer_rsc_0_7_i_radr_d),
      .accumulation_buffer_rsc_0_7_i_wadr_d(accumulation_buffer_rsc_0_7_i_wadr_d),
      .accumulation_buffer_rsc_0_7_i_d_d(accumulation_buffer_rsc_0_7_i_d_d),
      .accumulation_buffer_rsc_0_7_i_q_d(accumulation_buffer_rsc_0_7_i_q_d),
      .accumulation_buffer_rsc_0_8_i_radr_d(accumulation_buffer_rsc_0_8_i_radr_d),
      .accumulation_buffer_rsc_0_8_i_wadr_d(accumulation_buffer_rsc_0_8_i_wadr_d),
      .accumulation_buffer_rsc_0_8_i_d_d(accumulation_buffer_rsc_0_8_i_d_d),
      .accumulation_buffer_rsc_0_8_i_q_d(accumulation_buffer_rsc_0_8_i_q_d),
      .accumulation_buffer_rsc_0_9_i_radr_d(accumulation_buffer_rsc_0_9_i_radr_d),
      .accumulation_buffer_rsc_0_9_i_wadr_d(accumulation_buffer_rsc_0_9_i_wadr_d),
      .accumulation_buffer_rsc_0_9_i_d_d(accumulation_buffer_rsc_0_9_i_d_d),
      .accumulation_buffer_rsc_0_9_i_q_d(accumulation_buffer_rsc_0_9_i_q_d),
      .accumulation_buffer_rsc_0_10_i_radr_d(accumulation_buffer_rsc_0_10_i_radr_d),
      .accumulation_buffer_rsc_0_10_i_wadr_d(accumulation_buffer_rsc_0_10_i_wadr_d),
      .accumulation_buffer_rsc_0_10_i_d_d(accumulation_buffer_rsc_0_10_i_d_d),
      .accumulation_buffer_rsc_0_10_i_q_d(accumulation_buffer_rsc_0_10_i_q_d),
      .accumulation_buffer_rsc_0_11_i_radr_d(accumulation_buffer_rsc_0_11_i_radr_d),
      .accumulation_buffer_rsc_0_11_i_wadr_d(accumulation_buffer_rsc_0_11_i_wadr_d),
      .accumulation_buffer_rsc_0_11_i_d_d(accumulation_buffer_rsc_0_11_i_d_d),
      .accumulation_buffer_rsc_0_11_i_q_d(accumulation_buffer_rsc_0_11_i_q_d),
      .accumulation_buffer_rsc_0_12_i_radr_d(accumulation_buffer_rsc_0_12_i_radr_d),
      .accumulation_buffer_rsc_0_12_i_wadr_d(accumulation_buffer_rsc_0_12_i_wadr_d),
      .accumulation_buffer_rsc_0_12_i_d_d(accumulation_buffer_rsc_0_12_i_d_d),
      .accumulation_buffer_rsc_0_12_i_q_d(accumulation_buffer_rsc_0_12_i_q_d),
      .accumulation_buffer_rsc_0_13_i_radr_d(accumulation_buffer_rsc_0_13_i_radr_d),
      .accumulation_buffer_rsc_0_13_i_wadr_d(accumulation_buffer_rsc_0_13_i_wadr_d),
      .accumulation_buffer_rsc_0_13_i_d_d(accumulation_buffer_rsc_0_13_i_d_d),
      .accumulation_buffer_rsc_0_13_i_q_d(accumulation_buffer_rsc_0_13_i_q_d),
      .accumulation_buffer_rsc_0_14_i_radr_d(accumulation_buffer_rsc_0_14_i_radr_d),
      .accumulation_buffer_rsc_0_14_i_wadr_d(accumulation_buffer_rsc_0_14_i_wadr_d),
      .accumulation_buffer_rsc_0_14_i_d_d(accumulation_buffer_rsc_0_14_i_d_d),
      .accumulation_buffer_rsc_0_14_i_q_d(accumulation_buffer_rsc_0_14_i_q_d),
      .accumulation_buffer_rsc_0_15_i_radr_d(accumulation_buffer_rsc_0_15_i_radr_d),
      .accumulation_buffer_rsc_0_15_i_wadr_d(accumulation_buffer_rsc_0_15_i_wadr_d),
      .accumulation_buffer_rsc_0_15_i_d_d(accumulation_buffer_rsc_0_15_i_d_d),
      .accumulation_buffer_rsc_0_15_i_q_d(accumulation_buffer_rsc_0_15_i_q_d),
      .accumulation_buffer_rsc_0_0_i_we_d_pff(accumulation_buffer_rsc_0_0_i_we_d_iff),
      .accumulation_buffer_rsc_0_0_i_re_d_pff(accumulation_buffer_rsc_0_0_i_re_d_iff),
      .accumulation_buffer_rsc_0_1_i_we_d_pff(accumulation_buffer_rsc_0_1_i_we_d_iff),
      .accumulation_buffer_rsc_0_1_i_re_d_pff(accumulation_buffer_rsc_0_1_i_re_d_iff),
      .accumulation_buffer_rsc_0_2_i_we_d_pff(accumulation_buffer_rsc_0_2_i_we_d_iff),
      .accumulation_buffer_rsc_0_2_i_re_d_pff(accumulation_buffer_rsc_0_2_i_re_d_iff),
      .accumulation_buffer_rsc_0_3_i_we_d_pff(accumulation_buffer_rsc_0_3_i_we_d_iff),
      .accumulation_buffer_rsc_0_3_i_re_d_pff(accumulation_buffer_rsc_0_3_i_re_d_iff),
      .accumulation_buffer_rsc_0_4_i_we_d_pff(accumulation_buffer_rsc_0_4_i_we_d_iff),
      .accumulation_buffer_rsc_0_4_i_re_d_pff(accumulation_buffer_rsc_0_4_i_re_d_iff),
      .accumulation_buffer_rsc_0_5_i_we_d_pff(accumulation_buffer_rsc_0_5_i_we_d_iff),
      .accumulation_buffer_rsc_0_5_i_re_d_pff(accumulation_buffer_rsc_0_5_i_re_d_iff),
      .accumulation_buffer_rsc_0_6_i_we_d_pff(accumulation_buffer_rsc_0_6_i_we_d_iff),
      .accumulation_buffer_rsc_0_6_i_re_d_pff(accumulation_buffer_rsc_0_6_i_re_d_iff),
      .accumulation_buffer_rsc_0_7_i_we_d_pff(accumulation_buffer_rsc_0_7_i_we_d_iff),
      .accumulation_buffer_rsc_0_7_i_re_d_pff(accumulation_buffer_rsc_0_7_i_re_d_iff),
      .accumulation_buffer_rsc_0_8_i_we_d_pff(accumulation_buffer_rsc_0_8_i_we_d_iff),
      .accumulation_buffer_rsc_0_8_i_re_d_pff(accumulation_buffer_rsc_0_8_i_re_d_iff),
      .accumulation_buffer_rsc_0_9_i_we_d_pff(accumulation_buffer_rsc_0_9_i_we_d_iff),
      .accumulation_buffer_rsc_0_9_i_re_d_pff(accumulation_buffer_rsc_0_9_i_re_d_iff),
      .accumulation_buffer_rsc_0_10_i_we_d_pff(accumulation_buffer_rsc_0_10_i_we_d_iff),
      .accumulation_buffer_rsc_0_10_i_re_d_pff(accumulation_buffer_rsc_0_10_i_re_d_iff),
      .accumulation_buffer_rsc_0_11_i_we_d_pff(accumulation_buffer_rsc_0_11_i_we_d_iff),
      .accumulation_buffer_rsc_0_11_i_re_d_pff(accumulation_buffer_rsc_0_11_i_re_d_iff),
      .accumulation_buffer_rsc_0_12_i_we_d_pff(accumulation_buffer_rsc_0_12_i_we_d_iff),
      .accumulation_buffer_rsc_0_12_i_re_d_pff(accumulation_buffer_rsc_0_12_i_re_d_iff),
      .accumulation_buffer_rsc_0_13_i_we_d_pff(accumulation_buffer_rsc_0_13_i_we_d_iff),
      .accumulation_buffer_rsc_0_13_i_re_d_pff(accumulation_buffer_rsc_0_13_i_re_d_iff),
      .accumulation_buffer_rsc_0_14_i_we_d_pff(accumulation_buffer_rsc_0_14_i_we_d_iff),
      .accumulation_buffer_rsc_0_14_i_re_d_pff(accumulation_buffer_rsc_0_14_i_re_d_iff),
      .accumulation_buffer_rsc_0_15_i_we_d_pff(accumulation_buffer_rsc_0_15_i_we_d_iff),
      .accumulation_buffer_rsc_0_15_i_re_d_pff(accumulation_buffer_rsc_0_15_i_re_d_iff)
    );
  assign output_rsc_dat_value = output_rsc_dat;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16
// ------------------------------------------------------------------


module SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16 (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld,
      loopIndicesIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [47:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;


  // Interconnect Declarations
  wire [255:0] output_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE
      = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY
      = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX
      = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1
      = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1
      = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0
      = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0
      = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1
      = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1
      = paramsIn_rsc_dat[15:0];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx
      = loopIndicesIn_rsc_dat[47:32];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx
      = loopIndicesIn_rsc_dat[31:16];
  wire [15:0] nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx;
  assign nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx
      = loopIndicesIn_rsc_dat[15:0];
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat_value(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy),
      .weight_rsc_dat_value(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy),
      .output_rsc_dat_value(output_rsc_dat_value),
      .output_rsc_vld(output_rsc_vld),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .loopIndicesIn_rsc_dat_fy_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fy_idx[15:0]),
      .loopIndicesIn_rsc_dat_fx_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_fx_idx[15:0]),
      .loopIndicesIn_rsc_dat_ic1_idx(nl_SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16_struct_inst_loopIndicesIn_rsc_dat_ic1_idx[15:0]),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy)
    );
  assign output_rsc_dat = output_rsc_dat_value;
endmodule




//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_in_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_sync_v2 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0
    
    generate 
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data 
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd; 
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
    // synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
    // synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;       // experiment
 
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    // KH assign active = din_vld_int | dout_rdy; // (din_vld & ~din_rdy) | (dout_rdy & ~dout_vld);
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];
             
          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0)) 
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end
        
        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else 
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        if ( peak < count )
          peak = count;
        // synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT 
    generate
    if (ph_clk==1) 
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0) 
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif
   
endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock 
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;
   
    // synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
    // synopsys translate_on

    ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ../WeightDoubleBufferless_384comma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:04:07 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    WeightDoublefeSAqem_cns_bctl
// ------------------------------------------------------------------


module WeightDoublefeSAqem_cns_bctl (
  clk, arst_n, paramsIn_rsc_rdy_nweightDoubleBufferWriter, din_rsc_rdy_nweightDoubleBufferWriter,
      dout_rsc_wadr_nweightDoubleBufferWriter, dout_rsc_d_nweightDoubleBufferWriter,
      dout_rsc_we_nweightDoubleBufferWriter, dout_rsc_req_vz_nweightDoubleBufferWriter,
      paramsIn_rsc_rdy_nweightDoubleBufferReader, din_rsc_radr_nweightDoubleBufferReader,
      din_rsc_re_nweightDoubleBufferReader, din_rsc_q_nweightDoubleBufferReader,
      din_rsc_req_vz_nweightDoubleBufferReader, dout_rsc_vld_nweightDoubleBufferReader,
      paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud, din_rsc_rdy_nweightDoubleBufferWriter_bud,
      dout_rsc_rls_lz_nweightDoubleBufferWriter_bud, din_rsc_rls_lz_nweightDoubleBufferReader_bud,
      paramsIn_rsc_rdy_nweightDoubleBufferReader_bud, dout_rsc_vld_nweightDoubleBufferReader_bud,
      mem_cns_S0, mem_cns_R0, mem_cns_S1, mem_cns_R1, mem_cns_radr_shi0, mem_cns_radr_shi1,
      mem_cns_wadr_shi0, mem_cns_wadr_shi1, mem_cns_d_shi0, mem_cns_d_shi1, mem_cns_we_shi0,
      mem_cns_we_shi1, mem_cns_re_shi0, mem_cns_re_shi1, mem_cns_q_sho0, mem_cns_q_sho1,
      mem_cns_S0_pff, mem_cns_S1_pff
);
  input clk;
  input arst_n;
  output paramsIn_rsc_rdy_nweightDoubleBufferWriter;
  output din_rsc_rdy_nweightDoubleBufferWriter;
  input [8:0] dout_rsc_wadr_nweightDoubleBufferWriter;
  input [127:0] dout_rsc_d_nweightDoubleBufferWriter;
  input dout_rsc_we_nweightDoubleBufferWriter;
  output dout_rsc_req_vz_nweightDoubleBufferWriter;
  output paramsIn_rsc_rdy_nweightDoubleBufferReader;
  input [8:0] din_rsc_radr_nweightDoubleBufferReader;
  input din_rsc_re_nweightDoubleBufferReader;
  output [127:0] din_rsc_q_nweightDoubleBufferReader;
  output din_rsc_req_vz_nweightDoubleBufferReader;
  output dout_rsc_vld_nweightDoubleBufferReader;
  input paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  input din_rsc_rdy_nweightDoubleBufferWriter_bud;
  input dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  input din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  input paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  input dout_rsc_vld_nweightDoubleBufferReader_bud;
  output mem_cns_S0;
  input mem_cns_R0;
  output mem_cns_S1;
  input mem_cns_R1;
  output [8:0] mem_cns_radr_shi0;
  output [8:0] mem_cns_radr_shi1;
  output [8:0] mem_cns_wadr_shi0;
  output [8:0] mem_cns_wadr_shi1;
  output [127:0] mem_cns_d_shi0;
  output [127:0] mem_cns_d_shi1;
  output mem_cns_we_shi0;
  output mem_cns_we_shi1;
  output mem_cns_re_shi0;
  output mem_cns_re_shi1;
  input [127:0] mem_cns_q_sho0;
  input [127:0] mem_cns_q_sho1;
  output mem_cns_S0_pff;
  output mem_cns_S1_pff;


  // Interconnect Declarations
  wire mem_cns_PC0;
  reg mem_cns_ppidx;
  reg [1:0] mem_cns_ppown;
  wire mem_cns_PC1;
  reg mem_cns_ppidx_1;
  reg [1:0] mem_cns_ppown_1;
  wire [1:0] mem_acc_rmff;
  wire [3:0] nl_mem_acc_rmff;
  wire mem_xor_rmff;
  wire [1:0] mem_acc_1_rmff;
  wire [3:0] nl_mem_acc_1_rmff;
  wire mem_xor_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsc_rdy_nweightDoubleBufferWriter = paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  assign din_rsc_rdy_nweightDoubleBufferWriter = din_rsc_rdy_nweightDoubleBufferWriter_bud;
  assign paramsIn_rsc_rdy_nweightDoubleBufferReader = paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  assign dout_rsc_vld_nweightDoubleBufferReader = dout_rsc_vld_nweightDoubleBufferReader_bud;
  assign dout_rsc_req_vz_nweightDoubleBufferWriter = mem_cns_R0;
  assign din_rsc_req_vz_nweightDoubleBufferReader = mem_cns_R1;
  assign mem_xor_rmff = mem_cns_ppidx ^ mem_cns_PC0;
  assign nl_mem_acc_rmff = mem_cns_ppown + conv_u2u_1_2(mem_cns_PC0) + conv_s2u_1_2(mem_cns_PC1);
  assign mem_acc_rmff = nl_mem_acc_rmff[1:0];
  assign mem_cns_PC0 = mem_cns_S0 & dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  assign mem_xor_1_rmff = mem_cns_ppidx_1 ^ mem_cns_PC1;
  assign nl_mem_acc_1_rmff = mem_cns_ppown_1 + conv_u2u_1_2(mem_cns_PC1) + conv_s2u_1_2(mem_cns_PC0);
  assign mem_acc_1_rmff = nl_mem_acc_1_rmff[1:0];
  assign mem_cns_PC1 = mem_cns_S1 & din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  assign din_rsc_q_nweightDoubleBufferReader = MUX_v_128_2_2(mem_cns_q_sho0, mem_cns_q_sho1,
      mem_cns_ppidx_1);
  assign mem_cns_radr_shi0 = din_rsc_radr_nweightDoubleBufferReader;
  assign mem_cns_wadr_shi0 = dout_rsc_wadr_nweightDoubleBufferWriter;
  assign mem_cns_d_shi0 = dout_rsc_d_nweightDoubleBufferWriter;
  assign mem_cns_we_shi0 = dout_rsc_we_nweightDoubleBufferWriter & mem_cns_S0_pff
      & (~ mem_xor_rmff);
  assign mem_cns_S0 = ~((mem_cns_ppown==2'b10));
  assign mem_cns_S0_pff = ~((mem_acc_rmff==2'b10));
  assign mem_cns_re_shi0 = din_rsc_re_nweightDoubleBufferReader & mem_cns_S1_pff
      & (~ mem_xor_1_rmff);
  assign mem_cns_S1 = (mem_cns_ppown_1!=2'b00);
  assign mem_cns_S1_pff = (mem_acc_1_rmff!=2'b00);
  assign mem_cns_radr_shi1 = din_rsc_radr_nweightDoubleBufferReader;
  assign mem_cns_wadr_shi1 = dout_rsc_wadr_nweightDoubleBufferWriter;
  assign mem_cns_d_shi1 = dout_rsc_d_nweightDoubleBufferWriter;
  assign mem_cns_we_shi1 = dout_rsc_we_nweightDoubleBufferWriter & mem_cns_S0_pff
      & mem_xor_rmff;
  assign mem_cns_re_shi1 = din_rsc_re_nweightDoubleBufferReader & mem_cns_S1_pff
      & mem_xor_1_rmff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mem_cns_ppidx <= 1'b0;
      mem_cns_ppown <= 2'b00;
      mem_cns_ppidx_1 <= 1'b0;
      mem_cns_ppown_1 <= 2'b00;
    end
    else begin
      mem_cns_ppidx <= mem_xor_rmff;
      mem_cns_ppown <= mem_acc_rmff;
      mem_cns_ppidx_1 <= mem_xor_1_rmff;
      mem_cns_ppown_1 <= mem_acc_1_rmff;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier
// ------------------------------------------------------------------


module unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for WeightDoubleBuffer_384_16_16_run_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBuffer_384_16_16_run_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_staller
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_staller (
  run_wen, paramsIn_rsci_wen_comp, weightDoubleBufferWriterParams_cnsi_wen_comp,
      weightDoubleBufferReaderParams_cnsi_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input weightDoubleBufferWriterParams_cnsi_wen_comp;
  input weightDoubleBufferReaderParams_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & weightDoubleBufferWriterParams_cnsi_wen_comp
      & weightDoubleBufferReaderParams_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
    (
  clk, arst_n, weightDoubleBufferReaderParams_cnsi_oswt, weightDoubleBufferReaderParams_cnsi_wen_comp,
      weightDoubleBufferReaderParams_cnsi_biwt, weightDoubleBufferReaderParams_cnsi_bdwt,
      weightDoubleBufferReaderParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  output weightDoubleBufferReaderParams_cnsi_wen_comp;
  input weightDoubleBufferReaderParams_cnsi_biwt;
  input weightDoubleBufferReaderParams_cnsi_bdwt;
  output weightDoubleBufferReaderParams_cnsi_bcwt;
  reg weightDoubleBufferReaderParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferReaderParams_cnsi_wen_comp = (~ weightDoubleBufferReaderParams_cnsi_oswt)
      | weightDoubleBufferReaderParams_cnsi_biwt | weightDoubleBufferReaderParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weightDoubleBufferReaderParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      weightDoubleBufferReaderParams_cnsi_bcwt <= ~((~(weightDoubleBufferReaderParams_cnsi_bcwt
          | weightDoubleBufferReaderParams_cnsi_biwt)) | weightDoubleBufferReaderParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
    (
  run_wen, weightDoubleBufferReaderParams_cnsi_oswt, weightDoubleBufferReaderParams_cnsi_irdy,
      weightDoubleBufferReaderParams_cnsi_biwt, weightDoubleBufferReaderParams_cnsi_bdwt,
      weightDoubleBufferReaderParams_cnsi_bcwt, weightDoubleBufferReaderParams_cnsi_ivld_run_sct
);
  input run_wen;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  input weightDoubleBufferReaderParams_cnsi_irdy;
  output weightDoubleBufferReaderParams_cnsi_biwt;
  output weightDoubleBufferReaderParams_cnsi_bdwt;
  input weightDoubleBufferReaderParams_cnsi_bcwt;
  output weightDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire weightDoubleBufferReaderParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferReaderParams_cnsi_bdwt = weightDoubleBufferReaderParams_cnsi_oswt
      & run_wen;
  assign weightDoubleBufferReaderParams_cnsi_biwt = weightDoubleBufferReaderParams_cnsi_ogwt
      & weightDoubleBufferReaderParams_cnsi_irdy;
  assign weightDoubleBufferReaderParams_cnsi_ogwt = weightDoubleBufferReaderParams_cnsi_oswt
      & (~ weightDoubleBufferReaderParams_cnsi_bcwt);
  assign weightDoubleBufferReaderParams_cnsi_ivld_run_sct = weightDoubleBufferReaderParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
    (
  clk, arst_n, weightDoubleBufferWriterParams_cnsi_oswt, weightDoubleBufferWriterParams_cnsi_wen_comp,
      weightDoubleBufferWriterParams_cnsi_biwt, weightDoubleBufferWriterParams_cnsi_bdwt,
      weightDoubleBufferWriterParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  output weightDoubleBufferWriterParams_cnsi_wen_comp;
  input weightDoubleBufferWriterParams_cnsi_biwt;
  input weightDoubleBufferWriterParams_cnsi_bdwt;
  output weightDoubleBufferWriterParams_cnsi_bcwt;
  reg weightDoubleBufferWriterParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferWriterParams_cnsi_wen_comp = (~ weightDoubleBufferWriterParams_cnsi_oswt)
      | weightDoubleBufferWriterParams_cnsi_biwt | weightDoubleBufferWriterParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      weightDoubleBufferWriterParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      weightDoubleBufferWriterParams_cnsi_bcwt <= ~((~(weightDoubleBufferWriterParams_cnsi_bcwt
          | weightDoubleBufferWriterParams_cnsi_biwt)) | weightDoubleBufferWriterParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
    (
  run_wen, weightDoubleBufferWriterParams_cnsi_oswt, weightDoubleBufferWriterParams_cnsi_irdy,
      weightDoubleBufferWriterParams_cnsi_biwt, weightDoubleBufferWriterParams_cnsi_bdwt,
      weightDoubleBufferWriterParams_cnsi_bcwt, weightDoubleBufferWriterParams_cnsi_ivld_run_sct
);
  input run_wen;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  input weightDoubleBufferWriterParams_cnsi_irdy;
  output weightDoubleBufferWriterParams_cnsi_biwt;
  output weightDoubleBufferWriterParams_cnsi_bdwt;
  input weightDoubleBufferWriterParams_cnsi_bcwt;
  output weightDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire weightDoubleBufferWriterParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign weightDoubleBufferWriterParams_cnsi_bdwt = weightDoubleBufferWriterParams_cnsi_oswt
      & run_wen;
  assign weightDoubleBufferWriterParams_cnsi_biwt = weightDoubleBufferWriterParams_cnsi_ogwt
      & weightDoubleBufferWriterParams_cnsi_irdy;
  assign weightDoubleBufferWriterParams_cnsi_ogwt = weightDoubleBufferWriterParams_cnsi_oswt
      & (~ weightDoubleBufferWriterParams_cnsi_bcwt);
  assign weightDoubleBufferWriterParams_cnsi_ivld_run_sct = weightDoubleBufferWriterParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_384_384_128_5_gen
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_384_384_128_5_gen
    (
  we, d, wadr, wadr_d, d_d, we_d, port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [127:0] d;
  output [8:0] wadr;
  input [8:0] wadr_d;
  input [127:0] d_d;
  input we_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_2_tr0, while_while_C_0_tr0, while_while_C_0_tr1,
      while_while_for_for_C_0_tr0, while_while_for_C_1_tr0, while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input main_C_2_tr0;
  input while_while_C_0_tr0;
  input while_while_C_0_tr1;
  input while_while_for_for_C_0_tr0;
  input while_while_for_C_1_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for WeightDoubleBufferWriter_384_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    while_C_0 = 4'd4,
    while_while_C_0 = 4'd5,
    while_while_for_for_C_0 = 4'd6,
    while_while_for_C_0 = 4'd7,
    while_while_for_C_1 = 4'd8,
    while_while_C_1 = 4'd9,
    while_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBufferWriter_384_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 11'b00000001000;
        if ( main_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 11'b00000100000;
        if ( while_while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else if ( while_while_C_0_tr1 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_for_C_0 : begin
        fsm_output = 11'b00001000000;
        if ( while_while_for_for_C_0_tr0 ) begin
          state_var_NS = while_while_for_C_0;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = while_while_for_C_1;
      end
      while_while_for_C_1 : begin
        fsm_output = 11'b00100000000;
        if ( while_while_for_C_1_tr0 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_C_1 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 11'b10000000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_staller
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, din_rsci_wen_comp, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input din_rsci_wen_comp;
  input dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & din_rsci_wen_comp & dout_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
    (
  clk, arst_n, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt, dout_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;
  input dout_rsc_req_obj_biwt;
  input dout_rsc_req_obj_bdwt;
  output dout_rsc_req_obj_bcwt;
  reg dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_wen_comp = (~ dout_rsc_req_obj_oswt) | dout_rsc_req_obj_biwt
      | dout_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_bcwt <= ~((~(dout_rsc_req_obj_bcwt | dout_rsc_req_obj_biwt))
          | dout_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
    (
  run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_vd, dout_rsc_req_obj_biwt, dout_rsc_req_obj_bdwt,
      dout_rsc_req_obj_bcwt
);
  input run_wen;
  input dout_rsc_req_obj_oswt;
  input dout_rsc_req_obj_vd;
  output dout_rsc_req_obj_biwt;
  output dout_rsc_req_obj_bdwt;
  input dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_bdwt = dout_rsc_req_obj_oswt & run_wen;
  assign dout_rsc_req_obj_biwt = dout_rsc_req_obj_oswt & (~ dout_rsc_req_obj_bcwt)
      & dout_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
    (
  run_wten, dout_rsc_rls_obj_iswt0, dout_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input dout_rsc_rls_obj_iswt0;
  output dout_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_rls_obj_ld_run_sct = dout_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl (
  dout_rsci_we_d_run_sct_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_we_d_run_sct_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_we_d_run_sct_pff = dout_rsci_iswt0_pff & (~ run_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp (
  clk, arst_n, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt, din_rsci_biwt,
      din_rsci_bdwt, din_rsci_bcwt, din_rsci_idat
);
  input clk;
  input arst_n;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  output din_rsci_bcwt;
  reg din_rsci_bcwt;
  input [15:0] din_rsci_idat;


  // Interconnect Declarations
  reg [15:0] din_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_idat_mxwt = MUX_v_16_2_2(din_rsci_idat, din_rsci_idat_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_idat_bfwt <= din_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl (
  run_wen, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_bcwt, din_rsci_irdy_run_sct,
      din_rsci_ivld
);
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  input din_rsci_bcwt;
  output din_rsci_irdy_run_sct;
  input din_rsci_ivld;


  // Interconnect Declarations
  wire din_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_ivld;
  assign din_rsci_ogwt = din_rsci_oswt & (~ din_rsci_bcwt);
  assign din_rsci_irdy_run_sct = din_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [73:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [4:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [36:0] reg_paramsIn_rsci_idat_bfwt_ftd_12;
  reg [31:0] reg_paramsIn_rsci_idat_bfwt_ftd_45;
  wire [4:0] paramsIn_rsci_idat_mxwt_opt_116_112;
  wire [36:0] paramsIn_rsci_idat_mxwt_opt_100_64;
  wire [31:0] paramsIn_rsci_idat_mxwt_opt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_116_112 = MUX_v_5_2_2((paramsIn_rsci_idat[116:112]),
      reg_paramsIn_rsci_idat_bfwt_ftd, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_100_64 = MUX_v_37_2_2((paramsIn_rsci_idat[100:64]),
      reg_paramsIn_rsci_idat_bfwt_ftd_12, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_31_0 = MUX_v_32_2_2((paramsIn_rsci_idat[31:0]),
      reg_paramsIn_rsci_idat_bfwt_ftd_45, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {paramsIn_rsci_idat_mxwt_opt_116_112 , paramsIn_rsci_idat_mxwt_opt_100_64
      , paramsIn_rsci_idat_mxwt_opt_31_0};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 5'b00000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_opt_116_112;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= 37'b0000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= paramsIn_rsci_idat_mxwt_opt_100_64;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= paramsIn_rsci_idat_mxwt_opt_31_0;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [36:0] MUX_v_37_2_2;
    input [36:0] input_0;
    input [36:0] input_1;
    input [0:0] sel;
    reg [36:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_37_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_384_384_128_5_gen
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_384_384_128_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [127:0] q;
  output re;
  output [8:0] radr;
  input [8:0] radr_d;
  input re_d;
  output [127:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_2_tr0, while_while_C_0_tr0, while_while_for_C_0_tr0,
      while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input main_C_2_tr0;
  input while_while_C_0_tr0;
  input while_while_for_C_0_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for WeightDoubleBufferReader_384_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    while_C_0 = 4'd4,
    while_while_C_0 = 4'd5,
    while_while_for_C_0 = 4'd6,
    while_while_C_1 = 4'd7,
    while_C_1 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WeightDoubleBufferReader_384_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 9'b000001000;
        if ( main_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 9'b000010000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 9'b000100000;
        if ( while_while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 9'b001000000;
        if ( while_while_for_C_0_tr0 ) begin
          state_var_NS = while_while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_C_1 : begin
        fsm_output = 9'b010000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 9'b100000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_staller
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, dout_rsci_wen_comp, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input dout_rsci_wen_comp;
  input din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & dout_rsci_wen_comp & din_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
    (
  clk, arst_n, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt, din_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;
  input din_rsc_req_obj_biwt;
  input din_rsc_req_obj_bdwt;
  output din_rsc_req_obj_bcwt;
  reg din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_wen_comp = (~ din_rsc_req_obj_oswt) | din_rsc_req_obj_biwt
      | din_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_bcwt <= ~((~(din_rsc_req_obj_bcwt | din_rsc_req_obj_biwt))
          | din_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
    (
  run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_vd, din_rsc_req_obj_biwt, din_rsc_req_obj_bdwt,
      din_rsc_req_obj_bcwt
);
  input run_wen;
  input din_rsc_req_obj_oswt;
  input din_rsc_req_obj_vd;
  output din_rsc_req_obj_biwt;
  output din_rsc_req_obj_bdwt;
  input din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_bdwt = din_rsc_req_obj_oswt & run_wen;
  assign din_rsc_req_obj_biwt = din_rsc_req_obj_oswt & (~ din_rsc_req_obj_bcwt) &
      din_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
    (
  run_wten, din_rsc_rls_obj_iswt0, din_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input din_rsc_rls_obj_iswt0;
  output din_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_rls_obj_ld_run_sct = din_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp (
  clk, arst_n, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_bcwt
);
  input clk;
  input arst_n;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;
  output dout_rsci_bcwt;
  reg dout_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl (
  run_wen, dout_rsci_oswt, dout_rsci_irdy, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt,
      dout_rsci_ivld_run_sct
);
  input run_wen;
  input dout_rsci_oswt;
  input dout_rsci_irdy;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  input dout_rsci_bcwt;
  output dout_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dout_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_bdwt = dout_rsci_oswt & run_wen;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_irdy;
  assign dout_rsci_ogwt = dout_rsci_oswt & (~ dout_rsci_bcwt);
  assign dout_rsci_ivld_run_sct = dout_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp (
  clk, arst_n, din_rsci_q_d, din_rsci_q_d_mxwt, din_rsci_biwt, din_rsci_bdwt
);
  input clk;
  input arst_n;
  input [127:0] din_rsci_q_d;
  output [127:0] din_rsci_q_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [127:0] din_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_q_d_mxwt = MUX_v_128_2_2(din_rsci_q_d, din_rsci_q_d_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_q_d_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_q_d_bfwt <= din_rsci_q_d_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl (
  run_wen, run_wten, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_re_d_run_sct_pff,
      din_rsci_oswt_pff
);
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_re_d_run_sct_pff;
  input din_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = (~ run_wten) & din_rsci_oswt;
  assign din_rsci_re_d_run_sct_pff = din_rsci_oswt_pff & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [63:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [31:0] reg_paramsIn_rsci_idat_bfwt_ftd_33;
  wire [63:0] paramsIn_rsci_idat_mxwt_opt_127_64;
  wire [31:0] paramsIn_rsci_idat_mxwt_opt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_127_64 = MUX_v_64_2_2((paramsIn_rsci_idat[127:64]),
      reg_paramsIn_rsci_idat_bfwt_ftd, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt_opt_31_0 = MUX_v_32_2_2((paramsIn_rsci_idat[31:0]),
      reg_paramsIn_rsci_idat_bfwt_ftd_33, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {paramsIn_rsci_idat_mxwt_opt_127_64 , paramsIn_rsci_idat_mxwt_opt_31_0};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_opt_127_64;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_33 <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_33 <= paramsIn_rsci_idat_mxwt_opt_31_0;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi (
  clk, arst_n, weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy, run_wen, weightDoubleBufferReaderParams_cnsi_oswt,
      weightDoubleBufferReaderParams_cnsi_wen_comp, weightDoubleBufferReaderParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;
  input run_wen;
  input weightDoubleBufferReaderParams_cnsi_oswt;
  output weightDoubleBufferReaderParams_cnsi_wen_comp;
  input [143:0] weightDoubleBufferReaderParams_cnsi_idat;


  // Interconnect Declarations
  wire weightDoubleBufferReaderParams_cnsi_irdy;
  wire weightDoubleBufferReaderParams_cnsi_biwt;
  wire weightDoubleBufferReaderParams_cnsi_bdwt;
  wire weightDoubleBufferReaderParams_cnsi_bcwt;
  wire weightDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd19),
  .width(32'sd144)) weightDoubleBufferReaderParams_cnsi (
      .irdy(weightDoubleBufferReaderParams_cnsi_irdy),
      .ivld(weightDoubleBufferReaderParams_cnsi_ivld_run_sct),
      .idat(weightDoubleBufferReaderParams_cnsi_idat),
      .rdy(weightDoubleBufferReaderParams_cns_rdy),
      .vld(weightDoubleBufferReaderParams_cns_vld),
      .dat(weightDoubleBufferReaderParams_cns_dat)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weightDoubleBufferReaderParams_cnsi_oswt(weightDoubleBufferReaderParams_cnsi_oswt),
      .weightDoubleBufferReaderParams_cnsi_irdy(weightDoubleBufferReaderParams_cnsi_irdy),
      .weightDoubleBufferReaderParams_cnsi_biwt(weightDoubleBufferReaderParams_cnsi_biwt),
      .weightDoubleBufferReaderParams_cnsi_bdwt(weightDoubleBufferReaderParams_cnsi_bdwt),
      .weightDoubleBufferReaderParams_cnsi_bcwt(weightDoubleBufferReaderParams_cnsi_bcwt),
      .weightDoubleBufferReaderParams_cnsi_ivld_run_sct(weightDoubleBufferReaderParams_cnsi_ivld_run_sct)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_weightDoubleBufferReaderParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferReaderParams_cnsi_oswt(weightDoubleBufferReaderParams_cnsi_oswt),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_biwt(weightDoubleBufferReaderParams_cnsi_biwt),
      .weightDoubleBufferReaderParams_cnsi_bdwt(weightDoubleBufferReaderParams_cnsi_bdwt),
      .weightDoubleBufferReaderParams_cnsi_bcwt(weightDoubleBufferReaderParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi (
  clk, arst_n, weightDoubleBufferWriterParams_cns_dat, weightDoubleBufferWriterParams_cns_vld,
      weightDoubleBufferWriterParams_cns_rdy, run_wen, weightDoubleBufferWriterParams_cnsi_oswt,
      weightDoubleBufferWriterParams_cnsi_wen_comp, weightDoubleBufferWriterParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  input run_wen;
  input weightDoubleBufferWriterParams_cnsi_oswt;
  output weightDoubleBufferWriterParams_cnsi_wen_comp;
  input [143:0] weightDoubleBufferWriterParams_cnsi_idat;


  // Interconnect Declarations
  wire weightDoubleBufferWriterParams_cnsi_irdy;
  wire weightDoubleBufferWriterParams_cnsi_biwt;
  wire weightDoubleBufferWriterParams_cnsi_bdwt;
  wire weightDoubleBufferWriterParams_cnsi_bcwt;
  wire weightDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd18),
  .width(32'sd144)) weightDoubleBufferWriterParams_cnsi (
      .irdy(weightDoubleBufferWriterParams_cnsi_irdy),
      .ivld(weightDoubleBufferWriterParams_cnsi_ivld_run_sct),
      .idat(weightDoubleBufferWriterParams_cnsi_idat),
      .rdy(weightDoubleBufferWriterParams_cns_rdy),
      .vld(weightDoubleBufferWriterParams_cns_vld),
      .dat(weightDoubleBufferWriterParams_cns_dat)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .weightDoubleBufferWriterParams_cnsi_oswt(weightDoubleBufferWriterParams_cnsi_oswt),
      .weightDoubleBufferWriterParams_cnsi_irdy(weightDoubleBufferWriterParams_cnsi_irdy),
      .weightDoubleBufferWriterParams_cnsi_biwt(weightDoubleBufferWriterParams_cnsi_biwt),
      .weightDoubleBufferWriterParams_cnsi_bdwt(weightDoubleBufferWriterParams_cnsi_bdwt),
      .weightDoubleBufferWriterParams_cnsi_bcwt(weightDoubleBufferWriterParams_cnsi_bcwt),
      .weightDoubleBufferWriterParams_cnsi_ivld_run_sct(weightDoubleBufferWriterParams_cnsi_ivld_run_sct)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp
      WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_weightDoubleBufferWriterParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferWriterParams_cnsi_oswt(weightDoubleBufferWriterParams_cnsi_oswt),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_biwt(weightDoubleBufferWriterParams_cnsi_biwt),
      .weightDoubleBufferWriterParams_cnsi_bdwt(weightDoubleBufferWriterParams_cnsi_bdwt),
      .weightDoubleBufferWriterParams_cnsi_bcwt(weightDoubleBufferWriterParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd17),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj (
  clk, arst_n, dout_rsc_req_vz, run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input dout_rsc_req_vz;
  input run_wen;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_rsc_req_obj_vd;
  wire dout_rsc_req_obj_biwt;
  wire dout_rsc_req_obj_bdwt;
  wire dout_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) dout_rsc_req_obj (
      .vd(dout_rsc_req_obj_vd),
      .vz(dout_rsc_req_vz)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
      WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_vd(dout_rsc_req_obj_vd),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj (
  dout_rsc_rls_lz, run_wten, dout_rsc_rls_obj_iswt0
);
  output dout_rsc_rls_lz;
  input run_wten;
  input dout_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) dout_rsc_rls_obj (
      .ld(dout_rsc_rls_obj_ld_run_sct),
      .lz(dout_rsc_rls_lz)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
      WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(dout_rsc_rls_obj_iswt0),
      .dout_rsc_rls_obj_ld_run_sct(dout_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1 (
  dout_rsci_we_d_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_we_d_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;


  // Interconnect Declarations
  wire dout_rsci_we_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl_inst
      (
      .dout_rsci_we_d_run_sct_pff(dout_rsci_we_d_run_sct_iff),
      .dout_rsci_iswt0_pff(dout_rsci_iswt0_pff),
      .run_wten_pff(run_wten_pff)
    );
  assign dout_rsci_we_d_pff = dout_rsci_we_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_din_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_din_rsci (
  clk, arst_n, din_rsc_dat, din_rsc_vld, din_rsc_rdy, run_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_bcwt;
  wire din_rsci_irdy_run_sct;
  wire din_rsci_ivld;
  wire [15:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd16)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_irdy_run_sct),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_irdy_run_sct(din_rsci_irdy_run_sct),
      .din_rsci_ivld(din_rsci_ivld)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp WeightDoubleBufferWriter_384_16_16_run_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_idat(din_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [73:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [73:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj (
  clk, arst_n, din_rsc_req_vz, run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input din_rsc_req_vz;
  input run_wen;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_rsc_req_obj_vd;
  wire din_rsc_req_obj_biwt;
  wire din_rsc_req_obj_bdwt;
  wire din_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) din_rsc_req_obj (
      .vd(din_rsc_req_obj_vd),
      .vz(din_rsc_req_vz)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_vd(din_rsc_req_obj_vd),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj (
  din_rsc_rls_lz, run_wten, din_rsc_rls_obj_iswt0
);
  output din_rsc_rls_lz;
  input run_wten;
  input din_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) din_rsc_rls_obj (
      .ld(din_rsc_rls_obj_ld_run_sct),
      .lz(din_rsc_rls_lz)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(din_rsc_rls_obj_iswt0),
      .din_rsc_rls_obj_ld_run_sct(din_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_dout_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_dout_rsci (
  clk, arst_n, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, run_wen, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_idat
);
  input clk;
  input arst_n;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [127:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_irdy;
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_bcwt;
  wire dout_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd128)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_ivld_run_sct),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_irdy(dout_rsci_irdy),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt),
      .dout_rsci_ivld_run_sct(dout_rsci_ivld_run_sct)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp WeightDoubleBufferReader_384_16_16_run_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_din_rsci_1
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_din_rsci_1 (
  clk, arst_n, din_rsci_q_d, run_wen, run_wten, din_rsci_oswt, din_rsci_q_d_mxwt,
      din_rsci_re_d_pff, din_rsci_oswt_pff
);
  input clk;
  input arst_n;
  input [127:0] din_rsci_q_d;
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output [127:0] din_rsci_q_d_mxwt;
  output din_rsci_re_d_pff;
  input din_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_re_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_re_d_run_sct_pff(din_rsci_re_d_run_sct_iff),
      .din_rsci_oswt_pff(din_rsci_oswt_pff)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp WeightDoubleBufferReader_384_16_16_run_din_rsci_1_din_rsc_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_q_d(din_rsci_q_d),
      .din_rsci_q_d_mxwt(din_rsci_q_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt)
    );
  assign din_rsci_re_d_pff = din_rsci_re_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [95:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [95:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run_run
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, weightDoubleBufferWriterParams_cns_dat,
      weightDoubleBufferWriterParams_cns_vld, weightDoubleBufferWriterParams_cns_rdy,
      weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire weightDoubleBufferWriterParams_cnsi_wen_comp;
  wire weightDoubleBufferReaderParams_cnsi_wen_comp;
  wire [2:0] fsm_output;
  reg reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse;
  reg [143:0] reg_weightDoubleBufferReaderParams_cnsi_idat_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci WeightDoubleBuffer_384_16_16_run_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferWriterParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy),
      .run_wen(run_wen),
      .weightDoubleBufferWriterParams_cnsi_oswt(reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_idat(reg_weightDoubleBufferReaderParams_cnsi_idat_cse)
    );
  WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi WeightDoubleBuffer_384_16_16_run_run_weightDoubleBufferReaderParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy),
      .run_wen(run_wen),
      .weightDoubleBufferReaderParams_cnsi_oswt(reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_idat(reg_weightDoubleBufferReaderParams_cnsi_idat_cse)
    );
  WeightDoubleBuffer_384_16_16_run_run_staller WeightDoubleBuffer_384_16_16_run_run_staller_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .weightDoubleBufferWriterParams_cnsi_wen_comp(weightDoubleBufferWriterParams_cnsi_wen_comp),
      .weightDoubleBufferReaderParams_cnsi_wen_comp(weightDoubleBufferReaderParams_cnsi_wen_comp)
    );
  WeightDoubleBuffer_384_16_16_run_run_run_fsm WeightDoubleBuffer_384_16_16_run_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_weightDoubleBufferReaderParams_cnsi_idat_cse <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_weightDoubleBufferReaderParams_cnsi_idat_cse <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_weightDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= fsm_output[1];
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~ (fsm_output[1]);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_req_vz, dout_rsc_rls_lz, dout_rsci_wadr_d,
      dout_rsci_d_d, dout_rsci_we_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;
  output [8:0] dout_rsci_wadr_d;
  output [127:0] dout_rsci_d_d;
  output dout_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [73:0] paramsIn_rsci_idat_mxwt;
  wire din_rsci_wen_comp;
  wire [15:0] din_rsci_idat_mxwt;
  wire dout_rsc_req_obj_wen_comp;
  wire [10:0] fsm_output;
  wire [3:0] while_while_for_for_acc_1_tmp;
  wire [4:0] nl_while_while_for_for_acc_1_tmp;
  wire and_dcpl_3;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire or_dcpl_19;
  wire and_dcpl_10;
  wire or_dcpl_25;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_34;
  reg exit_while_while_for_sva;
  wire exit_while_sva_mx0;
  reg [2:0] while_while_for_for_oc0_idx_3_0_sva_2_0;
  reg [31:0] reg_paramsIn_crt_sva_116_0_ftd_21;
  reg reg_dout_rsc_req_obj_iswt0_cse;
  reg reg_dout_rsc_rls_obj_ld_run_psct_cse;
  reg reg_din_rsci_irdy_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire dout_rsci_we_d_iff;
  reg [4:0] while_current_buffer_size_8_4_sva;
  reg [8:0] while_while_for_idx_sva;
  reg [15:0] while_while_for_for_tmp_value_sva;
  reg [7:0] while_while_for_row_value_13_sva;
  reg [7:0] while_while_for_row_value_12_sva;
  reg [7:0] while_while_for_row_value_11_sva;
  reg [7:0] while_while_for_row_value_10_sva;
  reg [7:0] while_while_for_row_value_9_sva;
  reg [7:0] while_while_for_row_value_8_sva;
  reg [7:0] while_while_for_row_value_7_sva;
  reg [7:0] while_while_for_row_value_6_sva;
  reg [7:0] while_while_for_row_value_5_sva;
  reg [7:0] while_while_for_row_value_4_sva;
  reg [7:0] while_while_for_row_value_3_sva;
  reg [7:0] while_while_for_row_value_2_sva;
  reg [7:0] while_while_for_row_value_1_sva;
  reg [7:0] while_while_for_row_value_0_sva;
  reg [4:0] block_size_mul_psp_sva;
  wire [9:0] nl_block_size_mul_psp_sva;
  reg [63:0] total_blocks_lpi_3;
  reg [31:0] total_blocks_mul_2_itm;
  reg [47:0] total_blocks_mul_1_itm;
  wire [63:0] total_blocks_sva_1;
  wire [8:0] while_while_for_idx_sva_2;
  wire [9:0] nl_while_while_for_idx_sva_2;
  wire while_while_for_row_value_and_1_cse;
  wire while_while_for_row_value_and_cse;
  wire while_while_for_row_value_and_3_cse;
  wire while_while_for_row_value_and_2_cse;
  wire while_while_for_row_value_and_5_cse;
  wire while_while_for_row_value_and_4_cse;
  wire while_while_for_row_value_and_12_cse;
  wire operator_64_false_1_acc_1_itm_64_1;
  wire while_while_for_acc_2_itm_5_1;
  wire while_while_aelse_acc_itm_5_1;

  wire[63:0] while_while_acc_nl;
  wire[64:0] nl_while_while_acc_nl;
  wire[4:0] while_current_buffer_size_mux_nl;
  wire[4:0] while_while_acc_2_nl;
  wire[5:0] nl_while_while_acc_2_nl;
  wire[0:0] while_current_buffer_size_or_nl;
  wire[5:0] while_while_for_acc_3_nl;
  wire[7:0] nl_while_while_for_acc_3_nl;
  wire[8:0] while_while_for_idx_mux_nl;
  wire[0:0] or_nl;
  wire[0:0] not_60_nl;
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire[64:0] operator_64_false_1_acc_1_nl;
  wire[65:0] nl_operator_64_false_1_acc_1_nl;
  wire[5:0] while_while_for_acc_2_nl;
  wire[6:0] nl_while_while_for_acc_2_nl;
  wire[5:0] while_while_aelse_acc_nl;
  wire[6:0] nl_while_while_aelse_acc_nl;
  wire[5:0] while_while_aelse_acc_1_nl;
  wire[6:0] nl_while_while_aelse_acc_1_nl;
  wire[4:0] while_while_for_for_1_1_acc_4_nl;
  wire[5:0] nl_while_while_for_for_1_1_acc_4_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff
      = fsm_output[7];
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff
      = ~ run_wen;
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0
      = or_dcpl_19;
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1
      = and_dcpl_3 & (~ while_while_for_acc_2_itm_5_1);
  wire [0:0] nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0;
  assign nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0
      = while_while_for_for_acc_1_tmp[3];
  WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci WeightDoubleBufferWriter_384_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_din_rsci WeightDoubleBufferWriter_384_16_16_run_din_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .run_wen(run_wen),
      .din_rsci_oswt(reg_din_rsci_irdy_run_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1 WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst
      (
      .dout_rsci_we_d_pff(dout_rsci_we_d_iff),
      .dout_rsci_iswt0_pff(nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff[0:0]),
      .run_wten_pff(nl_WeightDoubleBufferWriter_384_16_16_run_dout_rsci_1_inst_run_wten_pff[0:0])
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj WeightDoubleBufferWriter_384_16_16_run_dout_rsc_rls_obj_inst
      (
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(reg_dout_rsc_rls_obj_ld_run_psct_cse)
    );
  WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj WeightDoubleBufferWriter_384_16_16_run_dout_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(reg_dout_rsc_req_obj_iswt0_cse),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferWriter_384_16_16_run_staller WeightDoubleBufferWriter_384_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferWriter_384_16_16_run_run_fsm WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_2_tr0(exit_while_sva_mx0),
      .while_while_C_0_tr0(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr0[0:0]),
      .while_while_C_0_tr1(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_C_0_tr1[0:0]),
      .while_while_for_for_C_0_tr0(nl_WeightDoubleBufferWriter_384_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0[0:0]),
      .while_while_for_C_1_tr0(exit_while_while_for_sva),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign while_while_for_row_value_and_cse = run_wen & (or_dcpl_7 | or_dcpl_6);
  assign while_while_for_row_value_and_1_cse = run_wen & (or_dcpl_4 | or_dcpl_9);
  assign while_while_for_row_value_and_2_cse = run_wen & (or_dcpl_7 | or_dcpl_9);
  assign while_while_for_row_value_and_3_cse = run_wen & (or_dcpl_4 | or_dcpl_6);
  assign while_while_for_row_value_and_4_cse = run_wen & (or_dcpl_7 | or_dcpl_3);
  assign while_while_for_row_value_and_5_cse = run_wen & (or_dcpl_4 | (while_while_for_for_acc_1_tmp[1:0]!=2'b11));
  assign while_while_for_row_value_and_12_cse = run_wen & (or_dcpl_4 | or_dcpl_3);
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ (readslicef_65_1_64((operator_64_false_acc_1_nl)))),
      (~ operator_64_false_1_acc_1_itm_64_1), fsm_output[10]);
  assign total_blocks_sva_1 = conv_u2u_64_64(total_blocks_mul_1_itm * (reg_paramsIn_crt_sva_116_0_ftd_21[15:0]));
  assign nl_while_while_for_idx_sva_2 = while_while_for_idx_sva + 9'b000000001;
  assign while_while_for_idx_sva_2 = nl_while_while_for_idx_sva_2[8:0];
  assign nl_while_while_for_for_acc_1_tmp = conv_u2s_3_4(while_while_for_for_oc0_idx_3_0_sva_2_0)
      + 4'b0001;
  assign while_while_for_for_acc_1_tmp = nl_while_while_for_for_acc_1_tmp[3:0];
  assign nl_operator_64_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_1_acc_1_nl = nl_operator_64_false_1_acc_1_nl[64:0];
  assign operator_64_false_1_acc_1_itm_64_1 = readslicef_65_1_64((operator_64_false_1_acc_1_nl));
  assign and_dcpl_3 = operator_64_false_1_acc_1_itm_64_1 & (~ while_while_aelse_acc_itm_5_1);
  assign or_dcpl_3 = (while_while_for_for_acc_1_tmp[1:0]!=2'b00);
  assign or_dcpl_4 = (while_while_for_for_acc_1_tmp[3:2]!=2'b00);
  assign or_dcpl_6 = (while_while_for_for_acc_1_tmp[1:0]!=2'b10);
  assign or_dcpl_7 = (while_while_for_for_acc_1_tmp[3:2]!=2'b01);
  assign or_dcpl_9 = (while_while_for_for_acc_1_tmp[1:0]!=2'b01);
  assign or_dcpl_19 = (~ operator_64_false_1_acc_1_itm_64_1) | while_while_aelse_acc_itm_5_1;
  assign and_dcpl_10 = ~((fsm_output[1:0]!=2'b00));
  assign or_dcpl_25 = (while_while_for_for_oc0_idx_3_0_sva_2_0!=3'b110);
  assign or_dcpl_26 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b00);
  assign or_dcpl_27 = or_dcpl_26 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_28 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b10);
  assign or_dcpl_29 = or_dcpl_28 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_30 = (while_while_for_for_oc0_idx_3_0_sva_2_0[2:1]!=2'b01);
  assign or_dcpl_31 = or_dcpl_30 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign or_dcpl_32 = or_dcpl_28 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign or_dcpl_33 = or_dcpl_30 | (~ (while_while_for_for_oc0_idx_3_0_sva_2_0[0]));
  assign or_dcpl_34 = or_dcpl_26 | (while_while_for_for_oc0_idx_3_0_sva_2_0[0]);
  assign nl_while_while_for_acc_2_nl = ({1'b1 , (~ block_size_mul_psp_sva)}) + 6'b000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[5:0];
  assign while_while_for_acc_2_itm_5_1 = readslicef_6_1_5((while_while_for_acc_2_nl));
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_5_6(~ while_current_buffer_size_8_4_sva)
      + conv_u2u_5_6(~ block_size_mul_psp_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[5:0];
  assign nl_while_while_aelse_acc_nl = conv_u2u_5_6(readslicef_6_5_1((while_while_aelse_acc_1_nl)))
      + 6'b101101;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[5:0];
  assign while_while_aelse_acc_itm_5_1 = readslicef_6_1_5((while_while_aelse_acc_nl));
  assign nl_while_while_for_for_1_1_acc_4_nl = while_current_buffer_size_8_4_sva
      + (while_while_for_idx_sva[8:4]);
  assign while_while_for_for_1_1_acc_4_nl = nl_while_while_for_for_1_1_acc_4_nl[4:0];
  assign dout_rsci_wadr_d = {(while_while_for_for_1_1_acc_4_nl) , (while_while_for_idx_sva[3:0])};
  assign dout_rsci_d_d = {while_while_for_for_tmp_value_sva , while_while_for_row_value_13_sva
      , while_while_for_row_value_12_sva , while_while_for_row_value_11_sva , while_while_for_row_value_10_sva
      , while_while_for_row_value_9_sva , while_while_for_row_value_8_sva , while_while_for_row_value_7_sva
      , while_while_for_row_value_6_sva , while_while_for_row_value_5_sva , while_while_for_row_value_4_sva
      , while_while_for_row_value_3_sva , while_while_for_row_value_2_sva , while_while_for_row_value_1_sva
      , while_while_for_row_value_0_sva};
  assign dout_rsci_we_d_pff = dout_rsci_we_d_iff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_din_rsci_irdy_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      total_blocks_mul_2_itm <= 32'b00000000000000000000000000000000;
      total_blocks_mul_1_itm <= 48'b000000000000000000000000000000000000000000000000;
      while_current_buffer_size_8_4_sva <= 5'b00000;
      exit_while_while_for_sva <= 1'b0;
      while_while_for_idx_sva <= 9'b000000000;
      while_while_for_for_oc0_idx_3_0_sva_2_0 <= 3'b000;
    end
    else if ( run_wen ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= ~(exit_while_sva_mx0 | (~((fsm_output[3])
          | (fsm_output[10]))));
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_19 & (fsm_output[5]);
      reg_din_rsci_irdy_run_psct_cse <= (and_dcpl_3 & while_while_for_acc_2_itm_5_1
          & (fsm_output[5])) | ((~ (while_while_for_for_acc_1_tmp[3])) & (fsm_output[6]))
          | ((~ exit_while_while_for_sva) & (fsm_output[8]));
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[3]) | (fsm_output[10])
          | (fsm_output[0]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      total_blocks_mul_2_itm <= conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16]) *
          (paramsIn_rsci_idat_mxwt[15:0]));
      total_blocks_mul_1_itm <= conv_u2u_48_48(total_blocks_mul_2_itm * (reg_paramsIn_crt_sva_116_0_ftd_21[31:16]));
      while_current_buffer_size_8_4_sva <= MUX_v_5_2_2(5'b00000, (while_current_buffer_size_mux_nl),
          (while_current_buffer_size_or_nl));
      exit_while_while_for_sva <= ~ (readslicef_6_1_5((while_while_for_acc_3_nl)));
      while_while_for_idx_sva <= MUX_v_9_2_2(9'b000000000, (while_while_for_idx_mux_nl),
          (not_60_nl));
      while_while_for_for_oc0_idx_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (while_while_for_for_acc_1_tmp[2:0]),
          (fsm_output[6]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_mul_psp_sva <= 5'b00000;
    end
    else if ( run_wen & (~ and_dcpl_10) ) begin
      block_size_mul_psp_sva <= nl_block_size_mul_psp_sva[4:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & ((fsm_output[2]) | (fsm_output[3]) | (fsm_output[9]) | (~
        and_dcpl_10)) ) begin
      total_blocks_lpi_3 <= MUX_v_64_2_2(total_blocks_sva_1, (while_while_acc_nl),
          fsm_output[9]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_13_sva <= 8'b00000000;
      while_while_for_row_value_12_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_cse ) begin
      while_while_for_row_value_13_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_13_sva, or_dcpl_25);
      while_while_for_row_value_12_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_row_value_12_sva, or_dcpl_25);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_3_sva <= 8'b00000000;
      while_while_for_row_value_2_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_1_cse ) begin
      while_while_for_row_value_3_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_3_sva, or_dcpl_27);
      while_while_for_row_value_2_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_2_sva,
          or_dcpl_27);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_11_sva <= 8'b00000000;
      while_while_for_row_value_10_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_2_cse ) begin
      while_while_for_row_value_11_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_11_sva, or_dcpl_29);
      while_while_for_row_value_10_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_row_value_10_sva, or_dcpl_29);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_5_sva <= 8'b00000000;
      while_while_for_row_value_4_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_3_cse ) begin
      while_while_for_row_value_5_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_5_sva, or_dcpl_31);
      while_while_for_row_value_4_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_4_sva,
          or_dcpl_31);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_9_sva <= 8'b00000000;
      while_while_for_row_value_8_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_4_cse ) begin
      while_while_for_row_value_9_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_9_sva, or_dcpl_32);
      while_while_for_row_value_8_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_8_sva,
          or_dcpl_32);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_7_sva <= 8'b00000000;
      while_while_for_row_value_6_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_5_cse ) begin
      while_while_for_row_value_7_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_7_sva, or_dcpl_33);
      while_while_for_row_value_6_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_6_sva,
          or_dcpl_33);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_row_value_1_sva <= 8'b00000000;
      while_while_for_row_value_0_sva <= 8'b00000000;
    end
    else if ( while_while_for_row_value_and_12_cse ) begin
      while_while_for_row_value_1_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_row_value_1_sva, or_dcpl_34);
      while_while_for_row_value_0_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]), while_while_for_row_value_0_sva,
          or_dcpl_34);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_tmp_value_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (while_while_for_for_acc_1_tmp[3]) ) begin
      while_while_for_for_tmp_value_sva <= din_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_crt_sva_116_0_ftd_21 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_paramsIn_crt_sva_116_0_ftd_21 <= paramsIn_rsci_idat_mxwt[63:32];
    end
  end
  assign nl_while_while_acc_2_nl = while_current_buffer_size_8_4_sva + block_size_mul_psp_sva;
  assign while_while_acc_2_nl = nl_while_while_acc_2_nl[4:0];
  assign while_current_buffer_size_mux_nl = MUX_v_5_2_2(while_current_buffer_size_8_4_sva,
      (while_while_acc_2_nl), fsm_output[9]);
  assign while_current_buffer_size_or_nl = (fsm_output[9:5]!=5'b00000);
  assign nl_while_while_for_acc_3_nl = ({1'b1 , (while_while_for_idx_sva_2[8:4])})
      + conv_u2u_5_6(~ block_size_mul_psp_sva) + 6'b000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[5:0];
  assign or_nl = (fsm_output[6]) | (fsm_output[8]);
  assign while_while_for_idx_mux_nl = MUX_v_9_2_2(while_while_for_idx_sva_2, while_while_for_idx_sva,
      or_nl);
  assign not_60_nl = ~ (fsm_output[5]);
  assign nl_block_size_mul_psp_sva  = (paramsIn_rsci_idat_mxwt[73:69]) * (paramsIn_rsci_idat_mxwt[68:64]);
  assign nl_while_while_acc_nl = total_blocks_lpi_3 + 64'b1111111111111111111111111111111111111111111111111111111111111111;
  assign while_while_acc_nl = nl_while_while_acc_nl[63:0];

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_6_5_1;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_6_5_1 = tmp[4:0];
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction


  function automatic [63:0] conv_u2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_64 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_req_vz,
      din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, din_rsci_radr_d,
      din_rsci_q_d, din_rsci_re_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  output [8:0] din_rsci_radr_d;
  input [127:0] din_rsci_q_d;
  output din_rsci_re_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [95:0] paramsIn_rsci_idat_mxwt;
  wire [127:0] din_rsci_q_d_mxwt;
  wire dout_rsci_wen_comp;
  reg [127:0] dout_rsci_idat;
  wire din_rsc_req_obj_wen_comp;
  wire [8:0] fsm_output;
  wire [4:0] while_while_for_for_acc_tmp;
  wire [5:0] nl_while_while_for_for_acc_tmp;
  wire or_dcpl;
  wire or_dcpl_4;
  wire or_dcpl_6;
  wire or_tmp_13;
  wire or_tmp_22;
  wire exit_while_sva_mx0;
  reg while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1;
  reg while_while_for_stage_0;
  reg while_while_for_stage_0_2;
  reg while_while_for_asn_3_itm_1;
  reg [63:0] reg_paramsIn_crt_sva_127_0_ftd;
  reg reg_din_rsc_req_obj_iswt0_cse;
  reg reg_din_rsc_rls_obj_ld_run_psct_cse;
  reg reg_dout_rsci_ivld_run_psct_cse;
  reg reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire din_rsci_re_d_iff;
  wire and_41_rmff;
  reg [4:0] while_block_count_4_0_sva;
  reg [4:0] block_size_mul_psp_sva;
  wire [31:0] total_blocks_mul_2_itm_mx1;
  wire [3:0] din_rsci_radr_d_run_3_0_mx1;
  reg [63:0] total_blocks_lpi_3;
  reg [4:0] while_current_buffer_size_8_4_sva;
  reg [31:0] total_blocks_mul_2_itm;
  reg [47:0] total_blocks_mul_1_itm;
  reg [3:0] while_while_for_for_r_idx_4_0_lpi_4_3_0;
  wire [63:0] total_blocks_sva_1;
  wire [31:0] while_while_for_wx_idx_sva_2;
  wire [32:0] nl_while_while_for_wx_idx_sva_2;
  wire while_while_for_acc_2_itm_32_1;
  wire operator_64_false_1_acc_1_itm_64_1;

  wire[4:0] block_size_mul_nl;
  wire[9:0] nl_block_size_mul_nl;
  wire[31:0] total_blocks_mux_nl;
  wire[31:0] total_blocks_mul_2_nl;
  wire[0:0] not_nl;
  wire[63:0] while_while_acc_1_nl;
  wire[64:0] nl_while_while_acc_1_nl;
  wire[4:0] while_while_acc_3_nl;
  wire[5:0] nl_while_while_acc_3_nl;
  wire[0:0] while_current_buffer_size_not_1_nl;
  wire[4:0] while_current_buffer_size_mux_1_nl;
  wire[4:0] while_while_acc_nl;
  wire[5:0] nl_while_while_acc_nl;
  wire[0:0] while_block_count_not_nl;
  wire[0:0] or_13_nl;
  wire[64:0] operator_64_false_acc_1_nl;
  wire[65:0] nl_operator_64_false_acc_1_nl;
  wire[32:0] while_while_for_acc_2_nl;
  wire[34:0] nl_while_while_for_acc_2_nl;
  wire[31:0] while_while_for_for_mux_2_nl;
  wire[31:0] while_while_for_mul_nl;
  wire[64:0] operator_64_false_1_acc_1_nl;
  wire[65:0] nl_operator_64_false_1_acc_1_nl;
  wire[5:0] while_while_aelse_acc_nl;
  wire[6:0] nl_while_while_aelse_acc_nl;
  wire[5:0] while_while_aelse_acc_1_nl;
  wire[6:0] nl_while_while_aelse_acc_1_nl;
  wire[4:0] while_while_for_for_address_acc_nl;
  wire[5:0] nl_while_while_for_for_address_acc_nl;
  wire[4:0] while_while_for_for_address_mul_nl;
  wire[9:0] nl_while_while_for_for_address_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0;
  assign nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0
      = or_dcpl_4;
  wire [0:0] nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0;
  assign nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0
      = ~(while_while_for_stage_0_2 | while_while_for_stage_0);
  WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci WeightDoubleBufferReader_384_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsci_1 WeightDoubleBufferReader_384_16_16_run_din_rsci_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_q_d(din_rsci_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .din_rsci_q_d_mxwt(din_rsci_q_d_mxwt),
      .din_rsci_re_d_pff(din_rsci_re_d_iff),
      .din_rsci_oswt_pff(and_41_rmff)
    );
  WeightDoubleBufferReader_384_16_16_run_dout_rsci WeightDoubleBufferReader_384_16_16_run_dout_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .run_wen(run_wen),
      .dout_rsci_oswt(reg_dout_rsci_ivld_run_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj WeightDoubleBufferReader_384_16_16_run_din_rsc_rls_obj_inst
      (
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(reg_din_rsc_rls_obj_ld_run_psct_cse)
    );
  WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj WeightDoubleBufferReader_384_16_16_run_din_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_vz(din_rsc_req_vz),
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(reg_din_rsc_req_obj_iswt0_cse),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferReader_384_16_16_run_staller WeightDoubleBufferReader_384_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  WeightDoubleBufferReader_384_16_16_run_run_fsm WeightDoubleBufferReader_384_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_2_tr0(exit_while_sva_mx0),
      .while_while_C_0_tr0(nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_C_0_tr0[0:0]),
      .while_while_for_C_0_tr0(nl_WeightDoubleBufferReader_384_16_16_run_run_fsm_inst_while_while_for_C_0_tr0[0:0]),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign and_41_rmff = or_dcpl & while_while_for_stage_0 & (fsm_output[6]);
  assign din_rsci_radr_d_run_3_0_mx1 = MUX_v_4_2_2(while_while_for_for_r_idx_4_0_lpi_4_3_0,
      (signext_4_1(~ while_while_for_acc_2_itm_32_1)), while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1);
  assign or_13_nl = or_dcpl_6 | (~ while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1);
  assign total_blocks_mul_2_itm_mx1 = MUX_v_32_2_2(while_while_for_wx_idx_sva_2,
      total_blocks_mul_2_itm, or_13_nl);
  assign nl_operator_64_false_acc_1_nl = ({1'b1 , (~ total_blocks_sva_1)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_acc_1_nl = nl_operator_64_false_acc_1_nl[64:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ (readslicef_65_1_64((operator_64_false_acc_1_nl)))),
      (~ operator_64_false_1_acc_1_itm_64_1), fsm_output[8]);
  assign total_blocks_sva_1 = conv_u2u_64_64(total_blocks_mul_1_itm * (reg_paramsIn_crt_sva_127_0_ftd[15:0]));
  assign nl_while_while_for_wx_idx_sva_2 = total_blocks_mul_2_itm + 32'b00000000000000000000000000000001;
  assign while_while_for_wx_idx_sva_2 = nl_while_while_for_wx_idx_sva_2[31:0];
  assign while_while_for_for_mux_2_nl = MUX_v_32_2_2(while_while_for_wx_idx_sva_2,
      total_blocks_mul_2_itm, or_dcpl_6);
  assign while_while_for_mul_nl = conv_u2u_32_32((reg_paramsIn_crt_sva_127_0_ftd[47:32])
      * (reg_paramsIn_crt_sva_127_0_ftd[63:48]));
  assign nl_while_while_for_acc_2_nl = ({1'b1 , (while_while_for_for_mux_2_nl)})
      + conv_u2u_32_33(~ (while_while_for_mul_nl)) + 33'b000000000000000000000000000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[32:0];
  assign while_while_for_acc_2_itm_32_1 = readslicef_33_1_32((while_while_for_acc_2_nl));
  assign nl_while_while_for_for_acc_tmp = conv_u2u_4_5(din_rsci_radr_d_run_3_0_mx1)
      + 5'b00001;
  assign while_while_for_for_acc_tmp = nl_while_while_for_for_acc_tmp[4:0];
  assign nl_operator_64_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign operator_64_false_1_acc_1_nl = nl_operator_64_false_1_acc_1_nl[64:0];
  assign operator_64_false_1_acc_1_itm_64_1 = readslicef_65_1_64((operator_64_false_1_acc_1_nl));
  assign or_dcpl = (~ while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1)
      | while_while_for_acc_2_itm_32_1;
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_5_6(~ while_current_buffer_size_8_4_sva)
      + conv_u2u_5_6(~ block_size_mul_psp_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[5:0];
  assign nl_while_while_aelse_acc_nl = conv_u2u_5_6(readslicef_6_5_1((while_while_aelse_acc_1_nl)))
      + 6'b101101;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[5:0];
  assign or_dcpl_4 = ~(operator_64_false_1_acc_1_itm_64_1 & (~ (readslicef_6_1_5((while_while_aelse_acc_nl)))));
  assign or_dcpl_6 = (~ while_while_for_stage_0_2) | while_while_for_asn_3_itm_1;
  assign or_tmp_13 = ~((fsm_output[1:0]!=2'b00));
  assign or_tmp_22 = ~((fsm_output[7:5]!=3'b000));
  assign nl_while_while_for_for_address_mul_nl = while_block_count_4_0_sva * block_size_mul_psp_sva;
  assign while_while_for_for_address_mul_nl = nl_while_while_for_for_address_mul_nl[4:0];
  assign nl_while_while_for_for_address_acc_nl = (while_while_for_for_address_mul_nl)
      + (total_blocks_mul_2_itm_mx1[4:0]);
  assign while_while_for_for_address_acc_nl = nl_while_while_for_for_address_acc_nl[4:0];
  assign din_rsci_radr_d = {(while_while_for_for_address_acc_nl) , din_rsci_radr_d_run_3_0_mx1};
  assign din_rsci_re_d_pff = din_rsci_re_d_iff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_din_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_din_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_dout_rsci_ivld_run_psct_cse <= 1'b0;
      reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      block_size_mul_psp_sva <= 5'b00000;
      total_blocks_mul_2_itm <= 32'b00000000000000000000000000000000;
      total_blocks_mul_1_itm <= 48'b000000000000000000000000000000000000000000000000;
      while_block_count_4_0_sva <= 5'b00000;
      while_while_for_stage_0 <= 1'b0;
      while_while_for_stage_0_2 <= 1'b0;
      while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1 <= 1'b0;
      reg_paramsIn_crt_sva_127_0_ftd <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_din_rsc_req_obj_iswt0_cse <= ~(exit_while_sva_mx0 | (~((fsm_output[3])
          | (fsm_output[8]))));
      reg_din_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_4 & (fsm_output[5]);
      reg_dout_rsci_ivld_run_psct_cse <= while_while_for_stage_0_2 & (~ while_while_for_asn_3_itm_1)
          & (fsm_output[6]);
      reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse <= and_41_rmff;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[3]) | (fsm_output[8])
          | (fsm_output[0]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      block_size_mul_psp_sva <= MUX_v_5_2_2((block_size_mul_nl), block_size_mul_psp_sva,
          or_tmp_13);
      total_blocks_mul_2_itm <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (total_blocks_mux_nl), (not_nl));
      total_blocks_mul_1_itm <= conv_u2u_48_48(total_blocks_mul_2_itm * (reg_paramsIn_crt_sva_127_0_ftd[31:16]));
      while_block_count_4_0_sva <= MUX_v_5_2_2(5'b00000, (while_current_buffer_size_mux_1_nl),
          (while_block_count_not_nl));
      while_while_for_stage_0 <= ~((~(while_while_for_stage_0 & or_dcpl)) & (fsm_output[6]));
      while_while_for_stage_0_2 <= while_while_for_stage_0 & (fsm_output[6]);
      while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1 <= (while_while_for_for_acc_tmp[4])
          | (~ (fsm_output[6]));
      reg_paramsIn_crt_sva_127_0_ftd <= MUX_v_64_2_2((paramsIn_rsci_idat_mxwt[95:32]),
          reg_paramsIn_crt_sva_127_0_ftd, or_tmp_13);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_idat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ (fsm_output[6])) | or_dcpl_6)) ) begin
      dout_rsci_idat <= din_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[5]) |
        (fsm_output[8]))) ) begin
      total_blocks_lpi_3 <= MUX_v_64_2_2(total_blocks_sva_1, (while_while_acc_1_nl),
          fsm_output[7]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_current_buffer_size_8_4_sva <= 5'b00000;
    end
    else if ( (fsm_output[6:5]==2'b00) & run_wen ) begin
      while_current_buffer_size_8_4_sva <= MUX_v_5_2_2(5'b00000, (while_while_acc_3_nl),
          (while_current_buffer_size_not_1_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_asn_3_itm_1 <= 1'b0;
    end
    else if ( run_wen & while_while_for_stage_0 ) begin
      while_while_for_asn_3_itm_1 <= (~ while_while_for_acc_2_itm_32_1) & while_while_for_for_r_idx_slc_while_while_for_for_r_idx_4_0_4_1_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_r_idx_4_0_lpi_4_3_0 <= 4'b0000;
    end
    else if ( run_wen & or_dcpl & while_while_for_stage_0 & (~ (while_while_for_for_acc_tmp[4]))
        ) begin
      while_while_for_for_r_idx_4_0_lpi_4_3_0 <= while_while_for_for_acc_tmp[3:0];
    end
  end
  assign nl_block_size_mul_nl = (paramsIn_rsci_idat_mxwt[84:80]) * (paramsIn_rsci_idat_mxwt[68:64]);
  assign block_size_mul_nl = nl_block_size_mul_nl[4:0];
  assign total_blocks_mul_2_nl = conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16])
      * (paramsIn_rsci_idat_mxwt[15:0]));
  assign total_blocks_mux_nl = MUX_v_32_2_2((total_blocks_mul_2_nl), total_blocks_mul_2_itm_mx1,
      fsm_output[6]);
  assign not_nl = ~ (fsm_output[5]);
  assign nl_while_while_acc_nl = while_block_count_4_0_sva + 5'b00001;
  assign while_while_acc_nl = nl_while_while_acc_nl[4:0];
  assign while_current_buffer_size_mux_1_nl = MUX_v_5_2_2(while_block_count_4_0_sva,
      (while_while_acc_nl), fsm_output[7]);
  assign while_block_count_not_nl = ~ or_tmp_22;
  assign nl_while_while_acc_1_nl = total_blocks_lpi_3 + 64'b1111111111111111111111111111111111111111111111111111111111111111;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[63:0];
  assign nl_while_while_acc_3_nl = while_current_buffer_size_8_4_sva + block_size_mul_psp_sva;
  assign while_while_acc_3_nl = nl_while_while_acc_3_nl[4:0];
  assign while_current_buffer_size_not_1_nl = ~ or_tmp_22;

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_65_1_64;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 64;
    readslicef_65_1_64 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_6_5_1;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_6_5_1 = tmp[4:0];
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [47:0] conv_u2u_48_48 ;
    input [47:0]  vector ;
  begin
    conv_u2u_48_48 = vector;
  end
  endfunction


  function automatic [63:0] conv_u2u_64_64 ;
    input [63:0]  vector ;
  begin
    conv_u2u_64_64 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_run
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, weightDoubleBufferWriterParams_cns_dat,
      weightDoubleBufferWriterParams_cns_vld, weightDoubleBufferWriterParams_cns_rdy,
      weightDoubleBufferReaderParams_cns_dat, weightDoubleBufferReaderParams_cns_vld,
      weightDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] weightDoubleBufferWriterParams_cns_dat;
  output weightDoubleBufferWriterParams_cns_vld;
  input weightDoubleBufferWriterParams_cns_rdy;
  output [143:0] weightDoubleBufferReaderParams_cns_dat;
  output weightDoubleBufferReaderParams_cns_vld;
  input weightDoubleBufferReaderParams_cns_rdy;



  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBuffer_384_16_16_run_run WeightDoubleBuffer_384_16_16_run_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferWriter_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBufferWriter_384_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_wadr, dout_rsc_d, dout_rsc_we, dout_rsc_req_vz,
      dout_rsc_rls_lz
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [8:0] dout_rsc_wadr;
  output [127:0] dout_rsc_d;
  output dout_rsc_we;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;


  // Interconnect Declarations
  wire [8:0] dout_rsci_wadr_d;
  wire [127:0] dout_rsci_d_d;
  wire dout_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferWriter_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_384_384_128_5_gen
      dout_rsci (
      .we(dout_rsc_we),
      .d(dout_rsc_d),
      .wadr(dout_rsc_wadr),
      .wadr_d(dout_rsci_wadr_d),
      .d_d(dout_rsci_d_d),
      .we_d(dout_rsci_we_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(dout_rsci_we_d_iff)
    );
  WeightDoubleBufferWriter_384_16_16_run WeightDoubleBufferWriter_384_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .dout_rsci_wadr_d(dout_rsci_wadr_d),
      .dout_rsci_d_d(dout_rsci_d_d),
      .dout_rsci_we_d_pff(dout_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBufferReader_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBufferReader_384_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_radr,
      din_rsc_re, din_rsc_q, din_rsc_req_vz, din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld,
      dout_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [8:0] din_rsc_radr;
  output din_rsc_re;
  input [127:0] din_rsc_q;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [8:0] din_rsci_radr_d;
  wire [127:0] din_rsci_q_d;
  wire din_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  WeightDoubleBufferReader_384_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_384_384_128_5_gen
      din_rsci (
      .q(din_rsc_q),
      .re(din_rsc_re),
      .radr(din_rsc_radr),
      .radr_d(din_rsci_radr_d),
      .re_d(din_rsci_re_d_iff),
      .q_d(din_rsci_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(din_rsci_re_d_iff)
    );
  WeightDoubleBufferReader_384_16_16_run WeightDoubleBufferReader_384_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_req_vz(din_rsc_req_vz),
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .din_rsci_radr_d(din_rsci_radr_d),
      .din_rsci_q_d(din_rsci_q_d),
      .din_rsci_re_d_pff(din_rsci_re_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16_struct
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16_struct (
  clk, arst_n, weights_in_rsc_dat_value, weights_in_rsc_vld, weights_in_rsc_rdy,
      weights_out_rsc_dat_value, weights_out_rsc_vld, weights_out_rsc_rdy, paramsIn_rsc_dat_STRIDE,
      paramsIn_rsc_dat_FY, paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1, paramsIn_rsc_dat_OC1,
      paramsIn_rsc_dat_OX0, paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1, paramsIn_rsc_dat_OY1,
      paramsIn_rsc_vld, paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] weights_in_rsc_dat_value;
  input weights_in_rsc_vld;
  output weights_in_rsc_rdy;
  output [127:0] weights_out_rsc_dat_value;
  output weights_out_rsc_vld;
  input weights_out_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBufferWriter;
  wire paramsIn_rsc_vld_nweightDoubleBufferWriter;
  wire paramsIn_rsc_rdy_nweightDoubleBufferWriter;
  wire din_rsc_rdy_nweightDoubleBufferWriter;
  wire [8:0] dout_rsc_wadr_nweightDoubleBufferWriter;
  wire [127:0] dout_rsc_d_nweightDoubleBufferWriter;
  wire dout_rsc_we_nweightDoubleBufferWriter;
  wire dout_rsc_req_vz_nweightDoubleBufferWriter;
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBufferReader;
  wire paramsIn_rsc_vld_nweightDoubleBufferReader;
  wire paramsIn_rsc_rdy_nweightDoubleBufferReader;
  wire [8:0] din_rsc_radr_nweightDoubleBufferReader;
  wire din_rsc_re_nweightDoubleBufferReader;
  wire [127:0] din_rsc_q_nweightDoubleBufferReader;
  wire din_rsc_req_vz_nweightDoubleBufferReader;
  wire [127:0] dout_rsc_dat_nweightDoubleBufferReader;
  wire dout_rsc_vld_nweightDoubleBufferReader;
  wire [143:0] weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst;
  wire weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst;
  wire [143:0] weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst;
  wire weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst;
  wire paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud;
  wire weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire din_rsc_rdy_nweightDoubleBufferWriter_bud;
  wire dout_rsc_rls_lz_nweightDoubleBufferWriter_bud;
  wire din_rsc_rls_lz_nweightDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nweightDoubleBufferReader_bud;
  wire weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire dout_rsc_vld_nweightDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud;
  wire weightDoubleBufferWriterParams_unc_2;
  wire weightDoubleBufferWriterParams_idle;
  wire mem_cns_R0;
  wire mem_cns_R1;
  wire [8:0] mem_cns_radr_shi0;
  wire [8:0] mem_cns_radr_shi1;
  wire [8:0] mem_cns_wadr_shi0;
  wire [8:0] mem_cns_wadr_shi1;
  wire [127:0] mem_cns_d_shi0;
  wire [127:0] mem_cns_d_shi1;
  wire mem_cns_we_shi0;
  wire mem_cns_we_shi1;
  wire mem_cns_re_shi0;
  wire mem_cns_re_shi1;
  wire [127:0] mem_cns_q_sho0;
  wire [127:0] mem_cns_q_sho1;
  wire weightDoubleBufferReaderParams_unc_2;
  wire weightDoubleBufferReaderParams_idle;
  wire mem_cns_S0_iff;
  wire mem_cns_S1_iff;
  wire mem_cns_S0_dmo;
  wire mem_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat = {paramsIn_rsc_dat_STRIDE
      , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1 , paramsIn_rsc_dat_OC1
      , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1 , paramsIn_rsc_dat_OY1};
  ccs_pipe_v5 #(.rscid(32'sd15),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferWriterParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .din_vld(weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .din(weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBufferWriter),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBufferWriter),
      .dout(paramsIn_rsc_dat_nweightDoubleBufferWriter),
      .sz(weightDoubleBufferWriterParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferWriterParams_idle)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd128),
  .addr_width(32'sd9),
  .depth(32'sd384)) mem_cns_comp (
      .radr(mem_cns_radr_shi0),
      .wadr(mem_cns_wadr_shi0),
      .d(mem_cns_d_shi0),
      .we(mem_cns_we_shi0),
      .re(mem_cns_re_shi0),
      .clk(clk),
      .q(mem_cns_q_sho0)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd128),
  .addr_width(32'sd9),
  .depth(32'sd384)) mem_cns_comp_1 (
      .radr(mem_cns_radr_shi1),
      .wadr(mem_cns_wadr_shi1),
      .d(mem_cns_d_shi1),
      .we(mem_cns_we_shi1),
      .re(mem_cns_re_shi1),
      .clk(clk),
      .q(mem_cns_q_sho1)
    );
  ccs_pipe_v5 #(.rscid(32'sd16),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferReaderParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .din_vld(weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .din(weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBufferReader),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBufferReader),
      .dout(paramsIn_rsc_dat_nweightDoubleBufferReader),
      .sz(weightDoubleBufferReaderParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferReaderParams_idle)
    );
  WeightDoubleBufferWriter_384_16_16 weightDoubleBufferWriter (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBufferWriter),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBufferWriter),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud),
      .din_rsc_dat(weights_in_rsc_dat_value),
      .din_rsc_vld(weights_in_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy_nweightDoubleBufferWriter_bud),
      .dout_rsc_wadr(dout_rsc_wadr_nweightDoubleBufferWriter),
      .dout_rsc_d(dout_rsc_d_nweightDoubleBufferWriter),
      .dout_rsc_we(dout_rsc_we_nweightDoubleBufferWriter),
      .dout_rsc_req_vz(dout_rsc_req_vz_nweightDoubleBufferWriter),
      .dout_rsc_rls_lz(dout_rsc_rls_lz_nweightDoubleBufferWriter_bud)
    );
  WeightDoubleBufferReader_384_16_16 weightDoubleBufferReader (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBufferReader),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBufferReader),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBufferReader_bud),
      .din_rsc_radr(din_rsc_radr_nweightDoubleBufferReader),
      .din_rsc_re(din_rsc_re_nweightDoubleBufferReader),
      .din_rsc_q(din_rsc_q_nweightDoubleBufferReader),
      .din_rsc_req_vz(din_rsc_req_vz_nweightDoubleBufferReader),
      .din_rsc_rls_lz(din_rsc_rls_lz_nweightDoubleBufferReader_bud),
      .dout_rsc_dat(dout_rsc_dat_nweightDoubleBufferReader),
      .dout_rsc_vld(dout_rsc_vld_nweightDoubleBufferReader_bud),
      .dout_rsc_rdy(weights_out_rsc_rdy)
    );
  WeightDoubleBuffer_384_16_16_run WeightDoubleBuffer_384_16_16_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(nl_WeightDoubleBuffer_384_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferWriterParams_cns_dat(weightDoubleBufferWriterParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferWriterParams_cns_vld(weightDoubleBufferWriterParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferWriterParams_cns_rdy(weightDoubleBufferWriterParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferReaderParams_cns_dat(weightDoubleBufferReaderParams_cns_dat_nWeightDoubleBuffer_384_16_16_run_inst),
      .weightDoubleBufferReaderParams_cns_vld(weightDoubleBufferReaderParams_cns_vld_nWeightDoubleBuffer_384_16_16_run_inst_bud),
      .weightDoubleBufferReaderParams_cns_rdy(weightDoubleBufferReaderParams_cns_rdy_nWeightDoubleBuffer_384_16_16_run_inst)
    );
  unreg_hier unreg (
      .in_0(mem_cns_S0_iff),
      .out_0(mem_cns_R0)
    );
  unreg_hier unreg_1 (
      .in_0(mem_cns_S1_iff),
      .out_0(mem_cns_R1)
    );
  WeightDoublefeSAqem_cns_bctl WeightDoublefeSAqem_cns_bctl_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_rdy_nweightDoubleBufferWriter(paramsIn_rsc_rdy_nweightDoubleBufferWriter),
      .din_rsc_rdy_nweightDoubleBufferWriter(din_rsc_rdy_nweightDoubleBufferWriter),
      .dout_rsc_wadr_nweightDoubleBufferWriter(dout_rsc_wadr_nweightDoubleBufferWriter),
      .dout_rsc_d_nweightDoubleBufferWriter(dout_rsc_d_nweightDoubleBufferWriter),
      .dout_rsc_we_nweightDoubleBufferWriter(dout_rsc_we_nweightDoubleBufferWriter),
      .dout_rsc_req_vz_nweightDoubleBufferWriter(dout_rsc_req_vz_nweightDoubleBufferWriter),
      .paramsIn_rsc_rdy_nweightDoubleBufferReader(paramsIn_rsc_rdy_nweightDoubleBufferReader),
      .din_rsc_radr_nweightDoubleBufferReader(din_rsc_radr_nweightDoubleBufferReader),
      .din_rsc_re_nweightDoubleBufferReader(din_rsc_re_nweightDoubleBufferReader),
      .din_rsc_q_nweightDoubleBufferReader(din_rsc_q_nweightDoubleBufferReader),
      .din_rsc_req_vz_nweightDoubleBufferReader(din_rsc_req_vz_nweightDoubleBufferReader),
      .dout_rsc_vld_nweightDoubleBufferReader(dout_rsc_vld_nweightDoubleBufferReader),
      .paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud(paramsIn_rsc_rdy_nweightDoubleBufferWriter_bud),
      .din_rsc_rdy_nweightDoubleBufferWriter_bud(din_rsc_rdy_nweightDoubleBufferWriter_bud),
      .dout_rsc_rls_lz_nweightDoubleBufferWriter_bud(dout_rsc_rls_lz_nweightDoubleBufferWriter_bud),
      .din_rsc_rls_lz_nweightDoubleBufferReader_bud(din_rsc_rls_lz_nweightDoubleBufferReader_bud),
      .paramsIn_rsc_rdy_nweightDoubleBufferReader_bud(paramsIn_rsc_rdy_nweightDoubleBufferReader_bud),
      .dout_rsc_vld_nweightDoubleBufferReader_bud(dout_rsc_vld_nweightDoubleBufferReader_bud),
      .mem_cns_S0(mem_cns_S0_dmo),
      .mem_cns_R0(mem_cns_R0),
      .mem_cns_S1(mem_cns_S1_dmo),
      .mem_cns_R1(mem_cns_R1),
      .mem_cns_radr_shi0(mem_cns_radr_shi0),
      .mem_cns_radr_shi1(mem_cns_radr_shi1),
      .mem_cns_wadr_shi0(mem_cns_wadr_shi0),
      .mem_cns_wadr_shi1(mem_cns_wadr_shi1),
      .mem_cns_d_shi0(mem_cns_d_shi0),
      .mem_cns_d_shi1(mem_cns_d_shi1),
      .mem_cns_we_shi0(mem_cns_we_shi0),
      .mem_cns_we_shi1(mem_cns_we_shi1),
      .mem_cns_re_shi0(mem_cns_re_shi0),
      .mem_cns_re_shi1(mem_cns_re_shi1),
      .mem_cns_q_sho0(mem_cns_q_sho0),
      .mem_cns_q_sho1(mem_cns_q_sho1),
      .mem_cns_S0_pff(mem_cns_S0_iff),
      .mem_cns_S1_pff(mem_cns_S1_iff)
    );
  assign weights_out_rsc_dat_value = dout_rsc_dat_nweightDoubleBufferReader;
  assign weights_in_rsc_rdy = din_rsc_rdy_nweightDoubleBufferWriter;
  assign weights_out_rsc_vld = dout_rsc_vld_nweightDoubleBufferReader;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nWeightDoubleBuffer_384_16_16_run_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WeightDoubleBuffer_384_16_16
// ------------------------------------------------------------------


module WeightDoubleBuffer_384_16_16 (
  clk, arst_n, weights_in_rsc_dat, weights_in_rsc_vld, weights_in_rsc_rdy, weights_out_rsc_dat,
      weights_out_rsc_vld, weights_out_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] weights_in_rsc_dat;
  input weights_in_rsc_vld;
  output weights_in_rsc_rdy;
  output [127:0] weights_out_rsc_dat;
  output weights_out_rsc_vld;
  input weights_out_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [127:0] weights_out_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1 = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1 = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0 = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0 = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1 = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1 = paramsIn_rsc_dat[15:0];
  WeightDoubleBuffer_384_16_16_struct WeightDoubleBuffer_384_16_16_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .weights_in_rsc_dat_value(weights_in_rsc_dat),
      .weights_in_rsc_vld(weights_in_rsc_vld),
      .weights_in_rsc_rdy(weights_in_rsc_rdy),
      .weights_out_rsc_dat_value(weights_out_rsc_dat_value),
      .weights_out_rsc_vld(weights_out_rsc_vld),
      .weights_out_rsc_rdy(weights_out_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_WeightDoubleBuffer_384_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy)
    );
  assign weights_out_rsc_dat = weights_out_rsc_dat_value;
endmodule




//------> ../InputDoubleBufferless_512comma_16comma_16greater_.v1/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:02:34 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBDjtfoem_cns_bctl
// ------------------------------------------------------------------


module InputDoubleBDjtfoem_cns_bctl (
  clk, arst_n, paramsIn_rsc_rdy_ninputDoubleBufferWriter, din_rsc_rdy_ninputDoubleBufferWriter,
      dout_rsc_wadr_ninputDoubleBufferWriter, dout_rsc_d_ninputDoubleBufferWriter,
      dout_rsc_we_ninputDoubleBufferWriter, dout_rsc_req_vz_ninputDoubleBufferWriter,
      paramsIn_rsc_rdy_ninputDoubleBufferReader, din_rsc_radr_ninputDoubleBufferReader,
      din_rsc_re_ninputDoubleBufferReader, din_rsc_q_ninputDoubleBufferReader, din_rsc_req_vz_ninputDoubleBufferReader,
      dout_rsc_vld_ninputDoubleBufferReader, paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud,
      din_rsc_rdy_ninputDoubleBufferWriter_bud, dout_rsc_rls_lz_ninputDoubleBufferWriter_bud,
      din_rsc_rls_lz_ninputDoubleBufferReader_bud, paramsIn_rsc_rdy_ninputDoubleBufferReader_bud,
      dout_rsc_vld_ninputDoubleBufferReader_bud, mem_cns_S0, mem_cns_R0, mem_cns_S1,
      mem_cns_R1, mem_cns_radr_shi0, mem_cns_radr_shi1, mem_cns_wadr_shi0, mem_cns_wadr_shi1,
      mem_cns_d_shi0, mem_cns_d_shi1, mem_cns_we_shi0, mem_cns_we_shi1, mem_cns_re_shi0,
      mem_cns_re_shi1, mem_cns_q_sho0, mem_cns_q_sho1, mem_cns_S0_pff, mem_cns_S1_pff
);
  input clk;
  input arst_n;
  output paramsIn_rsc_rdy_ninputDoubleBufferWriter;
  output din_rsc_rdy_ninputDoubleBufferWriter;
  input [8:0] dout_rsc_wadr_ninputDoubleBufferWriter;
  input [127:0] dout_rsc_d_ninputDoubleBufferWriter;
  input dout_rsc_we_ninputDoubleBufferWriter;
  output dout_rsc_req_vz_ninputDoubleBufferWriter;
  output paramsIn_rsc_rdy_ninputDoubleBufferReader;
  input [8:0] din_rsc_radr_ninputDoubleBufferReader;
  input din_rsc_re_ninputDoubleBufferReader;
  output [127:0] din_rsc_q_ninputDoubleBufferReader;
  output din_rsc_req_vz_ninputDoubleBufferReader;
  output dout_rsc_vld_ninputDoubleBufferReader;
  input paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  input din_rsc_rdy_ninputDoubleBufferWriter_bud;
  input dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  input din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  input paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  input dout_rsc_vld_ninputDoubleBufferReader_bud;
  output mem_cns_S0;
  input mem_cns_R0;
  output mem_cns_S1;
  input mem_cns_R1;
  output [8:0] mem_cns_radr_shi0;
  output [8:0] mem_cns_radr_shi1;
  output [8:0] mem_cns_wadr_shi0;
  output [8:0] mem_cns_wadr_shi1;
  output [127:0] mem_cns_d_shi0;
  output [127:0] mem_cns_d_shi1;
  output mem_cns_we_shi0;
  output mem_cns_we_shi1;
  output mem_cns_re_shi0;
  output mem_cns_re_shi1;
  input [127:0] mem_cns_q_sho0;
  input [127:0] mem_cns_q_sho1;
  output mem_cns_S0_pff;
  output mem_cns_S1_pff;


  // Interconnect Declarations
  wire mem_cns_PC0;
  reg mem_cns_ppidx;
  reg [1:0] mem_cns_ppown;
  wire mem_cns_PC1;
  reg mem_cns_ppidx_1;
  reg [1:0] mem_cns_ppown_1;
  wire [1:0] mem_acc_rmff;
  wire [3:0] nl_mem_acc_rmff;
  wire mem_xor_rmff;
  wire [1:0] mem_acc_1_rmff;
  wire [3:0] nl_mem_acc_1_rmff;
  wire mem_xor_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsc_rdy_ninputDoubleBufferWriter = paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  assign din_rsc_rdy_ninputDoubleBufferWriter = din_rsc_rdy_ninputDoubleBufferWriter_bud;
  assign paramsIn_rsc_rdy_ninputDoubleBufferReader = paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  assign dout_rsc_vld_ninputDoubleBufferReader = dout_rsc_vld_ninputDoubleBufferReader_bud;
  assign dout_rsc_req_vz_ninputDoubleBufferWriter = mem_cns_R0;
  assign din_rsc_req_vz_ninputDoubleBufferReader = mem_cns_R1;
  assign mem_xor_rmff = mem_cns_ppidx ^ mem_cns_PC0;
  assign nl_mem_acc_rmff = mem_cns_ppown + conv_u2u_1_2(mem_cns_PC0) + conv_s2u_1_2(mem_cns_PC1);
  assign mem_acc_rmff = nl_mem_acc_rmff[1:0];
  assign mem_cns_PC0 = mem_cns_S0 & dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  assign mem_xor_1_rmff = mem_cns_ppidx_1 ^ mem_cns_PC1;
  assign nl_mem_acc_1_rmff = mem_cns_ppown_1 + conv_u2u_1_2(mem_cns_PC1) + conv_s2u_1_2(mem_cns_PC0);
  assign mem_acc_1_rmff = nl_mem_acc_1_rmff[1:0];
  assign mem_cns_PC1 = mem_cns_S1 & din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  assign din_rsc_q_ninputDoubleBufferReader = MUX_v_128_2_2(mem_cns_q_sho0, mem_cns_q_sho1,
      mem_cns_ppidx_1);
  assign mem_cns_radr_shi0 = din_rsc_radr_ninputDoubleBufferReader;
  assign mem_cns_wadr_shi0 = dout_rsc_wadr_ninputDoubleBufferWriter;
  assign mem_cns_d_shi0 = dout_rsc_d_ninputDoubleBufferWriter;
  assign mem_cns_we_shi0 = dout_rsc_we_ninputDoubleBufferWriter & mem_cns_S0_pff
      & (~ mem_xor_rmff);
  assign mem_cns_S0 = ~((mem_cns_ppown==2'b10));
  assign mem_cns_S0_pff = ~((mem_acc_rmff==2'b10));
  assign mem_cns_re_shi0 = din_rsc_re_ninputDoubleBufferReader & mem_cns_S1_pff &
      (~ mem_xor_1_rmff);
  assign mem_cns_S1 = (mem_cns_ppown_1!=2'b00);
  assign mem_cns_S1_pff = (mem_acc_1_rmff!=2'b00);
  assign mem_cns_radr_shi1 = din_rsc_radr_ninputDoubleBufferReader;
  assign mem_cns_wadr_shi1 = dout_rsc_wadr_ninputDoubleBufferWriter;
  assign mem_cns_d_shi1 = dout_rsc_d_ninputDoubleBufferWriter;
  assign mem_cns_we_shi1 = dout_rsc_we_ninputDoubleBufferWriter & mem_cns_S0_pff
      & mem_xor_rmff;
  assign mem_cns_re_shi1 = din_rsc_re_ninputDoubleBufferReader & mem_cns_S1_pff &
      mem_xor_1_rmff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mem_cns_ppidx <= 1'b0;
      mem_cns_ppown <= 2'b00;
      mem_cns_ppidx_1 <= 1'b0;
      mem_cns_ppown_1 <= 2'b00;
    end
    else begin
      mem_cns_ppidx <= mem_xor_rmff;
      mem_cns_ppown <= mem_acc_rmff;
      mem_cns_ppidx_1 <= mem_xor_1_rmff;
      mem_cns_ppown_1 <= mem_acc_1_rmff;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    unreg_hier
// ------------------------------------------------------------------

/*
module unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule
*/
// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for InputDoubleBuffer_512_16_16_run_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBuffer_512_16_16_run_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_staller
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_staller (
  run_wen, paramsIn_rsci_wen_comp, inputDoubleBufferWriterParams_cnsi_wen_comp, inputDoubleBufferReaderParams_cnsi_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input inputDoubleBufferWriterParams_cnsi_wen_comp;
  input inputDoubleBufferReaderParams_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & inputDoubleBufferWriterParams_cnsi_wen_comp
      & inputDoubleBufferReaderParams_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
    (
  clk, arst_n, inputDoubleBufferReaderParams_cnsi_oswt, inputDoubleBufferReaderParams_cnsi_wen_comp,
      inputDoubleBufferReaderParams_cnsi_biwt, inputDoubleBufferReaderParams_cnsi_bdwt,
      inputDoubleBufferReaderParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  output inputDoubleBufferReaderParams_cnsi_wen_comp;
  input inputDoubleBufferReaderParams_cnsi_biwt;
  input inputDoubleBufferReaderParams_cnsi_bdwt;
  output inputDoubleBufferReaderParams_cnsi_bcwt;
  reg inputDoubleBufferReaderParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferReaderParams_cnsi_wen_comp = (~ inputDoubleBufferReaderParams_cnsi_oswt)
      | inputDoubleBufferReaderParams_cnsi_biwt | inputDoubleBufferReaderParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputDoubleBufferReaderParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      inputDoubleBufferReaderParams_cnsi_bcwt <= ~((~(inputDoubleBufferReaderParams_cnsi_bcwt
          | inputDoubleBufferReaderParams_cnsi_biwt)) | inputDoubleBufferReaderParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
    (
  run_wen, inputDoubleBufferReaderParams_cnsi_oswt, inputDoubleBufferReaderParams_cnsi_irdy,
      inputDoubleBufferReaderParams_cnsi_biwt, inputDoubleBufferReaderParams_cnsi_bdwt,
      inputDoubleBufferReaderParams_cnsi_bcwt, inputDoubleBufferReaderParams_cnsi_ivld_run_sct
);
  input run_wen;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  input inputDoubleBufferReaderParams_cnsi_irdy;
  output inputDoubleBufferReaderParams_cnsi_biwt;
  output inputDoubleBufferReaderParams_cnsi_bdwt;
  input inputDoubleBufferReaderParams_cnsi_bcwt;
  output inputDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire inputDoubleBufferReaderParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferReaderParams_cnsi_bdwt = inputDoubleBufferReaderParams_cnsi_oswt
      & run_wen;
  assign inputDoubleBufferReaderParams_cnsi_biwt = inputDoubleBufferReaderParams_cnsi_ogwt
      & inputDoubleBufferReaderParams_cnsi_irdy;
  assign inputDoubleBufferReaderParams_cnsi_ogwt = inputDoubleBufferReaderParams_cnsi_oswt
      & (~ inputDoubleBufferReaderParams_cnsi_bcwt);
  assign inputDoubleBufferReaderParams_cnsi_ivld_run_sct = inputDoubleBufferReaderParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
    (
  clk, arst_n, inputDoubleBufferWriterParams_cnsi_oswt, inputDoubleBufferWriterParams_cnsi_wen_comp,
      inputDoubleBufferWriterParams_cnsi_biwt, inputDoubleBufferWriterParams_cnsi_bdwt,
      inputDoubleBufferWriterParams_cnsi_bcwt
);
  input clk;
  input arst_n;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  output inputDoubleBufferWriterParams_cnsi_wen_comp;
  input inputDoubleBufferWriterParams_cnsi_biwt;
  input inputDoubleBufferWriterParams_cnsi_bdwt;
  output inputDoubleBufferWriterParams_cnsi_bcwt;
  reg inputDoubleBufferWriterParams_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferWriterParams_cnsi_wen_comp = (~ inputDoubleBufferWriterParams_cnsi_oswt)
      | inputDoubleBufferWriterParams_cnsi_biwt | inputDoubleBufferWriterParams_cnsi_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputDoubleBufferWriterParams_cnsi_bcwt <= 1'b0;
    end
    else begin
      inputDoubleBufferWriterParams_cnsi_bcwt <= ~((~(inputDoubleBufferWriterParams_cnsi_bcwt
          | inputDoubleBufferWriterParams_cnsi_biwt)) | inputDoubleBufferWriterParams_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
    (
  run_wen, inputDoubleBufferWriterParams_cnsi_oswt, inputDoubleBufferWriterParams_cnsi_irdy,
      inputDoubleBufferWriterParams_cnsi_biwt, inputDoubleBufferWriterParams_cnsi_bdwt,
      inputDoubleBufferWriterParams_cnsi_bcwt, inputDoubleBufferWriterParams_cnsi_ivld_run_sct
);
  input run_wen;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  input inputDoubleBufferWriterParams_cnsi_irdy;
  output inputDoubleBufferWriterParams_cnsi_biwt;
  output inputDoubleBufferWriterParams_cnsi_bdwt;
  input inputDoubleBufferWriterParams_cnsi_bcwt;
  output inputDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations
  wire inputDoubleBufferWriterParams_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputDoubleBufferWriterParams_cnsi_bdwt = inputDoubleBufferWriterParams_cnsi_oswt
      & run_wen;
  assign inputDoubleBufferWriterParams_cnsi_biwt = inputDoubleBufferWriterParams_cnsi_ogwt
      & inputDoubleBufferWriterParams_cnsi_irdy;
  assign inputDoubleBufferWriterParams_cnsi_ogwt = inputDoubleBufferWriterParams_cnsi_oswt
      & (~ inputDoubleBufferWriterParams_cnsi_bcwt);
  assign inputDoubleBufferWriterParams_cnsi_ivld_run_sct = inputDoubleBufferWriterParams_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_512_512_128_5_gen
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_512_512_128_5_gen
    (
  we, d, wadr, wadr_d, d_d, we_d, port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [127:0] d;
  output [8:0] wadr;
  input [8:0] wadr_d;
  input [127:0] d_d;
  input we_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_4_tr0, while_while_C_1_tr0, while_while_C_2_tr0,
      while_while_for_for_C_0_tr0, while_while_for_C_1_tr0, while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [14:0] fsm_output;
  reg [14:0] fsm_output;
  input main_C_4_tr0;
  input while_while_C_1_tr0;
  input while_while_C_2_tr0;
  input while_while_for_for_C_0_tr0;
  input while_while_for_C_1_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for InputDoubleBufferWriter_512_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    while_C_0 = 4'd6,
    while_while_C_0 = 4'd7,
    while_while_C_1 = 4'd8,
    while_while_C_2 = 4'd9,
    while_while_for_for_C_0 = 4'd10,
    while_while_for_C_0 = 4'd11,
    while_while_for_C_1 = 4'd12,
    while_while_C_3 = 4'd13,
    while_C_1 = 4'd14;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBufferWriter_512_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 15'b000000000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 15'b000000000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 15'b000000000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 15'b000000000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 15'b000000000100000;
        if ( main_C_4_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 15'b000000001000000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 15'b000000010000000;
        state_var_NS = while_while_C_1;
      end
      while_while_C_1 : begin
        fsm_output = 15'b000000100000000;
        if ( while_while_C_1_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_C_2;
        end
      end
      while_while_C_2 : begin
        fsm_output = 15'b000001000000000;
        if ( while_while_C_2_tr0 ) begin
          state_var_NS = while_while_C_3;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_for_C_0 : begin
        fsm_output = 15'b000010000000000;
        if ( while_while_for_for_C_0_tr0 ) begin
          state_var_NS = while_while_for_C_0;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 15'b000100000000000;
        state_var_NS = while_while_for_C_1;
      end
      while_while_for_C_1 : begin
        fsm_output = 15'b001000000000000;
        if ( while_while_for_C_1_tr0 ) begin
          state_var_NS = while_while_C_3;
        end
        else begin
          state_var_NS = while_while_for_for_C_0;
        end
      end
      while_while_C_3 : begin
        fsm_output = 15'b010000000000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 15'b100000000000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 15'b000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_staller
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, din_rsci_wen_comp, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input din_rsci_wen_comp;
  input dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & din_rsci_wen_comp & dout_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp
    (
  clk, arst_n, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp, dout_rsc_req_obj_biwt,
      dout_rsc_req_obj_bdwt, dout_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;
  input dout_rsc_req_obj_biwt;
  input dout_rsc_req_obj_bdwt;
  output dout_rsc_req_obj_bcwt;
  reg dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_wen_comp = (~ dout_rsc_req_obj_oswt) | dout_rsc_req_obj_biwt
      | dout_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      dout_rsc_req_obj_bcwt <= ~((~(dout_rsc_req_obj_bcwt | dout_rsc_req_obj_biwt))
          | dout_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl
    (
  run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_vd, dout_rsc_req_obj_biwt, dout_rsc_req_obj_bdwt,
      dout_rsc_req_obj_bcwt
);
  input run_wen;
  input dout_rsc_req_obj_oswt;
  input dout_rsc_req_obj_vd;
  output dout_rsc_req_obj_biwt;
  output dout_rsc_req_obj_bdwt;
  input dout_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_req_obj_bdwt = dout_rsc_req_obj_oswt & run_wen;
  assign dout_rsc_req_obj_biwt = dout_rsc_req_obj_oswt & (~ dout_rsc_req_obj_bcwt)
      & dout_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl
    (
  run_wten, dout_rsc_rls_obj_iswt0, dout_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input dout_rsc_rls_obj_iswt0;
  output dout_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsc_rls_obj_ld_run_sct = dout_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl (
  dout_rsci_we_d_run_sct_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_we_d_run_sct_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_we_d_run_sct_pff = dout_rsci_iswt0_pff & (~ run_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp (
  clk, arst_n, din_rsci_oswt, din_rsci_wen_comp, din_rsci_idat_mxwt, din_rsci_biwt,
      din_rsci_bdwt, din_rsci_bcwt, din_rsci_idat
);
  input clk;
  input arst_n;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;
  output din_rsci_bcwt;
  reg din_rsci_bcwt;
  input [15:0] din_rsci_idat;


  // Interconnect Declarations
  reg [15:0] din_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_wen_comp = (~ din_rsci_oswt) | din_rsci_biwt | din_rsci_bcwt;
  assign din_rsci_idat_mxwt = MUX_v_16_2_2(din_rsci_idat, din_rsci_idat_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_idat_bfwt <= din_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl (
  run_wen, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_bcwt, din_rsci_irdy_run_sct,
      din_rsci_ivld
);
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  input din_rsci_bcwt;
  output din_rsci_irdy_run_sct;
  input din_rsci_ivld;


  // Interconnect Declarations
  wire din_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = din_rsci_ogwt & din_rsci_ivld;
  assign din_rsci_ogwt = din_rsci_oswt & (~ din_rsci_bcwt);
  assign din_rsci_irdy_run_sct = din_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [136:0] paramsIn_rsci_idat_bfwt_136_0;
  wire [136:0] paramsIn_rsci_idat_mxwt_opt_136_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_136_0 = MUX_v_137_2_2((paramsIn_rsci_idat[136:0]),
      paramsIn_rsci_idat_bfwt_136_0, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_opt_136_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= paramsIn_rsci_idat_mxwt_opt_136_0;
    end
  end

  function automatic [136:0] MUX_v_137_2_2;
    input [136:0] input_0;
    input [136:0] input_1;
    input [0:0] sel;
    reg [136:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_137_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_512_512_128_5_gen
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_512_512_128_5_gen
    (
  q, re, radr, radr_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d
);
  input [127:0] q;
  output re;
  output [8:0] radr;
  input [8:0] radr_d;
  input re_d;
  output [127:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_1_tr0, while_while_C_1_tr0, while_while_for_C_0_tr0,
      while_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input main_C_1_tr0;
  input while_while_C_1_tr0;
  input while_while_for_C_0_tr0;
  input while_C_1_tr0;


  // FSM State Type Declaration for InputDoubleBufferReader_512_16_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    while_C_0 = 4'd3,
    while_while_C_0 = 4'd4,
    while_while_C_1 = 4'd5,
    while_while_for_C_0 = 4'd6,
    while_while_C_2 = 4'd7,
    while_C_1 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputDoubleBufferReader_512_16_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        if ( main_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      while_C_0 : begin
        fsm_output = 9'b000001000;
        state_var_NS = while_while_C_0;
      end
      while_while_C_0 : begin
        fsm_output = 9'b000010000;
        state_var_NS = while_while_C_1;
      end
      while_while_C_1 : begin
        fsm_output = 9'b000100000;
        if ( while_while_C_1_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_for_C_0 : begin
        fsm_output = 9'b001000000;
        if ( while_while_for_C_0_tr0 ) begin
          state_var_NS = while_while_C_2;
        end
        else begin
          state_var_NS = while_while_for_C_0;
        end
      end
      while_while_C_2 : begin
        fsm_output = 9'b010000000;
        state_var_NS = while_while_C_0;
      end
      while_C_1 : begin
        fsm_output = 9'b100000000;
        if ( while_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = while_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_staller
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_staller (
  clk, arst_n, run_wen, run_wten, paramsIn_rsci_wen_comp, dout_rsci_wen_comp, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  output run_wen;
  output run_wten;
  input paramsIn_rsci_wen_comp;
  input dout_rsci_wen_comp;
  input din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & dout_rsci_wen_comp & din_rsc_req_obj_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp
    (
  clk, arst_n, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp, din_rsc_req_obj_biwt,
      din_rsc_req_obj_bdwt, din_rsc_req_obj_bcwt
);
  input clk;
  input arst_n;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;
  input din_rsc_req_obj_biwt;
  input din_rsc_req_obj_bdwt;
  output din_rsc_req_obj_bcwt;
  reg din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_wen_comp = (~ din_rsc_req_obj_oswt) | din_rsc_req_obj_biwt
      | din_rsc_req_obj_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsc_req_obj_bcwt <= 1'b0;
    end
    else begin
      din_rsc_req_obj_bcwt <= ~((~(din_rsc_req_obj_bcwt | din_rsc_req_obj_biwt))
          | din_rsc_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl
    (
  run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_vd, din_rsc_req_obj_biwt, din_rsc_req_obj_bdwt,
      din_rsc_req_obj_bcwt
);
  input run_wen;
  input din_rsc_req_obj_oswt;
  input din_rsc_req_obj_vd;
  output din_rsc_req_obj_biwt;
  output din_rsc_req_obj_bdwt;
  input din_rsc_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_req_obj_bdwt = din_rsc_req_obj_oswt & run_wen;
  assign din_rsc_req_obj_biwt = din_rsc_req_obj_oswt & (~ din_rsc_req_obj_bcwt) &
      din_rsc_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl
    (
  run_wten, din_rsc_rls_obj_iswt0, din_rsc_rls_obj_ld_run_sct
);
  input run_wten;
  input din_rsc_rls_obj_iswt0;
  output din_rsc_rls_obj_ld_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsc_rls_obj_ld_run_sct = din_rsc_rls_obj_iswt0 & (~ run_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp (
  clk, arst_n, dout_rsci_oswt, dout_rsci_wen_comp, dout_rsci_biwt, dout_rsci_bdwt,
      dout_rsci_bcwt
);
  input clk;
  input arst_n;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input dout_rsci_biwt;
  input dout_rsci_bdwt;
  output dout_rsci_bcwt;
  reg dout_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_wen_comp = (~ dout_rsci_oswt) | dout_rsci_biwt | dout_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_bcwt <= 1'b0;
    end
    else begin
      dout_rsci_bcwt <= ~((~(dout_rsci_bcwt | dout_rsci_biwt)) | dout_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl (
  run_wen, dout_rsci_oswt, dout_rsci_irdy, dout_rsci_biwt, dout_rsci_bdwt, dout_rsci_bcwt,
      dout_rsci_ivld_run_sct
);
  input run_wen;
  input dout_rsci_oswt;
  input dout_rsci_irdy;
  output dout_rsci_biwt;
  output dout_rsci_bdwt;
  input dout_rsci_bcwt;
  output dout_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire dout_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign dout_rsci_bdwt = dout_rsci_oswt & run_wen;
  assign dout_rsci_biwt = dout_rsci_ogwt & dout_rsci_irdy;
  assign dout_rsci_ogwt = dout_rsci_oswt & (~ dout_rsci_bcwt);
  assign dout_rsci_ivld_run_sct = dout_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp (
  clk, arst_n, din_rsci_q_d, din_rsci_q_d_mxwt, din_rsci_biwt, din_rsci_bdwt
);
  input clk;
  input arst_n;
  input [127:0] din_rsci_q_d;
  output [127:0] din_rsci_q_d_mxwt;
  input din_rsci_biwt;
  input din_rsci_bdwt;


  // Interconnect Declarations
  reg din_rsci_bcwt;
  reg [127:0] din_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_q_d_mxwt = MUX_v_128_2_2(din_rsci_q_d, din_rsci_q_d_bfwt, din_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_bcwt <= 1'b0;
    end
    else begin
      din_rsci_bcwt <= ~((~(din_rsci_bcwt | din_rsci_biwt)) | din_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      din_rsci_q_d_bfwt <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ din_rsci_bcwt ) begin
      din_rsci_q_d_bfwt <= din_rsci_q_d_mxwt;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input [0:0] sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl (
  run_wen, run_wten, din_rsci_oswt, din_rsci_biwt, din_rsci_bdwt, din_rsci_re_d_run_sct_pff,
      din_rsci_oswt_pff
);
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output din_rsci_biwt;
  output din_rsci_bdwt;
  output din_rsci_re_d_run_sct_pff;
  input din_rsci_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign din_rsci_bdwt = din_rsci_oswt & run_wen;
  assign din_rsci_biwt = (~ run_wten) & din_rsci_oswt;
  assign din_rsci_re_d_run_sct_pff = din_rsci_oswt_pff & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [136:0] paramsIn_rsci_idat_bfwt_136_0;
  wire [136:0] paramsIn_rsci_idat_mxwt_opt_136_0;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_opt_136_0 = MUX_v_137_2_2((paramsIn_rsci_idat[136:0]),
      paramsIn_rsci_idat_bfwt_136_0, paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_opt_136_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt_136_0 <= paramsIn_rsci_idat_mxwt_opt_136_0;
    end
  end

  function automatic [136:0] MUX_v_137_2_2;
    input [136:0] input_0;
    input [136:0] input_1;
    input [0:0] sel;
    reg [136:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_137_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi (
  clk, arst_n, inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy, run_wen, inputDoubleBufferReaderParams_cnsi_oswt,
      inputDoubleBufferReaderParams_cnsi_wen_comp, inputDoubleBufferReaderParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;
  input run_wen;
  input inputDoubleBufferReaderParams_cnsi_oswt;
  output inputDoubleBufferReaderParams_cnsi_wen_comp;
  input [143:0] inputDoubleBufferReaderParams_cnsi_idat;


  // Interconnect Declarations
  wire inputDoubleBufferReaderParams_cnsi_irdy;
  wire inputDoubleBufferReaderParams_cnsi_biwt;
  wire inputDoubleBufferReaderParams_cnsi_bdwt;
  wire inputDoubleBufferReaderParams_cnsi_bcwt;
  wire inputDoubleBufferReaderParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd19),
  .width(32'sd144)) inputDoubleBufferReaderParams_cnsi (
      .irdy(inputDoubleBufferReaderParams_cnsi_irdy),
      .ivld(inputDoubleBufferReaderParams_cnsi_ivld_run_sct),
      .idat(inputDoubleBufferReaderParams_cnsi_idat),
      .rdy(inputDoubleBufferReaderParams_cns_rdy),
      .vld(inputDoubleBufferReaderParams_cns_vld),
      .dat(inputDoubleBufferReaderParams_cns_dat)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputDoubleBufferReaderParams_cnsi_oswt(inputDoubleBufferReaderParams_cnsi_oswt),
      .inputDoubleBufferReaderParams_cnsi_irdy(inputDoubleBufferReaderParams_cnsi_irdy),
      .inputDoubleBufferReaderParams_cnsi_biwt(inputDoubleBufferReaderParams_cnsi_biwt),
      .inputDoubleBufferReaderParams_cnsi_bdwt(inputDoubleBufferReaderParams_cnsi_bdwt),
      .inputDoubleBufferReaderParams_cnsi_bcwt(inputDoubleBufferReaderParams_cnsi_bcwt),
      .inputDoubleBufferReaderParams_cnsi_ivld_run_sct(inputDoubleBufferReaderParams_cnsi_ivld_run_sct)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inputDoubleBufferReaderParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferReaderParams_cnsi_oswt(inputDoubleBufferReaderParams_cnsi_oswt),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_biwt(inputDoubleBufferReaderParams_cnsi_biwt),
      .inputDoubleBufferReaderParams_cnsi_bdwt(inputDoubleBufferReaderParams_cnsi_bdwt),
      .inputDoubleBufferReaderParams_cnsi_bcwt(inputDoubleBufferReaderParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi (
  clk, arst_n, inputDoubleBufferWriterParams_cns_dat, inputDoubleBufferWriterParams_cns_vld,
      inputDoubleBufferWriterParams_cns_rdy, run_wen, inputDoubleBufferWriterParams_cnsi_oswt,
      inputDoubleBufferWriterParams_cnsi_wen_comp, inputDoubleBufferWriterParams_cnsi_idat
);
  input clk;
  input arst_n;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  input run_wen;
  input inputDoubleBufferWriterParams_cnsi_oswt;
  output inputDoubleBufferWriterParams_cnsi_wen_comp;
  input [143:0] inputDoubleBufferWriterParams_cnsi_idat;


  // Interconnect Declarations
  wire inputDoubleBufferWriterParams_cnsi_irdy;
  wire inputDoubleBufferWriterParams_cnsi_biwt;
  wire inputDoubleBufferWriterParams_cnsi_bdwt;
  wire inputDoubleBufferWriterParams_cnsi_bcwt;
  wire inputDoubleBufferWriterParams_cnsi_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd18),
  .width(32'sd144)) inputDoubleBufferWriterParams_cnsi (
      .irdy(inputDoubleBufferWriterParams_cnsi_irdy),
      .ivld(inputDoubleBufferWriterParams_cnsi_ivld_run_sct),
      .idat(inputDoubleBufferWriterParams_cnsi_idat),
      .rdy(inputDoubleBufferWriterParams_cns_rdy),
      .vld(inputDoubleBufferWriterParams_cns_vld),
      .dat(inputDoubleBufferWriterParams_cns_dat)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputDoubleBufferWriterParams_cnsi_oswt(inputDoubleBufferWriterParams_cnsi_oswt),
      .inputDoubleBufferWriterParams_cnsi_irdy(inputDoubleBufferWriterParams_cnsi_irdy),
      .inputDoubleBufferWriterParams_cnsi_biwt(inputDoubleBufferWriterParams_cnsi_biwt),
      .inputDoubleBufferWriterParams_cnsi_bdwt(inputDoubleBufferWriterParams_cnsi_bdwt),
      .inputDoubleBufferWriterParams_cnsi_bcwt(inputDoubleBufferWriterParams_cnsi_bcwt),
      .inputDoubleBufferWriterParams_cnsi_ivld_run_sct(inputDoubleBufferWriterParams_cnsi_ivld_run_sct)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp
      InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inputDoubleBufferWriterParams_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferWriterParams_cnsi_oswt(inputDoubleBufferWriterParams_cnsi_oswt),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_biwt(inputDoubleBufferWriterParams_cnsi_biwt),
      .inputDoubleBufferWriterParams_cnsi_bdwt(inputDoubleBufferWriterParams_cnsi_bdwt),
      .inputDoubleBufferWriterParams_cnsi_bcwt(inputDoubleBufferWriterParams_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd17),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj (
  clk, arst_n, dout_rsc_req_vz, run_wen, dout_rsc_req_obj_oswt, dout_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input dout_rsc_req_vz;
  input run_wen;
  input dout_rsc_req_obj_oswt;
  output dout_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire dout_rsc_req_obj_vd;
  wire dout_rsc_req_obj_biwt;
  wire dout_rsc_req_obj_bdwt;
  wire dout_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) dout_rsc_req_obj (
      .vd(dout_rsc_req_obj_vd),
      .vz(dout_rsc_req_vz)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_vd(dout_rsc_req_obj_vd),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_dout_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_obj_oswt(dout_rsc_req_obj_oswt),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp),
      .dout_rsc_req_obj_biwt(dout_rsc_req_obj_biwt),
      .dout_rsc_req_obj_bdwt(dout_rsc_req_obj_bdwt),
      .dout_rsc_req_obj_bcwt(dout_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj (
  dout_rsc_rls_lz, run_wten, dout_rsc_rls_obj_iswt0
);
  output dout_rsc_rls_lz;
  input run_wten;
  input dout_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire dout_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) dout_rsc_rls_obj (
      .ld(dout_rsc_rls_obj_ld_run_sct),
      .lz(dout_rsc_rls_lz)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_dout_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(dout_rsc_rls_obj_iswt0),
      .dout_rsc_rls_obj_ld_run_sct(dout_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_dout_rsci_1
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_dout_rsci_1 (
  dout_rsci_we_d_pff, dout_rsci_iswt0_pff, run_wten_pff
);
  output dout_rsci_we_d_pff;
  input dout_rsci_iswt0_pff;
  input run_wten_pff;


  // Interconnect Declarations
  wire dout_rsci_we_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_dout_rsc_wait_ctrl_inst
      (
      .dout_rsci_we_d_run_sct_pff(dout_rsci_we_d_run_sct_iff),
      .dout_rsci_iswt0_pff(dout_rsci_iswt0_pff),
      .run_wten_pff(run_wten_pff)
    );
  assign dout_rsci_we_d_pff = dout_rsci_we_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_din_rsci
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_din_rsci (
  clk, arst_n, din_rsc_dat, din_rsc_vld, din_rsc_rdy, run_wen, din_rsci_oswt, din_rsci_wen_comp,
      din_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input run_wen;
  input din_rsci_oswt;
  output din_rsci_wen_comp;
  output [15:0] din_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_bcwt;
  wire din_rsci_irdy_run_sct;
  wire din_rsci_ivld;
  wire [15:0] din_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd16)) din_rsci (
      .rdy(din_rsc_rdy),
      .vld(din_rsc_vld),
      .dat(din_rsc_dat),
      .irdy(din_rsci_irdy_run_sct),
      .ivld(din_rsci_ivld),
      .idat(din_rsci_idat)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_irdy_run_sct(din_rsci_irdy_run_sct),
      .din_rsci_ivld(din_rsci_ivld)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp InputDoubleBufferWriter_512_16_16_run_din_rsci_din_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_bcwt(din_rsci_bcwt),
      .din_rsci_idat(din_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [136:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj (
  clk, arst_n, din_rsc_req_vz, run_wen, din_rsc_req_obj_oswt, din_rsc_req_obj_wen_comp
);
  input clk;
  input arst_n;
  input din_rsc_req_vz;
  input run_wen;
  input din_rsc_req_obj_oswt;
  output din_rsc_req_obj_wen_comp;


  // Interconnect Declarations
  wire din_rsc_req_obj_vd;
  wire din_rsc_req_obj_biwt;
  wire din_rsc_req_obj_bdwt;
  wire din_rsc_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_sync_v2 #(.valid(32'sd1)) din_rsc_req_obj (
      .vd(din_rsc_req_obj_vd),
      .vz(din_rsc_req_vz)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_vd(din_rsc_req_obj_vd),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_din_rsc_req_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_obj_oswt(din_rsc_req_obj_oswt),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp),
      .din_rsc_req_obj_biwt(din_rsc_req_obj_biwt),
      .din_rsc_req_obj_bdwt(din_rsc_req_obj_bdwt),
      .din_rsc_req_obj_bcwt(din_rsc_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj (
  din_rsc_rls_lz, run_wten, din_rsc_rls_obj_iswt0
);
  output din_rsc_rls_lz;
  input run_wten;
  input din_rsc_rls_obj_iswt0;


  // Interconnect Declarations
  wire din_rsc_rls_obj_ld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) din_rsc_rls_obj (
      .ld(din_rsc_rls_obj_ld_run_sct),
      .lz(din_rsc_rls_lz)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_din_rsc_rls_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(din_rsc_rls_obj_iswt0),
      .din_rsc_rls_obj_ld_run_sct(din_rsc_rls_obj_ld_run_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_dout_rsci
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_dout_rsci (
  clk, arst_n, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, run_wen, dout_rsci_oswt,
      dout_rsci_wen_comp, dout_rsci_idat
);
  input clk;
  input arst_n;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  input run_wen;
  input dout_rsci_oswt;
  output dout_rsci_wen_comp;
  input [127:0] dout_rsci_idat;


  // Interconnect Declarations
  wire dout_rsci_irdy;
  wire dout_rsci_biwt;
  wire dout_rsci_bdwt;
  wire dout_rsci_bcwt;
  wire dout_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd128)) dout_rsci (
      .irdy(dout_rsci_irdy),
      .ivld(dout_rsci_ivld_run_sct),
      .idat(dout_rsci_idat),
      .rdy(dout_rsc_rdy),
      .vld(dout_rsc_vld),
      .dat(dout_rsc_dat)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_irdy(dout_rsci_irdy),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt),
      .dout_rsci_ivld_run_sct(dout_rsci_ivld_run_sct)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp InputDoubleBufferReader_512_16_16_run_dout_rsci_dout_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsci_oswt(dout_rsci_oswt),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_biwt(dout_rsci_biwt),
      .dout_rsci_bdwt(dout_rsci_bdwt),
      .dout_rsci_bcwt(dout_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_din_rsci_1
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_din_rsci_1 (
  clk, arst_n, din_rsci_q_d, run_wen, run_wten, din_rsci_oswt, din_rsci_q_d_mxwt,
      din_rsci_re_d_pff, din_rsci_oswt_pff
);
  input clk;
  input arst_n;
  input [127:0] din_rsci_q_d;
  input run_wen;
  input run_wten;
  input din_rsci_oswt;
  output [127:0] din_rsci_q_d_mxwt;
  output din_rsci_re_d_pff;
  input din_rsci_oswt_pff;


  // Interconnect Declarations
  wire din_rsci_biwt;
  wire din_rsci_bdwt;
  wire din_rsci_re_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(din_rsci_oswt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt),
      .din_rsci_re_d_run_sct_pff(din_rsci_re_d_run_sct_iff),
      .din_rsci_oswt_pff(din_rsci_oswt_pff)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp InputDoubleBufferReader_512_16_16_run_din_rsci_1_din_rsc_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_q_d(din_rsci_q_d),
      .din_rsci_q_d_mxwt(din_rsci_q_d_mxwt),
      .din_rsci_biwt(din_rsci_biwt),
      .din_rsci_bdwt(din_rsci_bdwt)
    );
  assign din_rsci_re_d_pff = din_rsci_re_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run_paramsIn_rsci
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [136:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;
  wire [136:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run_run
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, inputDoubleBufferWriterParams_cns_dat,
      inputDoubleBufferWriterParams_cns_vld, inputDoubleBufferWriterParams_cns_rdy,
      inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire inputDoubleBufferWriterParams_cnsi_wen_comp;
  wire inputDoubleBufferReaderParams_cnsi_wen_comp;
  wire [2:0] fsm_output;
  reg reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse;
  reg [143:0] reg_inputDoubleBufferReaderParams_cnsi_idat_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci InputDoubleBuffer_512_16_16_run_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferWriterParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy),
      .run_wen(run_wen),
      .inputDoubleBufferWriterParams_cnsi_oswt(reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_idat(reg_inputDoubleBufferReaderParams_cnsi_idat_cse)
    );
  InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi InputDoubleBuffer_512_16_16_run_run_inputDoubleBufferReaderParams_cnsi_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld),
      .inputDoubleBufferReaderParams_cns_rdy(inputDoubleBufferReaderParams_cns_rdy),
      .run_wen(run_wen),
      .inputDoubleBufferReaderParams_cnsi_oswt(reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_idat(reg_inputDoubleBufferReaderParams_cnsi_idat_cse)
    );
  InputDoubleBuffer_512_16_16_run_run_staller InputDoubleBuffer_512_16_16_run_run_staller_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .inputDoubleBufferWriterParams_cnsi_wen_comp(inputDoubleBufferWriterParams_cnsi_wen_comp),
      .inputDoubleBufferReaderParams_cnsi_wen_comp(inputDoubleBufferReaderParams_cnsi_wen_comp)
    );
  InputDoubleBuffer_512_16_16_run_run_run_fsm InputDoubleBuffer_512_16_16_run_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputDoubleBufferReaderParams_cnsi_idat_cse <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      reg_inputDoubleBufferReaderParams_cnsi_idat_cse <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_inputDoubleBufferReaderParams_cnsi_ivld_run_psct_cse <= fsm_output[1];
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~ (fsm_output[1]);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_req_vz, dout_rsc_rls_lz, dout_rsci_wadr_d,
      dout_rsci_d_d, dout_rsci_we_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;
  output [8:0] dout_rsci_wadr_d;
  wire [9:0] nl_dout_rsci_wadr_d;
  output [127:0] dout_rsci_d_d;
  output dout_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [136:0] paramsIn_rsci_idat_mxwt;
  wire din_rsci_wen_comp;
  wire [15:0] din_rsci_idat_mxwt;
  wire dout_rsc_req_obj_wen_comp;
  wire [14:0] fsm_output;
  wire [3:0] while_while_for_for_acc_1_tmp;
  wire [4:0] nl_while_while_for_for_acc_1_tmp;
  wire or_dcpl_7;
  wire or_dcpl_8;
  wire or_dcpl_10;
  wire or_dcpl_11;
  wire or_dcpl_13;
  wire or_dcpl_20;
  wire or_dcpl_21;
  wire and_dcpl_19;
  wire or_dcpl_25;
  wire or_dcpl_26;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_31;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_35;
  reg operator_32_false_1_slc_33_svs;
  wire exit_while_sva_mx0;
  reg [2:0] while_while_for_for_ic0_idx_3_0_sva_2_0;
  reg reg_dout_rsc_req_obj_iswt0_cse;
  reg reg_dout_rsc_rls_obj_ld_run_psct_cse;
  reg reg_din_rsci_irdy_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire dout_rsci_we_d_iff;
  reg [8:0] block_size_acc_itm;
  reg [8:0] operator_16_false_1_acc_itm;
  reg [15:0] while_while_for_for_tmp_value_sva;
  reg [7:0] while_while_for_column_value_13_sva;
  reg [7:0] while_while_for_column_value_12_sva;
  reg [7:0] while_while_for_column_value_11_sva;
  reg [7:0] while_while_for_column_value_10_sva;
  reg [7:0] while_while_for_column_value_9_sva;
  reg [7:0] while_while_for_column_value_8_sva;
  reg [7:0] while_while_for_column_value_7_sva;
  reg [7:0] while_while_for_column_value_6_sva;
  reg [7:0] while_while_for_column_value_5_sva;
  reg [7:0] while_while_for_column_value_4_sva;
  reg [7:0] while_while_for_column_value_3_sva;
  reg [7:0] while_while_for_column_value_2_sva;
  reg [7:0] while_while_for_column_value_1_sva;
  reg [7:0] while_while_for_column_value_0_sva;
  reg [8:0] block_size_sva;
  reg [31:0] total_blocks_lpi_3;
  reg [136:0] paramsIn_crt_sva_136_0;
  wire [8:0] while_while_for_idx_sva_2;
  wire [9:0] nl_while_while_for_idx_sva_2;
  wire while_while_for_column_value_and_cse;
  wire while_while_for_column_value_and_2_cse;
  wire while_while_for_column_value_and_1_cse;
  wire while_while_for_column_value_and_4_cse;
  wire while_while_for_column_value_and_3_cse;
  wire while_while_for_column_value_and_6_cse;
  wire while_while_for_column_value_and_5_cse;
  wire operator_32_false_1_acc_1_itm_32_1;
  wire while_while_for_acc_2_itm_9_1;

  wire[8:0] block_size_mux1h_1_nl;
  wire[8:0] block_size_acc_nl;
  wire[9:0] nl_block_size_acc_nl;
  wire[8:0] block_size_mul_2_nl;
  wire signed [18:0] nl_block_size_mul_2_nl;
  wire[8:0] operator_16_false_acc_nl;
  wire[9:0] nl_operator_16_false_acc_nl;
  wire[8:0] block_size_mul_1_nl;
  wire signed [18:0] nl_block_size_mul_1_nl;
  wire[8:0] while_while_acc_1_nl;
  wire[9:0] nl_while_while_acc_1_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_7_nl;
  wire[8:0] operator_16_false_1_mux1h_4_nl;
  wire[8:0] operator_16_false_1_acc_nl;
  wire[9:0] nl_operator_16_false_1_acc_nl;
  wire[9:0] while_while_aelse_acc_1_nl;
  wire[10:0] nl_while_while_aelse_acc_1_nl;
  wire[0:0] or_55_nl;
  wire[0:0] not_71_nl;
  wire[8:0] block_size_acc_1_nl;
  wire[9:0] nl_block_size_acc_1_nl;
  wire[8:0] block_size_mul_3_nl;
  wire signed [18:0] nl_block_size_mul_3_nl;
  wire[8:0] block_size_mul_nl;
  wire signed [18:0] nl_block_size_mul_nl;
  wire[31:0] total_blocks_mul_nl;
  wire[31:0] while_while_acc_nl;
  wire[32:0] nl_while_while_acc_nl;
  wire[9:0] while_while_for_acc_3_nl;
  wire[11:0] nl_while_while_for_acc_3_nl;
  wire[32:0] operator_32_false_1_acc_1_nl;
  wire[33:0] nl_operator_32_false_1_acc_1_nl;
  wire[9:0] while_while_aelse_acc_nl;
  wire[10:0] nl_while_while_aelse_acc_nl;
  wire[9:0] while_while_for_acc_2_nl;
  wire[10:0] nl_while_while_for_acc_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff;
  assign nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff
      = fsm_output[11];
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff;
  assign nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff =
      ~ run_wen;
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0;
  assign nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0
      = ~ while_while_for_acc_2_itm_9_1;
  wire [0:0] nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0;
  assign nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0
      = while_while_for_for_acc_1_tmp[3];
  InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci InputDoubleBufferWriter_512_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBufferWriter_512_16_16_run_din_rsci InputDoubleBufferWriter_512_16_16_run_din_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .run_wen(run_wen),
      .din_rsci_oswt(reg_din_rsci_irdy_run_psct_cse),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .din_rsci_idat_mxwt(din_rsci_idat_mxwt)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsci_1 InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst
      (
      .dout_rsci_we_d_pff(dout_rsci_we_d_iff),
      .dout_rsci_iswt0_pff(nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_dout_rsci_iswt0_pff[0:0]),
      .run_wten_pff(nl_InputDoubleBufferWriter_512_16_16_run_dout_rsci_1_inst_run_wten_pff[0:0])
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj InputDoubleBufferWriter_512_16_16_run_dout_rsc_rls_obj_inst
      (
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .run_wten(run_wten),
      .dout_rsc_rls_obj_iswt0(reg_dout_rsc_rls_obj_ld_run_psct_cse)
    );
  InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj InputDoubleBufferWriter_512_16_16_run_dout_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .run_wen(run_wen),
      .dout_rsc_req_obj_oswt(reg_dout_rsc_req_obj_iswt0_cse),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferWriter_512_16_16_run_staller InputDoubleBufferWriter_512_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .din_rsci_wen_comp(din_rsci_wen_comp),
      .dout_rsc_req_obj_wen_comp(dout_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferWriter_512_16_16_run_run_fsm InputDoubleBufferWriter_512_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_4_tr0(exit_while_sva_mx0),
      .while_while_C_1_tr0(or_dcpl_20),
      .while_while_C_2_tr0(nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_C_2_tr0[0:0]),
      .while_while_for_for_C_0_tr0(nl_InputDoubleBufferWriter_512_16_16_run_run_fsm_inst_while_while_for_for_C_0_tr0[0:0]),
      .while_while_for_C_1_tr0(operator_32_false_1_slc_33_svs),
      .while_C_1_tr0(exit_while_sva_mx0)
    );
  assign while_while_for_column_value_and_cse = run_wen & (or_dcpl_8 | or_dcpl_7);
  assign while_while_for_column_value_and_1_cse = run_wen & (or_dcpl_11 | or_dcpl_10);
  assign while_while_for_column_value_and_2_cse = run_wen & (or_dcpl_8 | or_dcpl_13);
  assign while_while_for_column_value_and_3_cse = run_wen & (or_dcpl_11 | or_dcpl_13);
  assign while_while_for_column_value_and_4_cse = run_wen & (or_dcpl_8 | or_dcpl_10);
  assign while_while_for_column_value_and_5_cse = run_wen & (or_dcpl_11 | or_dcpl_7);
  assign while_while_for_column_value_and_6_cse = run_wen & (or_dcpl_8 | (while_while_for_for_acc_1_tmp[1:0]!=2'b11));
  assign nl_while_while_for_idx_sva_2 = operator_16_false_1_acc_itm + 9'b000000001;
  assign while_while_for_idx_sva_2 = nl_while_while_for_idx_sva_2[8:0];
  assign exit_while_sva_mx0 = MUX_s_1_2_2((~ operator_32_false_1_slc_33_svs), (~
      operator_32_false_1_acc_1_itm_32_1), fsm_output[14]);
  assign nl_while_while_for_for_acc_1_tmp = conv_u2s_3_4(while_while_for_for_ic0_idx_3_0_sva_2_0)
      + 4'b0001;
  assign while_while_for_for_acc_1_tmp = nl_while_while_for_for_acc_1_tmp[3:0];
  assign nl_operator_32_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_1_acc_1_nl = nl_operator_32_false_1_acc_1_nl[32:0];
  assign operator_32_false_1_acc_1_itm_32_1 = readslicef_33_1_32((operator_32_false_1_acc_1_nl));
  assign or_dcpl_7 = (while_while_for_for_acc_1_tmp[1:0]!=2'b00);
  assign or_dcpl_8 = (while_while_for_for_acc_1_tmp[3:2]!=2'b00);
  assign or_dcpl_10 = (while_while_for_for_acc_1_tmp[1:0]!=2'b10);
  assign or_dcpl_11 = (while_while_for_for_acc_1_tmp[3:2]!=2'b01);
  assign or_dcpl_13 = (while_while_for_for_acc_1_tmp[1:0]!=2'b01);
  assign nl_while_while_aelse_acc_nl = conv_u2u_9_10(operator_16_false_1_acc_itm)
      + 10'b1100000001;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[9:0];
  assign or_dcpl_20 = (~ operator_32_false_1_slc_33_svs) | (readslicef_10_1_9((while_while_aelse_acc_nl)));
  assign or_dcpl_21 = (fsm_output[5]) | (fsm_output[14]);
  assign and_dcpl_19 = ~((fsm_output[0]) | (fsm_output[2]));
  assign or_dcpl_25 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b00);
  assign or_dcpl_26 = or_dcpl_25 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_27 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b10);
  assign or_dcpl_28 = or_dcpl_27 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_29 = (while_while_for_for_ic0_idx_3_0_sva_2_0[1:0]!=2'b01);
  assign or_dcpl_30 = or_dcpl_29 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_31 = or_dcpl_29 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_32 = or_dcpl_27 | (while_while_for_for_ic0_idx_3_0_sva_2_0[2]);
  assign or_dcpl_33 = or_dcpl_25 | (~ (while_while_for_for_ic0_idx_3_0_sva_2_0[2]));
  assign or_dcpl_35 = (while_while_for_for_ic0_idx_3_0_sva_2_0!=3'b011);
  assign nl_while_while_for_acc_2_nl = ({1'b1 , (~ block_size_sva)}) + 10'b0000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[9:0];
  assign while_while_for_acc_2_itm_9_1 = readslicef_10_1_9((while_while_for_acc_2_nl));
  assign nl_dout_rsci_wadr_d = block_size_acc_itm + operator_16_false_1_acc_itm;
  assign dout_rsci_wadr_d = nl_dout_rsci_wadr_d[8:0];
  assign dout_rsci_d_d = {while_while_for_for_tmp_value_sva , while_while_for_column_value_13_sva
      , while_while_for_column_value_12_sva , while_while_for_column_value_11_sva
      , while_while_for_column_value_10_sva , while_while_for_column_value_9_sva
      , while_while_for_column_value_8_sva , while_while_for_column_value_7_sva ,
      while_while_for_column_value_6_sva , while_while_for_column_value_5_sva , while_while_for_column_value_4_sva
      , while_while_for_column_value_3_sva , while_while_for_column_value_2_sva ,
      while_while_for_column_value_1_sva , while_while_for_column_value_0_sva};
  assign dout_rsci_we_d_pff = dout_rsci_we_d_iff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_din_rsci_irdy_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      block_size_acc_itm <= 9'b000000000;
      operator_16_false_1_acc_itm <= 9'b000000000;
      operator_32_false_1_slc_33_svs <= 1'b0;
      while_while_for_for_ic0_idx_3_0_sva_2_0 <= 3'b000;
    end
    else if ( run_wen ) begin
      reg_dout_rsc_req_obj_iswt0_cse <= (~ exit_while_sva_mx0) & or_dcpl_21;
      reg_dout_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_20 & (fsm_output[8]);
      reg_din_rsci_irdy_run_psct_cse <= (while_while_for_acc_2_itm_9_1 & (fsm_output[9]))
          | ((~ (while_while_for_for_acc_1_tmp[3])) & (fsm_output[10])) | ((~ operator_32_false_1_slc_33_svs)
          & (fsm_output[12]));
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[0]) | (fsm_output[5])
          | (fsm_output[14]))) | (~(exit_while_sva_mx0 | (fsm_output[0]))));
      block_size_acc_itm <= MUX_v_9_2_2(9'b000000000, (block_size_mux1h_1_nl), (nor_7_nl));
      operator_16_false_1_acc_itm <= MUX_v_9_2_2(9'b000000000, (operator_16_false_1_mux1h_4_nl),
          (not_71_nl));
      operator_32_false_1_slc_33_svs <= MUX_s_1_2_2(operator_32_false_1_acc_1_itm_32_1,
          (~ (readslicef_10_1_9((while_while_for_acc_3_nl)))), fsm_output[11]);
      while_while_for_for_ic0_idx_3_0_sva_2_0 <= MUX_v_3_2_2(3'b000, (while_while_for_for_acc_1_tmp[2:0]),
          (fsm_output[10]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_sva_136_0 <= 137'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      paramsIn_crt_sva_136_0 <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_sva <= 9'b000000000;
    end
    else if ( run_wen & ((~(and_dcpl_19 & (~ (fsm_output[1])))) | (fsm_output[5]))
        ) begin
      block_size_sva <= MUX_v_9_2_2((block_size_acc_1_nl), (block_size_mul_nl), fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & ((~ and_dcpl_19) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[13]))
        ) begin
      total_blocks_lpi_3 <= MUX_v_32_2_2((total_blocks_mul_nl), (while_while_acc_nl),
          fsm_output[13]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_1_sva <= 8'b00000000;
      while_while_for_column_value_0_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_cse ) begin
      while_while_for_column_value_1_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_1_sva, or_dcpl_26);
      while_while_for_column_value_0_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_0_sva, or_dcpl_26);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_13_sva <= 8'b00000000;
      while_while_for_column_value_12_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_1_cse ) begin
      while_while_for_column_value_13_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_13_sva, or_dcpl_28);
      while_while_for_column_value_12_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_12_sva, or_dcpl_28);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_3_sva <= 8'b00000000;
      while_while_for_column_value_2_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_2_cse ) begin
      while_while_for_column_value_3_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_3_sva, or_dcpl_30);
      while_while_for_column_value_2_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_2_sva, or_dcpl_30);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_11_sva <= 8'b00000000;
      while_while_for_column_value_10_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_3_cse ) begin
      while_while_for_column_value_11_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_11_sva, or_dcpl_31);
      while_while_for_column_value_10_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_10_sva, or_dcpl_31);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_5_sva <= 8'b00000000;
      while_while_for_column_value_4_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_4_cse ) begin
      while_while_for_column_value_5_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_5_sva, or_dcpl_32);
      while_while_for_column_value_4_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_4_sva, or_dcpl_32);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_9_sva <= 8'b00000000;
      while_while_for_column_value_8_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_5_cse ) begin
      while_while_for_column_value_9_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_9_sva, or_dcpl_33);
      while_while_for_column_value_8_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_8_sva, or_dcpl_33);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_column_value_7_sva <= 8'b00000000;
      while_while_for_column_value_6_sva <= 8'b00000000;
    end
    else if ( while_while_for_column_value_and_6_cse ) begin
      while_while_for_column_value_7_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[15:8]),
          while_while_for_column_value_7_sva, or_dcpl_35);
      while_while_for_column_value_6_sva <= MUX_v_8_2_2((din_rsci_idat_mxwt[7:0]),
          while_while_for_column_value_6_sva, or_dcpl_35);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_tmp_value_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (while_while_for_for_acc_1_tmp[3]) ) begin
      while_while_for_for_tmp_value_sva <= din_rsci_idat_mxwt;
    end
  end
  assign nl_operator_16_false_acc_nl = (paramsIn_rsci_idat_mxwt[56:48]) + 9'b111111111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[8:0];
  assign nl_block_size_mul_2_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[136:128]))
      * $signed((operator_16_false_acc_nl));
  assign block_size_mul_2_nl = nl_block_size_mul_2_nl[8:0];
  assign nl_block_size_acc_nl = (block_size_mul_2_nl) + (paramsIn_rsci_idat_mxwt[104:96]);
  assign block_size_acc_nl = nl_block_size_acc_nl[8:0];
  assign nl_block_size_mul_1_nl = $signed(conv_u2s_9_10(paramsIn_crt_sva_136_0[88:80]))
      * $signed(block_size_acc_itm);
  assign block_size_mul_1_nl = nl_block_size_mul_1_nl[8:0];
  assign nl_while_while_acc_1_nl = block_size_acc_itm + block_size_sva;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[8:0];
  assign nor_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[13]) | (fsm_output[5]) | (fsm_output[14]));
  assign block_size_mux1h_1_nl = MUX1HOT_v_9_4_2((block_size_acc_nl), (block_size_mul_1_nl),
      block_size_acc_itm, (while_while_acc_1_nl), {(fsm_output[1]) , (fsm_output[4])
      , (nor_nl) , (fsm_output[13])});
  assign nor_7_nl = ~((fsm_output[0]) | (fsm_output[6]) | or_dcpl_21);
  assign nl_operator_16_false_1_acc_nl = (paramsIn_rsci_idat_mxwt[40:32]) + 9'b111111111;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[8:0];
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_9_10(~ block_size_acc_itm) + conv_u2u_9_10(~
      block_size_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[9:0];
  assign or_55_nl = (fsm_output[10]) | (fsm_output[12]);
  assign operator_16_false_1_mux1h_4_nl = MUX1HOT_v_9_4_2((operator_16_false_1_acc_nl),
      (readslicef_10_9_1((while_while_aelse_acc_1_nl))), while_while_for_idx_sva_2,
      operator_16_false_1_acc_itm, {(fsm_output[1]) , (fsm_output[7]) , (fsm_output[11])
      , (or_55_nl)});
  assign not_71_nl = ~ (fsm_output[9]);
  assign nl_while_while_for_acc_3_nl = ({1'b1 , while_while_for_idx_sva_2}) + conv_u2u_9_10(~
      block_size_sva) + 10'b0000000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[9:0];
  assign nl_block_size_mul_3_nl = $signed(conv_u2s_9_10(paramsIn_crt_sva_136_0[136:128]))
      * $signed(operator_16_false_1_acc_itm);
  assign block_size_mul_3_nl = nl_block_size_mul_3_nl[8:0];
  assign nl_block_size_acc_1_nl = (block_size_mul_3_nl) + (paramsIn_crt_sva_136_0[120:112]);
  assign block_size_acc_1_nl = nl_block_size_acc_1_nl[8:0];
  assign nl_block_size_mul_nl = $signed(block_size_acc_itm) * $signed(conv_u2s_9_10(block_size_sva));
  assign block_size_mul_nl = nl_block_size_mul_nl[8:0];
  assign total_blocks_mul_nl = conv_u2u_32_32((paramsIn_crt_sva_136_0[31:16]) * (paramsIn_crt_sva_136_0[15:0]));
  assign nl_while_while_acc_nl = total_blocks_lpi_3 + 32'b11111111111111111111111111111111;
  assign while_while_acc_nl = nl_while_while_acc_nl[31:0];

  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_req_vz,
      din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld, dout_rsc_rdy, din_rsci_radr_d,
      din_rsci_q_d, din_rsci_re_d_pff
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;
  output [8:0] din_rsci_radr_d;
  wire [10:0] nl_din_rsci_radr_d;
  input [127:0] din_rsci_q_d;
  output din_rsci_re_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire paramsIn_rsci_wen_comp;
  wire [136:0] paramsIn_rsci_idat_mxwt;
  wire [127:0] din_rsci_q_d_mxwt;
  wire dout_rsci_wen_comp;
  reg [127:0] dout_rsci_idat;
  wire din_rsc_req_obj_wen_comp;
  wire [8:0] fsm_output;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire or_tmp_1;
  wire mux_tmp_2;
  wire mux_tmp_3;
  wire or_dcpl_8;
  wire and_dcpl_56;
  wire or_dcpl_23;
  wire or_dcpl_32;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_tmp_23;
  wire or_tmp_44;
  reg lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7;
  reg exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4;
  reg lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6;
  reg exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4;
  reg lfst_exitL_exit_while_while_for_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7;
  reg exitL_exitL_exit_while_while_for_for_for_for_lpi_2;
  reg lfst_exit_while_while_for_for_for_lpi_2;
  wire lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3;
  reg lfst_exitL_exit_while_while_for_for_for_lpi_2;
  wire exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6;
  reg exitL_exitL_exit_while_while_for_for_for_lpi_2;
  reg exitL_exit_while_while_for_for_sva;
  reg lfst_exit_while_while_for_for_lpi_2;
  reg while_while_for_for_asn_sft_lpi_4_dfm_st_1;
  reg exit_while_while_for_lpi_4_dfm_1;
  reg while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
  reg while_while_for_for_for_asn_sft_lpi_4_dfm_st_1;
  wire exit_while_while_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire exit_while_while_for_lpi_4_dfm_mx0w1;
  wire exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  wire while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  reg while_while_for_asn_4_itm_1;
  reg while_while_for_stage_0_2;
  reg while_while_for_stage_0_3;
  reg while_while_for_for_for_for_for_asn_sft_lpi_4;
  reg while_while_for_for_for_for_asn_sft_lpi_4;
  reg while_while_for_for_for_asn_sft_lpi_4;
  reg while_while_for_for_asn_sft_lpi_4;
  reg while_while_for_for_for_asn_sft_lpi_4_dfm_st_2;
  reg while_while_for_for_asn_sft_lpi_4_dfm_st_2;
  reg exit_while_while_for_lpi_4_dfm_st_2;
  reg while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_2;
  reg while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_2;
  reg while_while_for_for_for_for_for_for_not_mdf_sva_st_2;
  reg while_while_for_for_for_for_for_for_not_mdf_sva_st_1;
  wire [15:0] while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7;
  wire [15:0] while_while_for_for_for_for_for_x_idx_lpi_4_dfm_mx0w1;
  wire [15:0] while_while_for_for_for_for_wy_idx_lpi_4_dfm_6;
  wire lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0;
  wire and_93_m1c;
  reg [104:0] reg_paramsIn_crt_sva_136_0_ftd;
  reg reg_din_rsc_req_obj_iswt0_cse;
  reg reg_din_rsc_rls_obj_ld_run_psct_cse;
  reg reg_dout_rsci_ivld_run_psct_cse;
  reg reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire while_while_for_for_for_and_cse;
  reg reg_while_while_for_stage_0_cse;
  wire nor_12_cse;
  wire while_while_for_for_for_and_7_cse;
  wire while_while_for_for_for_for_and_3_cse;
  wire while_while_for_for_for_for_for_and_3_cse;
  wire while_while_aelse_while_while_aelse_and_cse;
  wire din_rsci_re_d_iff;
  wire and_103_rmff;
  reg [15:0] while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1;
  reg [8:0] while_while_for_for_for_for_for_for_slc_while_while_for_for_for_for_wy_idx_8_0_itm_1;
  reg [8:0] while_while_for_for_for_for_for_for_address_mul_itm_1;
  wire [17:0] nl_while_while_for_for_for_for_for_for_address_mul_itm_1;
  reg [8:0] operator_16_false_acc_itm;
  reg [8:0] while_while_for_for_for_for_for_for_address_mul_5_itm_1;
  wire signed [18:0] nl_while_while_for_for_for_for_for_for_address_mul_5_itm_1;
  reg [8:0] block_size_acc_cse_sva;
  reg [8:0] block_size_acc_1_cse_sva;
  wire [9:0] nl_block_size_acc_1_cse_sva;
  reg [8:0] block_size_sva;
  wire signed [17:0] nl_block_size_sva;
  reg [31:0] total_blocks_lpi_3;
  reg [8:0] while_current_buffer_size_sva;
  reg [8:0] while_block_count_8_0_sva;
  reg [15:0] while_while_for_for_co_idx_lpi_4;
  reg [15:0] while_while_for_for_for_wx_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_wy_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_for_x_idx_lpi_4;
  reg [15:0] while_while_for_for_for_for_for_for_y_idx_lpi_4;
  reg [15:0] while_while_for_koo_idx_sva;
  wire lfst_exit_while_while_for_for_lpi_2_mx0c1;
  wire [8:0] block_size_acc_cse_sva_1;
  wire [9:0] nl_block_size_acc_cse_sva_1;
  wire exit_while_while_for_for_lpi_4_dfm_mx1w0;
  wire while_while_for_for_for_or_tmp_1;
  wire while_while_for_for_or_3_tmp_1;
  wire exit_while_while_for_for_for_lpi_4_dfm_1;
  wire lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5;
  wire [15:0] while_while_for_for_for_wx_idx_lpi_4_dfm_5;
  wire [15:0] while_while_for_for_co_idx_lpi_4_dfm_1_mx0;
  wire exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
  wire exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
  wire while_while_for_and_1_cse;
  wire block_size_and_1_cse;
  wire mux_tmp;
  wire mux_tmp_9;
  wire and_184_cse;
  wire nor_32_cse;
  wire or_121_cse;
  wire and_181_cse;
  wire [15:0] while_while_for_for_for_for_for_acc_1_itm;
  wire [16:0] nl_while_while_for_for_for_for_for_acc_1_itm;
  wire while_while_for_for_for_while_while_for_for_for_nor_1_itm;
  wire while_while_for_for_for_for_for_for_acc_2_itm_16;
  wire while_while_for_for_for_for_for_acc_2_itm_16;
  wire while_while_for_for_for_for_acc_2_itm_16;
  wire while_while_for_for_for_acc_2_itm_16;
  wire while_while_for_for_acc_3_itm_16;
  wire while_while_for_acc_3_itm_16;
  wire operator_32_false_1_acc_1_itm_32_1;

  wire[8:0] block_size_mul_3_nl;
  wire signed [18:0] nl_block_size_mul_3_nl;
  wire[8:0] operator_16_false_1_acc_nl;
  wire[9:0] nl_operator_16_false_1_acc_nl;
  wire[8:0] operator_16_false_acc_nl;
  wire[9:0] nl_operator_16_false_acc_nl;
  wire[9:0] while_while_aelse_acc_1_nl;
  wire[10:0] nl_while_while_aelse_acc_1_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_1_nl;
  wire signed [17:0] nl_while_while_for_for_for_for_for_for_address_mul_1_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_2_nl;
  wire signed [18:0] nl_while_while_for_for_for_for_for_for_address_mul_2_nl;
  wire[31:0] total_blocks_mul_nl;
  wire[31:0] while_while_acc_1_nl;
  wire[32:0] nl_while_while_acc_1_nl;
  wire[8:0] block_size_mul_1_nl;
  wire signed [18:0] nl_block_size_mul_1_nl;
  wire[8:0] while_while_acc_2_nl;
  wire[9:0] nl_while_while_acc_2_nl;
  wire[0:0] while_current_buffer_size_not_1_nl;
  wire[8:0] while_while_acc_nl;
  wire[9:0] nl_while_while_acc_nl;
  wire[0:0] while_block_count_not_nl;
  wire[15:0] while_while_for_acc_2_nl;
  wire[16:0] nl_while_while_for_acc_2_nl;
  wire[0:0] while_while_for_mux_4_nl;
  wire[15:0] while_while_for_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_and_7_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] and_197_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_30_nl;
  wire[15:0] while_while_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_for_wx_idx_and_1_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] nor_41_nl;
  wire[0:0] nor_42_nl;
  wire[0:0] and_199_nl;
  wire[0:0] or_120_nl;
  wire[0:0] and_200_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] nor_9_nl;
  wire[15:0] while_while_for_for_acc_2_nl;
  wire[16:0] nl_while_while_for_for_acc_2_nl;
  wire[0:0] while_while_for_for_and_10_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_6_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_6_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_6_nl;
  wire[17:0] nl_while_while_for_for_for_for_for_for_address_mul_6_nl;
  wire[8:0] block_size_mul_2_nl;
  wire signed [18:0] nl_block_size_mul_2_nl;
  wire[15:0] while_while_for_for_for_for_for_x_idx_mux_nl;
  wire[0:0] while_while_for_for_for_for_for_x_idx_and_nl;
  wire[15:0] while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_mux1h_nl;
  wire[15:0] while_while_for_for_for_for_for_for_acc_1_nl;
  wire[16:0] nl_while_while_for_for_for_for_for_for_acc_1_nl;
  wire[0:0] while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_nl;
  wire[0:0] while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_1_nl;
  wire[0:0] while_while_for_for_for_for_for_for_y_idx_or_nl;
  wire[16:0] while_while_for_for_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_for_for_acc_2_nl;
  wire[0:0] or_48_nl;
  wire[0:0] or_56_nl;
  wire[16:0] while_while_for_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_for_acc_2_nl;
  wire[18:0] nl_while_while_for_for_for_acc_2_nl;
  wire[16:0] while_while_for_for_acc_3_nl;
  wire[18:0] nl_while_while_for_for_acc_3_nl;
  wire[0:0] while_while_for_for_mux_60_nl;
  wire[16:0] while_while_for_acc_3_nl;
  wire[18:0] nl_while_while_for_acc_3_nl;
  wire[32:0] operator_32_false_1_acc_1_nl;
  wire[33:0] nl_operator_32_false_1_acc_1_nl;
  wire[0:0] and_82_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] or_7_nl;
  wire[9:0] while_while_aelse_acc_nl;
  wire[10:0] nl_while_while_aelse_acc_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_acc_9_nl;
  wire[9:0] nl_while_while_for_for_for_for_for_for_address_acc_9_nl;
  wire[8:0] while_while_for_for_for_for_for_for_address_mul_8_nl;
  wire[17:0] nl_while_while_for_for_for_for_for_for_address_mul_8_nl;
  wire[0:0] nor_37_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_main_C_1_tr0;
  assign nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_main_C_1_tr0 = ~ operator_32_false_1_acc_1_itm_32_1;
  wire [0:0] nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0;
  assign nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0
      = ~(while_while_for_stage_0_2 | while_while_for_stage_0_3 | reg_while_while_for_stage_0_cse);
  wire [0:0] nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_C_1_tr0;
  assign nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_C_1_tr0 = ~
      operator_32_false_1_acc_1_itm_32_1;
  InputDoubleBufferReader_512_16_16_run_paramsIn_rsci InputDoubleBufferReader_512_16_16_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsci_1 InputDoubleBufferReader_512_16_16_run_din_rsci_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsci_q_d(din_rsci_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_rsci_oswt(reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse),
      .din_rsci_q_d_mxwt(din_rsci_q_d_mxwt),
      .din_rsci_re_d_pff(din_rsci_re_d_iff),
      .din_rsci_oswt_pff(and_103_rmff)
    );
  InputDoubleBufferReader_512_16_16_run_dout_rsci InputDoubleBufferReader_512_16_16_run_dout_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .run_wen(run_wen),
      .dout_rsci_oswt(reg_dout_rsci_ivld_run_psct_cse),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .dout_rsci_idat(dout_rsci_idat)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj InputDoubleBufferReader_512_16_16_run_din_rsc_rls_obj_inst
      (
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .run_wten(run_wten),
      .din_rsc_rls_obj_iswt0(reg_din_rsc_rls_obj_ld_run_psct_cse)
    );
  InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj InputDoubleBufferReader_512_16_16_run_din_rsc_req_obj_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .din_rsc_req_vz(din_rsc_req_vz),
      .run_wen(run_wen),
      .din_rsc_req_obj_oswt(reg_din_rsc_req_obj_iswt0_cse),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferReader_512_16_16_run_staller InputDoubleBufferReader_512_16_16_run_staller_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .dout_rsci_wen_comp(dout_rsci_wen_comp),
      .din_rsc_req_obj_wen_comp(din_rsc_req_obj_wen_comp)
    );
  InputDoubleBufferReader_512_16_16_run_run_fsm InputDoubleBufferReader_512_16_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_1_tr0(nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_main_C_1_tr0[0:0]),
      .while_while_C_1_tr0(or_dcpl_8),
      .while_while_for_C_0_tr0(nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_while_for_C_0_tr0[0:0]),
      .while_C_1_tr0(nl_InputDoubleBufferReader_512_16_16_run_run_fsm_inst_while_C_1_tr0[0:0])
    );
  assign and_103_rmff = and_dcpl_6 & nor_12_cse & (~(while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1
      | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_for_for_for_not_mdf_sva_st_1))
      & (fsm_output[6]);
  assign while_while_for_for_for_and_cse = run_wen & (~ or_tmp_23);
  assign while_while_for_for_for_and_7_cse = run_wen & (~(while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | or_tmp_23));
  assign while_while_for_for_for_for_and_3_cse = run_wen & (~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | or_tmp_23));
  assign while_while_for_for_for_for_for_and_3_cse = run_wen & (~(while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | or_tmp_23));
  assign block_size_and_1_cse = run_wen & ((fsm_output[2:0]!=3'b000));
  assign and_184_cse = (fsm_output[6:4]==3'b000) & run_wen;
  assign while_while_aelse_while_while_aelse_and_cse = reg_while_while_for_stage_0_cse
      & or_tmp_1;
  assign nor_12_cse = ~(while_while_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1);
  assign while_while_for_and_1_cse = run_wen & reg_while_while_for_stage_0_cse;
  assign nor_32_cse = ~(exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 |
      (~ lfst_exit_while_while_for_for_for_for_lpi_2));
  assign or_121_cse = (~ lfst_exit_while_while_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_lpi_2;
  assign and_93_m1c = (((~((~(((~ exitL_exitL_exit_while_while_for_for_for_for_lpi_2)
      & lfst_exit_while_while_for_for_for_lpi_2) | while_while_for_for_asn_sft_lpi_4))
      | exitL_exit_while_while_for_for_sva)) & (~ exitL_exitL_exit_while_while_for_for_for_lpi_2)
      & lfst_exit_while_while_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_lpi_2)
      | while_while_for_for_for_acc_2_itm_16) & reg_while_while_for_stage_0_cse;
  assign nl_block_size_mul_2_nl = $signed(conv_u2s_9_10(reg_paramsIn_crt_sva_136_0_ftd[104:96]))
      * $signed(operator_16_false_acc_itm);
  assign block_size_mul_2_nl = nl_block_size_mul_2_nl[8:0];
  assign nl_block_size_acc_cse_sva_1 = (block_size_mul_2_nl) + (reg_paramsIn_crt_sva_136_0_ftd[72:64]);
  assign block_size_acc_cse_sva_1 = nl_block_size_acc_cse_sva_1[8:0];
  assign exit_while_while_for_lpi_4_dfm_mx0w1 = (~ while_while_for_acc_3_itm_16)
      & exitL_exit_while_while_for_for_sva;
  assign exit_while_while_for_for_lpi_4_dfm_mx1w0 = (~ while_while_for_for_acc_3_itm_16)
      & exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6;
  assign while_while_for_for_for_for_for_x_idx_and_nl = while_while_for_for_for_while_while_for_for_for_nor_1_itm
      & (~ or_dcpl_23);
  assign while_while_for_for_for_for_for_x_idx_mux_nl = MUX_v_16_2_2(while_while_for_for_for_for_for_x_idx_lpi_4,
      while_while_for_for_for_for_for_acc_1_itm, while_while_for_for_for_for_for_x_idx_and_nl);
  assign while_while_for_for_for_for_for_x_idx_lpi_4_dfm_mx0w1 = MUX_v_16_2_2(16'b0000000000000000,
      (while_while_for_for_for_for_for_x_idx_mux_nl), lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4);
  assign nl_while_while_for_for_for_for_for_for_acc_1_nl = while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1
      + 16'b0000000000000001;
  assign while_while_for_for_for_for_for_for_acc_1_nl = nl_while_while_for_for_for_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_nl
      = ~(while_while_for_for_for_for_for_for_not_mdf_sva_st_1 | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1
      | while_while_for_for_for_or_tmp_1 | while_while_for_for_or_3_tmp_1 | or_dcpl_23);
  assign while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_1_nl
      = ~((~ while_while_for_for_for_for_for_for_not_mdf_sva_st_1) | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1
      | while_while_for_for_for_or_tmp_1 | while_while_for_for_or_3_tmp_1 | or_dcpl_23);
  assign while_while_for_for_for_for_for_for_y_idx_or_nl = while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1
      | while_while_for_for_for_or_tmp_1 | while_while_for_for_or_3_tmp_1 | or_dcpl_23;
  assign while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_mux1h_nl
      = MUX1HOT_v_16_3_2((while_while_for_for_for_for_for_for_acc_1_nl), while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1,
      while_while_for_for_for_for_for_for_y_idx_lpi_4, {(while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_nl)
      , (while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_nor_1_nl)
      , (while_while_for_for_for_for_for_for_y_idx_or_nl)});
  assign while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7 = MUX_v_16_2_2(16'b0000000000000000,
      (while_while_for_for_for_for_for_for_y_idx_while_while_for_for_for_for_for_for_y_idx_mux1h_nl),
      lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5);
  assign nl_while_while_for_for_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7})
      + conv_u2u_16_17(~ (reg_paramsIn_crt_sva_136_0_ftd[31:16])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_for_for_acc_2_itm_16 = readslicef_17_1_16((while_while_for_for_for_for_for_for_acc_2_nl));
  assign or_48_nl = or_dcpl_34 | (~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 | (~ lfst_exit_while_while_for_for_for_for_lpi_2)
      | (~ lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~ lfst_exit_while_while_for_for_for_for_for_lpi_2);
  assign while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_for_for_lpi_4_dfm_1, or_48_nl);
  assign or_56_nl = or_dcpl_32 | (~ lfst_exit_while_while_for_for_lpi_2) | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_for_lpi_2 | (~(lfst_exit_while_while_for_for_for_lpi_2
      & lfst_exitL_exit_while_while_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2))
      | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 | (~ lfst_exit_while_while_for_for_for_for_lpi_2);
  assign while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_for_lpi_4_dfm_1, or_56_nl);
  assign while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_for_lpi_4_dfm_1, or_dcpl_34);
  assign while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0 = MUX_s_1_2_2(while_while_for_for_asn_sft_lpi_4,
      exit_while_while_for_for_lpi_4_dfm_mx1w0, or_dcpl_33);
  assign while_while_for_for_for_or_tmp_1 = while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1
      | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1;
  assign nl_while_while_for_for_for_for_for_acc_1_itm = while_while_for_for_for_for_for_x_idx_lpi_4
      + 16'b0000000000000001;
  assign while_while_for_for_for_for_for_acc_1_itm = nl_while_while_for_for_for_for_for_acc_1_itm[15:0];
  assign while_while_for_for_for_while_while_for_for_for_nor_1_itm = ~((~ while_while_for_for_for_for_for_for_not_mdf_sva_st_1)
      | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_or_tmp_1
      | while_while_for_for_or_3_tmp_1);
  assign while_while_for_for_or_3_tmp_1 = while_while_for_for_asn_sft_lpi_4_dfm_st_1
      | exit_while_while_for_lpi_4_dfm_1;
  assign exit_while_while_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_acc_2_itm_16)
      & exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7;
  assign lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5 = lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7);
  assign nl_while_while_for_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_for_x_idx_lpi_4_dfm_mx0w1})
      + conv_u2u_16_17(~ (reg_paramsIn_crt_sva_136_0_ftd[15:0])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_for_acc_2_itm_16 = readslicef_17_1_16((while_while_for_for_for_for_for_acc_2_nl));
  assign exit_while_while_for_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_for_acc_2_itm_16)
      & exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7;
  assign exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_7 = exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4));
  assign lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4 = lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6);
  assign while_while_for_for_for_for_wy_idx_lpi_4_dfm_6 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_for_wy_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4);
  assign nl_while_while_for_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_for_wy_idx_lpi_4_dfm_6})
      + conv_u2u_16_17(~ (reg_paramsIn_crt_sva_136_0_ftd[95:80])) + 17'b00000000000000001;
  assign while_while_for_for_for_for_acc_2_nl = nl_while_while_for_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_for_acc_2_itm_16 = readslicef_17_1_16((while_while_for_for_for_for_acc_2_nl));
  assign exit_while_while_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_acc_2_itm_16)
      & exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6;
  assign exitL_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_6 = exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4));
  assign lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4 = lfst_exitL_exit_while_while_for_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7);
  assign nl_while_while_for_for_for_acc_2_nl = ({1'b1 , while_while_for_for_for_wx_idx_lpi_4_dfm_5})
      + conv_u2u_16_17(~ (reg_paramsIn_crt_sva_136_0_ftd[79:64])) + 17'b00000000000000001;
  assign while_while_for_for_for_acc_2_nl = nl_while_while_for_for_for_acc_2_nl[16:0];
  assign while_while_for_for_for_acc_2_itm_16 = readslicef_17_1_16((while_while_for_for_for_acc_2_nl));
  assign while_while_for_for_for_wx_idx_lpi_4_dfm_5 = MUX_v_16_2_2(16'b0000000000000000,
      while_while_for_for_for_wx_idx_lpi_4, lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3);
  assign exitL_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_7 = exitL_exitL_exit_while_while_for_for_for_for_lpi_2
      | (~(lfst_exit_while_while_for_for_for_lpi_2 & lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3));
  assign lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3 = lfst_exitL_exit_while_while_for_for_for_lpi_2
      & (~ exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6);
  assign nl_while_while_for_for_acc_3_nl = ({1'b1 , while_while_for_for_co_idx_lpi_4_dfm_1_mx0})
      + conv_u2u_16_17(~ (reg_paramsIn_crt_sva_136_0_ftd[63:48])) + 17'b00000000000000001;
  assign while_while_for_for_acc_3_nl = nl_while_while_for_for_acc_3_nl[16:0];
  assign while_while_for_for_acc_3_itm_16 = readslicef_17_1_16((while_while_for_for_acc_3_nl));
  assign while_while_for_for_co_idx_lpi_4_dfm_1_mx0 = MUX_v_16_2_2(while_while_for_for_co_idx_lpi_4,
      (signext_16_1(~ while_while_for_acc_3_itm_16)), exitL_exit_while_while_for_for_sva);
  assign while_while_for_for_mux_60_nl = MUX_s_1_2_2(lfst_exit_while_while_for_for_lpi_2,
      lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0, exitL_exit_while_while_for_for_sva);
  assign exitL_exitL_exit_while_while_for_for_for_lpi_4_dfm_6 = exitL_exitL_exit_while_while_for_for_for_lpi_2
      | (~ (while_while_for_for_mux_60_nl));
  assign lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0 = lfst_exit_while_while_for_for_lpi_2
      & (~ while_while_for_acc_3_itm_16);
  assign nl_while_while_for_acc_3_nl = ({1'b1 , while_while_for_koo_idx_sva}) + conv_u2u_16_17(~
      (reg_paramsIn_crt_sva_136_0_ftd[47:32])) + 17'b00000000000000001;
  assign while_while_for_acc_3_nl = nl_while_while_for_acc_3_nl[16:0];
  assign while_while_for_acc_3_itm_16 = readslicef_17_1_16((while_while_for_acc_3_nl));
  assign exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1 = (~ while_while_for_for_for_for_for_for_acc_2_itm_16)
      | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  assign exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1 = exit_while_while_for_for_for_for_for_lpi_4_dfm_1
      | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
  assign nl_operator_32_false_1_acc_1_nl = ({1'b1 , (~ total_blocks_lpi_3)}) + 33'b000000000000000000000000000000001;
  assign operator_32_false_1_acc_1_nl = nl_operator_32_false_1_acc_1_nl[32:0];
  assign operator_32_false_1_acc_1_itm_32_1 = readslicef_33_1_32((operator_32_false_1_acc_1_nl));
  assign and_dcpl_4 = ~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1);
  assign and_dcpl_6 = while_while_for_stage_0_2 & (~ while_while_for_asn_4_itm_1);
  assign and_dcpl_7 = and_dcpl_6 & (~ while_while_for_for_asn_sft_lpi_4_dfm_st_1);
  assign or_tmp_1 = while_while_for_acc_3_itm_16 | (~ exitL_exit_while_while_for_for_sva);
  assign and_82_nl = (~ exitL_exit_while_while_for_for_sva) & (~ exitL_exitL_exit_while_while_for_for_for_lpi_2)
      & lfst_exit_while_while_for_for_lpi_2;
  assign mux_tmp_2 = MUX_s_1_2_2((and_82_nl), or_tmp_1, while_while_for_for_acc_3_itm_16);
  assign and_181_cse = while_while_for_acc_3_itm_16 & exitL_exit_while_while_for_for_sva;
  assign nor_nl = ~(lfst_exitL_exit_while_while_for_for_for_lpi_2 | (~ lfst_exit_while_while_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_lpi_2 | exitL_exit_while_while_for_for_sva);
  assign or_7_nl = (~ lfst_exitL_exit_while_while_for_for_for_lpi_2) | (~ lfst_exit_while_while_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_lpi_2;
  assign mux_6_nl = MUX_s_1_2_2(and_181_cse, or_tmp_1, or_7_nl);
  assign mux_7_nl = MUX_s_1_2_2((nor_nl), (mux_6_nl), while_while_for_for_acc_3_itm_16);
  assign mux_tmp_3 = MUX_s_1_2_2(mux_tmp_2, (mux_7_nl), while_while_for_for_asn_sft_lpi_4);
  assign nl_while_while_aelse_acc_nl = conv_u2u_9_10(operator_16_false_acc_itm) +
      10'b1100000001;
  assign while_while_aelse_acc_nl = nl_while_while_aelse_acc_nl[9:0];
  assign or_dcpl_8 = ~(exit_while_while_for_lpi_4_dfm_1 & (~ (readslicef_10_1_9((while_while_aelse_acc_nl)))));
  assign and_dcpl_56 = ~((fsm_output[1:0]!=2'b00));
  assign or_dcpl_23 = (~ while_while_for_stage_0_2) | while_while_for_asn_4_itm_1;
  assign or_dcpl_32 = exitL_exit_while_while_for_for_sva | exitL_exitL_exit_while_while_for_for_for_lpi_2;
  assign or_dcpl_33 = or_dcpl_32 | (~ lfst_exit_while_while_for_for_lpi_2) | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2);
  assign or_dcpl_34 = or_dcpl_33 | or_121_cse | (~ lfst_exitL_exit_while_while_for_for_for_for_lpi_2);
  assign or_tmp_23 = (~ (fsm_output[6])) | exit_while_while_for_lpi_4_dfm_mx0w1 |
      (~ reg_while_while_for_stage_0_cse);
  assign or_tmp_44 = ~((fsm_output[7:4]!=4'b0000));
  assign lfst_exit_while_while_for_for_lpi_2_mx0c1 = exit_while_while_for_lpi_4_dfm_mx0w1
      & reg_while_while_for_stage_0_cse & (fsm_output[6]);
  assign nl_while_while_for_for_for_for_for_for_address_acc_9_nl = operator_16_false_acc_itm
      + while_while_for_for_for_for_for_for_address_mul_5_itm_1;
  assign while_while_for_for_for_for_for_for_address_acc_9_nl = nl_while_while_for_for_for_for_for_for_address_acc_9_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_8_nl = (reg_paramsIn_crt_sva_136_0_ftd[104:96])
      * (while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1[8:0]);
  assign while_while_for_for_for_for_for_for_address_mul_8_nl = nl_while_while_for_for_for_for_for_for_address_mul_8_nl[8:0];
  assign nl_din_rsci_radr_d = (while_while_for_for_for_for_for_for_address_acc_9_nl)
      + while_while_for_for_for_for_for_for_address_mul_itm_1 + (while_while_for_for_for_for_for_for_address_mul_8_nl)
      + while_while_for_for_for_for_for_for_slc_while_while_for_for_for_for_wy_idx_8_0_itm_1;
  assign din_rsci_radr_d = nl_din_rsci_radr_d[8:0];
  assign din_rsci_re_d_pff = din_rsci_re_d_iff;
  assign nor_37_nl = ~(while_while_for_for_asn_sft_lpi_4 | while_while_for_for_for_asn_sft_lpi_4);
  assign mux_tmp = MUX_s_1_2_2((nor_37_nl), while_while_for_acc_3_itm_16, exitL_exit_while_while_for_for_sva);
  assign mux_tmp_9 = MUX_s_1_2_2(and_181_cse, mux_tmp, while_while_for_for_for_for_acc_2_itm_16);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_din_rsc_req_obj_iswt0_cse <= 1'b0;
      reg_din_rsc_rls_obj_ld_run_psct_cse <= 1'b0;
      reg_dout_rsci_ivld_run_psct_cse <= 1'b0;
      reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      operator_16_false_acc_itm <= 9'b000000000;
      exit_while_while_for_lpi_4_dfm_1 <= 1'b0;
      reg_while_while_for_stage_0_cse <= 1'b0;
      exitL_exit_while_while_for_for_sva <= 1'b0;
      while_while_for_stage_0_2 <= 1'b0;
      while_while_for_stage_0_3 <= 1'b0;
      while_while_for_for_for_for_for_for_y_idx_lpi_4 <= 16'b0000000000000000;
      while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1 <= 16'b0000000000000000;
      while_while_for_for_for_for_for_for_not_mdf_sva_st_1 <= 1'b0;
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
      while_while_for_for_for_for_for_for_slc_while_while_for_for_for_for_wy_idx_8_0_itm_1
          <= 9'b000000000;
      while_while_for_for_for_for_for_for_address_mul_itm_1 <= 9'b000000000;
      while_while_for_for_for_for_for_for_address_mul_5_itm_1 <= 9'b000000000;
      reg_paramsIn_crt_sva_136_0_ftd <= 105'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_din_rsc_req_obj_iswt0_cse <= operator_32_false_1_acc_1_itm_32_1 & ((fsm_output[8])
          | (fsm_output[2]));
      reg_din_rsc_rls_obj_ld_run_psct_cse <= or_dcpl_8 & (fsm_output[5]);
      reg_dout_rsci_ivld_run_psct_cse <= while_while_for_stage_0_3 & (~ while_while_for_for_for_for_for_for_not_mdf_sva_st_2)
          & (~(while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_2 | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_2))
          & (~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_2 | while_while_for_for_asn_sft_lpi_4_dfm_st_2
          | exit_while_while_for_lpi_4_dfm_st_2)) & (fsm_output[6]);
      reg_din_rsci_port_0_r_ram_ir_internal_RMASK_B_d_run_psct_cse <= and_103_rmff;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[8]) | (fsm_output[2])
          | (fsm_output[0]))) | (~((~ operator_32_false_1_acc_1_itm_32_1) | (fsm_output[0]))));
      operator_16_false_acc_itm <= MUX1HOT_v_9_3_2((operator_16_false_acc_nl), (readslicef_10_9_1((while_while_aelse_acc_1_nl))),
          (while_while_for_for_for_for_for_for_address_mul_1_nl), {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[6])});
      exit_while_while_for_lpi_4_dfm_1 <= MUX_s_1_2_2(operator_32_false_1_acc_1_itm_32_1,
          exit_while_while_for_lpi_4_dfm_mx0w1, fsm_output[6]);
      reg_while_while_for_stage_0_cse <= while_while_aelse_while_while_aelse_and_cse
          | (~ (fsm_output[6]));
      exitL_exit_while_while_for_for_sva <= (while_while_for_mux_4_nl) | (~ (fsm_output[6]));
      while_while_for_stage_0_2 <= reg_while_while_for_stage_0_cse & (fsm_output[6]);
      while_while_for_stage_0_3 <= while_while_for_stage_0_2 & (fsm_output[6]);
      while_while_for_for_for_for_for_for_y_idx_lpi_4 <= 16'b0000000000000000;
      while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_1 <= while_while_for_for_for_for_for_for_y_idx_lpi_4_dfm_7;
      while_while_for_for_for_for_for_for_not_mdf_sva_st_1 <= ~ while_while_for_for_for_for_for_for_acc_2_itm_16;
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      while_while_for_for_for_for_for_for_slc_while_while_for_for_for_for_wy_idx_8_0_itm_1
          <= while_while_for_for_for_for_wy_idx_lpi_4_dfm_6[8:0];
      while_while_for_for_for_for_for_for_address_mul_itm_1 <= nl_while_while_for_for_for_for_for_for_address_mul_itm_1[8:0];
      while_while_for_for_for_for_for_for_address_mul_5_itm_1 <= nl_while_while_for_for_for_for_for_for_address_mul_5_itm_1[8:0];
      reg_paramsIn_crt_sva_136_0_ftd <= MUX_v_105_2_2((paramsIn_rsci_idat_mxwt[136:32]),
          reg_paramsIn_crt_sva_136_0_ftd, and_dcpl_56);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      dout_rsci_idat <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ (fsm_output[6])) | (~ while_while_for_stage_0_3) |
        while_while_for_for_for_for_for_for_not_mdf_sva_st_2 | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_2
        | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_2 | while_while_for_for_for_asn_sft_lpi_4_dfm_st_2
        | while_while_for_for_asn_sft_lpi_4_dfm_st_2 | exit_while_while_for_lpi_4_dfm_st_2))
        ) begin
      dout_rsci_idat <= din_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_lpi_2 <= 1'b0;
    end
    else if ( run_wen & ((or_tmp_1 & reg_while_while_for_stage_0_cse & (fsm_output[6]))
        | lfst_exit_while_while_for_for_lpi_2_mx0c1) ) begin
      lfst_exit_while_while_for_for_lpi_2 <= MUX_s_1_2_2((~ exit_while_while_for_for_lpi_4_dfm_mx1w0),
          lfst_exit_while_while_for_for_lpi_4_dfm_1_mx0w0, lfst_exit_while_while_for_for_lpi_2_mx0c1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exitL_exit_while_while_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_and_cse ) begin
      exitL_exitL_exit_while_while_for_for_for_lpi_2 <= exit_while_while_for_for_for_lpi_4_dfm_1
          | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      lfst_exitL_exit_while_while_for_for_for_lpi_2 <= ~(exit_while_while_for_for_for_lpi_4_dfm_1
          | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_and_7_cse ) begin
      lfst_exit_while_while_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_lpi_2 <= exit_while_while_for_for_for_for_lpi_4_dfm_1
          | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
      lfst_exitL_exit_while_while_for_for_for_for_lpi_2 <= ~(exit_while_while_for_for_for_for_lpi_4_dfm_1
          | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_for_and_3_cse ) begin
      lfst_exit_while_while_for_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
      lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2 <= ~ exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_while_while_for_for_for_for_for_lpi_2 <= 1'b0;
      exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= 1'b0;
      lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= 1'b0;
    end
    else if ( while_while_for_for_for_for_for_and_3_cse ) begin
      lfst_exit_while_while_for_for_for_for_for_lpi_2 <= ~ exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
      exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
      lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_2 <= ~ exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_acc_1_cse_sva <= 9'b000000000;
    end
    else if ( run_wen & (~ and_dcpl_56) ) begin
      block_size_acc_1_cse_sva <= nl_block_size_acc_1_cse_sva[8:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      total_blocks_lpi_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen & ((~ and_dcpl_56) | (fsm_output[7])) ) begin
      total_blocks_lpi_3 <= MUX_v_32_2_2((total_blocks_mul_nl), (while_while_acc_1_nl),
          fsm_output[7]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      block_size_sva <= 9'b000000000;
      block_size_acc_cse_sva <= 9'b000000000;
    end
    else if ( block_size_and_1_cse ) begin
      block_size_sva <= nl_block_size_sva[8:0];
      block_size_acc_cse_sva <= block_size_acc_cse_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_current_buffer_size_sva <= 9'b000000000;
      while_block_count_8_0_sva <= 9'b000000000;
    end
    else if ( and_184_cse ) begin
      while_current_buffer_size_sva <= MUX_v_9_2_2(9'b000000000, (while_while_acc_2_nl),
          (while_current_buffer_size_not_1_nl));
      while_block_count_8_0_sva <= MUX_v_9_2_2(9'b000000000, (while_while_acc_nl),
          (while_block_count_not_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_koo_idx_sva <= 16'b0000000000000000;
    end
    else if ( (~((~(((~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2
        | exitL_exit_while_while_for_for_sva) & reg_while_while_for_stage_0_cse &
        (~ while_while_for_for_acc_3_itm_16))) & (fsm_output[6]))) & run_wen ) begin
      while_while_for_koo_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, (while_while_for_acc_2_nl),
          (fsm_output[6]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_for_not_mdf_sva_st_2 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_7 & and_dcpl_4 & (~ while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1)
        ) begin
      while_while_for_for_for_for_for_for_not_mdf_sva_st_2 <= while_while_for_for_for_for_for_for_not_mdf_sva_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_2 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_7 & and_dcpl_4 ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_2 <= while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_2 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_6 & nor_12_cse ) begin
      while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_2 <= while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_2 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_7 ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_2 <= while_while_for_for_for_asn_sft_lpi_4_dfm_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_2 <= 1'b0;
    end
    else if ( run_wen & and_dcpl_6 ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_2 <= while_while_for_for_asn_sft_lpi_4_dfm_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_while_while_for_lpi_4_dfm_st_2 <= 1'b0;
    end
    else if ( run_wen & while_while_for_stage_0_2 ) begin
      exit_while_while_for_lpi_4_dfm_st_2 <= while_while_for_asn_4_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_x_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( (~(((~ while_while_for_stage_0_2) | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1
        | while_while_for_asn_4_itm_1 | (~ while_while_for_for_for_for_for_for_not_mdf_sva_st_1)
        | while_while_for_for_for_for_for_asn_sft_lpi_4_dfm_st_1 | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1
        | while_while_for_for_asn_sft_lpi_4_dfm_st_1 | exit_while_while_for_lpi_4_dfm_1)
        & (~(reg_while_while_for_stage_0_cse & ((~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2)
        | (~ lfst_exit_while_while_for_for_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_for_for_lpi_2
        | (~ lfst_exitL_exit_while_while_for_for_for_for_lpi_2) | (~ lfst_exit_while_while_for_for_for_lpi_2)
        | exitL_exitL_exit_while_while_for_for_for_for_lpi_2 | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2)
        | exitL_exitL_exit_while_while_for_for_for_lpi_2 | (~((~(exitL_exit_while_while_for_for_sva
        & while_while_for_acc_3_itm_16)) & lfst_exit_while_while_for_for_lpi_2)))))))
        & run_wen & (while_while_for_for_for_while_while_for_for_for_nor_1_itm |
        reg_while_while_for_stage_0_cse) ) begin
      while_while_for_for_for_for_for_x_idx_lpi_4 <= MUX_v_16_2_2(while_while_for_for_for_for_for_acc_1_itm,
          while_while_for_for_for_for_for_x_idx_lpi_4_dfm_mx0w1, reg_while_while_for_stage_0_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_3 & reg_while_while_for_stage_0_cse ) begin
      while_while_for_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_1 <= 1'b0;
    end
    else if ( run_wen & while_while_aelse_while_while_aelse_and_cse ) begin
      while_while_for_for_asn_sft_lpi_4_dfm_st_1 <= while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_asn_4_itm_1 <= 1'b0;
    end
    else if ( while_while_for_and_1_cse ) begin
      while_while_for_asn_4_itm_1 <= exit_while_while_for_lpi_4_dfm_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_for_for_lpi_4_dfm_5)
        | while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
        | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & reg_while_while_for_stage_0_cse
        ) begin
      while_while_for_for_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_for_lpi_4_dfm_4)
        | while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0 | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0)
        & reg_while_while_for_stage_0_cse ) begin
      while_while_for_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_for_wy_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( ((mux_20_nl) | (~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2
        | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2) | (~ lfst_exit_while_while_for_for_for_lpi_2)
        | exitL_exitL_exit_while_while_for_for_for_for_lpi_2 | (~ lfst_exitL_exit_while_while_for_for_for_for_lpi_2))
        & while_while_for_and_1_cse ) begin
      while_while_for_for_for_for_wy_idx_lpi_4 <= MUX_v_16_2_2(while_while_for_for_for_for_wy_idx_lpi_4_dfm_6,
          (while_while_for_for_for_for_acc_1_nl), while_while_for_for_and_7_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & ((~ lfst_exitL_exit_while_while_for_for_for_for_lpi_4_dfm_4)
        | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & reg_while_while_for_stage_0_cse
        ) begin
      while_while_for_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_for_lpi_4_dfm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_for_wx_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( (mux_25_nl) & while_while_for_and_1_cse ) begin
      while_while_for_for_for_wx_idx_lpi_4 <= MUX_v_16_2_2(while_while_for_for_for_wx_idx_lpi_4_dfm_5,
          (while_while_for_for_for_acc_1_nl), while_while_for_for_for_wx_idx_and_1_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_asn_sft_lpi_4 <= 1'b0;
    end
    else if ( run_wen & (mux_10_nl) & reg_while_while_for_stage_0_cse & (~ lfst_exitL_exit_while_while_for_for_for_lpi_4_dfm_3)
        ) begin
      while_while_for_for_asn_sft_lpi_4 <= exit_while_while_for_for_lpi_4_dfm_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      while_while_for_for_co_idx_lpi_4 <= 16'b0000000000000000;
    end
    else if ( run_wen & mux_tmp_2 & reg_while_while_for_stage_0_cse & (~((~ exitL_exit_while_while_for_for_sva)
        & and_93_m1c)) ) begin
      while_while_for_for_co_idx_lpi_4 <= MUX_v_16_2_2((while_while_for_for_acc_2_nl),
          (signext_16_1(~ while_while_for_acc_3_itm_16)), while_while_for_for_and_10_nl);
    end
  end
  assign nl_operator_16_false_acc_nl = (paramsIn_rsci_idat_mxwt[56:48]) + 9'b111111111;
  assign operator_16_false_acc_nl = nl_operator_16_false_acc_nl[8:0];
  assign nl_while_while_aelse_acc_1_nl = conv_u2u_9_10(~ while_current_buffer_size_sva)
      + conv_u2u_9_10(~ block_size_sva);
  assign while_while_aelse_acc_1_nl = nl_while_while_aelse_acc_1_nl[9:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_2_nl = $signed(conv_u2s_9_10(while_while_for_for_co_idx_lpi_4_dfm_1_mx0[8:0]))
      * $signed(block_size_acc_cse_sva);
  assign while_while_for_for_for_for_for_for_address_mul_2_nl = nl_while_while_for_for_for_for_for_for_address_mul_2_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_1_nl = $signed((while_while_for_for_for_for_for_for_address_mul_2_nl))
      * $signed(block_size_acc_1_cse_sva);
  assign while_while_for_for_for_for_for_for_address_mul_1_nl = nl_while_while_for_for_for_for_for_for_address_mul_1_nl[8:0];
  assign while_while_for_mux_4_nl = MUX_s_1_2_2(exitL_exit_while_while_for_for_sva,
      exit_while_while_for_for_lpi_4_dfm_mx1w0, reg_while_while_for_stage_0_cse);
  assign nl_while_while_for_for_for_for_for_for_address_mul_itm_1  = while_block_count_8_0_sva
      * block_size_sva;
  assign nl_while_while_for_for_for_for_for_for_address_mul_6_nl = (reg_paramsIn_crt_sva_136_0_ftd[104:96])
      * (while_while_for_for_for_for_for_x_idx_lpi_4_dfm_mx0w1[8:0]);
  assign while_while_for_for_for_for_for_for_address_mul_6_nl = nl_while_while_for_for_for_for_for_for_address_mul_6_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_acc_6_nl = (while_while_for_for_for_for_for_for_address_mul_6_nl)
      + (while_while_for_for_for_wx_idx_lpi_4_dfm_5[8:0]);
  assign while_while_for_for_for_for_for_for_address_acc_6_nl = nl_while_while_for_for_for_for_for_for_address_acc_6_nl[8:0];
  assign nl_while_while_for_for_for_for_for_for_address_mul_5_itm_1  = $signed(conv_u2s_9_10(while_while_for_for_for_for_for_for_address_acc_6_nl))
      * $signed(block_size_acc_cse_sva);
  assign nl_operator_16_false_1_acc_nl = (paramsIn_rsci_idat_mxwt[40:32]) + 9'b111111111;
  assign operator_16_false_1_acc_nl = nl_operator_16_false_1_acc_nl[8:0];
  assign nl_block_size_mul_3_nl = $signed(conv_u2s_9_10(paramsIn_rsci_idat_mxwt[136:128]))
      * $signed((operator_16_false_1_acc_nl));
  assign block_size_mul_3_nl = nl_block_size_mul_3_nl[8:0];
  assign nl_block_size_acc_1_cse_sva  = (block_size_mul_3_nl) + (paramsIn_rsci_idat_mxwt[120:112]);
  assign total_blocks_mul_nl = conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16]) *
      (paramsIn_rsci_idat_mxwt[15:0]));
  assign nl_while_while_acc_1_nl = total_blocks_lpi_3 + 32'b11111111111111111111111111111111;
  assign while_while_acc_1_nl = nl_while_while_acc_1_nl[31:0];
  assign nl_block_size_mul_1_nl = $signed(conv_u2s_9_10(reg_paramsIn_crt_sva_136_0_ftd[56:48]))
      * $signed(block_size_acc_cse_sva_1);
  assign block_size_mul_1_nl = nl_block_size_mul_1_nl[8:0];
  assign nl_block_size_sva  = $signed((block_size_mul_1_nl)) * $signed(block_size_acc_1_cse_sva);
  assign nl_while_while_acc_2_nl = while_current_buffer_size_sva + block_size_sva;
  assign while_while_acc_2_nl = nl_while_while_acc_2_nl[8:0];
  assign while_current_buffer_size_not_1_nl = ~ or_tmp_44;
  assign nl_while_while_acc_nl = while_block_count_8_0_sva + 9'b000000001;
  assign while_while_acc_nl = nl_while_while_acc_nl[8:0];
  assign while_block_count_not_nl = ~ or_tmp_44;
  assign nl_while_while_for_acc_2_nl = while_while_for_koo_idx_sva + 16'b0000000000000001;
  assign while_while_for_acc_2_nl = nl_while_while_for_acc_2_nl[15:0];
  assign nl_while_while_for_for_for_for_acc_1_nl = while_while_for_for_for_for_wy_idx_lpi_4_dfm_6
      + 16'b0000000000000001;
  assign while_while_for_for_for_for_acc_1_nl = nl_while_while_for_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_and_7_nl = exit_while_while_for_for_for_for_for_lpi_4_dfm_1
      & (~ while_while_for_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & (~(while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0)) & (~ exit_while_while_for_lpi_4_dfm_mx0w1);
  assign and_197_nl = while_while_for_for_for_for_asn_sft_lpi_4 & lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2;
  assign mux_17_nl = MUX_s_1_2_2(mux_tmp, and_181_cse, and_197_nl);
  assign mux_18_nl = MUX_s_1_2_2(mux_tmp_9, (mux_17_nl), nor_32_cse);
  assign mux_14_nl = MUX_s_1_2_2(mux_tmp, and_181_cse, lfst_exitL_exit_while_while_for_for_for_for_for_lpi_2);
  assign mux_16_nl = MUX_s_1_2_2(mux_tmp_9, (mux_14_nl), nor_32_cse);
  assign nor_30_nl = ~(exitL_exitL_exit_while_while_for_for_for_for_for_for_lpi_2
      | (~ lfst_exit_while_while_for_for_for_for_for_lpi_2));
  assign mux_19_nl = MUX_s_1_2_2((mux_18_nl), (mux_16_nl), nor_30_nl);
  assign mux_20_nl = MUX_s_1_2_2((mux_19_nl), and_181_cse, while_while_for_for_for_for_for_acc_2_itm_16);
  assign nl_while_while_for_for_for_acc_1_nl = while_while_for_for_for_wx_idx_lpi_4_dfm_5
      + 16'b0000000000000001;
  assign while_while_for_for_for_acc_1_nl = nl_while_while_for_for_for_acc_1_nl[15:0];
  assign while_while_for_for_for_wx_idx_and_1_nl = exit_while_while_for_for_for_for_lpi_4_dfm_1
      & (~ while_while_for_for_for_asn_sft_lpi_4_dfm_st_1_mx0) & (~(while_while_for_for_asn_sft_lpi_4_dfm_st_1_mx0
      | exit_while_while_for_lpi_4_dfm_mx0w1)) & reg_while_while_for_stage_0_cse;
  assign nor_40_nl = ~(while_while_for_for_asn_sft_lpi_4 | while_while_for_for_for_for_acc_2_itm_16);
  assign nor_41_nl = ~(while_while_for_for_for_asn_sft_lpi_4 | nor_32_cse | while_while_for_for_asn_sft_lpi_4
      | while_while_for_for_for_for_acc_2_itm_16);
  assign mux_21_nl = MUX_s_1_2_2((nor_40_nl), (nor_41_nl), lfst_exitL_exit_while_while_for_for_for_for_lpi_2);
  assign nor_42_nl = ~((~ while_while_for_for_for_acc_2_itm_16) | while_while_for_for_asn_sft_lpi_4
      | while_while_for_for_for_for_acc_2_itm_16);
  assign mux_22_nl = MUX_s_1_2_2((mux_21_nl), (nor_42_nl), or_121_cse);
  assign mux_23_nl = MUX_s_1_2_2(while_while_for_for_for_acc_2_itm_16, (mux_22_nl),
      lfst_exitL_exit_while_while_for_for_for_lpi_2);
  assign and_199_nl = while_while_for_for_acc_3_itm_16 & while_while_for_for_for_acc_2_itm_16;
  assign or_120_nl = (~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2;
  assign mux_24_nl = MUX_s_1_2_2((mux_23_nl), (and_199_nl), or_120_nl);
  assign and_200_nl = while_while_for_acc_3_itm_16 & while_while_for_for_acc_3_itm_16
      & while_while_for_for_for_acc_2_itm_16;
  assign mux_25_nl = MUX_s_1_2_2((mux_24_nl), (and_200_nl), exitL_exit_while_while_for_for_sva);
  assign nor_9_nl = ~(while_while_for_for_asn_sft_lpi_4 | (~ lfst_exit_while_while_for_for_for_lpi_2)
      | exitL_exitL_exit_while_while_for_for_for_for_lpi_2 | (~ lfst_exitL_exit_while_while_for_for_for_lpi_2)
      | (~ lfst_exit_while_while_for_for_lpi_2) | exitL_exitL_exit_while_while_for_for_for_lpi_2
      | exitL_exit_while_while_for_for_sva);
  assign mux_10_nl = MUX_s_1_2_2((nor_9_nl), mux_tmp_3, while_while_for_for_for_acc_2_itm_16);
  assign nl_while_while_for_for_acc_2_nl = while_while_for_for_co_idx_lpi_4_dfm_1_mx0
      + 16'b0000000000000001;
  assign while_while_for_for_acc_2_nl = nl_while_while_for_for_acc_2_nl[15:0];
  assign while_while_for_for_and_10_nl = exitL_exit_while_while_for_for_sva & and_93_m1c;

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [104:0] MUX_v_105_2_2;
    input [104:0] input_0;
    input [104:0] input_1;
    input [0:0] sel;
    reg [104:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_105_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_10_9_1;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_10_9_1 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] signext_16_1;
    input [0:0] vector;
  begin
    signext_16_1= {{15{vector[0]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [16:0] conv_u2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_run
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, inputDoubleBufferWriterParams_cns_dat,
      inputDoubleBufferWriterParams_cns_vld, inputDoubleBufferWriterParams_cns_rdy,
      inputDoubleBufferReaderParams_cns_dat, inputDoubleBufferReaderParams_cns_vld,
      inputDoubleBufferReaderParams_cns_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] inputDoubleBufferWriterParams_cns_dat;
  output inputDoubleBufferWriterParams_cns_vld;
  input inputDoubleBufferWriterParams_cns_rdy;
  output [143:0] inputDoubleBufferReaderParams_cns_dat;
  output inputDoubleBufferReaderParams_cns_vld;
  input inputDoubleBufferReaderParams_cns_rdy;



  // Interconnect Declarations for Component Instantiations 
  InputDoubleBuffer_512_16_16_run_run InputDoubleBuffer_512_16_16_run_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld),
      .inputDoubleBufferReaderParams_cns_rdy(inputDoubleBufferReaderParams_cns_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferWriter_512_16_16
// ------------------------------------------------------------------


module InputDoubleBufferWriter_512_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_dat,
      din_rsc_vld, din_rsc_rdy, dout_rsc_wadr, dout_rsc_d, dout_rsc_we, dout_rsc_req_vz,
      dout_rsc_rls_lz
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input [15:0] din_rsc_dat;
  input din_rsc_vld;
  output din_rsc_rdy;
  output [8:0] dout_rsc_wadr;
  output [127:0] dout_rsc_d;
  output dout_rsc_we;
  input dout_rsc_req_vz;
  output dout_rsc_rls_lz;


  // Interconnect Declarations
  wire [8:0] dout_rsci_wadr_d;
  wire [127:0] dout_rsci_d_d;
  wire dout_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferWriter_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_wport_3_128_9_512_512_128_5_gen
      dout_rsci (
      .we(dout_rsc_we),
      .d(dout_rsc_d),
      .wadr(dout_rsc_wadr),
      .wadr_d(dout_rsci_wadr_d),
      .d_d(dout_rsci_d_d),
      .we_d(dout_rsci_we_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(dout_rsci_we_d_iff)
    );
  InputDoubleBufferWriter_512_16_16_run InputDoubleBufferWriter_512_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_dat(din_rsc_dat),
      .din_rsc_vld(din_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy),
      .dout_rsc_req_vz(dout_rsc_req_vz),
      .dout_rsc_rls_lz(dout_rsc_rls_lz),
      .dout_rsci_wadr_d(dout_rsci_wadr_d),
      .dout_rsci_d_d(dout_rsci_d_d),
      .dout_rsci_we_d_pff(dout_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBufferReader_512_16_16
// ------------------------------------------------------------------


module InputDoubleBufferReader_512_16_16 (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, din_rsc_radr,
      din_rsc_re, din_rsc_q, din_rsc_req_vz, din_rsc_rls_lz, dout_rsc_dat, dout_rsc_vld,
      dout_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [8:0] din_rsc_radr;
  output din_rsc_re;
  input [127:0] din_rsc_q;
  input din_rsc_req_vz;
  output din_rsc_rls_lz;
  output [127:0] dout_rsc_dat;
  output dout_rsc_vld;
  input dout_rsc_rdy;


  // Interconnect Declarations
  wire [8:0] din_rsci_radr_d;
  wire [127:0] din_rsci_q_d;
  wire din_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  InputDoubleBufferReader_512_16_16_ccs_sample_mem_ccs_ram_sync_1R1W_rport_8_128_9_512_512_128_5_gen
      din_rsci (
      .q(din_rsc_q),
      .re(din_rsc_re),
      .radr(din_rsc_radr),
      .radr_d(din_rsci_radr_d),
      .re_d(din_rsci_re_d_iff),
      .q_d(din_rsci_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(din_rsci_re_d_iff)
    );
  InputDoubleBufferReader_512_16_16_run InputDoubleBufferReader_512_16_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .din_rsc_req_vz(din_rsc_req_vz),
      .din_rsc_rls_lz(din_rsc_rls_lz),
      .dout_rsc_dat(dout_rsc_dat),
      .dout_rsc_vld(dout_rsc_vld),
      .dout_rsc_rdy(dout_rsc_rdy),
      .din_rsci_radr_d(din_rsci_radr_d),
      .din_rsci_q_d(din_rsci_q_d),
      .din_rsci_re_d_pff(din_rsci_re_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16_struct
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16_struct (
  clk, arst_n, inputs_in_rsc_dat_value, inputs_in_rsc_vld, inputs_in_rsc_rdy, inputs_out_rsc_dat_value,
      inputs_out_rsc_vld, inputs_out_rsc_rdy, paramsIn_rsc_dat_STRIDE, paramsIn_rsc_dat_FY,
      paramsIn_rsc_dat_FX, paramsIn_rsc_dat_IC1, paramsIn_rsc_dat_OC1, paramsIn_rsc_dat_OX0,
      paramsIn_rsc_dat_OY0, paramsIn_rsc_dat_OX1, paramsIn_rsc_dat_OY1, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputs_in_rsc_dat_value;
  input inputs_in_rsc_vld;
  output inputs_in_rsc_rdy;
  output [127:0] inputs_out_rsc_dat_value;
  output inputs_out_rsc_vld;
  input inputs_out_rsc_rdy;
  input [15:0] paramsIn_rsc_dat_STRIDE;
  input [15:0] paramsIn_rsc_dat_FY;
  input [15:0] paramsIn_rsc_dat_FX;
  input [15:0] paramsIn_rsc_dat_IC1;
  input [15:0] paramsIn_rsc_dat_OC1;
  input [15:0] paramsIn_rsc_dat_OX0;
  input [15:0] paramsIn_rsc_dat_OY0;
  input [15:0] paramsIn_rsc_dat_OX1;
  input [15:0] paramsIn_rsc_dat_OY1;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] paramsIn_rsc_dat_ninputDoubleBufferWriter;
  wire paramsIn_rsc_vld_ninputDoubleBufferWriter;
  wire paramsIn_rsc_rdy_ninputDoubleBufferWriter;
  wire din_rsc_rdy_ninputDoubleBufferWriter;
  wire [8:0] dout_rsc_wadr_ninputDoubleBufferWriter;
  wire [127:0] dout_rsc_d_ninputDoubleBufferWriter;
  wire dout_rsc_we_ninputDoubleBufferWriter;
  wire dout_rsc_req_vz_ninputDoubleBufferWriter;
  wire paramsIn_rsc_rdy_ninputDoubleBufferReader;
  wire [8:0] din_rsc_radr_ninputDoubleBufferReader;
  wire din_rsc_re_ninputDoubleBufferReader;
  wire [127:0] din_rsc_q_ninputDoubleBufferReader;
  wire din_rsc_req_vz_ninputDoubleBufferReader;
  wire [127:0] dout_rsc_dat_ninputDoubleBufferReader;
  wire dout_rsc_vld_ninputDoubleBufferReader;
  wire [143:0] inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst;
  wire inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst;
  wire [143:0] inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst;
  wire paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud;
  wire inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire din_rsc_rdy_ninputDoubleBufferWriter_bud;
  wire dout_rsc_rls_lz_ninputDoubleBufferWriter_bud;
  wire din_rsc_rls_lz_ninputDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_ninputDoubleBufferReader_bud;
  wire inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire dout_rsc_vld_ninputDoubleBufferReader_bud;
  wire paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud;
  wire inputDoubleBufferWriterParams_unc_2;
  wire inputDoubleBufferWriterParams_idle;
  wire mem_cns_R0;
  wire mem_cns_R1;
  wire [8:0] mem_cns_radr_shi0;
  wire [8:0] mem_cns_radr_shi1;
  wire [8:0] mem_cns_wadr_shi0;
  wire [8:0] mem_cns_wadr_shi1;
  wire [127:0] mem_cns_d_shi0;
  wire [127:0] mem_cns_d_shi1;
  wire mem_cns_we_shi0;
  wire mem_cns_we_shi1;
  wire mem_cns_re_shi0;
  wire mem_cns_re_shi1;
  wire [127:0] mem_cns_q_sho0;
  wire [127:0] mem_cns_q_sho1;
  wire mem_cns_S0_iff;
  wire mem_cns_S1_iff;
  wire mem_cns_S0_dmo;
  wire mem_cns_S1_dmo;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat;
  assign nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat = {paramsIn_rsc_dat_STRIDE
      , paramsIn_rsc_dat_FY , paramsIn_rsc_dat_FX , paramsIn_rsc_dat_IC1 , paramsIn_rsc_dat_OC1
      , paramsIn_rsc_dat_OX0 , paramsIn_rsc_dat_OY0 , paramsIn_rsc_dat_OX1 , paramsIn_rsc_dat_OY1};
  ccs_pipe_v5 #(.rscid(32'sd15),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) inputDoubleBufferWriterParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst),
      .din_vld(inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .din(inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .dout_rdy(paramsIn_rsc_rdy_ninputDoubleBufferWriter),
      .dout_vld(paramsIn_rsc_vld_ninputDoubleBufferWriter),
      .dout(paramsIn_rsc_dat_ninputDoubleBufferWriter),
      .sz(inputDoubleBufferWriterParams_unc_2),
      .sz_req(1'b0),
      .is_idle(inputDoubleBufferWriterParams_idle)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd128),
  .addr_width(32'sd9),
  .depth(32'sd512)) mem_cns_comp (
      .radr(mem_cns_radr_shi0),
      .wadr(mem_cns_wadr_shi0),
      .d(mem_cns_d_shi0),
      .we(mem_cns_we_shi0),
      .re(mem_cns_re_shi0),
      .clk(clk),
      .q(mem_cns_q_sho0)
    );
  ccs_ram_sync_1R1W #(.data_width(32'sd128),
  .addr_width(32'sd9),
  .depth(32'sd512)) mem_cns_comp_1 (
      .radr(mem_cns_radr_shi1),
      .wadr(mem_cns_wadr_shi1),
      .d(mem_cns_d_shi1),
      .we(mem_cns_we_shi1),
      .re(mem_cns_re_shi1),
      .clk(clk),
      .q(mem_cns_q_sho1)
    );
  InputDoubleBufferWriter_512_16_16 inputDoubleBufferWriter (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_ninputDoubleBufferWriter),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_ninputDoubleBufferWriter),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud),
      .din_rsc_dat(inputs_in_rsc_dat_value),
      .din_rsc_vld(inputs_in_rsc_vld),
      .din_rsc_rdy(din_rsc_rdy_ninputDoubleBufferWriter_bud),
      .dout_rsc_wadr(dout_rsc_wadr_ninputDoubleBufferWriter),
      .dout_rsc_d(dout_rsc_d_ninputDoubleBufferWriter),
      .dout_rsc_we(dout_rsc_we_ninputDoubleBufferWriter),
      .dout_rsc_req_vz(dout_rsc_req_vz_ninputDoubleBufferWriter),
      .dout_rsc_rls_lz(dout_rsc_rls_lz_ninputDoubleBufferWriter_bud)
    );
  InputDoubleBufferReader_512_16_16 inputDoubleBufferReader (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .paramsIn_rsc_vld(inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBufferReader_bud),
      .din_rsc_radr(din_rsc_radr_ninputDoubleBufferReader),
      .din_rsc_re(din_rsc_re_ninputDoubleBufferReader),
      .din_rsc_q(din_rsc_q_ninputDoubleBufferReader),
      .din_rsc_req_vz(din_rsc_req_vz_ninputDoubleBufferReader),
      .din_rsc_rls_lz(din_rsc_rls_lz_ninputDoubleBufferReader_bud),
      .dout_rsc_dat(dout_rsc_dat_ninputDoubleBufferReader),
      .dout_rsc_vld(dout_rsc_vld_ninputDoubleBufferReader_bud),
      .dout_rsc_rdy(inputs_out_rsc_rdy)
    );
  InputDoubleBuffer_512_16_16_run InputDoubleBuffer_512_16_16_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(nl_InputDoubleBuffer_512_16_16_run_inst_paramsIn_rsc_dat[143:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferWriterParams_cns_dat(inputDoubleBufferWriterParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferWriterParams_cns_vld(inputDoubleBufferWriterParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferWriterParams_cns_rdy(inputDoubleBufferWriterParams_cns_rdy_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferReaderParams_cns_dat(inputDoubleBufferReaderParams_cns_dat_nInputDoubleBuffer_512_16_16_run_inst),
      .inputDoubleBufferReaderParams_cns_vld(inputDoubleBufferReaderParams_cns_vld_nInputDoubleBuffer_512_16_16_run_inst_bud),
      .inputDoubleBufferReaderParams_cns_rdy(paramsIn_rsc_rdy_ninputDoubleBufferReader)
    );
  unreg_hier unreg (
      .in_0(mem_cns_S0_iff),
      .out_0(mem_cns_R0)
    );
  unreg_hier unreg_1 (
      .in_0(mem_cns_S1_iff),
      .out_0(mem_cns_R1)
    );
  InputDoubleBDjtfoem_cns_bctl InputDoubleBDjtfoem_cns_bctl_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_rdy_ninputDoubleBufferWriter(paramsIn_rsc_rdy_ninputDoubleBufferWriter),
      .din_rsc_rdy_ninputDoubleBufferWriter(din_rsc_rdy_ninputDoubleBufferWriter),
      .dout_rsc_wadr_ninputDoubleBufferWriter(dout_rsc_wadr_ninputDoubleBufferWriter),
      .dout_rsc_d_ninputDoubleBufferWriter(dout_rsc_d_ninputDoubleBufferWriter),
      .dout_rsc_we_ninputDoubleBufferWriter(dout_rsc_we_ninputDoubleBufferWriter),
      .dout_rsc_req_vz_ninputDoubleBufferWriter(dout_rsc_req_vz_ninputDoubleBufferWriter),
      .paramsIn_rsc_rdy_ninputDoubleBufferReader(paramsIn_rsc_rdy_ninputDoubleBufferReader),
      .din_rsc_radr_ninputDoubleBufferReader(din_rsc_radr_ninputDoubleBufferReader),
      .din_rsc_re_ninputDoubleBufferReader(din_rsc_re_ninputDoubleBufferReader),
      .din_rsc_q_ninputDoubleBufferReader(din_rsc_q_ninputDoubleBufferReader),
      .din_rsc_req_vz_ninputDoubleBufferReader(din_rsc_req_vz_ninputDoubleBufferReader),
      .dout_rsc_vld_ninputDoubleBufferReader(dout_rsc_vld_ninputDoubleBufferReader),
      .paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud(paramsIn_rsc_rdy_ninputDoubleBufferWriter_bud),
      .din_rsc_rdy_ninputDoubleBufferWriter_bud(din_rsc_rdy_ninputDoubleBufferWriter_bud),
      .dout_rsc_rls_lz_ninputDoubleBufferWriter_bud(dout_rsc_rls_lz_ninputDoubleBufferWriter_bud),
      .din_rsc_rls_lz_ninputDoubleBufferReader_bud(din_rsc_rls_lz_ninputDoubleBufferReader_bud),
      .paramsIn_rsc_rdy_ninputDoubleBufferReader_bud(paramsIn_rsc_rdy_ninputDoubleBufferReader_bud),
      .dout_rsc_vld_ninputDoubleBufferReader_bud(dout_rsc_vld_ninputDoubleBufferReader_bud),
      .mem_cns_S0(mem_cns_S0_dmo),
      .mem_cns_R0(mem_cns_R0),
      .mem_cns_S1(mem_cns_S1_dmo),
      .mem_cns_R1(mem_cns_R1),
      .mem_cns_radr_shi0(mem_cns_radr_shi0),
      .mem_cns_radr_shi1(mem_cns_radr_shi1),
      .mem_cns_wadr_shi0(mem_cns_wadr_shi0),
      .mem_cns_wadr_shi1(mem_cns_wadr_shi1),
      .mem_cns_d_shi0(mem_cns_d_shi0),
      .mem_cns_d_shi1(mem_cns_d_shi1),
      .mem_cns_we_shi0(mem_cns_we_shi0),
      .mem_cns_we_shi1(mem_cns_we_shi1),
      .mem_cns_re_shi0(mem_cns_re_shi0),
      .mem_cns_re_shi1(mem_cns_re_shi1),
      .mem_cns_q_sho0(mem_cns_q_sho0),
      .mem_cns_q_sho1(mem_cns_q_sho1),
      .mem_cns_S0_pff(mem_cns_S0_iff),
      .mem_cns_S1_pff(mem_cns_S1_iff)
    );
  assign inputs_out_rsc_dat_value = dout_rsc_dat_ninputDoubleBufferReader;
  assign inputs_in_rsc_rdy = din_rsc_rdy_ninputDoubleBufferWriter;
  assign inputs_out_rsc_vld = dout_rsc_vld_ninputDoubleBufferReader;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nInputDoubleBuffer_512_16_16_run_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputDoubleBuffer_512_16_16
// ------------------------------------------------------------------


module InputDoubleBuffer_512_16_16 (
  clk, arst_n, inputs_in_rsc_dat, inputs_in_rsc_vld, inputs_in_rsc_rdy, inputs_out_rsc_dat,
      inputs_out_rsc_vld, inputs_out_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputs_in_rsc_dat;
  input inputs_in_rsc_vld;
  output inputs_in_rsc_rdy;
  output [127:0] inputs_out_rsc_dat;
  output inputs_out_rsc_vld;
  input inputs_out_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [127:0] inputs_out_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE = paramsIn_rsc_dat[143:128];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY = paramsIn_rsc_dat[127:112];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX = paramsIn_rsc_dat[111:96];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1 = paramsIn_rsc_dat[95:80];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1 = paramsIn_rsc_dat[79:64];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0 = paramsIn_rsc_dat[63:48];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0 = paramsIn_rsc_dat[47:32];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1 = paramsIn_rsc_dat[31:16];
  wire [15:0] nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1;
  assign nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1 = paramsIn_rsc_dat[15:0];
  InputDoubleBuffer_512_16_16_struct InputDoubleBuffer_512_16_16_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputs_in_rsc_dat_value(inputs_in_rsc_dat),
      .inputs_in_rsc_vld(inputs_in_rsc_vld),
      .inputs_in_rsc_rdy(inputs_in_rsc_rdy),
      .inputs_out_rsc_dat_value(inputs_out_rsc_dat_value),
      .inputs_out_rsc_vld(inputs_out_rsc_vld),
      .inputs_out_rsc_rdy(inputs_out_rsc_rdy),
      .paramsIn_rsc_dat_STRIDE(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_STRIDE[15:0]),
      .paramsIn_rsc_dat_FY(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FY[15:0]),
      .paramsIn_rsc_dat_FX(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_FX[15:0]),
      .paramsIn_rsc_dat_IC1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_IC1[15:0]),
      .paramsIn_rsc_dat_OC1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OC1[15:0]),
      .paramsIn_rsc_dat_OX0(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX0[15:0]),
      .paramsIn_rsc_dat_OY0(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY0[15:0]),
      .paramsIn_rsc_dat_OX1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OX1[15:0]),
      .paramsIn_rsc_dat_OY1(nl_InputDoubleBuffer_512_16_16_struct_inst_paramsIn_rsc_dat_OY1[15:0]),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy)
    );
  assign inputs_out_rsc_dat = inputs_out_rsc_dat_value;
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   skavya@caddy09
//  Generated date: Thu Feb 20 23:21:09 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ParamsDeserializer_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;


  // FSM State Type Declaration for ParamsDeserializer_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8,
    main_C_8 = 4'd9,
    main_C_9 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ParamsDeserializer_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 11'b00000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_staller
// ------------------------------------------------------------------


module ParamsDeserializer_run_staller (
  run_wen, inputChannel_rsci_wen_comp, outputChannel1_rsci_wen_comp, outputChannel2_rsci_wen_comp,
      outputChannel3_rsci_wen_comp
);
  output run_wen;
  input inputChannel_rsci_wen_comp;
  input outputChannel1_rsci_wen_comp;
  input outputChannel2_rsci_wen_comp;
  input outputChannel3_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = inputChannel_rsci_wen_comp & outputChannel1_rsci_wen_comp & outputChannel2_rsci_wen_comp
      & outputChannel3_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp (
  clk, arst_n, outputChannel3_rsci_oswt, outputChannel3_rsci_wen_comp, outputChannel3_rsci_biwt,
      outputChannel3_rsci_bdwt, outputChannel3_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel3_rsci_oswt;
  output outputChannel3_rsci_wen_comp;
  input outputChannel3_rsci_biwt;
  input outputChannel3_rsci_bdwt;
  output outputChannel3_rsci_bcwt;
  reg outputChannel3_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel3_rsci_wen_comp = (~ outputChannel3_rsci_oswt) | outputChannel3_rsci_biwt
      | outputChannel3_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel3_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel3_rsci_bcwt <= ~((~(outputChannel3_rsci_bcwt | outputChannel3_rsci_biwt))
          | outputChannel3_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl (
  run_wen, outputChannel3_rsci_oswt, outputChannel3_rsci_irdy, outputChannel3_rsci_biwt,
      outputChannel3_rsci_bdwt, outputChannel3_rsci_bcwt, outputChannel3_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel3_rsci_oswt;
  input outputChannel3_rsci_irdy;
  output outputChannel3_rsci_biwt;
  output outputChannel3_rsci_bdwt;
  input outputChannel3_rsci_bcwt;
  output outputChannel3_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel3_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel3_rsci_bdwt = outputChannel3_rsci_oswt & run_wen;
  assign outputChannel3_rsci_biwt = outputChannel3_rsci_ogwt & outputChannel3_rsci_irdy;
  assign outputChannel3_rsci_ogwt = outputChannel3_rsci_oswt & (~ outputChannel3_rsci_bcwt);
  assign outputChannel3_rsci_ivld_run_sct = outputChannel3_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp (
  clk, arst_n, outputChannel2_rsci_oswt, outputChannel2_rsci_wen_comp, outputChannel2_rsci_biwt,
      outputChannel2_rsci_bdwt, outputChannel2_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel2_rsci_oswt;
  output outputChannel2_rsci_wen_comp;
  input outputChannel2_rsci_biwt;
  input outputChannel2_rsci_bdwt;
  output outputChannel2_rsci_bcwt;
  reg outputChannel2_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel2_rsci_wen_comp = (~ outputChannel2_rsci_oswt) | outputChannel2_rsci_biwt
      | outputChannel2_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel2_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel2_rsci_bcwt <= ~((~(outputChannel2_rsci_bcwt | outputChannel2_rsci_biwt))
          | outputChannel2_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl (
  run_wen, outputChannel2_rsci_oswt, outputChannel2_rsci_irdy, outputChannel2_rsci_biwt,
      outputChannel2_rsci_bdwt, outputChannel2_rsci_bcwt, outputChannel2_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel2_rsci_oswt;
  input outputChannel2_rsci_irdy;
  output outputChannel2_rsci_biwt;
  output outputChannel2_rsci_bdwt;
  input outputChannel2_rsci_bcwt;
  output outputChannel2_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel2_rsci_bdwt = outputChannel2_rsci_oswt & run_wen;
  assign outputChannel2_rsci_biwt = outputChannel2_rsci_ogwt & outputChannel2_rsci_irdy;
  assign outputChannel2_rsci_ogwt = outputChannel2_rsci_oswt & (~ outputChannel2_rsci_bcwt);
  assign outputChannel2_rsci_ivld_run_sct = outputChannel2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp (
  clk, arst_n, outputChannel1_rsci_oswt, outputChannel1_rsci_wen_comp, outputChannel1_rsci_biwt,
      outputChannel1_rsci_bdwt, outputChannel1_rsci_bcwt
);
  input clk;
  input arst_n;
  input outputChannel1_rsci_oswt;
  output outputChannel1_rsci_wen_comp;
  input outputChannel1_rsci_biwt;
  input outputChannel1_rsci_bdwt;
  output outputChannel1_rsci_bcwt;
  reg outputChannel1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign outputChannel1_rsci_wen_comp = (~ outputChannel1_rsci_oswt) | outputChannel1_rsci_biwt
      | outputChannel1_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      outputChannel1_rsci_bcwt <= 1'b0;
    end
    else begin
      outputChannel1_rsci_bcwt <= ~((~(outputChannel1_rsci_bcwt | outputChannel1_rsci_biwt))
          | outputChannel1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl (
  run_wen, outputChannel1_rsci_oswt, outputChannel1_rsci_irdy, outputChannel1_rsci_biwt,
      outputChannel1_rsci_bdwt, outputChannel1_rsci_bcwt, outputChannel1_rsci_ivld_run_sct
);
  input run_wen;
  input outputChannel1_rsci_oswt;
  input outputChannel1_rsci_irdy;
  output outputChannel1_rsci_biwt;
  output outputChannel1_rsci_bdwt;
  input outputChannel1_rsci_bcwt;
  output outputChannel1_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire outputChannel1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign outputChannel1_rsci_bdwt = outputChannel1_rsci_oswt & run_wen;
  assign outputChannel1_rsci_biwt = outputChannel1_rsci_ogwt & outputChannel1_rsci_irdy;
  assign outputChannel1_rsci_ogwt = outputChannel1_rsci_oswt & (~ outputChannel1_rsci_bcwt);
  assign outputChannel1_rsci_ivld_run_sct = outputChannel1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp (
  clk, arst_n, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt,
      inputChannel_rsci_biwt, inputChannel_rsci_bdwt, inputChannel_rsci_bcwt, inputChannel_rsci_idat
);
  input clk;
  input arst_n;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [15:0] inputChannel_rsci_idat_mxwt;
  input inputChannel_rsci_biwt;
  input inputChannel_rsci_bdwt;
  output inputChannel_rsci_bcwt;
  reg inputChannel_rsci_bcwt;
  input [15:0] inputChannel_rsci_idat;


  // Interconnect Declarations
  reg [15:0] inputChannel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_wen_comp = (~ inputChannel_rsci_oswt) | inputChannel_rsci_biwt
      | inputChannel_rsci_bcwt;
  assign inputChannel_rsci_idat_mxwt = MUX_v_16_2_2(inputChannel_rsci_idat, inputChannel_rsci_idat_bfwt,
      inputChannel_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      inputChannel_rsci_bcwt <= ~((~(inputChannel_rsci_bcwt | inputChannel_rsci_biwt))
          | inputChannel_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_idat_bfwt <= 16'b0000000000000000;
    end
    else if ( ~ inputChannel_rsci_bcwt ) begin
      inputChannel_rsci_idat_bfwt <= inputChannel_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl (
  run_wen, inputChannel_rsci_oswt, inputChannel_rsci_biwt, inputChannel_rsci_bdwt,
      inputChannel_rsci_bcwt, inputChannel_rsci_irdy_run_sct, inputChannel_rsci_ivld
);
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_biwt;
  output inputChannel_rsci_bdwt;
  input inputChannel_rsci_bcwt;
  output inputChannel_rsci_irdy_run_sct;
  input inputChannel_rsci_ivld;


  // Interconnect Declarations
  wire inputChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_bdwt = inputChannel_rsci_oswt & run_wen;
  assign inputChannel_rsci_biwt = inputChannel_rsci_ogwt & inputChannel_rsci_ivld;
  assign inputChannel_rsci_ogwt = inputChannel_rsci_oswt & (~ inputChannel_rsci_bcwt);
  assign inputChannel_rsci_irdy_run_sct = inputChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller (
  run_wen, inputChannel_rsci_wen_comp, serialOutChannel_rsci_wen_comp
);
  output run_wen;
  input inputChannel_rsci_wen_comp;
  input serialOutChannel_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = inputChannel_rsci_wen_comp & serialOutChannel_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
    (
  clk, arst_n, serialOutChannel_rsci_oswt, serialOutChannel_rsci_wen_comp, serialOutChannel_rsci_biwt,
      serialOutChannel_rsci_bdwt, serialOutChannel_rsci_bcwt
);
  input clk;
  input arst_n;
  input serialOutChannel_rsci_oswt;
  output serialOutChannel_rsci_wen_comp;
  input serialOutChannel_rsci_biwt;
  input serialOutChannel_rsci_bdwt;
  output serialOutChannel_rsci_bcwt;
  reg serialOutChannel_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign serialOutChannel_rsci_wen_comp = (~ serialOutChannel_rsci_oswt) | serialOutChannel_rsci_biwt
      | serialOutChannel_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      serialOutChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      serialOutChannel_rsci_bcwt <= ~((~(serialOutChannel_rsci_bcwt | serialOutChannel_rsci_biwt))
          | serialOutChannel_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
    (
  run_wen, serialOutChannel_rsci_oswt, serialOutChannel_rsci_irdy, serialOutChannel_rsci_biwt,
      serialOutChannel_rsci_bdwt, serialOutChannel_rsci_bcwt, serialOutChannel_rsci_ivld_run_sct
);
  input run_wen;
  input serialOutChannel_rsci_oswt;
  input serialOutChannel_rsci_irdy;
  output serialOutChannel_rsci_biwt;
  output serialOutChannel_rsci_bdwt;
  input serialOutChannel_rsci_bcwt;
  output serialOutChannel_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire serialOutChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign serialOutChannel_rsci_bdwt = serialOutChannel_rsci_oswt & run_wen;
  assign serialOutChannel_rsci_biwt = serialOutChannel_rsci_ogwt & serialOutChannel_rsci_irdy;
  assign serialOutChannel_rsci_ogwt = serialOutChannel_rsci_oswt & (~ serialOutChannel_rsci_bcwt);
  assign serialOutChannel_rsci_ivld_run_sct = serialOutChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
    (
  clk, arst_n, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt,
      inputChannel_rsci_biwt, inputChannel_rsci_bdwt, inputChannel_rsci_bcwt, inputChannel_rsci_idat
);
  input clk;
  input arst_n;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [255:0] inputChannel_rsci_idat_mxwt;
  input inputChannel_rsci_biwt;
  input inputChannel_rsci_bdwt;
  output inputChannel_rsci_bcwt;
  reg inputChannel_rsci_bcwt;
  input [255:0] inputChannel_rsci_idat;


  // Interconnect Declarations
  reg [255:0] inputChannel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_wen_comp = (~ inputChannel_rsci_oswt) | inputChannel_rsci_biwt
      | inputChannel_rsci_bcwt;
  assign inputChannel_rsci_idat_mxwt = MUX_v_256_2_2(inputChannel_rsci_idat, inputChannel_rsci_idat_bfwt,
      inputChannel_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      inputChannel_rsci_bcwt <= ~((~(inputChannel_rsci_bcwt | inputChannel_rsci_biwt))
          | inputChannel_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_idat_bfwt <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ inputChannel_rsci_bcwt ) begin
      inputChannel_rsci_idat_bfwt <= inputChannel_rsci_idat_mxwt;
    end
  end

  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
    (
  run_wen, inputChannel_rsci_oswt, inputChannel_rsci_biwt, inputChannel_rsci_bdwt,
      inputChannel_rsci_bcwt, inputChannel_rsci_irdy_run_sct, inputChannel_rsci_ivld
);
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_biwt;
  output inputChannel_rsci_bdwt;
  input inputChannel_rsci_bcwt;
  output inputChannel_rsci_irdy_run_sct;
  input inputChannel_rsci_ivld;


  // Interconnect Declarations
  wire inputChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_bdwt = inputChannel_rsci_oswt & run_wen;
  assign inputChannel_rsci_biwt = inputChannel_rsci_ogwt & inputChannel_rsci_ivld;
  assign inputChannel_rsci_ogwt = inputChannel_rsci_oswt & (~ inputChannel_rsci_bcwt);
  assign inputChannel_rsci_irdy_run_sct = inputChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module SystolicArrayLooper_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, main_C_1_tr0, xy_o_C_0_tr0, OC2_C_0_tr0, co_C_0_tr0,
      winx_C_0_tr0, winy_C_0_tr0, winx_C_1_tr0, co_C_1_tr0, OC2_C_1_tr0, xy_o_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [11:0] fsm_output;
  reg [11:0] fsm_output;
  input main_C_1_tr0;
  input xy_o_C_0_tr0;
  input OC2_C_0_tr0;
  input co_C_0_tr0;
  input winx_C_0_tr0;
  input winy_C_0_tr0;
  input winx_C_1_tr0;
  input co_C_1_tr0;
  input OC2_C_1_tr0;
  input xy_o_C_1_tr0;


  // FSM State Type Declaration for SystolicArrayLooper_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    xy_o_C_0 = 4'd3,
    OC2_C_0 = 4'd4,
    co_C_0 = 4'd5,
    winx_C_0 = 4'd6,
    winy_C_0 = 4'd7,
    winx_C_1 = 4'd8,
    co_C_1 = 4'd9,
    OC2_C_1 = 4'd10,
    xy_o_C_1 = 4'd11;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SystolicArrayLooper_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 12'b000000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 12'b000000000100;
        if ( main_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = xy_o_C_0;
        end
      end
      xy_o_C_0 : begin
        fsm_output = 12'b000000001000;
        if ( xy_o_C_0_tr0 ) begin
          state_var_NS = xy_o_C_1;
        end
        else begin
          state_var_NS = OC2_C_0;
        end
      end
      OC2_C_0 : begin
        fsm_output = 12'b000000010000;
        if ( OC2_C_0_tr0 ) begin
          state_var_NS = OC2_C_1;
        end
        else begin
          state_var_NS = co_C_0;
        end
      end
      co_C_0 : begin
        fsm_output = 12'b000000100000;
        if ( co_C_0_tr0 ) begin
          state_var_NS = co_C_1;
        end
        else begin
          state_var_NS = winx_C_0;
        end
      end
      winx_C_0 : begin
        fsm_output = 12'b000001000000;
        if ( winx_C_0_tr0 ) begin
          state_var_NS = winx_C_1;
        end
        else begin
          state_var_NS = winy_C_0;
        end
      end
      winy_C_0 : begin
        fsm_output = 12'b000010000000;
        if ( winy_C_0_tr0 ) begin
          state_var_NS = winx_C_1;
        end
        else begin
          state_var_NS = winy_C_0;
        end
      end
      winx_C_1 : begin
        fsm_output = 12'b000100000000;
        if ( winx_C_1_tr0 ) begin
          state_var_NS = co_C_1;
        end
        else begin
          state_var_NS = winx_C_0;
        end
      end
      co_C_1 : begin
        fsm_output = 12'b001000000000;
        if ( co_C_1_tr0 ) begin
          state_var_NS = OC2_C_1;
        end
        else begin
          state_var_NS = co_C_0;
        end
      end
      OC2_C_1 : begin
        fsm_output = 12'b010000000000;
        if ( OC2_C_1_tr0 ) begin
          state_var_NS = xy_o_C_1;
        end
        else begin
          state_var_NS = OC2_C_0;
        end
      end
      xy_o_C_1 : begin
        fsm_output = 12'b100000000000;
        if ( xy_o_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = xy_o_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 12'b000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_staller
// ------------------------------------------------------------------


module SystolicArrayLooper_run_staller (
  run_wen, paramsIn_rsci_wen_comp, paramsOut_rsci_wen_comp, loopIndicesOut_rsci_wen_comp
);
  output run_wen;
  input paramsIn_rsci_wen_comp;
  input paramsOut_rsci_wen_comp;
  input loopIndicesOut_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = paramsIn_rsci_wen_comp & paramsOut_rsci_wen_comp & loopIndicesOut_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp (
  clk, arst_n, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input loopIndicesOut_rsci_biwt;
  input loopIndicesOut_rsci_bdwt;
  output loopIndicesOut_rsci_bcwt;
  reg loopIndicesOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_wen_comp = (~ loopIndicesOut_rsci_oswt) | loopIndicesOut_rsci_biwt
      | loopIndicesOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_bcwt <= 1'b0;
    end
    else begin
      loopIndicesOut_rsci_bcwt <= ~((~(loopIndicesOut_rsci_bcwt | loopIndicesOut_rsci_biwt))
          | loopIndicesOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl (
  run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_irdy, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt, loopIndicesOut_rsci_ivld_run_sct
);
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  input loopIndicesOut_rsci_irdy;
  output loopIndicesOut_rsci_biwt;
  output loopIndicesOut_rsci_bdwt;
  input loopIndicesOut_rsci_bcwt;
  output loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_bdwt = loopIndicesOut_rsci_oswt & run_wen;
  assign loopIndicesOut_rsci_biwt = loopIndicesOut_rsci_ogwt & loopIndicesOut_rsci_irdy;
  assign loopIndicesOut_rsci_ogwt = loopIndicesOut_rsci_oswt & (~ loopIndicesOut_rsci_bcwt);
  assign loopIndicesOut_rsci_ivld_run_sct = loopIndicesOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp (
  clk, arst_n, paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_biwt,
      paramsOut_rsci_bdwt, paramsOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input paramsOut_rsci_biwt;
  input paramsOut_rsci_bdwt;
  output paramsOut_rsci_bcwt;
  reg paramsOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_wen_comp = (~ paramsOut_rsci_oswt) | paramsOut_rsci_biwt
      | paramsOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsOut_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsOut_rsci_bcwt <= ~((~(paramsOut_rsci_bcwt | paramsOut_rsci_biwt)) | paramsOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl (
  run_wen, paramsOut_rsci_oswt, paramsOut_rsci_irdy, paramsOut_rsci_biwt, paramsOut_rsci_bdwt,
      paramsOut_rsci_bcwt, paramsOut_rsci_ivld_run_sct
);
  input run_wen;
  input paramsOut_rsci_oswt;
  input paramsOut_rsci_irdy;
  output paramsOut_rsci_biwt;
  output paramsOut_rsci_bdwt;
  input paramsOut_rsci_bcwt;
  output paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire paramsOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_bdwt = paramsOut_rsci_oswt & run_wen;
  assign paramsOut_rsci_biwt = paramsOut_rsci_ogwt & paramsOut_rsci_irdy;
  assign paramsOut_rsci_ogwt = paramsOut_rsci_oswt & (~ paramsOut_rsci_bcwt);
  assign paramsOut_rsci_ivld_run_sct = paramsOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [143:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_144_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [143:0] MUX_v_144_2_2;
    input [143:0] input_0;
    input [143:0] input_1;
    input [0:0] sel;
    reg [143:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_144_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel3_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel3_rsci (
  clk, arst_n, outputChannel3_rsc_dat, outputChannel3_rsc_vld, outputChannel3_rsc_rdy,
      run_wen, outputChannel3_rsci_oswt, outputChannel3_rsci_wen_comp, outputChannel3_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;
  input run_wen;
  input outputChannel3_rsci_oswt;
  output outputChannel3_rsci_wen_comp;
  input [143:0] outputChannel3_rsci_idat;


  // Interconnect Declarations
  wire outputChannel3_rsci_irdy;
  wire outputChannel3_rsci_biwt;
  wire outputChannel3_rsci_bdwt;
  wire outputChannel3_rsci_bcwt;
  wire outputChannel3_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd144)) outputChannel3_rsci (
      .irdy(outputChannel3_rsci_irdy),
      .ivld(outputChannel3_rsci_ivld_run_sct),
      .idat(outputChannel3_rsci_idat),
      .rdy(outputChannel3_rsc_rdy),
      .vld(outputChannel3_rsc_vld),
      .dat(outputChannel3_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel3_rsci_oswt(outputChannel3_rsci_oswt),
      .outputChannel3_rsci_irdy(outputChannel3_rsci_irdy),
      .outputChannel3_rsci_biwt(outputChannel3_rsci_biwt),
      .outputChannel3_rsci_bdwt(outputChannel3_rsci_bdwt),
      .outputChannel3_rsci_bcwt(outputChannel3_rsci_bcwt),
      .outputChannel3_rsci_ivld_run_sct(outputChannel3_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp ParamsDeserializer_run_outputChannel3_rsci_outputChannel3_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel3_rsci_oswt(outputChannel3_rsci_oswt),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp),
      .outputChannel3_rsci_biwt(outputChannel3_rsci_biwt),
      .outputChannel3_rsci_bdwt(outputChannel3_rsci_bdwt),
      .outputChannel3_rsci_bcwt(outputChannel3_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel2_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel2_rsci (
  clk, arst_n, outputChannel2_rsc_dat, outputChannel2_rsc_vld, outputChannel2_rsc_rdy,
      run_wen, outputChannel2_rsci_oswt, outputChannel2_rsci_wen_comp, outputChannel2_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  input run_wen;
  input outputChannel2_rsci_oswt;
  output outputChannel2_rsci_wen_comp;
  input [143:0] outputChannel2_rsci_idat;


  // Interconnect Declarations
  wire outputChannel2_rsci_irdy;
  wire outputChannel2_rsci_biwt;
  wire outputChannel2_rsci_bdwt;
  wire outputChannel2_rsci_bcwt;
  wire outputChannel2_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd144)) outputChannel2_rsci (
      .irdy(outputChannel2_rsci_irdy),
      .ivld(outputChannel2_rsci_ivld_run_sct),
      .idat(outputChannel2_rsci_idat),
      .rdy(outputChannel2_rsc_rdy),
      .vld(outputChannel2_rsc_vld),
      .dat(outputChannel2_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel2_rsci_oswt(outputChannel2_rsci_oswt),
      .outputChannel2_rsci_irdy(outputChannel2_rsci_irdy),
      .outputChannel2_rsci_biwt(outputChannel2_rsci_biwt),
      .outputChannel2_rsci_bdwt(outputChannel2_rsci_bdwt),
      .outputChannel2_rsci_bcwt(outputChannel2_rsci_bcwt),
      .outputChannel2_rsci_ivld_run_sct(outputChannel2_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp ParamsDeserializer_run_outputChannel2_rsci_outputChannel2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel2_rsci_oswt(outputChannel2_rsci_oswt),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel2_rsci_biwt(outputChannel2_rsci_biwt),
      .outputChannel2_rsci_bdwt(outputChannel2_rsci_bdwt),
      .outputChannel2_rsci_bcwt(outputChannel2_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_outputChannel1_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_outputChannel1_rsci (
  clk, arst_n, outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy,
      run_wen, outputChannel1_rsci_oswt, outputChannel1_rsci_wen_comp, outputChannel1_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  input run_wen;
  input outputChannel1_rsci_oswt;
  output outputChannel1_rsci_wen_comp;
  input [143:0] outputChannel1_rsci_idat;


  // Interconnect Declarations
  wire outputChannel1_rsci_irdy;
  wire outputChannel1_rsci_biwt;
  wire outputChannel1_rsci_bdwt;
  wire outputChannel1_rsci_bcwt;
  wire outputChannel1_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd144)) outputChannel1_rsci (
      .irdy(outputChannel1_rsci_irdy),
      .ivld(outputChannel1_rsci_ivld_run_sct),
      .idat(outputChannel1_rsci_idat),
      .rdy(outputChannel1_rsc_rdy),
      .vld(outputChannel1_rsc_vld),
      .dat(outputChannel1_rsc_dat)
    );
  ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .outputChannel1_rsci_oswt(outputChannel1_rsci_oswt),
      .outputChannel1_rsci_irdy(outputChannel1_rsci_irdy),
      .outputChannel1_rsci_biwt(outputChannel1_rsci_biwt),
      .outputChannel1_rsci_bdwt(outputChannel1_rsci_bdwt),
      .outputChannel1_rsci_bcwt(outputChannel1_rsci_bcwt),
      .outputChannel1_rsci_ivld_run_sct(outputChannel1_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp ParamsDeserializer_run_outputChannel1_rsci_outputChannel1_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel1_rsci_oswt(outputChannel1_rsci_oswt),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel1_rsci_biwt(outputChannel1_rsci_biwt),
      .outputChannel1_rsci_bdwt(outputChannel1_rsci_bdwt),
      .outputChannel1_rsci_bcwt(outputChannel1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      run_wen, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [15:0] inputChannel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire inputChannel_rsci_biwt;
  wire inputChannel_rsci_bdwt;
  wire inputChannel_rsci_bcwt;
  wire inputChannel_rsci_irdy_run_sct;
  wire inputChannel_rsci_ivld;
  wire [15:0] inputChannel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd16)) inputChannel_rsci (
      .rdy(inputChannel_rsc_rdy),
      .vld(inputChannel_rsc_vld),
      .dat(inputChannel_rsc_dat),
      .irdy(inputChannel_rsci_irdy_run_sct),
      .ivld(inputChannel_rsci_ivld),
      .idat(inputChannel_rsci_idat)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_irdy_run_sct(inputChannel_rsci_irdy_run_sct),
      .inputChannel_rsci_ivld(inputChannel_rsci_ivld)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_idat(inputChannel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci (
  clk, arst_n, serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy,
      run_wen, serialOutChannel_rsci_oswt, serialOutChannel_rsci_wen_comp, serialOutChannel_rsci_idat
);
  input clk;
  input arst_n;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;
  input run_wen;
  input serialOutChannel_rsci_oswt;
  output serialOutChannel_rsci_wen_comp;
  input [15:0] serialOutChannel_rsci_idat;


  // Interconnect Declarations
  wire serialOutChannel_rsci_irdy;
  wire serialOutChannel_rsci_biwt;
  wire serialOutChannel_rsci_bdwt;
  wire serialOutChannel_rsci_bcwt;
  wire serialOutChannel_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd6),
  .width(32'sd16)) serialOutChannel_rsci (
      .irdy(serialOutChannel_rsci_irdy),
      .ivld(serialOutChannel_rsci_ivld_run_sct),
      .idat(serialOutChannel_rsci_idat),
      .rdy(serialOutChannel_rsc_rdy),
      .vld(serialOutChannel_rsc_vld),
      .dat(serialOutChannel_rsc_dat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .serialOutChannel_rsci_oswt(serialOutChannel_rsci_oswt),
      .serialOutChannel_rsci_irdy(serialOutChannel_rsci_irdy),
      .serialOutChannel_rsci_biwt(serialOutChannel_rsci_biwt),
      .serialOutChannel_rsci_bdwt(serialOutChannel_rsci_bdwt),
      .serialOutChannel_rsci_bcwt(serialOutChannel_rsci_bcwt),
      .serialOutChannel_rsci_ivld_run_sct(serialOutChannel_rsci_ivld_run_sct)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_serialOutChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .serialOutChannel_rsci_oswt(serialOutChannel_rsci_oswt),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp),
      .serialOutChannel_rsci_biwt(serialOutChannel_rsci_biwt),
      .serialOutChannel_rsci_bdwt(serialOutChannel_rsci_bdwt),
      .serialOutChannel_rsci_bcwt(serialOutChannel_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      run_wen, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [255:0] inputChannel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire inputChannel_rsci_biwt;
  wire inputChannel_rsci_bdwt;
  wire inputChannel_rsci_bcwt;
  wire inputChannel_rsci_irdy_run_sct;
  wire inputChannel_rsci_ivld;
  wire [255:0] inputChannel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd256)) inputChannel_rsci (
      .rdy(inputChannel_rsc_rdy),
      .vld(inputChannel_rsc_vld),
      .dat(inputChannel_rsc_dat),
      .irdy(inputChannel_rsci_irdy_run_sct),
      .ivld(inputChannel_rsci_ivld),
      .idat(inputChannel_rsci_idat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_irdy_run_sct(inputChannel_rsci_irdy_run_sct),
      .inputChannel_rsci_ivld(inputChannel_rsci_ivld)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp
      Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inputChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_idat(inputChannel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_loopIndicesOut_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_loopIndicesOut_rsci (
  clk, arst_n, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld, loopIndicesOut_rsc_rdy,
      run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_idat
);
  input clk;
  input arst_n;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input [47:0] loopIndicesOut_rsci_idat;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_irdy;
  wire loopIndicesOut_rsci_biwt;
  wire loopIndicesOut_rsci_bdwt;
  wire loopIndicesOut_rsci_bcwt;
  wire loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd158),
  .width(32'sd48)) loopIndicesOut_rsci (
      .irdy(loopIndicesOut_rsci_irdy),
      .ivld(loopIndicesOut_rsci_ivld_run_sct),
      .idat(loopIndicesOut_rsci_idat),
      .rdy(loopIndicesOut_rsc_rdy),
      .vld(loopIndicesOut_rsc_vld),
      .dat(loopIndicesOut_rsc_dat)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_irdy(loopIndicesOut_rsci_irdy),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt),
      .loopIndicesOut_rsci_ivld_run_sct(loopIndicesOut_rsci_ivld_run_sct)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp SystolicArrayLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsOut_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsOut_rsci (
  clk, arst_n, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy, run_wen,
      paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_idat
);
  input clk;
  input arst_n;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  input run_wen;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input [143:0] paramsOut_rsci_idat;


  // Interconnect Declarations
  wire paramsOut_rsci_irdy;
  wire paramsOut_rsci_biwt;
  wire paramsOut_rsci_bdwt;
  wire paramsOut_rsci_bcwt;
  wire paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd157),
  .width(32'sd144)) paramsOut_rsci (
      .irdy(paramsOut_rsci_irdy),
      .ivld(paramsOut_rsci_ivld_run_sct),
      .idat(paramsOut_rsci_idat),
      .rdy(paramsOut_rsc_rdy),
      .vld(paramsOut_rsc_vld),
      .dat(paramsOut_rsc_dat)
    );
  SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_irdy(paramsOut_rsci_irdy),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt),
      .paramsOut_rsci_ivld_run_sct(paramsOut_rsci_ivld_run_sct)
    );
  SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp SystolicArrayLooper_run_paramsOut_rsci_paramsOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run_paramsIn_rsci
// ------------------------------------------------------------------


module SystolicArrayLooper_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [143:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [143:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd156),
  .width(32'sd144)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp SystolicArrayLooper_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run
// ------------------------------------------------------------------


module ParamsDeserializer_run (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy, outputChannel2_rsc_dat,
      outputChannel2_rsc_vld, outputChannel2_rsc_rdy, outputChannel3_rsc_dat, outputChannel3_rsc_vld,
      outputChannel3_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire inputChannel_rsci_wen_comp;
  wire [15:0] inputChannel_rsci_idat_mxwt;
  wire outputChannel1_rsci_wen_comp;
  wire outputChannel2_rsci_wen_comp;
  wire outputChannel3_rsci_wen_comp;
  wire [10:0] fsm_output;
  wire outputChannel3_and_cse;
  reg reg_outputChannel3_rsci_ivld_run_psct_cse;
  reg reg_inputChannel_rsci_irdy_run_psct_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_15_0_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_31_16_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_47_32_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_63_48_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_79_64_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_95_80_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_111_96_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_127_112_cse;
  reg [15:0] reg_outputChannel3_rsci_idat_143_128_cse;
  reg [15:0] params_OY1_sva;
  reg [15:0] params_OX1_sva;
  reg [15:0] params_OY0_sva;
  reg [15:0] params_OX0_sva;
  reg [15:0] params_OC1_sva;
  reg [15:0] params_IC1_sva;
  reg [15:0] params_FX_sva;
  reg [15:0] params_FY_sva;


  // Interconnect Declarations for Component Instantiations 
  wire [143:0] nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  wire [143:0] nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  wire [143:0] nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat;
  assign nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat
      = {reg_outputChannel3_rsci_idat_143_128_cse , reg_outputChannel3_rsci_idat_127_112_cse
      , reg_outputChannel3_rsci_idat_111_96_cse , reg_outputChannel3_rsci_idat_95_80_cse
      , reg_outputChannel3_rsci_idat_79_64_cse , reg_outputChannel3_rsci_idat_63_48_cse
      , reg_outputChannel3_rsci_idat_47_32_cse , reg_outputChannel3_rsci_idat_31_16_cse
      , reg_outputChannel3_rsci_idat_15_0_cse};
  ParamsDeserializer_run_inputChannel_rsci ParamsDeserializer_run_inputChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(reg_inputChannel_rsci_irdy_run_psct_cse),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt)
    );
  ParamsDeserializer_run_outputChannel1_rsci ParamsDeserializer_run_outputChannel1_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel1_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel1_rsci_idat(nl_ParamsDeserializer_run_outputChannel1_rsci_inst_outputChannel1_rsci_idat[143:0])
    );
  ParamsDeserializer_run_outputChannel2_rsci ParamsDeserializer_run_outputChannel2_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel2_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel2_rsci_idat(nl_ParamsDeserializer_run_outputChannel2_rsci_inst_outputChannel2_rsci_idat[143:0])
    );
  ParamsDeserializer_run_outputChannel3_rsci ParamsDeserializer_run_outputChannel3_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy),
      .run_wen(run_wen),
      .outputChannel3_rsci_oswt(reg_outputChannel3_rsci_ivld_run_psct_cse),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp),
      .outputChannel3_rsci_idat(nl_ParamsDeserializer_run_outputChannel3_rsci_inst_outputChannel3_rsci_idat[143:0])
    );
  ParamsDeserializer_run_staller ParamsDeserializer_run_staller_inst (
      .run_wen(run_wen),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .outputChannel1_rsci_wen_comp(outputChannel1_rsci_wen_comp),
      .outputChannel2_rsci_wen_comp(outputChannel2_rsci_wen_comp),
      .outputChannel3_rsci_wen_comp(outputChannel3_rsci_wen_comp)
    );
  ParamsDeserializer_run_run_fsm ParamsDeserializer_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign outputChannel3_and_cse = run_wen & (fsm_output[9]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_outputChannel3_rsci_idat_15_0_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_31_16_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_47_32_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_63_48_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_79_64_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_95_80_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_111_96_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_127_112_cse <= 16'b0000000000000000;
      reg_outputChannel3_rsci_idat_143_128_cse <= 16'b0000000000000000;
    end
    else if ( outputChannel3_and_cse ) begin
      reg_outputChannel3_rsci_idat_15_0_cse <= params_OY1_sva;
      reg_outputChannel3_rsci_idat_31_16_cse <= params_OX1_sva;
      reg_outputChannel3_rsci_idat_47_32_cse <= params_OY0_sva;
      reg_outputChannel3_rsci_idat_63_48_cse <= params_OX0_sva;
      reg_outputChannel3_rsci_idat_79_64_cse <= params_OC1_sva;
      reg_outputChannel3_rsci_idat_95_80_cse <= params_IC1_sva;
      reg_outputChannel3_rsci_idat_111_96_cse <= params_FX_sva;
      reg_outputChannel3_rsci_idat_127_112_cse <= params_FY_sva;
      reg_outputChannel3_rsci_idat_143_128_cse <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_outputChannel3_rsci_ivld_run_psct_cse <= 1'b0;
      reg_inputChannel_rsci_irdy_run_psct_cse <= 1'b0;
      params_FY_sva <= 16'b0000000000000000;
    end
    else if ( run_wen ) begin
      reg_outputChannel3_rsci_ivld_run_psct_cse <= fsm_output[9];
      reg_inputChannel_rsci_irdy_run_psct_cse <= ~ (fsm_output[9]);
      params_FY_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OY1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[1]) ) begin
      params_OY1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OX1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      params_OX1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OY0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[3]) ) begin
      params_OY0_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OX0_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[4]) ) begin
      params_OX0_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_OC1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[5]) ) begin
      params_OC1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_IC1_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[6]) ) begin
      params_IC1_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_FX_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & (fsm_output[7]) ) begin
      params_FX_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16_run
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16_run (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire inputChannel_rsci_wen_comp;
  wire [255:0] inputChannel_rsci_idat_mxwt;
  wire serialOutChannel_rsci_wen_comp;
  reg [15:0] serialOutChannel_rsci_idat;
  wire [1:0] fsm_output;
  reg exitL_exit_for_sva;
  wire [4:0] for_i_4_0_sva_3;
  wire [5:0] nl_for_i_4_0_sva_3;
  reg reg_inputChannel_rsci_oswt_cse;
  reg reg_serialOutChannel_rsci_ivld_run_psct_cse;
  wire serialOutChannel_and_cse;
  reg [255:0] input_value_lpi_1_dfm;
  wire [255:0] input_value_lpi_1_dfm_mx0;
  wire [3:0] for_i_4_0_lpi_1_dfm_3_0_1;
  reg [3:0] for_i_4_0_sva_1_3_0;

  wire[0:0] for_not_nl;

  // Interconnect Declarations for Component Instantiations 
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inputChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(reg_inputChannel_rsci_oswt_cse),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_serialOutChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld),
      .serialOutChannel_rsc_rdy(serialOutChannel_rsc_rdy),
      .run_wen(run_wen),
      .serialOutChannel_rsci_oswt(reg_serialOutChannel_rsci_ivld_run_psct_cse),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp),
      .serialOutChannel_rsci_idat(serialOutChannel_rsci_idat)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_staller_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .serialOutChannel_rsci_wen_comp(serialOutChannel_rsci_wen_comp)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign serialOutChannel_and_cse = run_wen & (~ (fsm_output[0]));
  assign input_value_lpi_1_dfm_mx0 = MUX_v_256_2_2(input_value_lpi_1_dfm, inputChannel_rsci_idat_mxwt,
      exitL_exit_for_sva);
  assign nl_for_i_4_0_sva_3 = conv_u2s_4_5(for_i_4_0_lpi_1_dfm_3_0_1) + 5'b00001;
  assign for_i_4_0_sva_3 = nl_for_i_4_0_sva_3[4:0];
  assign for_not_nl = ~ exitL_exit_for_sva;
  assign for_i_4_0_lpi_1_dfm_3_0_1 = MUX_v_4_2_2(4'b0000, for_i_4_0_sva_1_3_0, (for_not_nl));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_inputChannel_rsci_oswt_cse <= 1'b0;
      reg_serialOutChannel_rsci_ivld_run_psct_cse <= 1'b0;
      for_i_4_0_sva_1_3_0 <= 4'b0000;
    end
    else if ( run_wen ) begin
      reg_inputChannel_rsci_oswt_cse <= ~((~ (for_i_4_0_sva_3[4])) & (fsm_output[1]));
      reg_serialOutChannel_rsci_ivld_run_psct_cse <= fsm_output[1];
      for_i_4_0_sva_1_3_0 <= for_i_4_0_sva_3[3:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      serialOutChannel_rsci_idat <= 16'b0000000000000000;
      exitL_exit_for_sva <= 1'b1;
    end
    else if ( serialOutChannel_and_cse ) begin
      serialOutChannel_rsci_idat <= MUX_v_16_16_2((input_value_lpi_1_dfm_mx0[15:0]),
          (input_value_lpi_1_dfm_mx0[31:16]), (input_value_lpi_1_dfm_mx0[47:32]),
          (input_value_lpi_1_dfm_mx0[63:48]), (input_value_lpi_1_dfm_mx0[79:64]),
          (input_value_lpi_1_dfm_mx0[95:80]), (input_value_lpi_1_dfm_mx0[111:96]),
          (input_value_lpi_1_dfm_mx0[127:112]), (input_value_lpi_1_dfm_mx0[143:128]),
          (input_value_lpi_1_dfm_mx0[159:144]), (input_value_lpi_1_dfm_mx0[175:160]),
          (input_value_lpi_1_dfm_mx0[191:176]), (input_value_lpi_1_dfm_mx0[207:192]),
          (input_value_lpi_1_dfm_mx0[223:208]), (input_value_lpi_1_dfm_mx0[239:224]),
          (input_value_lpi_1_dfm_mx0[255:240]), for_i_4_0_lpi_1_dfm_3_0_1);
      exitL_exit_for_sva <= for_i_4_0_sva_3[4];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      input_value_lpi_1_dfm <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (~ (for_i_4_0_sva_3[4])) & run_wen & exitL_exit_for_sva ) begin
      input_value_lpi_1_dfm <= input_value_lpi_1_dfm_mx0;
    end
  end

  function automatic [15:0] MUX_v_16_16_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_16_16_2 = result;
  end
  endfunction


  function automatic [255:0] MUX_v_256_2_2;
    input [255:0] input_0;
    input [255:0] input_1;
    input [0:0] sel;
    reg [255:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_256_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper_run
// ------------------------------------------------------------------


module SystolicArrayLooper_run (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat,
      paramsOut_rsc_vld, paramsOut_rsc_rdy, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld,
      loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire paramsIn_rsci_wen_comp;
  wire [143:0] paramsIn_rsci_idat_mxwt;
  wire paramsOut_rsci_wen_comp;
  reg [143:0] paramsOut_rsci_idat;
  wire loopIndicesOut_rsci_wen_comp;
  reg [15:0] loopIndicesOut_rsci_idat_47_32;
  reg [15:0] loopIndicesOut_rsci_idat_31_16;
  reg [15:0] loopIndicesOut_rsci_idat_15_0;
  wire [11:0] fsm_output;
  wire loopIndicesOut_and_cse;
  reg reg_loopIndicesOut_rsci_ivld_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
  wire [15:0] z_out_1;
  wire [16:0] nl_z_out_1;
  reg [143:0] paramsIn_crt_sva;
  reg [15:0] xy_o_p_sva;
  reg [15:0] OC2_koo_idx_sva;
  reg [15:0] co_c_idx_sva;
  reg [15:0] winx_wx_idx_sva;
  reg [31:0] xy_o_mul_1_itm;
  wire loopIndicesOut_rsci_idat_47_32_mx0c0;
  wire xy_o_and_cse;
  wire [16:0] z_out_32_16;

  wire[0:0] loopIndicesOut_not_1_nl;
  wire[33:0] acc_nl;
  wire[34:0] nl_acc_nl;
  wire[0:0] xy_o_xy_o_or_16_nl;
  wire[0:0] xy_o_xy_o_or_17_nl;
  wire[0:0] xy_o_xy_o_or_18_nl;
  wire[0:0] xy_o_xy_o_or_19_nl;
  wire[0:0] xy_o_xy_o_or_20_nl;
  wire[0:0] xy_o_xy_o_or_21_nl;
  wire[0:0] xy_o_xy_o_or_22_nl;
  wire[0:0] xy_o_xy_o_or_23_nl;
  wire[0:0] xy_o_xy_o_or_24_nl;
  wire[0:0] xy_o_xy_o_or_25_nl;
  wire[0:0] xy_o_xy_o_or_26_nl;
  wire[0:0] xy_o_xy_o_or_27_nl;
  wire[0:0] xy_o_xy_o_or_28_nl;
  wire[0:0] xy_o_xy_o_or_29_nl;
  wire[0:0] xy_o_xy_o_or_30_nl;
  wire[0:0] xy_o_xy_o_or_31_nl;
  wire[15:0] xy_o_mux1h_3_nl;
  wire[0:0] xy_o_or_3_nl;
  wire[0:0] xy_o_or_4_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_16_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_17_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_18_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_19_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_20_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_21_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_22_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_23_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_24_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_25_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_26_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_27_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_28_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_29_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_30_nl;
  wire[0:0] xy_o_xy_o_xy_o_nor_31_nl;
  wire[15:0] xy_o_mux1h_4_nl;
  wire[0:0] xy_o_or_5_nl;
  wire[15:0] winy_mux1h_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat;
  assign nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat
      = {loopIndicesOut_rsci_idat_47_32 , loopIndicesOut_rsci_idat_31_16 , loopIndicesOut_rsci_idat_15_0};
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_main_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_main_C_1_tr0 = ~ (z_out_32_16[16]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0 = ~ (z_out_32_16[0]);
  wire [0:0] nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0;
  assign nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0 = ~ (z_out_32_16[16]);
  SystolicArrayLooper_run_paramsIn_rsci SystolicArrayLooper_run_paramsIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  SystolicArrayLooper_run_paramsOut_rsci SystolicArrayLooper_run_paramsOut_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_idat(paramsOut_rsci_idat)
    );
  SystolicArrayLooper_run_loopIndicesOut_rsci SystolicArrayLooper_run_loopIndicesOut_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_idat(nl_SystolicArrayLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat[47:0])
    );
  SystolicArrayLooper_run_staller SystolicArrayLooper_run_staller_inst (
      .run_wen(run_wen),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp)
    );
  SystolicArrayLooper_run_run_fsm SystolicArrayLooper_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .main_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_main_C_1_tr0[0:0]),
      .xy_o_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_0_tr0[0:0]),
      .OC2_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_0_tr0[0:0]),
      .co_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_co_C_0_tr0[0:0]),
      .winx_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_0_tr0[0:0]),
      .winy_C_0_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winy_C_0_tr0[0:0]),
      .winx_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_winx_C_1_tr0[0:0]),
      .co_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_co_C_1_tr0[0:0]),
      .OC2_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_OC2_C_1_tr0[0:0]),
      .xy_o_C_1_tr0(nl_SystolicArrayLooper_run_run_fsm_inst_xy_o_C_1_tr0[0:0])
    );
  assign reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm = (z_out_32_16[0])
      & ((fsm_output[7:6]!=2'b00));
  assign loopIndicesOut_and_cse = run_wen & reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
  assign xy_o_and_cse = run_wen & ((fsm_output[1:0]!=2'b00));
  assign loopIndicesOut_rsci_idat_47_32_mx0c0 = (z_out_32_16[0]) & (fsm_output[6]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_15_0 <= 16'b0000000000000000;
      loopIndicesOut_rsci_idat_31_16 <= 16'b0000000000000000;
      paramsOut_rsci_idat <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( loopIndicesOut_and_cse ) begin
      loopIndicesOut_rsci_idat_15_0 <= co_c_idx_sva;
      loopIndicesOut_rsci_idat_31_16 <= winx_wx_idx_sva;
      paramsOut_rsci_idat <= paramsIn_crt_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( run_wen & (loopIndicesOut_rsci_idat_47_32_mx0c0 | ((z_out_32_16[0])
        & (fsm_output[7]))) ) begin
      loopIndicesOut_rsci_idat_47_32 <= MUX_v_16_2_2(16'b0000000000000000, z_out_1,
          (loopIndicesOut_not_1_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= reg_loopIndicesOut_rsci_idat_15_loopIndicesOut_nor_itm;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((~((fsm_output[0]) | (fsm_output[2])
          | (fsm_output[11]))) | (~((~ (z_out_32_16[16])) | (fsm_output[0]))));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      xy_o_mul_1_itm <= 32'b00000000000000000000000000000000;
      paramsIn_crt_sva <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( xy_o_and_cse ) begin
      xy_o_mul_1_itm <= conv_u2u_32_32((paramsIn_rsci_idat_mxwt[31:16]) * (paramsIn_rsci_idat_mxwt[15:0]));
      paramsIn_crt_sva <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      xy_o_p_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[11]) | (fsm_output[2])) ) begin
      xy_o_p_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[11]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      OC2_koo_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[10]) | (fsm_output[3])) ) begin
      OC2_koo_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[10]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      co_c_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[9]) | (fsm_output[4])) ) begin
      co_c_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[9]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      winx_wx_idx_sva <= 16'b0000000000000000;
    end
    else if ( run_wen & ((fsm_output[8]) | (fsm_output[5])) ) begin
      winx_wx_idx_sva <= MUX_v_16_2_2(16'b0000000000000000, z_out_1, (fsm_output[8]));
    end
  end
  assign loopIndicesOut_not_1_nl = ~ loopIndicesOut_rsci_idat_47_32_mx0c0;
  assign xy_o_xy_o_or_16_nl = (~((xy_o_mul_1_itm[31]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_17_nl = (~((xy_o_mul_1_itm[30]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_18_nl = (~((xy_o_mul_1_itm[29]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_19_nl = (~((xy_o_mul_1_itm[28]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_20_nl = (~((xy_o_mul_1_itm[27]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_21_nl = (~((xy_o_mul_1_itm[26]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_22_nl = (~((xy_o_mul_1_itm[25]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_23_nl = (~((xy_o_mul_1_itm[24]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_24_nl = (~((xy_o_mul_1_itm[23]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_25_nl = (~((xy_o_mul_1_itm[22]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_26_nl = (~((xy_o_mul_1_itm[21]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_27_nl = (~((xy_o_mul_1_itm[20]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_28_nl = (~((xy_o_mul_1_itm[19]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_29_nl = (~((xy_o_mul_1_itm[18]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_30_nl = (~((xy_o_mul_1_itm[17]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_xy_o_or_31_nl = (~((xy_o_mul_1_itm[16]) | (fsm_output[11]))) | (fsm_output[10:3]!=8'b00000000);
  assign xy_o_or_3_nl = (fsm_output[11:7]!=5'b00000);
  assign xy_o_mux1h_3_nl = MUX1HOT_v_16_6_2((~ (xy_o_mul_1_itm[15:0])), z_out_1,
      (~ (paramsIn_crt_sva[79:64])), (~ (paramsIn_crt_sva[95:80])), (~ (paramsIn_crt_sva[111:96])),
      (~ (paramsIn_crt_sva[127:112])), {(fsm_output[2]) , (xy_o_or_3_nl) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign xy_o_or_4_nl = (~((fsm_output[6:2]!=5'b00000))) | (fsm_output[11:7]!=5'b00000);
  assign xy_o_xy_o_xy_o_nor_16_nl = ~((xy_o_mul_1_itm[31]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_17_nl = ~((xy_o_mul_1_itm[30]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_18_nl = ~((xy_o_mul_1_itm[29]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_19_nl = ~((xy_o_mul_1_itm[28]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_20_nl = ~((xy_o_mul_1_itm[27]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_21_nl = ~((xy_o_mul_1_itm[26]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_22_nl = ~((xy_o_mul_1_itm[25]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_23_nl = ~((xy_o_mul_1_itm[24]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_24_nl = ~((xy_o_mul_1_itm[23]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_25_nl = ~((xy_o_mul_1_itm[22]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_26_nl = ~((xy_o_mul_1_itm[21]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_27_nl = ~((xy_o_mul_1_itm[20]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_28_nl = ~((xy_o_mul_1_itm[19]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_29_nl = ~((xy_o_mul_1_itm[18]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_30_nl = ~((xy_o_mul_1_itm[17]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_xy_o_xy_o_nor_31_nl = ~((xy_o_mul_1_itm[16]) | (fsm_output[10:2]!=9'b000000000));
  assign xy_o_or_5_nl = (fsm_output[6:2]!=5'b00000);
  assign xy_o_mux1h_4_nl = MUX1HOT_v_16_6_2(16'b0000000000000001, (~ (xy_o_mul_1_itm[15:0])),
      (~ (paramsIn_crt_sva[79:64])), (~ (paramsIn_crt_sva[95:80])), (~ (paramsIn_crt_sva[111:96])),
      (~ (paramsIn_crt_sva[127:112])), {(xy_o_or_5_nl) , (fsm_output[11]) , (fsm_output[10])
      , (fsm_output[9]) , (fsm_output[8]) , (fsm_output[7])});
  assign nl_acc_nl = ({1'b1 , (xy_o_xy_o_or_16_nl) , (xy_o_xy_o_or_17_nl) , (xy_o_xy_o_or_18_nl)
      , (xy_o_xy_o_or_19_nl) , (xy_o_xy_o_or_20_nl) , (xy_o_xy_o_or_21_nl) , (xy_o_xy_o_or_22_nl)
      , (xy_o_xy_o_or_23_nl) , (xy_o_xy_o_or_24_nl) , (xy_o_xy_o_or_25_nl) , (xy_o_xy_o_or_26_nl)
      , (xy_o_xy_o_or_27_nl) , (xy_o_xy_o_or_28_nl) , (xy_o_xy_o_or_29_nl) , (xy_o_xy_o_or_30_nl)
      , (xy_o_xy_o_or_31_nl) , (xy_o_mux1h_3_nl) , (xy_o_or_4_nl)}) + conv_u2u_33_34({(xy_o_xy_o_xy_o_nor_16_nl)
      , (xy_o_xy_o_xy_o_nor_17_nl) , (xy_o_xy_o_xy_o_nor_18_nl) , (xy_o_xy_o_xy_o_nor_19_nl)
      , (xy_o_xy_o_xy_o_nor_20_nl) , (xy_o_xy_o_xy_o_nor_21_nl) , (xy_o_xy_o_xy_o_nor_22_nl)
      , (xy_o_xy_o_xy_o_nor_23_nl) , (xy_o_xy_o_xy_o_nor_24_nl) , (xy_o_xy_o_xy_o_nor_25_nl)
      , (xy_o_xy_o_xy_o_nor_26_nl) , (xy_o_xy_o_xy_o_nor_27_nl) , (xy_o_xy_o_xy_o_nor_28_nl)
      , (xy_o_xy_o_xy_o_nor_29_nl) , (xy_o_xy_o_xy_o_nor_30_nl) , (xy_o_xy_o_xy_o_nor_31_nl)
      , (xy_o_mux1h_4_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[33:0];
  assign z_out_32_16 = readslicef_34_17_17((acc_nl));
  assign winy_mux1h_1_nl = MUX1HOT_v_16_5_2(loopIndicesOut_rsci_idat_47_32, xy_o_p_sva,
      OC2_koo_idx_sva, co_c_idx_sva, winx_wx_idx_sva, {(fsm_output[7]) , (fsm_output[11])
      , (fsm_output[10]) , (fsm_output[9]) , (fsm_output[8])});
  assign nl_z_out_1 = (winy_mux1h_1_nl) + 16'b0000000000000001;
  assign z_out_1 = nl_z_out_1[15:0];

  function automatic [15:0] MUX1HOT_v_16_5_2;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [4:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    MUX1HOT_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_6_2;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [5:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    result = result | ( input_3 & {16{sel[3]}});
    result = result | ( input_4 & {16{sel[4]}});
    result = result | ( input_5 & {16{sel[5]}});
    MUX1HOT_v_16_6_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [16:0] readslicef_34_17_17;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 17;
    readslicef_34_17_17 = tmp[16:0];
  end
  endfunction


  function automatic [31:0] conv_u2u_32_32 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_32 = vector;
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer
// ------------------------------------------------------------------


module ParamsDeserializer (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      outputChannel1_rsc_dat, outputChannel1_rsc_vld, outputChannel1_rsc_rdy, outputChannel2_rsc_dat,
      outputChannel2_rsc_vld, outputChannel2_rsc_rdy, outputChannel3_rsc_dat, outputChannel3_rsc_vld,
      outputChannel3_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [143:0] outputChannel1_rsc_dat;
  output outputChannel1_rsc_vld;
  input outputChannel1_rsc_rdy;
  output [143:0] outputChannel2_rsc_dat;
  output outputChannel2_rsc_vld;
  input outputChannel2_rsc_rdy;
  output [143:0] outputChannel3_rsc_dat;
  output outputChannel3_rsc_vld;
  input outputChannel3_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ParamsDeserializer_run ParamsDeserializer_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Serializer_PackedInt_16UL_16UL_ODTYPE_16
// ------------------------------------------------------------------


module Serializer_PackedInt_16UL_16UL_ODTYPE_16 (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      serialOutChannel_rsc_dat, serialOutChannel_rsc_vld, serialOutChannel_rsc_rdy
);
  input clk;
  input arst_n;
  input [255:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [15:0] serialOutChannel_rsc_dat;
  output serialOutChannel_rsc_vld;
  input serialOutChannel_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  Serializer_PackedInt_16UL_16UL_ODTYPE_16_run Serializer_PackedInt_16UL_16UL_ODTYPE_16_run_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld),
      .serialOutChannel_rsc_rdy(serialOutChannel_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayLooper
// ------------------------------------------------------------------


module SystolicArrayLooper (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat,
      paramsOut_rsc_vld, paramsOut_rsc_rdy, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld,
      loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [143:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [47:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  SystolicArrayLooper_run SystolicArrayLooper_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16
// ------------------------------------------------------------------


module SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16 (
  clk, arst_n, input_rsc_dat, input_rsc_vld, input_rsc_rdy, weight_rsc_dat, weight_rsc_vld,
      weight_rsc_rdy, output_rsc_dat, output_rsc_vld, output_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [127:0] input_rsc_dat;
  input input_rsc_vld;
  output input_rsc_rdy;
  input [127:0] weight_rsc_dat;
  input weight_rsc_vld;
  output weight_rsc_rdy;
  output [255:0] output_rsc_dat;
  output output_rsc_vld;
  input output_rsc_rdy;
  input [143:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [255:0] output_rsc_dat_nsystolicArrayCore;
  wire [143:0] paramsIn_rsc_dat_nsystolicArrayCore;
  wire paramsIn_rsc_vld_nsystolicArrayCore;
  wire [47:0] loopIndicesIn_rsc_dat_nsystolicArrayCore;
  wire loopIndicesIn_rsc_vld_nsystolicArrayCore;
  wire [143:0] paramsOut_rsc_dat_nsystolicArrayLooper;
  wire paramsOut_rsc_rdy_nsystolicArrayLooper;
  wire [47:0] loopIndicesOut_rsc_dat_nsystolicArrayLooper;
  wire loopIndicesOut_rsc_rdy_nsystolicArrayLooper;
  wire input_rsc_rdy_nsystolicArrayCore_bud;
  wire weight_rsc_rdy_nsystolicArrayCore_bud;
  wire output_rsc_vld_nsystolicArrayCore_bud;
  wire paramsIn_rsc_rdy_nsystolicArrayCore_bud;
  wire paramsOut_rsc_vld_nsystolicArrayLooper_bud;
  wire loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud;
  wire loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud;
  wire paramsIn_rsc_rdy_nsystolicArrayLooper_bud;
  wire paramsChannel_unc_2;
  wire paramsChannel_idle;
  wire loopIndicesChannel_unc_2;
  wire loopIndicesChannel_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd163),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) paramsChannel_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(paramsOut_rsc_rdy_nsystolicArrayLooper),
      .din_vld(paramsOut_rsc_vld_nsystolicArrayLooper_bud),
      .din(paramsOut_rsc_dat_nsystolicArrayLooper),
      .dout_rdy(paramsIn_rsc_rdy_nsystolicArrayCore_bud),
      .dout_vld(paramsIn_rsc_vld_nsystolicArrayCore),
      .dout(paramsIn_rsc_dat_nsystolicArrayCore),
      .sz(paramsChannel_unc_2),
      .sz_req(1'b0),
      .is_idle(paramsChannel_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd164),
  .width(32'sd48),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) loopIndicesChannel_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(loopIndicesOut_rsc_rdy_nsystolicArrayLooper),
      .din_vld(loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud),
      .din(loopIndicesOut_rsc_dat_nsystolicArrayLooper),
      .dout_rdy(loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud),
      .dout_vld(loopIndicesIn_rsc_vld_nsystolicArrayCore),
      .dout(loopIndicesIn_rsc_dat_nsystolicArrayCore),
      .sz(loopIndicesChannel_unc_2),
      .sz_req(1'b0),
      .is_idle(loopIndicesChannel_idle)
    );
  SystolicArrayCore_IDTYPE_WDTYPE_ODTYPE_16_16 systolicArrayCore (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_vld(input_rsc_vld),
      .input_rsc_rdy(input_rsc_rdy_nsystolicArrayCore_bud),
      .weight_rsc_dat(weight_rsc_dat),
      .weight_rsc_vld(weight_rsc_vld),
      .weight_rsc_rdy(weight_rsc_rdy_nsystolicArrayCore_bud),
      .output_rsc_dat(output_rsc_dat_nsystolicArrayCore),
      .output_rsc_vld(output_rsc_vld_nsystolicArrayCore_bud),
      .output_rsc_rdy(output_rsc_rdy),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nsystolicArrayCore),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nsystolicArrayCore),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArrayCore_bud),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat_nsystolicArrayCore),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld_nsystolicArrayCore),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy_nsystolicArrayCore_bud)
    );
  SystolicArrayLooper systolicArrayLooper_1 (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArrayLooper_bud),
      .paramsOut_rsc_dat(paramsOut_rsc_dat_nsystolicArrayLooper),
      .paramsOut_rsc_vld(paramsOut_rsc_vld_nsystolicArrayLooper_bud),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy_nsystolicArrayLooper),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat_nsystolicArrayLooper),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld_nsystolicArrayLooper_bud),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy_nsystolicArrayLooper)
    );
  assign input_rsc_rdy = input_rsc_rdy_nsystolicArrayCore_bud;
  assign weight_rsc_rdy = weight_rsc_rdy_nsystolicArrayCore_bud;
  assign output_rsc_vld = output_rsc_vld_nsystolicArrayCore_bud;
  assign output_rsc_dat = output_rsc_dat_nsystolicArrayCore;
  assign paramsIn_rsc_rdy = paramsIn_rsc_rdy_nsystolicArrayLooper_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Conv
// ------------------------------------------------------------------


module Conv (
  clk, arst_n, input_serial_rsc_dat, input_serial_rsc_vld, input_serial_rsc_rdy,
      weight_serial_rsc_dat, weight_serial_rsc_vld, weight_serial_rsc_rdy, output_serial_rsc_dat,
      output_serial_rsc_vld, output_serial_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy
);
  input clk;
  input arst_n;
  input [15:0] input_serial_rsc_dat;
  input input_serial_rsc_vld;
  output input_serial_rsc_rdy;
  input [15:0] weight_serial_rsc_dat;
  input weight_serial_rsc_vld;
  output weight_serial_rsc_rdy;
  output [15:0] output_serial_rsc_dat;
  output output_serial_rsc_vld;
  input output_serial_rsc_rdy;
  input [15:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;


  // Interconnect Declarations
  wire [143:0] outputChannel1_rsc_dat_nparamsDeserializer;
  wire outputChannel1_rsc_rdy_nparamsDeserializer;
  wire [143:0] outputChannel2_rsc_dat_nparamsDeserializer;
  wire outputChannel2_rsc_rdy_nparamsDeserializer;
  wire [143:0] outputChannel3_rsc_dat_nparamsDeserializer;
  wire outputChannel3_rsc_rdy_nparamsDeserializer;
  wire [255:0] inputChannel_rsc_dat_noutputSerializer;
  wire inputChannel_rsc_vld_noutputSerializer;
  wire [15:0] serialOutChannel_rsc_dat_noutputSerializer;
  wire [127:0] inputs_out_rsc_dat_ninputDoubleBuffer;
  wire inputs_out_rsc_rdy_ninputDoubleBuffer;
  wire [143:0] paramsIn_rsc_dat_ninputDoubleBuffer;
  wire paramsIn_rsc_vld_ninputDoubleBuffer;
  wire [127:0] weights_out_rsc_dat_nweightDoubleBuffer;
  wire weights_out_rsc_rdy_nweightDoubleBuffer;
  wire [143:0] paramsIn_rsc_dat_nweightDoubleBuffer;
  wire paramsIn_rsc_vld_nweightDoubleBuffer;
  wire [127:0] input_rsc_dat_nsystolicArray;
  wire input_rsc_vld_nsystolicArray;
  wire [127:0] weight_rsc_dat_nsystolicArray;
  wire weight_rsc_vld_nsystolicArray;
  wire [255:0] output_rsc_dat_nsystolicArray;
  wire output_rsc_rdy_nsystolicArray;
  wire [143:0] paramsIn_rsc_dat_nsystolicArray;
  wire paramsIn_rsc_vld_nsystolicArray;
  wire inputChannel_rsc_rdy_nparamsDeserializer_bud;
  wire outputChannel1_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_ninputDoubleBuffer_bud;
  wire outputChannel2_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_nweightDoubleBuffer_bud;
  wire outputChannel3_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_nsystolicArray_bud;
  wire inputChannel_rsc_rdy_noutputSerializer_bud;
  wire output_rsc_vld_nsystolicArray_bud;
  wire serialOutChannel_rsc_vld_noutputSerializer_bud;
  wire inputs_in_rsc_rdy_ninputDoubleBuffer_bud;
  wire inputs_out_rsc_vld_ninputDoubleBuffer_bud;
  wire input_rsc_rdy_nsystolicArray_bud;
  wire weights_in_rsc_rdy_nweightDoubleBuffer_bud;
  wire weights_out_rsc_vld_nweightDoubleBuffer_bud;
  wire weight_rsc_rdy_nsystolicArray_bud;
  wire inputDoubleBufferParams_unc_2;
  wire inputDoubleBufferParams_idle;
  wire weightDoubleBufferParams_unc_2;
  wire weightDoubleBufferParams_idle;
  wire systolicArrayParams_unc_2;
  wire systolicArrayParams_idle;
  wire output_unc_2;
  wire output_idle;
  wire input_out_unc_2;
  wire input_out_idle;
  wire weight_out_unc_2;
  wire weight_out_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd169),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) inputDoubleBufferParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel1_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel1_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel1_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_ninputDoubleBuffer_bud),
      .dout_vld(paramsIn_rsc_vld_ninputDoubleBuffer),
      .dout(paramsIn_rsc_dat_ninputDoubleBuffer),
      .sz(inputDoubleBufferParams_unc_2),
      .sz_req(1'b0),
      .is_idle(inputDoubleBufferParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd170),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weightDoubleBufferParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel2_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel2_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel2_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_nweightDoubleBuffer_bud),
      .dout_vld(paramsIn_rsc_vld_nweightDoubleBuffer),
      .dout(paramsIn_rsc_dat_nweightDoubleBuffer),
      .sz(weightDoubleBufferParams_unc_2),
      .sz_req(1'b0),
      .is_idle(weightDoubleBufferParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd174),
  .width(32'sd144),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) systolicArrayParams_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(outputChannel3_rsc_rdy_nparamsDeserializer),
      .din_vld(outputChannel3_rsc_vld_nparamsDeserializer_bud),
      .din(outputChannel3_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_nsystolicArray_bud),
      .dout_vld(paramsIn_rsc_vld_nsystolicArray),
      .dout(paramsIn_rsc_dat_nsystolicArray),
      .sz(systolicArrayParams_unc_2),
      .sz_req(1'b0),
      .is_idle(systolicArrayParams_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd173),
  .width(32'sd256),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) output_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(output_rsc_rdy_nsystolicArray),
      .din_vld(output_rsc_vld_nsystolicArray_bud),
      .din(output_rsc_dat_nsystolicArray),
      .dout_rdy(inputChannel_rsc_rdy_noutputSerializer_bud),
      .dout_vld(inputChannel_rsc_vld_noutputSerializer),
      .dout(inputChannel_rsc_dat_noutputSerializer),
      .sz(output_unc_2),
      .sz_req(1'b0),
      .is_idle(output_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd171),
  .width(32'sd128),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) input_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(inputs_out_rsc_rdy_ninputDoubleBuffer),
      .din_vld(inputs_out_rsc_vld_ninputDoubleBuffer_bud),
      .din(inputs_out_rsc_dat_ninputDoubleBuffer),
      .dout_rdy(input_rsc_rdy_nsystolicArray_bud),
      .dout_vld(input_rsc_vld_nsystolicArray),
      .dout(input_rsc_dat_nsystolicArray),
      .sz(input_out_unc_2),
      .sz_req(1'b0),
      .is_idle(input_out_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd172),
  .width(32'sd128),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) weight_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(weights_out_rsc_rdy_nweightDoubleBuffer),
      .din_vld(weights_out_rsc_vld_nweightDoubleBuffer_bud),
      .din(weights_out_rsc_dat_nweightDoubleBuffer),
      .dout_rdy(weight_rsc_rdy_nsystolicArray_bud),
      .dout_vld(weight_rsc_vld_nsystolicArray),
      .dout(weight_rsc_dat_nsystolicArray),
      .sz(weight_out_unc_2),
      .sz_req(1'b0),
      .is_idle(weight_out_idle)
    );
  ParamsDeserializer paramsDeserializer_1 (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(paramsIn_rsc_dat),
      .inputChannel_rsc_vld(paramsIn_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy_nparamsDeserializer_bud),
      .outputChannel1_rsc_dat(outputChannel1_rsc_dat_nparamsDeserializer),
      .outputChannel1_rsc_vld(outputChannel1_rsc_vld_nparamsDeserializer_bud),
      .outputChannel1_rsc_rdy(outputChannel1_rsc_rdy_nparamsDeserializer),
      .outputChannel2_rsc_dat(outputChannel2_rsc_dat_nparamsDeserializer),
      .outputChannel2_rsc_vld(outputChannel2_rsc_vld_nparamsDeserializer_bud),
      .outputChannel2_rsc_rdy(outputChannel2_rsc_rdy_nparamsDeserializer),
      .outputChannel3_rsc_dat(outputChannel3_rsc_dat_nparamsDeserializer),
      .outputChannel3_rsc_vld(outputChannel3_rsc_vld_nparamsDeserializer_bud),
      .outputChannel3_rsc_rdy(outputChannel3_rsc_rdy_nparamsDeserializer)
    );
  Serializer_PackedInt_16UL_16UL_ODTYPE_16 outputSerializer (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat_noutputSerializer),
      .inputChannel_rsc_vld(inputChannel_rsc_vld_noutputSerializer),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy_noutputSerializer_bud),
      .serialOutChannel_rsc_dat(serialOutChannel_rsc_dat_noutputSerializer),
      .serialOutChannel_rsc_vld(serialOutChannel_rsc_vld_noutputSerializer_bud),
      .serialOutChannel_rsc_rdy(output_serial_rsc_rdy)
    );
  InputDoubleBuffer_512_16_16 inputDoubleBuffer (
      .clk(clk),
      .arst_n(arst_n),
      .inputs_in_rsc_dat(input_serial_rsc_dat),
      .inputs_in_rsc_vld(input_serial_rsc_vld),
      .inputs_in_rsc_rdy(inputs_in_rsc_rdy_ninputDoubleBuffer_bud),
      .inputs_out_rsc_dat(inputs_out_rsc_dat_ninputDoubleBuffer),
      .inputs_out_rsc_vld(inputs_out_rsc_vld_ninputDoubleBuffer_bud),
      .inputs_out_rsc_rdy(inputs_out_rsc_rdy_ninputDoubleBuffer),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_ninputDoubleBuffer),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_ninputDoubleBuffer),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_ninputDoubleBuffer_bud)
    );
  WeightDoubleBuffer_384_16_16 weightDoubleBuffer (
      .clk(clk),
      .arst_n(arst_n),
      .weights_in_rsc_dat(weight_serial_rsc_dat),
      .weights_in_rsc_vld(weight_serial_rsc_vld),
      .weights_in_rsc_rdy(weights_in_rsc_rdy_nweightDoubleBuffer_bud),
      .weights_out_rsc_dat(weights_out_rsc_dat_nweightDoubleBuffer),
      .weights_out_rsc_vld(weights_out_rsc_vld_nweightDoubleBuffer_bud),
      .weights_out_rsc_rdy(weights_out_rsc_rdy_nweightDoubleBuffer),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nweightDoubleBuffer),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nweightDoubleBuffer),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nweightDoubleBuffer_bud)
    );
  SystolicArrayWrapper_IDTYPE_WDTYPE_ODTYPE_16_16 systolicArray (
      .clk(clk),
      .arst_n(arst_n),
      .input_rsc_dat(input_rsc_dat_nsystolicArray),
      .input_rsc_vld(input_rsc_vld_nsystolicArray),
      .input_rsc_rdy(input_rsc_rdy_nsystolicArray_bud),
      .weight_rsc_dat(weight_rsc_dat_nsystolicArray),
      .weight_rsc_vld(weight_rsc_vld_nsystolicArray),
      .weight_rsc_rdy(weight_rsc_rdy_nsystolicArray_bud),
      .output_rsc_dat(output_rsc_dat_nsystolicArray),
      .output_rsc_vld(output_rsc_vld_nsystolicArray_bud),
      .output_rsc_rdy(output_rsc_rdy_nsystolicArray),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nsystolicArray),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nsystolicArray),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nsystolicArray_bud)
    );
  assign paramsIn_rsc_rdy = inputChannel_rsc_rdy_nparamsDeserializer_bud;
  assign output_serial_rsc_vld = serialOutChannel_rsc_vld_noutputSerializer_bud;
  assign output_serial_rsc_dat = serialOutChannel_rsc_dat_noutputSerializer;
  assign input_serial_rsc_rdy = inputs_in_rsc_rdy_ninputDoubleBuffer_bud;
  assign weight_serial_rsc_rdy = weights_in_rsc_rdy_nweightDoubleBuffer_bud;
endmodule



