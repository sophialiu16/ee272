module accum_double_buffer
#(
  parameter DATA_WIDTH = 64,
  parameter BANK_ADDR_WIDTH = 32 // There are two banks
)(
  input clk,
  input rst_n,
  input switch_banks,
  input ren_out,
  input ren_sys_arr,
  input [BANK_ADDR_WIDTH - 1 : 0] radr_out,
  input [BANK_ADDR_WIDTH - 1 : 0] radr_sys_arr,
  output [DATA_WIDTH - 1 : 0] rdata_out,
  output [DATA_WIDTH - 1 : 0] rdata_sys_arr,
  input wen,
  input [BANK_ADDR_WIDTH - 1 : 0] wadr,
  input [DATA_WIDTH - 1 : 0] wdata
);

  // Internally keeps track of which bank is being used for reading and which
  // for writing using some state
  logic systolic_bank;

  logic wen0, ren0, wen1, ren1;

  ram_sync_1r1w #(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(BANK_ADDR_WIDTH),
    .DEPTH(128) //todo
  )
  ram0 (
    .clk(clk),
    .wen(wen0),
    .wadr(wadr),
    .wdata(wdata),
    .ren(ren0),
    .radr(radr),
    .rdata(rdata0)
  );

   ram_sync_1r1w #(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(BANK_ADDR_WIDTH),
    .DEPTH(128) //todo
  )
  ram1 (
    .clk(clk),
    .wen(wen1),
    .wadr(wadr),
    .wdata(wdata),
    .ren(ren1),
    .radr(radr),
    .rdata(rdata1)
  );

  always_ff @(posedge clk) begin
    if (~rst_n) begin
      systolic_bank <= 0;
      rdata_sys_arr <= 0;
    end
    else if begin

      if (ren_sys_arr) begin
        if (systolic_bank) begin
          rdata_sys_arr <= rdata1;
          ren1 <= systolic_bank;
        end else begin
          rdata_sys_arr <= rdata0;
          ren0 <= ~systolic_bank;
        end
     end else begin
       rdata_sys_arr <= 0;
     end
      
      if (ren_out) begin 
        if (systolic_bank) begin
          rdata_out <= rdata0;
          ren0 <= systolic_bank;
        end else begin
          rdata_out <= rdata1;
          ren1 <= ~systolic_bank;
        end
      end

      if (wen) begin
        wen0 <= ~systolic_bank;
        wen1 <= systolic_bank;
      end

      if (switch_banks) begin
         systolic_bank <= ~systolic_bank;
      end
    end // end reset
  end // end always_ff

endmodule

