module double_buffer
#(
  parameter DATA_WIDTH = 64,
  parameter BANK_ADDR_WIDTH = 32 // There are two banks
)(
  input clk,
  input rst_n,
  input switch_banks,
  input ren,
  input [BANK_ADDR_WIDTH - 1 : 0] radr,
  output [DATA_WIDTH - 1 : 0] rdata,
  input wen,
  input [BANK_ADDR_WIDTH - 1 : 0] wadr,
  input [DATA_WIDTH - 1 : 0] wdata
);

  // Internally keeps track of which bank is being used for reading and which
  // for writing using some state
  logic read_bank;
  logic [DATA_WIDTH - 1 : 0] buffers [1 : 0][BANK_ADDR_WIDTH - 1 : 0]
  
  logic wen0, ren0, wen1, ren1;
  
  ram_sync_1r1w #(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(BANK_ADDR_WIDTH),
    .DEPTH(128) //todo
  ) 
  ram0 (
    .clk(clk),
    .wen(wen0),
    .wadr(wadr),
    .wdata(wdata),
    .ren(ren0),
    .radr(radr),
    .rdata(rdata0)
  );
  
   ram_sync_1r1w #(
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(BANK_ADDR_WIDTH),
    .DEPTH(128) //todo
  ) 
  ram1 (
    .clk(clk),
    .wen(wen1),
    .wadr(wadr),
    .wdata(wdata),
    .ren(ren1),
    .radr(radr),
    .rdata(rdata1)
  );
  
  always_ff @(posedge clk) begin
    if (~rst_n) begin
      read_bank <= 0;
    end
    else if begin

      if (ren) begin
        ren0 <= ~read_bank;
        ren1 <= read_bank;
        if (read_bank) begin
          rdata <= rdata1;
        end else begin 
          rdata <= rdata0;
        end
     end

      if (wen) begin
        if (~read_bank) begin
          wen0 <= 0;
          wen1 <= 1;
        end
        buffers[~read_bank][wadr] <= wdata;
      end

      if (switch_banks) begin
        read_bank <= ~read_bank;
      end
    end // end reset
  end // end always_ff

endmodule
~

