**************************************************
* OpenRAM generated memory.
* Words: 512
* Data bits: 128
* Banks: 1
* Column mux: 2:1
**************************************************
* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
*
.subckt dff D Q clk vdd gnd
*
MM21 Q a_66_6# gnd gnd NMOS_VTG L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd NMOS_VTG L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd PMOS_VTG L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd PMOS_VTG L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd PMOS_VTG L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd PMOS_VTG L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.SUBCKT row_addr_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 8 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r1_c0 din_1 dout_1 clk vdd gnd dff
Xdff_r2_c0 din_2 dout_2 clk vdd gnd dff
Xdff_r3_c0 din_3 dout_3 clk vdd gnd dff
Xdff_r4_c0 din_4 dout_4 clk vdd gnd dff
Xdff_r5_c0 din_5 dout_5 clk vdd gnd dff
Xdff_r6_c0 din_6 dout_6 clk vdd gnd dff
Xdff_r7_c0 din_7 dout_7 clk vdd gnd dff
.ENDS row_addr_dff

.SUBCKT col_addr_dff din_0 dout_0 clk vdd gnd
* INPUT : din_0 
* OUTPUT: dout_0 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
.ENDS col_addr_dff

.SUBCKT data_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38 dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46 dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54 dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62 dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70 dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78 dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86 dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94 dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102 dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109 dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116 dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123 dout_124 dout_125 dout_126 dout_127 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 128
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
Xdff_r0_c3 din_3 dout_3 clk vdd gnd dff
Xdff_r0_c4 din_4 dout_4 clk vdd gnd dff
Xdff_r0_c5 din_5 dout_5 clk vdd gnd dff
Xdff_r0_c6 din_6 dout_6 clk vdd gnd dff
Xdff_r0_c7 din_7 dout_7 clk vdd gnd dff
Xdff_r0_c8 din_8 dout_8 clk vdd gnd dff
Xdff_r0_c9 din_9 dout_9 clk vdd gnd dff
Xdff_r0_c10 din_10 dout_10 clk vdd gnd dff
Xdff_r0_c11 din_11 dout_11 clk vdd gnd dff
Xdff_r0_c12 din_12 dout_12 clk vdd gnd dff
Xdff_r0_c13 din_13 dout_13 clk vdd gnd dff
Xdff_r0_c14 din_14 dout_14 clk vdd gnd dff
Xdff_r0_c15 din_15 dout_15 clk vdd gnd dff
Xdff_r0_c16 din_16 dout_16 clk vdd gnd dff
Xdff_r0_c17 din_17 dout_17 clk vdd gnd dff
Xdff_r0_c18 din_18 dout_18 clk vdd gnd dff
Xdff_r0_c19 din_19 dout_19 clk vdd gnd dff
Xdff_r0_c20 din_20 dout_20 clk vdd gnd dff
Xdff_r0_c21 din_21 dout_21 clk vdd gnd dff
Xdff_r0_c22 din_22 dout_22 clk vdd gnd dff
Xdff_r0_c23 din_23 dout_23 clk vdd gnd dff
Xdff_r0_c24 din_24 dout_24 clk vdd gnd dff
Xdff_r0_c25 din_25 dout_25 clk vdd gnd dff
Xdff_r0_c26 din_26 dout_26 clk vdd gnd dff
Xdff_r0_c27 din_27 dout_27 clk vdd gnd dff
Xdff_r0_c28 din_28 dout_28 clk vdd gnd dff
Xdff_r0_c29 din_29 dout_29 clk vdd gnd dff
Xdff_r0_c30 din_30 dout_30 clk vdd gnd dff
Xdff_r0_c31 din_31 dout_31 clk vdd gnd dff
Xdff_r0_c32 din_32 dout_32 clk vdd gnd dff
Xdff_r0_c33 din_33 dout_33 clk vdd gnd dff
Xdff_r0_c34 din_34 dout_34 clk vdd gnd dff
Xdff_r0_c35 din_35 dout_35 clk vdd gnd dff
Xdff_r0_c36 din_36 dout_36 clk vdd gnd dff
Xdff_r0_c37 din_37 dout_37 clk vdd gnd dff
Xdff_r0_c38 din_38 dout_38 clk vdd gnd dff
Xdff_r0_c39 din_39 dout_39 clk vdd gnd dff
Xdff_r0_c40 din_40 dout_40 clk vdd gnd dff
Xdff_r0_c41 din_41 dout_41 clk vdd gnd dff
Xdff_r0_c42 din_42 dout_42 clk vdd gnd dff
Xdff_r0_c43 din_43 dout_43 clk vdd gnd dff
Xdff_r0_c44 din_44 dout_44 clk vdd gnd dff
Xdff_r0_c45 din_45 dout_45 clk vdd gnd dff
Xdff_r0_c46 din_46 dout_46 clk vdd gnd dff
Xdff_r0_c47 din_47 dout_47 clk vdd gnd dff
Xdff_r0_c48 din_48 dout_48 clk vdd gnd dff
Xdff_r0_c49 din_49 dout_49 clk vdd gnd dff
Xdff_r0_c50 din_50 dout_50 clk vdd gnd dff
Xdff_r0_c51 din_51 dout_51 clk vdd gnd dff
Xdff_r0_c52 din_52 dout_52 clk vdd gnd dff
Xdff_r0_c53 din_53 dout_53 clk vdd gnd dff
Xdff_r0_c54 din_54 dout_54 clk vdd gnd dff
Xdff_r0_c55 din_55 dout_55 clk vdd gnd dff
Xdff_r0_c56 din_56 dout_56 clk vdd gnd dff
Xdff_r0_c57 din_57 dout_57 clk vdd gnd dff
Xdff_r0_c58 din_58 dout_58 clk vdd gnd dff
Xdff_r0_c59 din_59 dout_59 clk vdd gnd dff
Xdff_r0_c60 din_60 dout_60 clk vdd gnd dff
Xdff_r0_c61 din_61 dout_61 clk vdd gnd dff
Xdff_r0_c62 din_62 dout_62 clk vdd gnd dff
Xdff_r0_c63 din_63 dout_63 clk vdd gnd dff
Xdff_r0_c64 din_64 dout_64 clk vdd gnd dff
Xdff_r0_c65 din_65 dout_65 clk vdd gnd dff
Xdff_r0_c66 din_66 dout_66 clk vdd gnd dff
Xdff_r0_c67 din_67 dout_67 clk vdd gnd dff
Xdff_r0_c68 din_68 dout_68 clk vdd gnd dff
Xdff_r0_c69 din_69 dout_69 clk vdd gnd dff
Xdff_r0_c70 din_70 dout_70 clk vdd gnd dff
Xdff_r0_c71 din_71 dout_71 clk vdd gnd dff
Xdff_r0_c72 din_72 dout_72 clk vdd gnd dff
Xdff_r0_c73 din_73 dout_73 clk vdd gnd dff
Xdff_r0_c74 din_74 dout_74 clk vdd gnd dff
Xdff_r0_c75 din_75 dout_75 clk vdd gnd dff
Xdff_r0_c76 din_76 dout_76 clk vdd gnd dff
Xdff_r0_c77 din_77 dout_77 clk vdd gnd dff
Xdff_r0_c78 din_78 dout_78 clk vdd gnd dff
Xdff_r0_c79 din_79 dout_79 clk vdd gnd dff
Xdff_r0_c80 din_80 dout_80 clk vdd gnd dff
Xdff_r0_c81 din_81 dout_81 clk vdd gnd dff
Xdff_r0_c82 din_82 dout_82 clk vdd gnd dff
Xdff_r0_c83 din_83 dout_83 clk vdd gnd dff
Xdff_r0_c84 din_84 dout_84 clk vdd gnd dff
Xdff_r0_c85 din_85 dout_85 clk vdd gnd dff
Xdff_r0_c86 din_86 dout_86 clk vdd gnd dff
Xdff_r0_c87 din_87 dout_87 clk vdd gnd dff
Xdff_r0_c88 din_88 dout_88 clk vdd gnd dff
Xdff_r0_c89 din_89 dout_89 clk vdd gnd dff
Xdff_r0_c90 din_90 dout_90 clk vdd gnd dff
Xdff_r0_c91 din_91 dout_91 clk vdd gnd dff
Xdff_r0_c92 din_92 dout_92 clk vdd gnd dff
Xdff_r0_c93 din_93 dout_93 clk vdd gnd dff
Xdff_r0_c94 din_94 dout_94 clk vdd gnd dff
Xdff_r0_c95 din_95 dout_95 clk vdd gnd dff
Xdff_r0_c96 din_96 dout_96 clk vdd gnd dff
Xdff_r0_c97 din_97 dout_97 clk vdd gnd dff
Xdff_r0_c98 din_98 dout_98 clk vdd gnd dff
Xdff_r0_c99 din_99 dout_99 clk vdd gnd dff
Xdff_r0_c100 din_100 dout_100 clk vdd gnd dff
Xdff_r0_c101 din_101 dout_101 clk vdd gnd dff
Xdff_r0_c102 din_102 dout_102 clk vdd gnd dff
Xdff_r0_c103 din_103 dout_103 clk vdd gnd dff
Xdff_r0_c104 din_104 dout_104 clk vdd gnd dff
Xdff_r0_c105 din_105 dout_105 clk vdd gnd dff
Xdff_r0_c106 din_106 dout_106 clk vdd gnd dff
Xdff_r0_c107 din_107 dout_107 clk vdd gnd dff
Xdff_r0_c108 din_108 dout_108 clk vdd gnd dff
Xdff_r0_c109 din_109 dout_109 clk vdd gnd dff
Xdff_r0_c110 din_110 dout_110 clk vdd gnd dff
Xdff_r0_c111 din_111 dout_111 clk vdd gnd dff
Xdff_r0_c112 din_112 dout_112 clk vdd gnd dff
Xdff_r0_c113 din_113 dout_113 clk vdd gnd dff
Xdff_r0_c114 din_114 dout_114 clk vdd gnd dff
Xdff_r0_c115 din_115 dout_115 clk vdd gnd dff
Xdff_r0_c116 din_116 dout_116 clk vdd gnd dff
Xdff_r0_c117 din_117 dout_117 clk vdd gnd dff
Xdff_r0_c118 din_118 dout_118 clk vdd gnd dff
Xdff_r0_c119 din_119 dout_119 clk vdd gnd dff
Xdff_r0_c120 din_120 dout_120 clk vdd gnd dff
Xdff_r0_c121 din_121 dout_121 clk vdd gnd dff
Xdff_r0_c122 din_122 dout_122 clk vdd gnd dff
Xdff_r0_c123 din_123 dout_123 clk vdd gnd dff
Xdff_r0_c124 din_124 dout_124 clk vdd gnd dff
Xdff_r0_c125 din_125 dout_125 clk vdd gnd dff
Xdff_r0_c126 din_126 dout_126 clk vdd gnd dff
Xdff_r0_c127 din_127 dout_127 clk vdd gnd dff
.ENDS data_dff

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT precharge_1 bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos1 bl en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos2 br en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS precharge_1

.SUBCKT precharge_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 bl_256 br_256 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* INPUT : en_bar 
* POWER : vdd 
* cols: 257 size: 1 bl: bl br: br
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_1
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_1
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_1
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_1
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_1
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_1
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_1
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_1
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_1
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_1
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_1
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_1
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_1
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_1
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_1
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_1
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_1
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_1
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_1
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_1
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_1
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_1
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_1
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_1
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_1
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_1
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_1
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_1
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_1
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_1
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_1
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_1
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_1
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_1
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_1
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_1
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_1
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_1
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_1
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_1
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_1
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_1
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_1
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_1
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_1
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_1
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_1
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_1
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_1
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_1
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_1
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_1
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_1
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_1
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_1
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_1
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_1
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_1
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_1
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_1
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_1
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_1
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_1
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_1
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_1
Xpre_column_65 bl_65 br_65 en_bar vdd precharge_1
Xpre_column_66 bl_66 br_66 en_bar vdd precharge_1
Xpre_column_67 bl_67 br_67 en_bar vdd precharge_1
Xpre_column_68 bl_68 br_68 en_bar vdd precharge_1
Xpre_column_69 bl_69 br_69 en_bar vdd precharge_1
Xpre_column_70 bl_70 br_70 en_bar vdd precharge_1
Xpre_column_71 bl_71 br_71 en_bar vdd precharge_1
Xpre_column_72 bl_72 br_72 en_bar vdd precharge_1
Xpre_column_73 bl_73 br_73 en_bar vdd precharge_1
Xpre_column_74 bl_74 br_74 en_bar vdd precharge_1
Xpre_column_75 bl_75 br_75 en_bar vdd precharge_1
Xpre_column_76 bl_76 br_76 en_bar vdd precharge_1
Xpre_column_77 bl_77 br_77 en_bar vdd precharge_1
Xpre_column_78 bl_78 br_78 en_bar vdd precharge_1
Xpre_column_79 bl_79 br_79 en_bar vdd precharge_1
Xpre_column_80 bl_80 br_80 en_bar vdd precharge_1
Xpre_column_81 bl_81 br_81 en_bar vdd precharge_1
Xpre_column_82 bl_82 br_82 en_bar vdd precharge_1
Xpre_column_83 bl_83 br_83 en_bar vdd precharge_1
Xpre_column_84 bl_84 br_84 en_bar vdd precharge_1
Xpre_column_85 bl_85 br_85 en_bar vdd precharge_1
Xpre_column_86 bl_86 br_86 en_bar vdd precharge_1
Xpre_column_87 bl_87 br_87 en_bar vdd precharge_1
Xpre_column_88 bl_88 br_88 en_bar vdd precharge_1
Xpre_column_89 bl_89 br_89 en_bar vdd precharge_1
Xpre_column_90 bl_90 br_90 en_bar vdd precharge_1
Xpre_column_91 bl_91 br_91 en_bar vdd precharge_1
Xpre_column_92 bl_92 br_92 en_bar vdd precharge_1
Xpre_column_93 bl_93 br_93 en_bar vdd precharge_1
Xpre_column_94 bl_94 br_94 en_bar vdd precharge_1
Xpre_column_95 bl_95 br_95 en_bar vdd precharge_1
Xpre_column_96 bl_96 br_96 en_bar vdd precharge_1
Xpre_column_97 bl_97 br_97 en_bar vdd precharge_1
Xpre_column_98 bl_98 br_98 en_bar vdd precharge_1
Xpre_column_99 bl_99 br_99 en_bar vdd precharge_1
Xpre_column_100 bl_100 br_100 en_bar vdd precharge_1
Xpre_column_101 bl_101 br_101 en_bar vdd precharge_1
Xpre_column_102 bl_102 br_102 en_bar vdd precharge_1
Xpre_column_103 bl_103 br_103 en_bar vdd precharge_1
Xpre_column_104 bl_104 br_104 en_bar vdd precharge_1
Xpre_column_105 bl_105 br_105 en_bar vdd precharge_1
Xpre_column_106 bl_106 br_106 en_bar vdd precharge_1
Xpre_column_107 bl_107 br_107 en_bar vdd precharge_1
Xpre_column_108 bl_108 br_108 en_bar vdd precharge_1
Xpre_column_109 bl_109 br_109 en_bar vdd precharge_1
Xpre_column_110 bl_110 br_110 en_bar vdd precharge_1
Xpre_column_111 bl_111 br_111 en_bar vdd precharge_1
Xpre_column_112 bl_112 br_112 en_bar vdd precharge_1
Xpre_column_113 bl_113 br_113 en_bar vdd precharge_1
Xpre_column_114 bl_114 br_114 en_bar vdd precharge_1
Xpre_column_115 bl_115 br_115 en_bar vdd precharge_1
Xpre_column_116 bl_116 br_116 en_bar vdd precharge_1
Xpre_column_117 bl_117 br_117 en_bar vdd precharge_1
Xpre_column_118 bl_118 br_118 en_bar vdd precharge_1
Xpre_column_119 bl_119 br_119 en_bar vdd precharge_1
Xpre_column_120 bl_120 br_120 en_bar vdd precharge_1
Xpre_column_121 bl_121 br_121 en_bar vdd precharge_1
Xpre_column_122 bl_122 br_122 en_bar vdd precharge_1
Xpre_column_123 bl_123 br_123 en_bar vdd precharge_1
Xpre_column_124 bl_124 br_124 en_bar vdd precharge_1
Xpre_column_125 bl_125 br_125 en_bar vdd precharge_1
Xpre_column_126 bl_126 br_126 en_bar vdd precharge_1
Xpre_column_127 bl_127 br_127 en_bar vdd precharge_1
Xpre_column_128 bl_128 br_128 en_bar vdd precharge_1
Xpre_column_129 bl_129 br_129 en_bar vdd precharge_1
Xpre_column_130 bl_130 br_130 en_bar vdd precharge_1
Xpre_column_131 bl_131 br_131 en_bar vdd precharge_1
Xpre_column_132 bl_132 br_132 en_bar vdd precharge_1
Xpre_column_133 bl_133 br_133 en_bar vdd precharge_1
Xpre_column_134 bl_134 br_134 en_bar vdd precharge_1
Xpre_column_135 bl_135 br_135 en_bar vdd precharge_1
Xpre_column_136 bl_136 br_136 en_bar vdd precharge_1
Xpre_column_137 bl_137 br_137 en_bar vdd precharge_1
Xpre_column_138 bl_138 br_138 en_bar vdd precharge_1
Xpre_column_139 bl_139 br_139 en_bar vdd precharge_1
Xpre_column_140 bl_140 br_140 en_bar vdd precharge_1
Xpre_column_141 bl_141 br_141 en_bar vdd precharge_1
Xpre_column_142 bl_142 br_142 en_bar vdd precharge_1
Xpre_column_143 bl_143 br_143 en_bar vdd precharge_1
Xpre_column_144 bl_144 br_144 en_bar vdd precharge_1
Xpre_column_145 bl_145 br_145 en_bar vdd precharge_1
Xpre_column_146 bl_146 br_146 en_bar vdd precharge_1
Xpre_column_147 bl_147 br_147 en_bar vdd precharge_1
Xpre_column_148 bl_148 br_148 en_bar vdd precharge_1
Xpre_column_149 bl_149 br_149 en_bar vdd precharge_1
Xpre_column_150 bl_150 br_150 en_bar vdd precharge_1
Xpre_column_151 bl_151 br_151 en_bar vdd precharge_1
Xpre_column_152 bl_152 br_152 en_bar vdd precharge_1
Xpre_column_153 bl_153 br_153 en_bar vdd precharge_1
Xpre_column_154 bl_154 br_154 en_bar vdd precharge_1
Xpre_column_155 bl_155 br_155 en_bar vdd precharge_1
Xpre_column_156 bl_156 br_156 en_bar vdd precharge_1
Xpre_column_157 bl_157 br_157 en_bar vdd precharge_1
Xpre_column_158 bl_158 br_158 en_bar vdd precharge_1
Xpre_column_159 bl_159 br_159 en_bar vdd precharge_1
Xpre_column_160 bl_160 br_160 en_bar vdd precharge_1
Xpre_column_161 bl_161 br_161 en_bar vdd precharge_1
Xpre_column_162 bl_162 br_162 en_bar vdd precharge_1
Xpre_column_163 bl_163 br_163 en_bar vdd precharge_1
Xpre_column_164 bl_164 br_164 en_bar vdd precharge_1
Xpre_column_165 bl_165 br_165 en_bar vdd precharge_1
Xpre_column_166 bl_166 br_166 en_bar vdd precharge_1
Xpre_column_167 bl_167 br_167 en_bar vdd precharge_1
Xpre_column_168 bl_168 br_168 en_bar vdd precharge_1
Xpre_column_169 bl_169 br_169 en_bar vdd precharge_1
Xpre_column_170 bl_170 br_170 en_bar vdd precharge_1
Xpre_column_171 bl_171 br_171 en_bar vdd precharge_1
Xpre_column_172 bl_172 br_172 en_bar vdd precharge_1
Xpre_column_173 bl_173 br_173 en_bar vdd precharge_1
Xpre_column_174 bl_174 br_174 en_bar vdd precharge_1
Xpre_column_175 bl_175 br_175 en_bar vdd precharge_1
Xpre_column_176 bl_176 br_176 en_bar vdd precharge_1
Xpre_column_177 bl_177 br_177 en_bar vdd precharge_1
Xpre_column_178 bl_178 br_178 en_bar vdd precharge_1
Xpre_column_179 bl_179 br_179 en_bar vdd precharge_1
Xpre_column_180 bl_180 br_180 en_bar vdd precharge_1
Xpre_column_181 bl_181 br_181 en_bar vdd precharge_1
Xpre_column_182 bl_182 br_182 en_bar vdd precharge_1
Xpre_column_183 bl_183 br_183 en_bar vdd precharge_1
Xpre_column_184 bl_184 br_184 en_bar vdd precharge_1
Xpre_column_185 bl_185 br_185 en_bar vdd precharge_1
Xpre_column_186 bl_186 br_186 en_bar vdd precharge_1
Xpre_column_187 bl_187 br_187 en_bar vdd precharge_1
Xpre_column_188 bl_188 br_188 en_bar vdd precharge_1
Xpre_column_189 bl_189 br_189 en_bar vdd precharge_1
Xpre_column_190 bl_190 br_190 en_bar vdd precharge_1
Xpre_column_191 bl_191 br_191 en_bar vdd precharge_1
Xpre_column_192 bl_192 br_192 en_bar vdd precharge_1
Xpre_column_193 bl_193 br_193 en_bar vdd precharge_1
Xpre_column_194 bl_194 br_194 en_bar vdd precharge_1
Xpre_column_195 bl_195 br_195 en_bar vdd precharge_1
Xpre_column_196 bl_196 br_196 en_bar vdd precharge_1
Xpre_column_197 bl_197 br_197 en_bar vdd precharge_1
Xpre_column_198 bl_198 br_198 en_bar vdd precharge_1
Xpre_column_199 bl_199 br_199 en_bar vdd precharge_1
Xpre_column_200 bl_200 br_200 en_bar vdd precharge_1
Xpre_column_201 bl_201 br_201 en_bar vdd precharge_1
Xpre_column_202 bl_202 br_202 en_bar vdd precharge_1
Xpre_column_203 bl_203 br_203 en_bar vdd precharge_1
Xpre_column_204 bl_204 br_204 en_bar vdd precharge_1
Xpre_column_205 bl_205 br_205 en_bar vdd precharge_1
Xpre_column_206 bl_206 br_206 en_bar vdd precharge_1
Xpre_column_207 bl_207 br_207 en_bar vdd precharge_1
Xpre_column_208 bl_208 br_208 en_bar vdd precharge_1
Xpre_column_209 bl_209 br_209 en_bar vdd precharge_1
Xpre_column_210 bl_210 br_210 en_bar vdd precharge_1
Xpre_column_211 bl_211 br_211 en_bar vdd precharge_1
Xpre_column_212 bl_212 br_212 en_bar vdd precharge_1
Xpre_column_213 bl_213 br_213 en_bar vdd precharge_1
Xpre_column_214 bl_214 br_214 en_bar vdd precharge_1
Xpre_column_215 bl_215 br_215 en_bar vdd precharge_1
Xpre_column_216 bl_216 br_216 en_bar vdd precharge_1
Xpre_column_217 bl_217 br_217 en_bar vdd precharge_1
Xpre_column_218 bl_218 br_218 en_bar vdd precharge_1
Xpre_column_219 bl_219 br_219 en_bar vdd precharge_1
Xpre_column_220 bl_220 br_220 en_bar vdd precharge_1
Xpre_column_221 bl_221 br_221 en_bar vdd precharge_1
Xpre_column_222 bl_222 br_222 en_bar vdd precharge_1
Xpre_column_223 bl_223 br_223 en_bar vdd precharge_1
Xpre_column_224 bl_224 br_224 en_bar vdd precharge_1
Xpre_column_225 bl_225 br_225 en_bar vdd precharge_1
Xpre_column_226 bl_226 br_226 en_bar vdd precharge_1
Xpre_column_227 bl_227 br_227 en_bar vdd precharge_1
Xpre_column_228 bl_228 br_228 en_bar vdd precharge_1
Xpre_column_229 bl_229 br_229 en_bar vdd precharge_1
Xpre_column_230 bl_230 br_230 en_bar vdd precharge_1
Xpre_column_231 bl_231 br_231 en_bar vdd precharge_1
Xpre_column_232 bl_232 br_232 en_bar vdd precharge_1
Xpre_column_233 bl_233 br_233 en_bar vdd precharge_1
Xpre_column_234 bl_234 br_234 en_bar vdd precharge_1
Xpre_column_235 bl_235 br_235 en_bar vdd precharge_1
Xpre_column_236 bl_236 br_236 en_bar vdd precharge_1
Xpre_column_237 bl_237 br_237 en_bar vdd precharge_1
Xpre_column_238 bl_238 br_238 en_bar vdd precharge_1
Xpre_column_239 bl_239 br_239 en_bar vdd precharge_1
Xpre_column_240 bl_240 br_240 en_bar vdd precharge_1
Xpre_column_241 bl_241 br_241 en_bar vdd precharge_1
Xpre_column_242 bl_242 br_242 en_bar vdd precharge_1
Xpre_column_243 bl_243 br_243 en_bar vdd precharge_1
Xpre_column_244 bl_244 br_244 en_bar vdd precharge_1
Xpre_column_245 bl_245 br_245 en_bar vdd precharge_1
Xpre_column_246 bl_246 br_246 en_bar vdd precharge_1
Xpre_column_247 bl_247 br_247 en_bar vdd precharge_1
Xpre_column_248 bl_248 br_248 en_bar vdd precharge_1
Xpre_column_249 bl_249 br_249 en_bar vdd precharge_1
Xpre_column_250 bl_250 br_250 en_bar vdd precharge_1
Xpre_column_251 bl_251 br_251 en_bar vdd precharge_1
Xpre_column_252 bl_252 br_252 en_bar vdd precharge_1
Xpre_column_253 bl_253 br_253 en_bar vdd precharge_1
Xpre_column_254 bl_254 br_254 en_bar vdd precharge_1
Xpre_column_255 bl_255 br_255 en_bar vdd precharge_1
Xpre_column_256 bl_256 br_256 en_bar vdd precharge_1
.ENDS precharge_array_0

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sense_amp_array_0 data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14 data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18 bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31 br_31 data_32 bl_32 br_32 data_33 bl_33 br_33 data_34 bl_34 br_34 data_35 bl_35 br_35 data_36 bl_36 br_36 data_37 bl_37 br_37 data_38 bl_38 br_38 data_39 bl_39 br_39 data_40 bl_40 br_40 data_41 bl_41 br_41 data_42 bl_42 br_42 data_43 bl_43 br_43 data_44 bl_44 br_44 data_45 bl_45 br_45 data_46 bl_46 br_46 data_47 bl_47 br_47 data_48 bl_48 br_48 data_49 bl_49 br_49 data_50 bl_50 br_50 data_51 bl_51 br_51 data_52 bl_52 br_52 data_53 bl_53 br_53 data_54 bl_54 br_54 data_55 bl_55 br_55 data_56 bl_56 br_56 data_57 bl_57 br_57 data_58 bl_58 br_58 data_59 bl_59 br_59 data_60 bl_60 br_60 data_61 bl_61 br_61 data_62 bl_62 br_62 data_63 bl_63 br_63 data_64 bl_64 br_64 data_65 bl_65 br_65 data_66 bl_66 br_66 data_67 bl_67 br_67 data_68 bl_68 br_68 data_69 bl_69 br_69 data_70 bl_70 br_70 data_71 bl_71 br_71 data_72 bl_72 br_72 data_73 bl_73 br_73 data_74 bl_74 br_74 data_75 bl_75 br_75 data_76 bl_76 br_76 data_77 bl_77 br_77 data_78 bl_78 br_78 data_79 bl_79 br_79 data_80 bl_80 br_80 data_81 bl_81 br_81 data_82 bl_82 br_82 data_83 bl_83 br_83 data_84 bl_84 br_84 data_85 bl_85 br_85 data_86 bl_86 br_86 data_87 bl_87 br_87 data_88 bl_88 br_88 data_89 bl_89 br_89 data_90 bl_90 br_90 data_91 bl_91 br_91 data_92 bl_92 br_92 data_93 bl_93 br_93 data_94 bl_94 br_94 data_95 bl_95 br_95 data_96 bl_96 br_96 data_97 bl_97 br_97 data_98 bl_98 br_98 data_99 bl_99 br_99 data_100 bl_100 br_100 data_101 bl_101 br_101 data_102 bl_102 br_102 data_103 bl_103 br_103 data_104 bl_104 br_104 data_105 bl_105 br_105 data_106 bl_106 br_106 data_107 bl_107 br_107 data_108 bl_108 br_108 data_109 bl_109 br_109 data_110 bl_110 br_110 data_111 bl_111 br_111 data_112 bl_112 br_112 data_113 bl_113 br_113 data_114 bl_114 br_114 data_115 bl_115 br_115 data_116 bl_116 br_116 data_117 bl_117 br_117 data_118 bl_118 br_118 data_119 bl_119 br_119 data_120 bl_120 br_120 data_121 bl_121 br_121 data_122 bl_122 br_122 data_123 bl_123 br_123 data_124 bl_124 br_124 data_125 bl_125 br_125 data_126 bl_126 br_126 data_127 bl_127 br_127 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* OUTPUT: data_32 
* INPUT : bl_32 
* INPUT : br_32 
* OUTPUT: data_33 
* INPUT : bl_33 
* INPUT : br_33 
* OUTPUT: data_34 
* INPUT : bl_34 
* INPUT : br_34 
* OUTPUT: data_35 
* INPUT : bl_35 
* INPUT : br_35 
* OUTPUT: data_36 
* INPUT : bl_36 
* INPUT : br_36 
* OUTPUT: data_37 
* INPUT : bl_37 
* INPUT : br_37 
* OUTPUT: data_38 
* INPUT : bl_38 
* INPUT : br_38 
* OUTPUT: data_39 
* INPUT : bl_39 
* INPUT : br_39 
* OUTPUT: data_40 
* INPUT : bl_40 
* INPUT : br_40 
* OUTPUT: data_41 
* INPUT : bl_41 
* INPUT : br_41 
* OUTPUT: data_42 
* INPUT : bl_42 
* INPUT : br_42 
* OUTPUT: data_43 
* INPUT : bl_43 
* INPUT : br_43 
* OUTPUT: data_44 
* INPUT : bl_44 
* INPUT : br_44 
* OUTPUT: data_45 
* INPUT : bl_45 
* INPUT : br_45 
* OUTPUT: data_46 
* INPUT : bl_46 
* INPUT : br_46 
* OUTPUT: data_47 
* INPUT : bl_47 
* INPUT : br_47 
* OUTPUT: data_48 
* INPUT : bl_48 
* INPUT : br_48 
* OUTPUT: data_49 
* INPUT : bl_49 
* INPUT : br_49 
* OUTPUT: data_50 
* INPUT : bl_50 
* INPUT : br_50 
* OUTPUT: data_51 
* INPUT : bl_51 
* INPUT : br_51 
* OUTPUT: data_52 
* INPUT : bl_52 
* INPUT : br_52 
* OUTPUT: data_53 
* INPUT : bl_53 
* INPUT : br_53 
* OUTPUT: data_54 
* INPUT : bl_54 
* INPUT : br_54 
* OUTPUT: data_55 
* INPUT : bl_55 
* INPUT : br_55 
* OUTPUT: data_56 
* INPUT : bl_56 
* INPUT : br_56 
* OUTPUT: data_57 
* INPUT : bl_57 
* INPUT : br_57 
* OUTPUT: data_58 
* INPUT : bl_58 
* INPUT : br_58 
* OUTPUT: data_59 
* INPUT : bl_59 
* INPUT : br_59 
* OUTPUT: data_60 
* INPUT : bl_60 
* INPUT : br_60 
* OUTPUT: data_61 
* INPUT : bl_61 
* INPUT : br_61 
* OUTPUT: data_62 
* INPUT : bl_62 
* INPUT : br_62 
* OUTPUT: data_63 
* INPUT : bl_63 
* INPUT : br_63 
* OUTPUT: data_64 
* INPUT : bl_64 
* INPUT : br_64 
* OUTPUT: data_65 
* INPUT : bl_65 
* INPUT : br_65 
* OUTPUT: data_66 
* INPUT : bl_66 
* INPUT : br_66 
* OUTPUT: data_67 
* INPUT : bl_67 
* INPUT : br_67 
* OUTPUT: data_68 
* INPUT : bl_68 
* INPUT : br_68 
* OUTPUT: data_69 
* INPUT : bl_69 
* INPUT : br_69 
* OUTPUT: data_70 
* INPUT : bl_70 
* INPUT : br_70 
* OUTPUT: data_71 
* INPUT : bl_71 
* INPUT : br_71 
* OUTPUT: data_72 
* INPUT : bl_72 
* INPUT : br_72 
* OUTPUT: data_73 
* INPUT : bl_73 
* INPUT : br_73 
* OUTPUT: data_74 
* INPUT : bl_74 
* INPUT : br_74 
* OUTPUT: data_75 
* INPUT : bl_75 
* INPUT : br_75 
* OUTPUT: data_76 
* INPUT : bl_76 
* INPUT : br_76 
* OUTPUT: data_77 
* INPUT : bl_77 
* INPUT : br_77 
* OUTPUT: data_78 
* INPUT : bl_78 
* INPUT : br_78 
* OUTPUT: data_79 
* INPUT : bl_79 
* INPUT : br_79 
* OUTPUT: data_80 
* INPUT : bl_80 
* INPUT : br_80 
* OUTPUT: data_81 
* INPUT : bl_81 
* INPUT : br_81 
* OUTPUT: data_82 
* INPUT : bl_82 
* INPUT : br_82 
* OUTPUT: data_83 
* INPUT : bl_83 
* INPUT : br_83 
* OUTPUT: data_84 
* INPUT : bl_84 
* INPUT : br_84 
* OUTPUT: data_85 
* INPUT : bl_85 
* INPUT : br_85 
* OUTPUT: data_86 
* INPUT : bl_86 
* INPUT : br_86 
* OUTPUT: data_87 
* INPUT : bl_87 
* INPUT : br_87 
* OUTPUT: data_88 
* INPUT : bl_88 
* INPUT : br_88 
* OUTPUT: data_89 
* INPUT : bl_89 
* INPUT : br_89 
* OUTPUT: data_90 
* INPUT : bl_90 
* INPUT : br_90 
* OUTPUT: data_91 
* INPUT : bl_91 
* INPUT : br_91 
* OUTPUT: data_92 
* INPUT : bl_92 
* INPUT : br_92 
* OUTPUT: data_93 
* INPUT : bl_93 
* INPUT : br_93 
* OUTPUT: data_94 
* INPUT : bl_94 
* INPUT : br_94 
* OUTPUT: data_95 
* INPUT : bl_95 
* INPUT : br_95 
* OUTPUT: data_96 
* INPUT : bl_96 
* INPUT : br_96 
* OUTPUT: data_97 
* INPUT : bl_97 
* INPUT : br_97 
* OUTPUT: data_98 
* INPUT : bl_98 
* INPUT : br_98 
* OUTPUT: data_99 
* INPUT : bl_99 
* INPUT : br_99 
* OUTPUT: data_100 
* INPUT : bl_100 
* INPUT : br_100 
* OUTPUT: data_101 
* INPUT : bl_101 
* INPUT : br_101 
* OUTPUT: data_102 
* INPUT : bl_102 
* INPUT : br_102 
* OUTPUT: data_103 
* INPUT : bl_103 
* INPUT : br_103 
* OUTPUT: data_104 
* INPUT : bl_104 
* INPUT : br_104 
* OUTPUT: data_105 
* INPUT : bl_105 
* INPUT : br_105 
* OUTPUT: data_106 
* INPUT : bl_106 
* INPUT : br_106 
* OUTPUT: data_107 
* INPUT : bl_107 
* INPUT : br_107 
* OUTPUT: data_108 
* INPUT : bl_108 
* INPUT : br_108 
* OUTPUT: data_109 
* INPUT : bl_109 
* INPUT : br_109 
* OUTPUT: data_110 
* INPUT : bl_110 
* INPUT : br_110 
* OUTPUT: data_111 
* INPUT : bl_111 
* INPUT : br_111 
* OUTPUT: data_112 
* INPUT : bl_112 
* INPUT : br_112 
* OUTPUT: data_113 
* INPUT : bl_113 
* INPUT : br_113 
* OUTPUT: data_114 
* INPUT : bl_114 
* INPUT : br_114 
* OUTPUT: data_115 
* INPUT : bl_115 
* INPUT : br_115 
* OUTPUT: data_116 
* INPUT : bl_116 
* INPUT : br_116 
* OUTPUT: data_117 
* INPUT : bl_117 
* INPUT : br_117 
* OUTPUT: data_118 
* INPUT : bl_118 
* INPUT : br_118 
* OUTPUT: data_119 
* INPUT : bl_119 
* INPUT : br_119 
* OUTPUT: data_120 
* INPUT : bl_120 
* INPUT : br_120 
* OUTPUT: data_121 
* INPUT : bl_121 
* INPUT : br_121 
* OUTPUT: data_122 
* INPUT : bl_122 
* INPUT : br_122 
* OUTPUT: data_123 
* INPUT : bl_123 
* INPUT : br_123 
* OUTPUT: data_124 
* INPUT : bl_124 
* INPUT : br_124 
* OUTPUT: data_125 
* INPUT : bl_125 
* INPUT : br_125 
* OUTPUT: data_126 
* INPUT : bl_126 
* INPUT : br_126 
* OUTPUT: data_127 
* INPUT : bl_127 
* INPUT : br_127 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 2
Xsa_d0 bl_0 br_0 data_0 en vdd gnd sense_amp
Xsa_d1 bl_1 br_1 data_1 en vdd gnd sense_amp
Xsa_d2 bl_2 br_2 data_2 en vdd gnd sense_amp
Xsa_d3 bl_3 br_3 data_3 en vdd gnd sense_amp
Xsa_d4 bl_4 br_4 data_4 en vdd gnd sense_amp
Xsa_d5 bl_5 br_5 data_5 en vdd gnd sense_amp
Xsa_d6 bl_6 br_6 data_6 en vdd gnd sense_amp
Xsa_d7 bl_7 br_7 data_7 en vdd gnd sense_amp
Xsa_d8 bl_8 br_8 data_8 en vdd gnd sense_amp
Xsa_d9 bl_9 br_9 data_9 en vdd gnd sense_amp
Xsa_d10 bl_10 br_10 data_10 en vdd gnd sense_amp
Xsa_d11 bl_11 br_11 data_11 en vdd gnd sense_amp
Xsa_d12 bl_12 br_12 data_12 en vdd gnd sense_amp
Xsa_d13 bl_13 br_13 data_13 en vdd gnd sense_amp
Xsa_d14 bl_14 br_14 data_14 en vdd gnd sense_amp
Xsa_d15 bl_15 br_15 data_15 en vdd gnd sense_amp
Xsa_d16 bl_16 br_16 data_16 en vdd gnd sense_amp
Xsa_d17 bl_17 br_17 data_17 en vdd gnd sense_amp
Xsa_d18 bl_18 br_18 data_18 en vdd gnd sense_amp
Xsa_d19 bl_19 br_19 data_19 en vdd gnd sense_amp
Xsa_d20 bl_20 br_20 data_20 en vdd gnd sense_amp
Xsa_d21 bl_21 br_21 data_21 en vdd gnd sense_amp
Xsa_d22 bl_22 br_22 data_22 en vdd gnd sense_amp
Xsa_d23 bl_23 br_23 data_23 en vdd gnd sense_amp
Xsa_d24 bl_24 br_24 data_24 en vdd gnd sense_amp
Xsa_d25 bl_25 br_25 data_25 en vdd gnd sense_amp
Xsa_d26 bl_26 br_26 data_26 en vdd gnd sense_amp
Xsa_d27 bl_27 br_27 data_27 en vdd gnd sense_amp
Xsa_d28 bl_28 br_28 data_28 en vdd gnd sense_amp
Xsa_d29 bl_29 br_29 data_29 en vdd gnd sense_amp
Xsa_d30 bl_30 br_30 data_30 en vdd gnd sense_amp
Xsa_d31 bl_31 br_31 data_31 en vdd gnd sense_amp
Xsa_d32 bl_32 br_32 data_32 en vdd gnd sense_amp
Xsa_d33 bl_33 br_33 data_33 en vdd gnd sense_amp
Xsa_d34 bl_34 br_34 data_34 en vdd gnd sense_amp
Xsa_d35 bl_35 br_35 data_35 en vdd gnd sense_amp
Xsa_d36 bl_36 br_36 data_36 en vdd gnd sense_amp
Xsa_d37 bl_37 br_37 data_37 en vdd gnd sense_amp
Xsa_d38 bl_38 br_38 data_38 en vdd gnd sense_amp
Xsa_d39 bl_39 br_39 data_39 en vdd gnd sense_amp
Xsa_d40 bl_40 br_40 data_40 en vdd gnd sense_amp
Xsa_d41 bl_41 br_41 data_41 en vdd gnd sense_amp
Xsa_d42 bl_42 br_42 data_42 en vdd gnd sense_amp
Xsa_d43 bl_43 br_43 data_43 en vdd gnd sense_amp
Xsa_d44 bl_44 br_44 data_44 en vdd gnd sense_amp
Xsa_d45 bl_45 br_45 data_45 en vdd gnd sense_amp
Xsa_d46 bl_46 br_46 data_46 en vdd gnd sense_amp
Xsa_d47 bl_47 br_47 data_47 en vdd gnd sense_amp
Xsa_d48 bl_48 br_48 data_48 en vdd gnd sense_amp
Xsa_d49 bl_49 br_49 data_49 en vdd gnd sense_amp
Xsa_d50 bl_50 br_50 data_50 en vdd gnd sense_amp
Xsa_d51 bl_51 br_51 data_51 en vdd gnd sense_amp
Xsa_d52 bl_52 br_52 data_52 en vdd gnd sense_amp
Xsa_d53 bl_53 br_53 data_53 en vdd gnd sense_amp
Xsa_d54 bl_54 br_54 data_54 en vdd gnd sense_amp
Xsa_d55 bl_55 br_55 data_55 en vdd gnd sense_amp
Xsa_d56 bl_56 br_56 data_56 en vdd gnd sense_amp
Xsa_d57 bl_57 br_57 data_57 en vdd gnd sense_amp
Xsa_d58 bl_58 br_58 data_58 en vdd gnd sense_amp
Xsa_d59 bl_59 br_59 data_59 en vdd gnd sense_amp
Xsa_d60 bl_60 br_60 data_60 en vdd gnd sense_amp
Xsa_d61 bl_61 br_61 data_61 en vdd gnd sense_amp
Xsa_d62 bl_62 br_62 data_62 en vdd gnd sense_amp
Xsa_d63 bl_63 br_63 data_63 en vdd gnd sense_amp
Xsa_d64 bl_64 br_64 data_64 en vdd gnd sense_amp
Xsa_d65 bl_65 br_65 data_65 en vdd gnd sense_amp
Xsa_d66 bl_66 br_66 data_66 en vdd gnd sense_amp
Xsa_d67 bl_67 br_67 data_67 en vdd gnd sense_amp
Xsa_d68 bl_68 br_68 data_68 en vdd gnd sense_amp
Xsa_d69 bl_69 br_69 data_69 en vdd gnd sense_amp
Xsa_d70 bl_70 br_70 data_70 en vdd gnd sense_amp
Xsa_d71 bl_71 br_71 data_71 en vdd gnd sense_amp
Xsa_d72 bl_72 br_72 data_72 en vdd gnd sense_amp
Xsa_d73 bl_73 br_73 data_73 en vdd gnd sense_amp
Xsa_d74 bl_74 br_74 data_74 en vdd gnd sense_amp
Xsa_d75 bl_75 br_75 data_75 en vdd gnd sense_amp
Xsa_d76 bl_76 br_76 data_76 en vdd gnd sense_amp
Xsa_d77 bl_77 br_77 data_77 en vdd gnd sense_amp
Xsa_d78 bl_78 br_78 data_78 en vdd gnd sense_amp
Xsa_d79 bl_79 br_79 data_79 en vdd gnd sense_amp
Xsa_d80 bl_80 br_80 data_80 en vdd gnd sense_amp
Xsa_d81 bl_81 br_81 data_81 en vdd gnd sense_amp
Xsa_d82 bl_82 br_82 data_82 en vdd gnd sense_amp
Xsa_d83 bl_83 br_83 data_83 en vdd gnd sense_amp
Xsa_d84 bl_84 br_84 data_84 en vdd gnd sense_amp
Xsa_d85 bl_85 br_85 data_85 en vdd gnd sense_amp
Xsa_d86 bl_86 br_86 data_86 en vdd gnd sense_amp
Xsa_d87 bl_87 br_87 data_87 en vdd gnd sense_amp
Xsa_d88 bl_88 br_88 data_88 en vdd gnd sense_amp
Xsa_d89 bl_89 br_89 data_89 en vdd gnd sense_amp
Xsa_d90 bl_90 br_90 data_90 en vdd gnd sense_amp
Xsa_d91 bl_91 br_91 data_91 en vdd gnd sense_amp
Xsa_d92 bl_92 br_92 data_92 en vdd gnd sense_amp
Xsa_d93 bl_93 br_93 data_93 en vdd gnd sense_amp
Xsa_d94 bl_94 br_94 data_94 en vdd gnd sense_amp
Xsa_d95 bl_95 br_95 data_95 en vdd gnd sense_amp
Xsa_d96 bl_96 br_96 data_96 en vdd gnd sense_amp
Xsa_d97 bl_97 br_97 data_97 en vdd gnd sense_amp
Xsa_d98 bl_98 br_98 data_98 en vdd gnd sense_amp
Xsa_d99 bl_99 br_99 data_99 en vdd gnd sense_amp
Xsa_d100 bl_100 br_100 data_100 en vdd gnd sense_amp
Xsa_d101 bl_101 br_101 data_101 en vdd gnd sense_amp
Xsa_d102 bl_102 br_102 data_102 en vdd gnd sense_amp
Xsa_d103 bl_103 br_103 data_103 en vdd gnd sense_amp
Xsa_d104 bl_104 br_104 data_104 en vdd gnd sense_amp
Xsa_d105 bl_105 br_105 data_105 en vdd gnd sense_amp
Xsa_d106 bl_106 br_106 data_106 en vdd gnd sense_amp
Xsa_d107 bl_107 br_107 data_107 en vdd gnd sense_amp
Xsa_d108 bl_108 br_108 data_108 en vdd gnd sense_amp
Xsa_d109 bl_109 br_109 data_109 en vdd gnd sense_amp
Xsa_d110 bl_110 br_110 data_110 en vdd gnd sense_amp
Xsa_d111 bl_111 br_111 data_111 en vdd gnd sense_amp
Xsa_d112 bl_112 br_112 data_112 en vdd gnd sense_amp
Xsa_d113 bl_113 br_113 data_113 en vdd gnd sense_amp
Xsa_d114 bl_114 br_114 data_114 en vdd gnd sense_amp
Xsa_d115 bl_115 br_115 data_115 en vdd gnd sense_amp
Xsa_d116 bl_116 br_116 data_116 en vdd gnd sense_amp
Xsa_d117 bl_117 br_117 data_117 en vdd gnd sense_amp
Xsa_d118 bl_118 br_118 data_118 en vdd gnd sense_amp
Xsa_d119 bl_119 br_119 data_119 en vdd gnd sense_amp
Xsa_d120 bl_120 br_120 data_120 en vdd gnd sense_amp
Xsa_d121 bl_121 br_121 data_121 en vdd gnd sense_amp
Xsa_d122 bl_122 br_122 data_122 en vdd gnd sense_amp
Xsa_d123 bl_123 br_123 data_123 en vdd gnd sense_amp
Xsa_d124 bl_124 br_124 data_124 en vdd gnd sense_amp
Xsa_d125 bl_125 br_125 data_125 en vdd gnd sense_amp
Xsa_d126 bl_126 br_126 data_126 en vdd gnd sense_amp
Xsa_d127 bl_127 br_127 data_127 en vdd gnd sense_amp
.ENDS sense_amp_array_0

* ptx M{0} {1} nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT single_level_column_mux_0 bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Mmux_tx1 bl sel bl_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mmux_tx2 br sel br_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
.ENDS single_level_column_mux_0

.SUBCKT single_level_column_mux_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 sel_0 sel_1 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 bl_out_32 br_out_32 bl_out_33 br_out_33 bl_out_34 br_out_34 bl_out_35 br_out_35 bl_out_36 br_out_36 bl_out_37 br_out_37 bl_out_38 br_out_38 bl_out_39 br_out_39 bl_out_40 br_out_40 bl_out_41 br_out_41 bl_out_42 br_out_42 bl_out_43 br_out_43 bl_out_44 br_out_44 bl_out_45 br_out_45 bl_out_46 br_out_46 bl_out_47 br_out_47 bl_out_48 br_out_48 bl_out_49 br_out_49 bl_out_50 br_out_50 bl_out_51 br_out_51 bl_out_52 br_out_52 bl_out_53 br_out_53 bl_out_54 br_out_54 bl_out_55 br_out_55 bl_out_56 br_out_56 bl_out_57 br_out_57 bl_out_58 br_out_58 bl_out_59 br_out_59 bl_out_60 br_out_60 bl_out_61 br_out_61 bl_out_62 br_out_62 bl_out_63 br_out_63 bl_out_64 br_out_64 bl_out_65 br_out_65 bl_out_66 br_out_66 bl_out_67 br_out_67 bl_out_68 br_out_68 bl_out_69 br_out_69 bl_out_70 br_out_70 bl_out_71 br_out_71 bl_out_72 br_out_72 bl_out_73 br_out_73 bl_out_74 br_out_74 bl_out_75 br_out_75 bl_out_76 br_out_76 bl_out_77 br_out_77 bl_out_78 br_out_78 bl_out_79 br_out_79 bl_out_80 br_out_80 bl_out_81 br_out_81 bl_out_82 br_out_82 bl_out_83 br_out_83 bl_out_84 br_out_84 bl_out_85 br_out_85 bl_out_86 br_out_86 bl_out_87 br_out_87 bl_out_88 br_out_88 bl_out_89 br_out_89 bl_out_90 br_out_90 bl_out_91 br_out_91 bl_out_92 br_out_92 bl_out_93 br_out_93 bl_out_94 br_out_94 bl_out_95 br_out_95 bl_out_96 br_out_96 bl_out_97 br_out_97 bl_out_98 br_out_98 bl_out_99 br_out_99 bl_out_100 br_out_100 bl_out_101 br_out_101 bl_out_102 br_out_102 bl_out_103 br_out_103 bl_out_104 br_out_104 bl_out_105 br_out_105 bl_out_106 br_out_106 bl_out_107 br_out_107 bl_out_108 br_out_108 bl_out_109 br_out_109 bl_out_110 br_out_110 bl_out_111 br_out_111 bl_out_112 br_out_112 bl_out_113 br_out_113 bl_out_114 br_out_114 bl_out_115 br_out_115 bl_out_116 br_out_116 bl_out_117 br_out_117 bl_out_118 br_out_118 bl_out_119 br_out_119 bl_out_120 br_out_120 bl_out_121 br_out_121 bl_out_122 br_out_122 bl_out_123 br_out_123 bl_out_124 br_out_124 bl_out_125 br_out_125 bl_out_126 br_out_126 bl_out_127 br_out_127 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : bl_out_32 
* INOUT : br_out_32 
* INOUT : bl_out_33 
* INOUT : br_out_33 
* INOUT : bl_out_34 
* INOUT : br_out_34 
* INOUT : bl_out_35 
* INOUT : br_out_35 
* INOUT : bl_out_36 
* INOUT : br_out_36 
* INOUT : bl_out_37 
* INOUT : br_out_37 
* INOUT : bl_out_38 
* INOUT : br_out_38 
* INOUT : bl_out_39 
* INOUT : br_out_39 
* INOUT : bl_out_40 
* INOUT : br_out_40 
* INOUT : bl_out_41 
* INOUT : br_out_41 
* INOUT : bl_out_42 
* INOUT : br_out_42 
* INOUT : bl_out_43 
* INOUT : br_out_43 
* INOUT : bl_out_44 
* INOUT : br_out_44 
* INOUT : bl_out_45 
* INOUT : br_out_45 
* INOUT : bl_out_46 
* INOUT : br_out_46 
* INOUT : bl_out_47 
* INOUT : br_out_47 
* INOUT : bl_out_48 
* INOUT : br_out_48 
* INOUT : bl_out_49 
* INOUT : br_out_49 
* INOUT : bl_out_50 
* INOUT : br_out_50 
* INOUT : bl_out_51 
* INOUT : br_out_51 
* INOUT : bl_out_52 
* INOUT : br_out_52 
* INOUT : bl_out_53 
* INOUT : br_out_53 
* INOUT : bl_out_54 
* INOUT : br_out_54 
* INOUT : bl_out_55 
* INOUT : br_out_55 
* INOUT : bl_out_56 
* INOUT : br_out_56 
* INOUT : bl_out_57 
* INOUT : br_out_57 
* INOUT : bl_out_58 
* INOUT : br_out_58 
* INOUT : bl_out_59 
* INOUT : br_out_59 
* INOUT : bl_out_60 
* INOUT : br_out_60 
* INOUT : bl_out_61 
* INOUT : br_out_61 
* INOUT : bl_out_62 
* INOUT : br_out_62 
* INOUT : bl_out_63 
* INOUT : br_out_63 
* INOUT : bl_out_64 
* INOUT : br_out_64 
* INOUT : bl_out_65 
* INOUT : br_out_65 
* INOUT : bl_out_66 
* INOUT : br_out_66 
* INOUT : bl_out_67 
* INOUT : br_out_67 
* INOUT : bl_out_68 
* INOUT : br_out_68 
* INOUT : bl_out_69 
* INOUT : br_out_69 
* INOUT : bl_out_70 
* INOUT : br_out_70 
* INOUT : bl_out_71 
* INOUT : br_out_71 
* INOUT : bl_out_72 
* INOUT : br_out_72 
* INOUT : bl_out_73 
* INOUT : br_out_73 
* INOUT : bl_out_74 
* INOUT : br_out_74 
* INOUT : bl_out_75 
* INOUT : br_out_75 
* INOUT : bl_out_76 
* INOUT : br_out_76 
* INOUT : bl_out_77 
* INOUT : br_out_77 
* INOUT : bl_out_78 
* INOUT : br_out_78 
* INOUT : bl_out_79 
* INOUT : br_out_79 
* INOUT : bl_out_80 
* INOUT : br_out_80 
* INOUT : bl_out_81 
* INOUT : br_out_81 
* INOUT : bl_out_82 
* INOUT : br_out_82 
* INOUT : bl_out_83 
* INOUT : br_out_83 
* INOUT : bl_out_84 
* INOUT : br_out_84 
* INOUT : bl_out_85 
* INOUT : br_out_85 
* INOUT : bl_out_86 
* INOUT : br_out_86 
* INOUT : bl_out_87 
* INOUT : br_out_87 
* INOUT : bl_out_88 
* INOUT : br_out_88 
* INOUT : bl_out_89 
* INOUT : br_out_89 
* INOUT : bl_out_90 
* INOUT : br_out_90 
* INOUT : bl_out_91 
* INOUT : br_out_91 
* INOUT : bl_out_92 
* INOUT : br_out_92 
* INOUT : bl_out_93 
* INOUT : br_out_93 
* INOUT : bl_out_94 
* INOUT : br_out_94 
* INOUT : bl_out_95 
* INOUT : br_out_95 
* INOUT : bl_out_96 
* INOUT : br_out_96 
* INOUT : bl_out_97 
* INOUT : br_out_97 
* INOUT : bl_out_98 
* INOUT : br_out_98 
* INOUT : bl_out_99 
* INOUT : br_out_99 
* INOUT : bl_out_100 
* INOUT : br_out_100 
* INOUT : bl_out_101 
* INOUT : br_out_101 
* INOUT : bl_out_102 
* INOUT : br_out_102 
* INOUT : bl_out_103 
* INOUT : br_out_103 
* INOUT : bl_out_104 
* INOUT : br_out_104 
* INOUT : bl_out_105 
* INOUT : br_out_105 
* INOUT : bl_out_106 
* INOUT : br_out_106 
* INOUT : bl_out_107 
* INOUT : br_out_107 
* INOUT : bl_out_108 
* INOUT : br_out_108 
* INOUT : bl_out_109 
* INOUT : br_out_109 
* INOUT : bl_out_110 
* INOUT : br_out_110 
* INOUT : bl_out_111 
* INOUT : br_out_111 
* INOUT : bl_out_112 
* INOUT : br_out_112 
* INOUT : bl_out_113 
* INOUT : br_out_113 
* INOUT : bl_out_114 
* INOUT : br_out_114 
* INOUT : bl_out_115 
* INOUT : br_out_115 
* INOUT : bl_out_116 
* INOUT : br_out_116 
* INOUT : bl_out_117 
* INOUT : br_out_117 
* INOUT : bl_out_118 
* INOUT : br_out_118 
* INOUT : bl_out_119 
* INOUT : br_out_119 
* INOUT : bl_out_120 
* INOUT : br_out_120 
* INOUT : bl_out_121 
* INOUT : br_out_121 
* INOUT : bl_out_122 
* INOUT : br_out_122 
* INOUT : bl_out_123 
* INOUT : br_out_123 
* INOUT : bl_out_124 
* INOUT : br_out_124 
* INOUT : bl_out_125 
* INOUT : br_out_125 
* INOUT : bl_out_126 
* INOUT : br_out_126 
* INOUT : bl_out_127 
* INOUT : br_out_127 
* INOUT : gnd 
* cols: 256 word_size: 128 bl: bl br: br
XXMUX0 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd single_level_column_mux_0
XXMUX1 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd single_level_column_mux_0
XXMUX2 bl_2 br_2 bl_out_1 br_out_1 sel_0 gnd single_level_column_mux_0
XXMUX3 bl_3 br_3 bl_out_1 br_out_1 sel_1 gnd single_level_column_mux_0
XXMUX4 bl_4 br_4 bl_out_2 br_out_2 sel_0 gnd single_level_column_mux_0
XXMUX5 bl_5 br_5 bl_out_2 br_out_2 sel_1 gnd single_level_column_mux_0
XXMUX6 bl_6 br_6 bl_out_3 br_out_3 sel_0 gnd single_level_column_mux_0
XXMUX7 bl_7 br_7 bl_out_3 br_out_3 sel_1 gnd single_level_column_mux_0
XXMUX8 bl_8 br_8 bl_out_4 br_out_4 sel_0 gnd single_level_column_mux_0
XXMUX9 bl_9 br_9 bl_out_4 br_out_4 sel_1 gnd single_level_column_mux_0
XXMUX10 bl_10 br_10 bl_out_5 br_out_5 sel_0 gnd single_level_column_mux_0
XXMUX11 bl_11 br_11 bl_out_5 br_out_5 sel_1 gnd single_level_column_mux_0
XXMUX12 bl_12 br_12 bl_out_6 br_out_6 sel_0 gnd single_level_column_mux_0
XXMUX13 bl_13 br_13 bl_out_6 br_out_6 sel_1 gnd single_level_column_mux_0
XXMUX14 bl_14 br_14 bl_out_7 br_out_7 sel_0 gnd single_level_column_mux_0
XXMUX15 bl_15 br_15 bl_out_7 br_out_7 sel_1 gnd single_level_column_mux_0
XXMUX16 bl_16 br_16 bl_out_8 br_out_8 sel_0 gnd single_level_column_mux_0
XXMUX17 bl_17 br_17 bl_out_8 br_out_8 sel_1 gnd single_level_column_mux_0
XXMUX18 bl_18 br_18 bl_out_9 br_out_9 sel_0 gnd single_level_column_mux_0
XXMUX19 bl_19 br_19 bl_out_9 br_out_9 sel_1 gnd single_level_column_mux_0
XXMUX20 bl_20 br_20 bl_out_10 br_out_10 sel_0 gnd single_level_column_mux_0
XXMUX21 bl_21 br_21 bl_out_10 br_out_10 sel_1 gnd single_level_column_mux_0
XXMUX22 bl_22 br_22 bl_out_11 br_out_11 sel_0 gnd single_level_column_mux_0
XXMUX23 bl_23 br_23 bl_out_11 br_out_11 sel_1 gnd single_level_column_mux_0
XXMUX24 bl_24 br_24 bl_out_12 br_out_12 sel_0 gnd single_level_column_mux_0
XXMUX25 bl_25 br_25 bl_out_12 br_out_12 sel_1 gnd single_level_column_mux_0
XXMUX26 bl_26 br_26 bl_out_13 br_out_13 sel_0 gnd single_level_column_mux_0
XXMUX27 bl_27 br_27 bl_out_13 br_out_13 sel_1 gnd single_level_column_mux_0
XXMUX28 bl_28 br_28 bl_out_14 br_out_14 sel_0 gnd single_level_column_mux_0
XXMUX29 bl_29 br_29 bl_out_14 br_out_14 sel_1 gnd single_level_column_mux_0
XXMUX30 bl_30 br_30 bl_out_15 br_out_15 sel_0 gnd single_level_column_mux_0
XXMUX31 bl_31 br_31 bl_out_15 br_out_15 sel_1 gnd single_level_column_mux_0
XXMUX32 bl_32 br_32 bl_out_16 br_out_16 sel_0 gnd single_level_column_mux_0
XXMUX33 bl_33 br_33 bl_out_16 br_out_16 sel_1 gnd single_level_column_mux_0
XXMUX34 bl_34 br_34 bl_out_17 br_out_17 sel_0 gnd single_level_column_mux_0
XXMUX35 bl_35 br_35 bl_out_17 br_out_17 sel_1 gnd single_level_column_mux_0
XXMUX36 bl_36 br_36 bl_out_18 br_out_18 sel_0 gnd single_level_column_mux_0
XXMUX37 bl_37 br_37 bl_out_18 br_out_18 sel_1 gnd single_level_column_mux_0
XXMUX38 bl_38 br_38 bl_out_19 br_out_19 sel_0 gnd single_level_column_mux_0
XXMUX39 bl_39 br_39 bl_out_19 br_out_19 sel_1 gnd single_level_column_mux_0
XXMUX40 bl_40 br_40 bl_out_20 br_out_20 sel_0 gnd single_level_column_mux_0
XXMUX41 bl_41 br_41 bl_out_20 br_out_20 sel_1 gnd single_level_column_mux_0
XXMUX42 bl_42 br_42 bl_out_21 br_out_21 sel_0 gnd single_level_column_mux_0
XXMUX43 bl_43 br_43 bl_out_21 br_out_21 sel_1 gnd single_level_column_mux_0
XXMUX44 bl_44 br_44 bl_out_22 br_out_22 sel_0 gnd single_level_column_mux_0
XXMUX45 bl_45 br_45 bl_out_22 br_out_22 sel_1 gnd single_level_column_mux_0
XXMUX46 bl_46 br_46 bl_out_23 br_out_23 sel_0 gnd single_level_column_mux_0
XXMUX47 bl_47 br_47 bl_out_23 br_out_23 sel_1 gnd single_level_column_mux_0
XXMUX48 bl_48 br_48 bl_out_24 br_out_24 sel_0 gnd single_level_column_mux_0
XXMUX49 bl_49 br_49 bl_out_24 br_out_24 sel_1 gnd single_level_column_mux_0
XXMUX50 bl_50 br_50 bl_out_25 br_out_25 sel_0 gnd single_level_column_mux_0
XXMUX51 bl_51 br_51 bl_out_25 br_out_25 sel_1 gnd single_level_column_mux_0
XXMUX52 bl_52 br_52 bl_out_26 br_out_26 sel_0 gnd single_level_column_mux_0
XXMUX53 bl_53 br_53 bl_out_26 br_out_26 sel_1 gnd single_level_column_mux_0
XXMUX54 bl_54 br_54 bl_out_27 br_out_27 sel_0 gnd single_level_column_mux_0
XXMUX55 bl_55 br_55 bl_out_27 br_out_27 sel_1 gnd single_level_column_mux_0
XXMUX56 bl_56 br_56 bl_out_28 br_out_28 sel_0 gnd single_level_column_mux_0
XXMUX57 bl_57 br_57 bl_out_28 br_out_28 sel_1 gnd single_level_column_mux_0
XXMUX58 bl_58 br_58 bl_out_29 br_out_29 sel_0 gnd single_level_column_mux_0
XXMUX59 bl_59 br_59 bl_out_29 br_out_29 sel_1 gnd single_level_column_mux_0
XXMUX60 bl_60 br_60 bl_out_30 br_out_30 sel_0 gnd single_level_column_mux_0
XXMUX61 bl_61 br_61 bl_out_30 br_out_30 sel_1 gnd single_level_column_mux_0
XXMUX62 bl_62 br_62 bl_out_31 br_out_31 sel_0 gnd single_level_column_mux_0
XXMUX63 bl_63 br_63 bl_out_31 br_out_31 sel_1 gnd single_level_column_mux_0
XXMUX64 bl_64 br_64 bl_out_32 br_out_32 sel_0 gnd single_level_column_mux_0
XXMUX65 bl_65 br_65 bl_out_32 br_out_32 sel_1 gnd single_level_column_mux_0
XXMUX66 bl_66 br_66 bl_out_33 br_out_33 sel_0 gnd single_level_column_mux_0
XXMUX67 bl_67 br_67 bl_out_33 br_out_33 sel_1 gnd single_level_column_mux_0
XXMUX68 bl_68 br_68 bl_out_34 br_out_34 sel_0 gnd single_level_column_mux_0
XXMUX69 bl_69 br_69 bl_out_34 br_out_34 sel_1 gnd single_level_column_mux_0
XXMUX70 bl_70 br_70 bl_out_35 br_out_35 sel_0 gnd single_level_column_mux_0
XXMUX71 bl_71 br_71 bl_out_35 br_out_35 sel_1 gnd single_level_column_mux_0
XXMUX72 bl_72 br_72 bl_out_36 br_out_36 sel_0 gnd single_level_column_mux_0
XXMUX73 bl_73 br_73 bl_out_36 br_out_36 sel_1 gnd single_level_column_mux_0
XXMUX74 bl_74 br_74 bl_out_37 br_out_37 sel_0 gnd single_level_column_mux_0
XXMUX75 bl_75 br_75 bl_out_37 br_out_37 sel_1 gnd single_level_column_mux_0
XXMUX76 bl_76 br_76 bl_out_38 br_out_38 sel_0 gnd single_level_column_mux_0
XXMUX77 bl_77 br_77 bl_out_38 br_out_38 sel_1 gnd single_level_column_mux_0
XXMUX78 bl_78 br_78 bl_out_39 br_out_39 sel_0 gnd single_level_column_mux_0
XXMUX79 bl_79 br_79 bl_out_39 br_out_39 sel_1 gnd single_level_column_mux_0
XXMUX80 bl_80 br_80 bl_out_40 br_out_40 sel_0 gnd single_level_column_mux_0
XXMUX81 bl_81 br_81 bl_out_40 br_out_40 sel_1 gnd single_level_column_mux_0
XXMUX82 bl_82 br_82 bl_out_41 br_out_41 sel_0 gnd single_level_column_mux_0
XXMUX83 bl_83 br_83 bl_out_41 br_out_41 sel_1 gnd single_level_column_mux_0
XXMUX84 bl_84 br_84 bl_out_42 br_out_42 sel_0 gnd single_level_column_mux_0
XXMUX85 bl_85 br_85 bl_out_42 br_out_42 sel_1 gnd single_level_column_mux_0
XXMUX86 bl_86 br_86 bl_out_43 br_out_43 sel_0 gnd single_level_column_mux_0
XXMUX87 bl_87 br_87 bl_out_43 br_out_43 sel_1 gnd single_level_column_mux_0
XXMUX88 bl_88 br_88 bl_out_44 br_out_44 sel_0 gnd single_level_column_mux_0
XXMUX89 bl_89 br_89 bl_out_44 br_out_44 sel_1 gnd single_level_column_mux_0
XXMUX90 bl_90 br_90 bl_out_45 br_out_45 sel_0 gnd single_level_column_mux_0
XXMUX91 bl_91 br_91 bl_out_45 br_out_45 sel_1 gnd single_level_column_mux_0
XXMUX92 bl_92 br_92 bl_out_46 br_out_46 sel_0 gnd single_level_column_mux_0
XXMUX93 bl_93 br_93 bl_out_46 br_out_46 sel_1 gnd single_level_column_mux_0
XXMUX94 bl_94 br_94 bl_out_47 br_out_47 sel_0 gnd single_level_column_mux_0
XXMUX95 bl_95 br_95 bl_out_47 br_out_47 sel_1 gnd single_level_column_mux_0
XXMUX96 bl_96 br_96 bl_out_48 br_out_48 sel_0 gnd single_level_column_mux_0
XXMUX97 bl_97 br_97 bl_out_48 br_out_48 sel_1 gnd single_level_column_mux_0
XXMUX98 bl_98 br_98 bl_out_49 br_out_49 sel_0 gnd single_level_column_mux_0
XXMUX99 bl_99 br_99 bl_out_49 br_out_49 sel_1 gnd single_level_column_mux_0
XXMUX100 bl_100 br_100 bl_out_50 br_out_50 sel_0 gnd single_level_column_mux_0
XXMUX101 bl_101 br_101 bl_out_50 br_out_50 sel_1 gnd single_level_column_mux_0
XXMUX102 bl_102 br_102 bl_out_51 br_out_51 sel_0 gnd single_level_column_mux_0
XXMUX103 bl_103 br_103 bl_out_51 br_out_51 sel_1 gnd single_level_column_mux_0
XXMUX104 bl_104 br_104 bl_out_52 br_out_52 sel_0 gnd single_level_column_mux_0
XXMUX105 bl_105 br_105 bl_out_52 br_out_52 sel_1 gnd single_level_column_mux_0
XXMUX106 bl_106 br_106 bl_out_53 br_out_53 sel_0 gnd single_level_column_mux_0
XXMUX107 bl_107 br_107 bl_out_53 br_out_53 sel_1 gnd single_level_column_mux_0
XXMUX108 bl_108 br_108 bl_out_54 br_out_54 sel_0 gnd single_level_column_mux_0
XXMUX109 bl_109 br_109 bl_out_54 br_out_54 sel_1 gnd single_level_column_mux_0
XXMUX110 bl_110 br_110 bl_out_55 br_out_55 sel_0 gnd single_level_column_mux_0
XXMUX111 bl_111 br_111 bl_out_55 br_out_55 sel_1 gnd single_level_column_mux_0
XXMUX112 bl_112 br_112 bl_out_56 br_out_56 sel_0 gnd single_level_column_mux_0
XXMUX113 bl_113 br_113 bl_out_56 br_out_56 sel_1 gnd single_level_column_mux_0
XXMUX114 bl_114 br_114 bl_out_57 br_out_57 sel_0 gnd single_level_column_mux_0
XXMUX115 bl_115 br_115 bl_out_57 br_out_57 sel_1 gnd single_level_column_mux_0
XXMUX116 bl_116 br_116 bl_out_58 br_out_58 sel_0 gnd single_level_column_mux_0
XXMUX117 bl_117 br_117 bl_out_58 br_out_58 sel_1 gnd single_level_column_mux_0
XXMUX118 bl_118 br_118 bl_out_59 br_out_59 sel_0 gnd single_level_column_mux_0
XXMUX119 bl_119 br_119 bl_out_59 br_out_59 sel_1 gnd single_level_column_mux_0
XXMUX120 bl_120 br_120 bl_out_60 br_out_60 sel_0 gnd single_level_column_mux_0
XXMUX121 bl_121 br_121 bl_out_60 br_out_60 sel_1 gnd single_level_column_mux_0
XXMUX122 bl_122 br_122 bl_out_61 br_out_61 sel_0 gnd single_level_column_mux_0
XXMUX123 bl_123 br_123 bl_out_61 br_out_61 sel_1 gnd single_level_column_mux_0
XXMUX124 bl_124 br_124 bl_out_62 br_out_62 sel_0 gnd single_level_column_mux_0
XXMUX125 bl_125 br_125 bl_out_62 br_out_62 sel_1 gnd single_level_column_mux_0
XXMUX126 bl_126 br_126 bl_out_63 br_out_63 sel_0 gnd single_level_column_mux_0
XXMUX127 bl_127 br_127 bl_out_63 br_out_63 sel_1 gnd single_level_column_mux_0
XXMUX128 bl_128 br_128 bl_out_64 br_out_64 sel_0 gnd single_level_column_mux_0
XXMUX129 bl_129 br_129 bl_out_64 br_out_64 sel_1 gnd single_level_column_mux_0
XXMUX130 bl_130 br_130 bl_out_65 br_out_65 sel_0 gnd single_level_column_mux_0
XXMUX131 bl_131 br_131 bl_out_65 br_out_65 sel_1 gnd single_level_column_mux_0
XXMUX132 bl_132 br_132 bl_out_66 br_out_66 sel_0 gnd single_level_column_mux_0
XXMUX133 bl_133 br_133 bl_out_66 br_out_66 sel_1 gnd single_level_column_mux_0
XXMUX134 bl_134 br_134 bl_out_67 br_out_67 sel_0 gnd single_level_column_mux_0
XXMUX135 bl_135 br_135 bl_out_67 br_out_67 sel_1 gnd single_level_column_mux_0
XXMUX136 bl_136 br_136 bl_out_68 br_out_68 sel_0 gnd single_level_column_mux_0
XXMUX137 bl_137 br_137 bl_out_68 br_out_68 sel_1 gnd single_level_column_mux_0
XXMUX138 bl_138 br_138 bl_out_69 br_out_69 sel_0 gnd single_level_column_mux_0
XXMUX139 bl_139 br_139 bl_out_69 br_out_69 sel_1 gnd single_level_column_mux_0
XXMUX140 bl_140 br_140 bl_out_70 br_out_70 sel_0 gnd single_level_column_mux_0
XXMUX141 bl_141 br_141 bl_out_70 br_out_70 sel_1 gnd single_level_column_mux_0
XXMUX142 bl_142 br_142 bl_out_71 br_out_71 sel_0 gnd single_level_column_mux_0
XXMUX143 bl_143 br_143 bl_out_71 br_out_71 sel_1 gnd single_level_column_mux_0
XXMUX144 bl_144 br_144 bl_out_72 br_out_72 sel_0 gnd single_level_column_mux_0
XXMUX145 bl_145 br_145 bl_out_72 br_out_72 sel_1 gnd single_level_column_mux_0
XXMUX146 bl_146 br_146 bl_out_73 br_out_73 sel_0 gnd single_level_column_mux_0
XXMUX147 bl_147 br_147 bl_out_73 br_out_73 sel_1 gnd single_level_column_mux_0
XXMUX148 bl_148 br_148 bl_out_74 br_out_74 sel_0 gnd single_level_column_mux_0
XXMUX149 bl_149 br_149 bl_out_74 br_out_74 sel_1 gnd single_level_column_mux_0
XXMUX150 bl_150 br_150 bl_out_75 br_out_75 sel_0 gnd single_level_column_mux_0
XXMUX151 bl_151 br_151 bl_out_75 br_out_75 sel_1 gnd single_level_column_mux_0
XXMUX152 bl_152 br_152 bl_out_76 br_out_76 sel_0 gnd single_level_column_mux_0
XXMUX153 bl_153 br_153 bl_out_76 br_out_76 sel_1 gnd single_level_column_mux_0
XXMUX154 bl_154 br_154 bl_out_77 br_out_77 sel_0 gnd single_level_column_mux_0
XXMUX155 bl_155 br_155 bl_out_77 br_out_77 sel_1 gnd single_level_column_mux_0
XXMUX156 bl_156 br_156 bl_out_78 br_out_78 sel_0 gnd single_level_column_mux_0
XXMUX157 bl_157 br_157 bl_out_78 br_out_78 sel_1 gnd single_level_column_mux_0
XXMUX158 bl_158 br_158 bl_out_79 br_out_79 sel_0 gnd single_level_column_mux_0
XXMUX159 bl_159 br_159 bl_out_79 br_out_79 sel_1 gnd single_level_column_mux_0
XXMUX160 bl_160 br_160 bl_out_80 br_out_80 sel_0 gnd single_level_column_mux_0
XXMUX161 bl_161 br_161 bl_out_80 br_out_80 sel_1 gnd single_level_column_mux_0
XXMUX162 bl_162 br_162 bl_out_81 br_out_81 sel_0 gnd single_level_column_mux_0
XXMUX163 bl_163 br_163 bl_out_81 br_out_81 sel_1 gnd single_level_column_mux_0
XXMUX164 bl_164 br_164 bl_out_82 br_out_82 sel_0 gnd single_level_column_mux_0
XXMUX165 bl_165 br_165 bl_out_82 br_out_82 sel_1 gnd single_level_column_mux_0
XXMUX166 bl_166 br_166 bl_out_83 br_out_83 sel_0 gnd single_level_column_mux_0
XXMUX167 bl_167 br_167 bl_out_83 br_out_83 sel_1 gnd single_level_column_mux_0
XXMUX168 bl_168 br_168 bl_out_84 br_out_84 sel_0 gnd single_level_column_mux_0
XXMUX169 bl_169 br_169 bl_out_84 br_out_84 sel_1 gnd single_level_column_mux_0
XXMUX170 bl_170 br_170 bl_out_85 br_out_85 sel_0 gnd single_level_column_mux_0
XXMUX171 bl_171 br_171 bl_out_85 br_out_85 sel_1 gnd single_level_column_mux_0
XXMUX172 bl_172 br_172 bl_out_86 br_out_86 sel_0 gnd single_level_column_mux_0
XXMUX173 bl_173 br_173 bl_out_86 br_out_86 sel_1 gnd single_level_column_mux_0
XXMUX174 bl_174 br_174 bl_out_87 br_out_87 sel_0 gnd single_level_column_mux_0
XXMUX175 bl_175 br_175 bl_out_87 br_out_87 sel_1 gnd single_level_column_mux_0
XXMUX176 bl_176 br_176 bl_out_88 br_out_88 sel_0 gnd single_level_column_mux_0
XXMUX177 bl_177 br_177 bl_out_88 br_out_88 sel_1 gnd single_level_column_mux_0
XXMUX178 bl_178 br_178 bl_out_89 br_out_89 sel_0 gnd single_level_column_mux_0
XXMUX179 bl_179 br_179 bl_out_89 br_out_89 sel_1 gnd single_level_column_mux_0
XXMUX180 bl_180 br_180 bl_out_90 br_out_90 sel_0 gnd single_level_column_mux_0
XXMUX181 bl_181 br_181 bl_out_90 br_out_90 sel_1 gnd single_level_column_mux_0
XXMUX182 bl_182 br_182 bl_out_91 br_out_91 sel_0 gnd single_level_column_mux_0
XXMUX183 bl_183 br_183 bl_out_91 br_out_91 sel_1 gnd single_level_column_mux_0
XXMUX184 bl_184 br_184 bl_out_92 br_out_92 sel_0 gnd single_level_column_mux_0
XXMUX185 bl_185 br_185 bl_out_92 br_out_92 sel_1 gnd single_level_column_mux_0
XXMUX186 bl_186 br_186 bl_out_93 br_out_93 sel_0 gnd single_level_column_mux_0
XXMUX187 bl_187 br_187 bl_out_93 br_out_93 sel_1 gnd single_level_column_mux_0
XXMUX188 bl_188 br_188 bl_out_94 br_out_94 sel_0 gnd single_level_column_mux_0
XXMUX189 bl_189 br_189 bl_out_94 br_out_94 sel_1 gnd single_level_column_mux_0
XXMUX190 bl_190 br_190 bl_out_95 br_out_95 sel_0 gnd single_level_column_mux_0
XXMUX191 bl_191 br_191 bl_out_95 br_out_95 sel_1 gnd single_level_column_mux_0
XXMUX192 bl_192 br_192 bl_out_96 br_out_96 sel_0 gnd single_level_column_mux_0
XXMUX193 bl_193 br_193 bl_out_96 br_out_96 sel_1 gnd single_level_column_mux_0
XXMUX194 bl_194 br_194 bl_out_97 br_out_97 sel_0 gnd single_level_column_mux_0
XXMUX195 bl_195 br_195 bl_out_97 br_out_97 sel_1 gnd single_level_column_mux_0
XXMUX196 bl_196 br_196 bl_out_98 br_out_98 sel_0 gnd single_level_column_mux_0
XXMUX197 bl_197 br_197 bl_out_98 br_out_98 sel_1 gnd single_level_column_mux_0
XXMUX198 bl_198 br_198 bl_out_99 br_out_99 sel_0 gnd single_level_column_mux_0
XXMUX199 bl_199 br_199 bl_out_99 br_out_99 sel_1 gnd single_level_column_mux_0
XXMUX200 bl_200 br_200 bl_out_100 br_out_100 sel_0 gnd single_level_column_mux_0
XXMUX201 bl_201 br_201 bl_out_100 br_out_100 sel_1 gnd single_level_column_mux_0
XXMUX202 bl_202 br_202 bl_out_101 br_out_101 sel_0 gnd single_level_column_mux_0
XXMUX203 bl_203 br_203 bl_out_101 br_out_101 sel_1 gnd single_level_column_mux_0
XXMUX204 bl_204 br_204 bl_out_102 br_out_102 sel_0 gnd single_level_column_mux_0
XXMUX205 bl_205 br_205 bl_out_102 br_out_102 sel_1 gnd single_level_column_mux_0
XXMUX206 bl_206 br_206 bl_out_103 br_out_103 sel_0 gnd single_level_column_mux_0
XXMUX207 bl_207 br_207 bl_out_103 br_out_103 sel_1 gnd single_level_column_mux_0
XXMUX208 bl_208 br_208 bl_out_104 br_out_104 sel_0 gnd single_level_column_mux_0
XXMUX209 bl_209 br_209 bl_out_104 br_out_104 sel_1 gnd single_level_column_mux_0
XXMUX210 bl_210 br_210 bl_out_105 br_out_105 sel_0 gnd single_level_column_mux_0
XXMUX211 bl_211 br_211 bl_out_105 br_out_105 sel_1 gnd single_level_column_mux_0
XXMUX212 bl_212 br_212 bl_out_106 br_out_106 sel_0 gnd single_level_column_mux_0
XXMUX213 bl_213 br_213 bl_out_106 br_out_106 sel_1 gnd single_level_column_mux_0
XXMUX214 bl_214 br_214 bl_out_107 br_out_107 sel_0 gnd single_level_column_mux_0
XXMUX215 bl_215 br_215 bl_out_107 br_out_107 sel_1 gnd single_level_column_mux_0
XXMUX216 bl_216 br_216 bl_out_108 br_out_108 sel_0 gnd single_level_column_mux_0
XXMUX217 bl_217 br_217 bl_out_108 br_out_108 sel_1 gnd single_level_column_mux_0
XXMUX218 bl_218 br_218 bl_out_109 br_out_109 sel_0 gnd single_level_column_mux_0
XXMUX219 bl_219 br_219 bl_out_109 br_out_109 sel_1 gnd single_level_column_mux_0
XXMUX220 bl_220 br_220 bl_out_110 br_out_110 sel_0 gnd single_level_column_mux_0
XXMUX221 bl_221 br_221 bl_out_110 br_out_110 sel_1 gnd single_level_column_mux_0
XXMUX222 bl_222 br_222 bl_out_111 br_out_111 sel_0 gnd single_level_column_mux_0
XXMUX223 bl_223 br_223 bl_out_111 br_out_111 sel_1 gnd single_level_column_mux_0
XXMUX224 bl_224 br_224 bl_out_112 br_out_112 sel_0 gnd single_level_column_mux_0
XXMUX225 bl_225 br_225 bl_out_112 br_out_112 sel_1 gnd single_level_column_mux_0
XXMUX226 bl_226 br_226 bl_out_113 br_out_113 sel_0 gnd single_level_column_mux_0
XXMUX227 bl_227 br_227 bl_out_113 br_out_113 sel_1 gnd single_level_column_mux_0
XXMUX228 bl_228 br_228 bl_out_114 br_out_114 sel_0 gnd single_level_column_mux_0
XXMUX229 bl_229 br_229 bl_out_114 br_out_114 sel_1 gnd single_level_column_mux_0
XXMUX230 bl_230 br_230 bl_out_115 br_out_115 sel_0 gnd single_level_column_mux_0
XXMUX231 bl_231 br_231 bl_out_115 br_out_115 sel_1 gnd single_level_column_mux_0
XXMUX232 bl_232 br_232 bl_out_116 br_out_116 sel_0 gnd single_level_column_mux_0
XXMUX233 bl_233 br_233 bl_out_116 br_out_116 sel_1 gnd single_level_column_mux_0
XXMUX234 bl_234 br_234 bl_out_117 br_out_117 sel_0 gnd single_level_column_mux_0
XXMUX235 bl_235 br_235 bl_out_117 br_out_117 sel_1 gnd single_level_column_mux_0
XXMUX236 bl_236 br_236 bl_out_118 br_out_118 sel_0 gnd single_level_column_mux_0
XXMUX237 bl_237 br_237 bl_out_118 br_out_118 sel_1 gnd single_level_column_mux_0
XXMUX238 bl_238 br_238 bl_out_119 br_out_119 sel_0 gnd single_level_column_mux_0
XXMUX239 bl_239 br_239 bl_out_119 br_out_119 sel_1 gnd single_level_column_mux_0
XXMUX240 bl_240 br_240 bl_out_120 br_out_120 sel_0 gnd single_level_column_mux_0
XXMUX241 bl_241 br_241 bl_out_120 br_out_120 sel_1 gnd single_level_column_mux_0
XXMUX242 bl_242 br_242 bl_out_121 br_out_121 sel_0 gnd single_level_column_mux_0
XXMUX243 bl_243 br_243 bl_out_121 br_out_121 sel_1 gnd single_level_column_mux_0
XXMUX244 bl_244 br_244 bl_out_122 br_out_122 sel_0 gnd single_level_column_mux_0
XXMUX245 bl_245 br_245 bl_out_122 br_out_122 sel_1 gnd single_level_column_mux_0
XXMUX246 bl_246 br_246 bl_out_123 br_out_123 sel_0 gnd single_level_column_mux_0
XXMUX247 bl_247 br_247 bl_out_123 br_out_123 sel_1 gnd single_level_column_mux_0
XXMUX248 bl_248 br_248 bl_out_124 br_out_124 sel_0 gnd single_level_column_mux_0
XXMUX249 bl_249 br_249 bl_out_124 br_out_124 sel_1 gnd single_level_column_mux_0
XXMUX250 bl_250 br_250 bl_out_125 br_out_125 sel_0 gnd single_level_column_mux_0
XXMUX251 bl_251 br_251 bl_out_125 br_out_125 sel_1 gnd single_level_column_mux_0
XXMUX252 bl_252 br_252 bl_out_126 br_out_126 sel_0 gnd single_level_column_mux_0
XXMUX253 bl_253 br_253 bl_out_126 br_out_126 sel_1 gnd single_level_column_mux_0
XXMUX254 bl_254 br_254 bl_out_127 br_out_127 sel_0 gnd single_level_column_mux_0
XXMUX255 bl_255 br_255 bl_out_127 br_out_127 sel_1 gnd single_level_column_mux_0
.ENDS single_level_column_mux_array_0

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT write_driver_array_0 data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9 data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17 data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25 data_26 data_27 data_28 data_29 data_30 data_31 data_32 data_33 data_34 data_35 data_36 data_37 data_38 data_39 data_40 data_41 data_42 data_43 data_44 data_45 data_46 data_47 data_48 data_49 data_50 data_51 data_52 data_53 data_54 data_55 data_56 data_57 data_58 data_59 data_60 data_61 data_62 data_63 data_64 data_65 data_66 data_67 data_68 data_69 data_70 data_71 data_72 data_73 data_74 data_75 data_76 data_77 data_78 data_79 data_80 data_81 data_82 data_83 data_84 data_85 data_86 data_87 data_88 data_89 data_90 data_91 data_92 data_93 data_94 data_95 data_96 data_97 data_98 data_99 data_100 data_101 data_102 data_103 data_104 data_105 data_106 data_107 data_108 data_109 data_110 data_111 data_112 data_113 data_114 data_115 data_116 data_117 data_118 data_119 data_120 data_121 data_122 data_123 data_124 data_125 data_126 data_127 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 en vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* INPUT : data_32 
* INPUT : data_33 
* INPUT : data_34 
* INPUT : data_35 
* INPUT : data_36 
* INPUT : data_37 
* INPUT : data_38 
* INPUT : data_39 
* INPUT : data_40 
* INPUT : data_41 
* INPUT : data_42 
* INPUT : data_43 
* INPUT : data_44 
* INPUT : data_45 
* INPUT : data_46 
* INPUT : data_47 
* INPUT : data_48 
* INPUT : data_49 
* INPUT : data_50 
* INPUT : data_51 
* INPUT : data_52 
* INPUT : data_53 
* INPUT : data_54 
* INPUT : data_55 
* INPUT : data_56 
* INPUT : data_57 
* INPUT : data_58 
* INPUT : data_59 
* INPUT : data_60 
* INPUT : data_61 
* INPUT : data_62 
* INPUT : data_63 
* INPUT : data_64 
* INPUT : data_65 
* INPUT : data_66 
* INPUT : data_67 
* INPUT : data_68 
* INPUT : data_69 
* INPUT : data_70 
* INPUT : data_71 
* INPUT : data_72 
* INPUT : data_73 
* INPUT : data_74 
* INPUT : data_75 
* INPUT : data_76 
* INPUT : data_77 
* INPUT : data_78 
* INPUT : data_79 
* INPUT : data_80 
* INPUT : data_81 
* INPUT : data_82 
* INPUT : data_83 
* INPUT : data_84 
* INPUT : data_85 
* INPUT : data_86 
* INPUT : data_87 
* INPUT : data_88 
* INPUT : data_89 
* INPUT : data_90 
* INPUT : data_91 
* INPUT : data_92 
* INPUT : data_93 
* INPUT : data_94 
* INPUT : data_95 
* INPUT : data_96 
* INPUT : data_97 
* INPUT : data_98 
* INPUT : data_99 
* INPUT : data_100 
* INPUT : data_101 
* INPUT : data_102 
* INPUT : data_103 
* INPUT : data_104 
* INPUT : data_105 
* INPUT : data_106 
* INPUT : data_107 
* INPUT : data_108 
* INPUT : data_109 
* INPUT : data_110 
* INPUT : data_111 
* INPUT : data_112 
* INPUT : data_113 
* INPUT : data_114 
* INPUT : data_115 
* INPUT : data_116 
* INPUT : data_117 
* INPUT : data_118 
* INPUT : data_119 
* INPUT : data_120 
* INPUT : data_121 
* INPUT : data_122 
* INPUT : data_123 
* INPUT : data_124 
* INPUT : data_125 
* INPUT : data_126 
* INPUT : data_127 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 128
Xwrite_driver0 data_0 bl_0 br_0 en vdd gnd write_driver
Xwrite_driver2 data_1 bl_1 br_1 en vdd gnd write_driver
Xwrite_driver4 data_2 bl_2 br_2 en vdd gnd write_driver
Xwrite_driver6 data_3 bl_3 br_3 en vdd gnd write_driver
Xwrite_driver8 data_4 bl_4 br_4 en vdd gnd write_driver
Xwrite_driver10 data_5 bl_5 br_5 en vdd gnd write_driver
Xwrite_driver12 data_6 bl_6 br_6 en vdd gnd write_driver
Xwrite_driver14 data_7 bl_7 br_7 en vdd gnd write_driver
Xwrite_driver16 data_8 bl_8 br_8 en vdd gnd write_driver
Xwrite_driver18 data_9 bl_9 br_9 en vdd gnd write_driver
Xwrite_driver20 data_10 bl_10 br_10 en vdd gnd write_driver
Xwrite_driver22 data_11 bl_11 br_11 en vdd gnd write_driver
Xwrite_driver24 data_12 bl_12 br_12 en vdd gnd write_driver
Xwrite_driver26 data_13 bl_13 br_13 en vdd gnd write_driver
Xwrite_driver28 data_14 bl_14 br_14 en vdd gnd write_driver
Xwrite_driver30 data_15 bl_15 br_15 en vdd gnd write_driver
Xwrite_driver32 data_16 bl_16 br_16 en vdd gnd write_driver
Xwrite_driver34 data_17 bl_17 br_17 en vdd gnd write_driver
Xwrite_driver36 data_18 bl_18 br_18 en vdd gnd write_driver
Xwrite_driver38 data_19 bl_19 br_19 en vdd gnd write_driver
Xwrite_driver40 data_20 bl_20 br_20 en vdd gnd write_driver
Xwrite_driver42 data_21 bl_21 br_21 en vdd gnd write_driver
Xwrite_driver44 data_22 bl_22 br_22 en vdd gnd write_driver
Xwrite_driver46 data_23 bl_23 br_23 en vdd gnd write_driver
Xwrite_driver48 data_24 bl_24 br_24 en vdd gnd write_driver
Xwrite_driver50 data_25 bl_25 br_25 en vdd gnd write_driver
Xwrite_driver52 data_26 bl_26 br_26 en vdd gnd write_driver
Xwrite_driver54 data_27 bl_27 br_27 en vdd gnd write_driver
Xwrite_driver56 data_28 bl_28 br_28 en vdd gnd write_driver
Xwrite_driver58 data_29 bl_29 br_29 en vdd gnd write_driver
Xwrite_driver60 data_30 bl_30 br_30 en vdd gnd write_driver
Xwrite_driver62 data_31 bl_31 br_31 en vdd gnd write_driver
Xwrite_driver64 data_32 bl_32 br_32 en vdd gnd write_driver
Xwrite_driver66 data_33 bl_33 br_33 en vdd gnd write_driver
Xwrite_driver68 data_34 bl_34 br_34 en vdd gnd write_driver
Xwrite_driver70 data_35 bl_35 br_35 en vdd gnd write_driver
Xwrite_driver72 data_36 bl_36 br_36 en vdd gnd write_driver
Xwrite_driver74 data_37 bl_37 br_37 en vdd gnd write_driver
Xwrite_driver76 data_38 bl_38 br_38 en vdd gnd write_driver
Xwrite_driver78 data_39 bl_39 br_39 en vdd gnd write_driver
Xwrite_driver80 data_40 bl_40 br_40 en vdd gnd write_driver
Xwrite_driver82 data_41 bl_41 br_41 en vdd gnd write_driver
Xwrite_driver84 data_42 bl_42 br_42 en vdd gnd write_driver
Xwrite_driver86 data_43 bl_43 br_43 en vdd gnd write_driver
Xwrite_driver88 data_44 bl_44 br_44 en vdd gnd write_driver
Xwrite_driver90 data_45 bl_45 br_45 en vdd gnd write_driver
Xwrite_driver92 data_46 bl_46 br_46 en vdd gnd write_driver
Xwrite_driver94 data_47 bl_47 br_47 en vdd gnd write_driver
Xwrite_driver96 data_48 bl_48 br_48 en vdd gnd write_driver
Xwrite_driver98 data_49 bl_49 br_49 en vdd gnd write_driver
Xwrite_driver100 data_50 bl_50 br_50 en vdd gnd write_driver
Xwrite_driver102 data_51 bl_51 br_51 en vdd gnd write_driver
Xwrite_driver104 data_52 bl_52 br_52 en vdd gnd write_driver
Xwrite_driver106 data_53 bl_53 br_53 en vdd gnd write_driver
Xwrite_driver108 data_54 bl_54 br_54 en vdd gnd write_driver
Xwrite_driver110 data_55 bl_55 br_55 en vdd gnd write_driver
Xwrite_driver112 data_56 bl_56 br_56 en vdd gnd write_driver
Xwrite_driver114 data_57 bl_57 br_57 en vdd gnd write_driver
Xwrite_driver116 data_58 bl_58 br_58 en vdd gnd write_driver
Xwrite_driver118 data_59 bl_59 br_59 en vdd gnd write_driver
Xwrite_driver120 data_60 bl_60 br_60 en vdd gnd write_driver
Xwrite_driver122 data_61 bl_61 br_61 en vdd gnd write_driver
Xwrite_driver124 data_62 bl_62 br_62 en vdd gnd write_driver
Xwrite_driver126 data_63 bl_63 br_63 en vdd gnd write_driver
Xwrite_driver128 data_64 bl_64 br_64 en vdd gnd write_driver
Xwrite_driver130 data_65 bl_65 br_65 en vdd gnd write_driver
Xwrite_driver132 data_66 bl_66 br_66 en vdd gnd write_driver
Xwrite_driver134 data_67 bl_67 br_67 en vdd gnd write_driver
Xwrite_driver136 data_68 bl_68 br_68 en vdd gnd write_driver
Xwrite_driver138 data_69 bl_69 br_69 en vdd gnd write_driver
Xwrite_driver140 data_70 bl_70 br_70 en vdd gnd write_driver
Xwrite_driver142 data_71 bl_71 br_71 en vdd gnd write_driver
Xwrite_driver144 data_72 bl_72 br_72 en vdd gnd write_driver
Xwrite_driver146 data_73 bl_73 br_73 en vdd gnd write_driver
Xwrite_driver148 data_74 bl_74 br_74 en vdd gnd write_driver
Xwrite_driver150 data_75 bl_75 br_75 en vdd gnd write_driver
Xwrite_driver152 data_76 bl_76 br_76 en vdd gnd write_driver
Xwrite_driver154 data_77 bl_77 br_77 en vdd gnd write_driver
Xwrite_driver156 data_78 bl_78 br_78 en vdd gnd write_driver
Xwrite_driver158 data_79 bl_79 br_79 en vdd gnd write_driver
Xwrite_driver160 data_80 bl_80 br_80 en vdd gnd write_driver
Xwrite_driver162 data_81 bl_81 br_81 en vdd gnd write_driver
Xwrite_driver164 data_82 bl_82 br_82 en vdd gnd write_driver
Xwrite_driver166 data_83 bl_83 br_83 en vdd gnd write_driver
Xwrite_driver168 data_84 bl_84 br_84 en vdd gnd write_driver
Xwrite_driver170 data_85 bl_85 br_85 en vdd gnd write_driver
Xwrite_driver172 data_86 bl_86 br_86 en vdd gnd write_driver
Xwrite_driver174 data_87 bl_87 br_87 en vdd gnd write_driver
Xwrite_driver176 data_88 bl_88 br_88 en vdd gnd write_driver
Xwrite_driver178 data_89 bl_89 br_89 en vdd gnd write_driver
Xwrite_driver180 data_90 bl_90 br_90 en vdd gnd write_driver
Xwrite_driver182 data_91 bl_91 br_91 en vdd gnd write_driver
Xwrite_driver184 data_92 bl_92 br_92 en vdd gnd write_driver
Xwrite_driver186 data_93 bl_93 br_93 en vdd gnd write_driver
Xwrite_driver188 data_94 bl_94 br_94 en vdd gnd write_driver
Xwrite_driver190 data_95 bl_95 br_95 en vdd gnd write_driver
Xwrite_driver192 data_96 bl_96 br_96 en vdd gnd write_driver
Xwrite_driver194 data_97 bl_97 br_97 en vdd gnd write_driver
Xwrite_driver196 data_98 bl_98 br_98 en vdd gnd write_driver
Xwrite_driver198 data_99 bl_99 br_99 en vdd gnd write_driver
Xwrite_driver200 data_100 bl_100 br_100 en vdd gnd write_driver
Xwrite_driver202 data_101 bl_101 br_101 en vdd gnd write_driver
Xwrite_driver204 data_102 bl_102 br_102 en vdd gnd write_driver
Xwrite_driver206 data_103 bl_103 br_103 en vdd gnd write_driver
Xwrite_driver208 data_104 bl_104 br_104 en vdd gnd write_driver
Xwrite_driver210 data_105 bl_105 br_105 en vdd gnd write_driver
Xwrite_driver212 data_106 bl_106 br_106 en vdd gnd write_driver
Xwrite_driver214 data_107 bl_107 br_107 en vdd gnd write_driver
Xwrite_driver216 data_108 bl_108 br_108 en vdd gnd write_driver
Xwrite_driver218 data_109 bl_109 br_109 en vdd gnd write_driver
Xwrite_driver220 data_110 bl_110 br_110 en vdd gnd write_driver
Xwrite_driver222 data_111 bl_111 br_111 en vdd gnd write_driver
Xwrite_driver224 data_112 bl_112 br_112 en vdd gnd write_driver
Xwrite_driver226 data_113 bl_113 br_113 en vdd gnd write_driver
Xwrite_driver228 data_114 bl_114 br_114 en vdd gnd write_driver
Xwrite_driver230 data_115 bl_115 br_115 en vdd gnd write_driver
Xwrite_driver232 data_116 bl_116 br_116 en vdd gnd write_driver
Xwrite_driver234 data_117 bl_117 br_117 en vdd gnd write_driver
Xwrite_driver236 data_118 bl_118 br_118 en vdd gnd write_driver
Xwrite_driver238 data_119 bl_119 br_119 en vdd gnd write_driver
Xwrite_driver240 data_120 bl_120 br_120 en vdd gnd write_driver
Xwrite_driver242 data_121 bl_121 br_121 en vdd gnd write_driver
Xwrite_driver244 data_122 bl_122 br_122 en vdd gnd write_driver
Xwrite_driver246 data_123 bl_123 br_123 en vdd gnd write_driver
Xwrite_driver248 data_124 bl_124 br_124 en vdd gnd write_driver
Xwrite_driver250 data_125 bl_125 br_125 en vdd gnd write_driver
Xwrite_driver252 data_126 bl_126 br_126 en vdd gnd write_driver
Xwrite_driver254 data_127 bl_127 br_127 en vdd gnd write_driver
.ENDS write_driver_array_0

.SUBCKT port_data_0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 dout_32 dout_33 dout_34 dout_35 dout_36 dout_37 dout_38 dout_39 dout_40 dout_41 dout_42 dout_43 dout_44 dout_45 dout_46 dout_47 dout_48 dout_49 dout_50 dout_51 dout_52 dout_53 dout_54 dout_55 dout_56 dout_57 dout_58 dout_59 dout_60 dout_61 dout_62 dout_63 dout_64 dout_65 dout_66 dout_67 dout_68 dout_69 dout_70 dout_71 dout_72 dout_73 dout_74 dout_75 dout_76 dout_77 dout_78 dout_79 dout_80 dout_81 dout_82 dout_83 dout_84 dout_85 dout_86 dout_87 dout_88 dout_89 dout_90 dout_91 dout_92 dout_93 dout_94 dout_95 dout_96 dout_97 dout_98 dout_99 dout_100 dout_101 dout_102 dout_103 dout_104 dout_105 dout_106 dout_107 dout_108 dout_109 dout_110 dout_111 dout_112 dout_113 dout_114 dout_115 dout_116 dout_117 dout_118 dout_119 dout_120 dout_121 dout_122 dout_123 dout_124 dout_125 dout_126 dout_127 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 sel_0 sel_1 s_en p_en_bar w_en vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* OUTPUT: dout_32 
* OUTPUT: dout_33 
* OUTPUT: dout_34 
* OUTPUT: dout_35 
* OUTPUT: dout_36 
* OUTPUT: dout_37 
* OUTPUT: dout_38 
* OUTPUT: dout_39 
* OUTPUT: dout_40 
* OUTPUT: dout_41 
* OUTPUT: dout_42 
* OUTPUT: dout_43 
* OUTPUT: dout_44 
* OUTPUT: dout_45 
* OUTPUT: dout_46 
* OUTPUT: dout_47 
* OUTPUT: dout_48 
* OUTPUT: dout_49 
* OUTPUT: dout_50 
* OUTPUT: dout_51 
* OUTPUT: dout_52 
* OUTPUT: dout_53 
* OUTPUT: dout_54 
* OUTPUT: dout_55 
* OUTPUT: dout_56 
* OUTPUT: dout_57 
* OUTPUT: dout_58 
* OUTPUT: dout_59 
* OUTPUT: dout_60 
* OUTPUT: dout_61 
* OUTPUT: dout_62 
* OUTPUT: dout_63 
* OUTPUT: dout_64 
* OUTPUT: dout_65 
* OUTPUT: dout_66 
* OUTPUT: dout_67 
* OUTPUT: dout_68 
* OUTPUT: dout_69 
* OUTPUT: dout_70 
* OUTPUT: dout_71 
* OUTPUT: dout_72 
* OUTPUT: dout_73 
* OUTPUT: dout_74 
* OUTPUT: dout_75 
* OUTPUT: dout_76 
* OUTPUT: dout_77 
* OUTPUT: dout_78 
* OUTPUT: dout_79 
* OUTPUT: dout_80 
* OUTPUT: dout_81 
* OUTPUT: dout_82 
* OUTPUT: dout_83 
* OUTPUT: dout_84 
* OUTPUT: dout_85 
* OUTPUT: dout_86 
* OUTPUT: dout_87 
* OUTPUT: dout_88 
* OUTPUT: dout_89 
* OUTPUT: dout_90 
* OUTPUT: dout_91 
* OUTPUT: dout_92 
* OUTPUT: dout_93 
* OUTPUT: dout_94 
* OUTPUT: dout_95 
* OUTPUT: dout_96 
* OUTPUT: dout_97 
* OUTPUT: dout_98 
* OUTPUT: dout_99 
* OUTPUT: dout_100 
* OUTPUT: dout_101 
* OUTPUT: dout_102 
* OUTPUT: dout_103 
* OUTPUT: dout_104 
* OUTPUT: dout_105 
* OUTPUT: dout_106 
* OUTPUT: dout_107 
* OUTPUT: dout_108 
* OUTPUT: dout_109 
* OUTPUT: dout_110 
* OUTPUT: dout_111 
* OUTPUT: dout_112 
* OUTPUT: dout_113 
* OUTPUT: dout_114 
* OUTPUT: dout_115 
* OUTPUT: dout_116 
* OUTPUT: dout_117 
* OUTPUT: dout_118 
* OUTPUT: dout_119 
* OUTPUT: dout_120 
* OUTPUT: dout_121 
* OUTPUT: dout_122 
* OUTPUT: dout_123 
* OUTPUT: dout_124 
* OUTPUT: dout_125 
* OUTPUT: dout_126 
* OUTPUT: dout_127 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : din_32 
* INPUT : din_33 
* INPUT : din_34 
* INPUT : din_35 
* INPUT : din_36 
* INPUT : din_37 
* INPUT : din_38 
* INPUT : din_39 
* INPUT : din_40 
* INPUT : din_41 
* INPUT : din_42 
* INPUT : din_43 
* INPUT : din_44 
* INPUT : din_45 
* INPUT : din_46 
* INPUT : din_47 
* INPUT : din_48 
* INPUT : din_49 
* INPUT : din_50 
* INPUT : din_51 
* INPUT : din_52 
* INPUT : din_53 
* INPUT : din_54 
* INPUT : din_55 
* INPUT : din_56 
* INPUT : din_57 
* INPUT : din_58 
* INPUT : din_59 
* INPUT : din_60 
* INPUT : din_61 
* INPUT : din_62 
* INPUT : din_63 
* INPUT : din_64 
* INPUT : din_65 
* INPUT : din_66 
* INPUT : din_67 
* INPUT : din_68 
* INPUT : din_69 
* INPUT : din_70 
* INPUT : din_71 
* INPUT : din_72 
* INPUT : din_73 
* INPUT : din_74 
* INPUT : din_75 
* INPUT : din_76 
* INPUT : din_77 
* INPUT : din_78 
* INPUT : din_79 
* INPUT : din_80 
* INPUT : din_81 
* INPUT : din_82 
* INPUT : din_83 
* INPUT : din_84 
* INPUT : din_85 
* INPUT : din_86 
* INPUT : din_87 
* INPUT : din_88 
* INPUT : din_89 
* INPUT : din_90 
* INPUT : din_91 
* INPUT : din_92 
* INPUT : din_93 
* INPUT : din_94 
* INPUT : din_95 
* INPUT : din_96 
* INPUT : din_97 
* INPUT : din_98 
* INPUT : din_99 
* INPUT : din_100 
* INPUT : din_101 
* INPUT : din_102 
* INPUT : din_103 
* INPUT : din_104 
* INPUT : din_105 
* INPUT : din_106 
* INPUT : din_107 
* INPUT : din_108 
* INPUT : din_109 
* INPUT : din_110 
* INPUT : din_111 
* INPUT : din_112 
* INPUT : din_113 
* INPUT : din_114 
* INPUT : din_115 
* INPUT : din_116 
* INPUT : din_117 
* INPUT : din_118 
* INPUT : din_119 
* INPUT : din_120 
* INPUT : din_121 
* INPUT : din_122 
* INPUT : din_123 
* INPUT : din_124 
* INPUT : din_125 
* INPUT : din_126 
* INPUT : din_127 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 p_en_bar vdd precharge_array_0
Xsense_amp_array0 dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2 br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5 bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7 dout_8 bl_out_8 br_out_8 dout_9 bl_out_9 br_out_9 dout_10 bl_out_10 br_out_10 dout_11 bl_out_11 br_out_11 dout_12 bl_out_12 br_out_12 dout_13 bl_out_13 br_out_13 dout_14 bl_out_14 br_out_14 dout_15 bl_out_15 br_out_15 dout_16 bl_out_16 br_out_16 dout_17 bl_out_17 br_out_17 dout_18 bl_out_18 br_out_18 dout_19 bl_out_19 br_out_19 dout_20 bl_out_20 br_out_20 dout_21 bl_out_21 br_out_21 dout_22 bl_out_22 br_out_22 dout_23 bl_out_23 br_out_23 dout_24 bl_out_24 br_out_24 dout_25 bl_out_25 br_out_25 dout_26 bl_out_26 br_out_26 dout_27 bl_out_27 br_out_27 dout_28 bl_out_28 br_out_28 dout_29 bl_out_29 br_out_29 dout_30 bl_out_30 br_out_30 dout_31 bl_out_31 br_out_31 dout_32 bl_out_32 br_out_32 dout_33 bl_out_33 br_out_33 dout_34 bl_out_34 br_out_34 dout_35 bl_out_35 br_out_35 dout_36 bl_out_36 br_out_36 dout_37 bl_out_37 br_out_37 dout_38 bl_out_38 br_out_38 dout_39 bl_out_39 br_out_39 dout_40 bl_out_40 br_out_40 dout_41 bl_out_41 br_out_41 dout_42 bl_out_42 br_out_42 dout_43 bl_out_43 br_out_43 dout_44 bl_out_44 br_out_44 dout_45 bl_out_45 br_out_45 dout_46 bl_out_46 br_out_46 dout_47 bl_out_47 br_out_47 dout_48 bl_out_48 br_out_48 dout_49 bl_out_49 br_out_49 dout_50 bl_out_50 br_out_50 dout_51 bl_out_51 br_out_51 dout_52 bl_out_52 br_out_52 dout_53 bl_out_53 br_out_53 dout_54 bl_out_54 br_out_54 dout_55 bl_out_55 br_out_55 dout_56 bl_out_56 br_out_56 dout_57 bl_out_57 br_out_57 dout_58 bl_out_58 br_out_58 dout_59 bl_out_59 br_out_59 dout_60 bl_out_60 br_out_60 dout_61 bl_out_61 br_out_61 dout_62 bl_out_62 br_out_62 dout_63 bl_out_63 br_out_63 dout_64 bl_out_64 br_out_64 dout_65 bl_out_65 br_out_65 dout_66 bl_out_66 br_out_66 dout_67 bl_out_67 br_out_67 dout_68 bl_out_68 br_out_68 dout_69 bl_out_69 br_out_69 dout_70 bl_out_70 br_out_70 dout_71 bl_out_71 br_out_71 dout_72 bl_out_72 br_out_72 dout_73 bl_out_73 br_out_73 dout_74 bl_out_74 br_out_74 dout_75 bl_out_75 br_out_75 dout_76 bl_out_76 br_out_76 dout_77 bl_out_77 br_out_77 dout_78 bl_out_78 br_out_78 dout_79 bl_out_79 br_out_79 dout_80 bl_out_80 br_out_80 dout_81 bl_out_81 br_out_81 dout_82 bl_out_82 br_out_82 dout_83 bl_out_83 br_out_83 dout_84 bl_out_84 br_out_84 dout_85 bl_out_85 br_out_85 dout_86 bl_out_86 br_out_86 dout_87 bl_out_87 br_out_87 dout_88 bl_out_88 br_out_88 dout_89 bl_out_89 br_out_89 dout_90 bl_out_90 br_out_90 dout_91 bl_out_91 br_out_91 dout_92 bl_out_92 br_out_92 dout_93 bl_out_93 br_out_93 dout_94 bl_out_94 br_out_94 dout_95 bl_out_95 br_out_95 dout_96 bl_out_96 br_out_96 dout_97 bl_out_97 br_out_97 dout_98 bl_out_98 br_out_98 dout_99 bl_out_99 br_out_99 dout_100 bl_out_100 br_out_100 dout_101 bl_out_101 br_out_101 dout_102 bl_out_102 br_out_102 dout_103 bl_out_103 br_out_103 dout_104 bl_out_104 br_out_104 dout_105 bl_out_105 br_out_105 dout_106 bl_out_106 br_out_106 dout_107 bl_out_107 br_out_107 dout_108 bl_out_108 br_out_108 dout_109 bl_out_109 br_out_109 dout_110 bl_out_110 br_out_110 dout_111 bl_out_111 br_out_111 dout_112 bl_out_112 br_out_112 dout_113 bl_out_113 br_out_113 dout_114 bl_out_114 br_out_114 dout_115 bl_out_115 br_out_115 dout_116 bl_out_116 br_out_116 dout_117 bl_out_117 br_out_117 dout_118 bl_out_118 br_out_118 dout_119 bl_out_119 br_out_119 dout_120 bl_out_120 br_out_120 dout_121 bl_out_121 br_out_121 dout_122 bl_out_122 br_out_122 dout_123 bl_out_123 br_out_123 dout_124 bl_out_124 br_out_124 dout_125 bl_out_125 br_out_125 dout_126 bl_out_126 br_out_126 dout_127 bl_out_127 br_out_127 s_en vdd gnd sense_amp_array_0
Xwrite_driver_array0 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 din_32 din_33 din_34 din_35 din_36 din_37 din_38 din_39 din_40 din_41 din_42 din_43 din_44 din_45 din_46 din_47 din_48 din_49 din_50 din_51 din_52 din_53 din_54 din_55 din_56 din_57 din_58 din_59 din_60 din_61 din_62 din_63 din_64 din_65 din_66 din_67 din_68 din_69 din_70 din_71 din_72 din_73 din_74 din_75 din_76 din_77 din_78 din_79 din_80 din_81 din_82 din_83 din_84 din_85 din_86 din_87 din_88 din_89 din_90 din_91 din_92 din_93 din_94 din_95 din_96 din_97 din_98 din_99 din_100 din_101 din_102 din_103 din_104 din_105 din_106 din_107 din_108 din_109 din_110 din_111 din_112 din_113 din_114 din_115 din_116 din_117 din_118 din_119 din_120 din_121 din_122 din_123 din_124 din_125 din_126 din_127 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 bl_out_32 br_out_32 bl_out_33 br_out_33 bl_out_34 br_out_34 bl_out_35 br_out_35 bl_out_36 br_out_36 bl_out_37 br_out_37 bl_out_38 br_out_38 bl_out_39 br_out_39 bl_out_40 br_out_40 bl_out_41 br_out_41 bl_out_42 br_out_42 bl_out_43 br_out_43 bl_out_44 br_out_44 bl_out_45 br_out_45 bl_out_46 br_out_46 bl_out_47 br_out_47 bl_out_48 br_out_48 bl_out_49 br_out_49 bl_out_50 br_out_50 bl_out_51 br_out_51 bl_out_52 br_out_52 bl_out_53 br_out_53 bl_out_54 br_out_54 bl_out_55 br_out_55 bl_out_56 br_out_56 bl_out_57 br_out_57 bl_out_58 br_out_58 bl_out_59 br_out_59 bl_out_60 br_out_60 bl_out_61 br_out_61 bl_out_62 br_out_62 bl_out_63 br_out_63 bl_out_64 br_out_64 bl_out_65 br_out_65 bl_out_66 br_out_66 bl_out_67 br_out_67 bl_out_68 br_out_68 bl_out_69 br_out_69 bl_out_70 br_out_70 bl_out_71 br_out_71 bl_out_72 br_out_72 bl_out_73 br_out_73 bl_out_74 br_out_74 bl_out_75 br_out_75 bl_out_76 br_out_76 bl_out_77 br_out_77 bl_out_78 br_out_78 bl_out_79 br_out_79 bl_out_80 br_out_80 bl_out_81 br_out_81 bl_out_82 br_out_82 bl_out_83 br_out_83 bl_out_84 br_out_84 bl_out_85 br_out_85 bl_out_86 br_out_86 bl_out_87 br_out_87 bl_out_88 br_out_88 bl_out_89 br_out_89 bl_out_90 br_out_90 bl_out_91 br_out_91 bl_out_92 br_out_92 bl_out_93 br_out_93 bl_out_94 br_out_94 bl_out_95 br_out_95 bl_out_96 br_out_96 bl_out_97 br_out_97 bl_out_98 br_out_98 bl_out_99 br_out_99 bl_out_100 br_out_100 bl_out_101 br_out_101 bl_out_102 br_out_102 bl_out_103 br_out_103 bl_out_104 br_out_104 bl_out_105 br_out_105 bl_out_106 br_out_106 bl_out_107 br_out_107 bl_out_108 br_out_108 bl_out_109 br_out_109 bl_out_110 br_out_110 bl_out_111 br_out_111 bl_out_112 br_out_112 bl_out_113 br_out_113 bl_out_114 br_out_114 bl_out_115 br_out_115 bl_out_116 br_out_116 bl_out_117 br_out_117 bl_out_118 br_out_118 bl_out_119 br_out_119 bl_out_120 br_out_120 bl_out_121 br_out_121 bl_out_122 br_out_122 bl_out_123 br_out_123 bl_out_124 br_out_124 bl_out_125 br_out_125 bl_out_126 br_out_126 bl_out_127 br_out_127 w_en vdd gnd write_driver_array_0
Xcolumn_mux_array0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 sel_0 sel_1 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 bl_out_32 br_out_32 bl_out_33 br_out_33 bl_out_34 br_out_34 bl_out_35 br_out_35 bl_out_36 br_out_36 bl_out_37 br_out_37 bl_out_38 br_out_38 bl_out_39 br_out_39 bl_out_40 br_out_40 bl_out_41 br_out_41 bl_out_42 br_out_42 bl_out_43 br_out_43 bl_out_44 br_out_44 bl_out_45 br_out_45 bl_out_46 br_out_46 bl_out_47 br_out_47 bl_out_48 br_out_48 bl_out_49 br_out_49 bl_out_50 br_out_50 bl_out_51 br_out_51 bl_out_52 br_out_52 bl_out_53 br_out_53 bl_out_54 br_out_54 bl_out_55 br_out_55 bl_out_56 br_out_56 bl_out_57 br_out_57 bl_out_58 br_out_58 bl_out_59 br_out_59 bl_out_60 br_out_60 bl_out_61 br_out_61 bl_out_62 br_out_62 bl_out_63 br_out_63 bl_out_64 br_out_64 bl_out_65 br_out_65 bl_out_66 br_out_66 bl_out_67 br_out_67 bl_out_68 br_out_68 bl_out_69 br_out_69 bl_out_70 br_out_70 bl_out_71 br_out_71 bl_out_72 br_out_72 bl_out_73 br_out_73 bl_out_74 br_out_74 bl_out_75 br_out_75 bl_out_76 br_out_76 bl_out_77 br_out_77 bl_out_78 br_out_78 bl_out_79 br_out_79 bl_out_80 br_out_80 bl_out_81 br_out_81 bl_out_82 br_out_82 bl_out_83 br_out_83 bl_out_84 br_out_84 bl_out_85 br_out_85 bl_out_86 br_out_86 bl_out_87 br_out_87 bl_out_88 br_out_88 bl_out_89 br_out_89 bl_out_90 br_out_90 bl_out_91 br_out_91 bl_out_92 br_out_92 bl_out_93 br_out_93 bl_out_94 br_out_94 bl_out_95 br_out_95 bl_out_96 br_out_96 bl_out_97 br_out_97 bl_out_98 br_out_98 bl_out_99 br_out_99 bl_out_100 br_out_100 bl_out_101 br_out_101 bl_out_102 br_out_102 bl_out_103 br_out_103 bl_out_104 br_out_104 bl_out_105 br_out_105 bl_out_106 br_out_106 bl_out_107 br_out_107 bl_out_108 br_out_108 bl_out_109 br_out_109 bl_out_110 br_out_110 bl_out_111 br_out_111 bl_out_112 br_out_112 bl_out_113 br_out_113 bl_out_114 br_out_114 bl_out_115 br_out_115 bl_out_116 br_out_116 bl_out_117 br_out_117 bl_out_118 br_out_118 bl_out_119 br_out_119 bl_out_120 br_out_120 bl_out_121 br_out_121 bl_out_122 br_out_122 bl_out_123 br_out_123 bl_out_124 br_out_124 bl_out_125 br_out_125 bl_out_126 br_out_126 bl_out_127 br_out_127 gnd single_level_column_mux_array_0
.ENDS port_data_0

* ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_0

* ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT pnand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_0

.SUBCKT pnand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_0

.SUBCKT hierarchical_predecode2x4_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
XXpre2x4_nand_0 inbar_0 inbar_1 Z_0 vdd gnd pnand2_0
XXpre2x4_nand_1 in_0 inbar_1 Z_1 vdd gnd pnand2_0
XXpre2x4_nand_2 inbar_0 in_1 Z_2 vdd gnd pnand2_0
XXpre2x4_nand_3 in_0 in_1 Z_3 vdd gnd pnand2_0
.ENDS hierarchical_predecode2x4_0

.SUBCKT hierarchical_predecode3x8_0 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
Xpre_nand_inv_4 Z_4 out_4 vdd gnd pinv_0
Xpre_nand_inv_5 Z_5 out_5 vdd gnd pinv_0
Xpre_nand_inv_6 Z_6 out_6 vdd gnd pinv_0
Xpre_nand_inv_7 Z_7 out_7 vdd gnd pinv_0
XXpre3x8_nand_0 inbar_0 inbar_1 inbar_2 Z_0 vdd gnd pnand3_0
XXpre3x8_nand_1 in_0 inbar_1 inbar_2 Z_1 vdd gnd pnand3_0
XXpre3x8_nand_2 inbar_0 in_1 inbar_2 Z_2 vdd gnd pnand3_0
XXpre3x8_nand_3 in_0 in_1 inbar_2 Z_3 vdd gnd pnand3_0
XXpre3x8_nand_4 inbar_0 inbar_1 in_2 Z_4 vdd gnd pnand3_0
XXpre3x8_nand_5 in_0 inbar_1 in_2 Z_5 vdd gnd pnand3_0
XXpre3x8_nand_6 inbar_0 in_1 in_2 Z_6 vdd gnd pnand3_0
XXpre3x8_nand_7 in_0 in_1 in_2 Z_7 vdd gnd pnand3_0
.ENDS hierarchical_predecode3x8_0

.SUBCKT hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 decode_0 decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64 decode_65 decode_66 decode_67 decode_68 decode_69 decode_70 decode_71 decode_72 decode_73 decode_74 decode_75 decode_76 decode_77 decode_78 decode_79 decode_80 decode_81 decode_82 decode_83 decode_84 decode_85 decode_86 decode_87 decode_88 decode_89 decode_90 decode_91 decode_92 decode_93 decode_94 decode_95 decode_96 decode_97 decode_98 decode_99 decode_100 decode_101 decode_102 decode_103 decode_104 decode_105 decode_106 decode_107 decode_108 decode_109 decode_110 decode_111 decode_112 decode_113 decode_114 decode_115 decode_116 decode_117 decode_118 decode_119 decode_120 decode_121 decode_122 decode_123 decode_124 decode_125 decode_126 decode_127 decode_128 decode_129 decode_130 decode_131 decode_132 decode_133 decode_134 decode_135 decode_136 decode_137 decode_138 decode_139 decode_140 decode_141 decode_142 decode_143 decode_144 decode_145 decode_146 decode_147 decode_148 decode_149 decode_150 decode_151 decode_152 decode_153 decode_154 decode_155 decode_156 decode_157 decode_158 decode_159 decode_160 decode_161 decode_162 decode_163 decode_164 decode_165 decode_166 decode_167 decode_168 decode_169 decode_170 decode_171 decode_172 decode_173 decode_174 decode_175 decode_176 decode_177 decode_178 decode_179 decode_180 decode_181 decode_182 decode_183 decode_184 decode_185 decode_186 decode_187 decode_188 decode_189 decode_190 decode_191 decode_192 decode_193 decode_194 decode_195 decode_196 decode_197 decode_198 decode_199 decode_200 decode_201 decode_202 decode_203 decode_204 decode_205 decode_206 decode_207 decode_208 decode_209 decode_210 decode_211 decode_212 decode_213 decode_214 decode_215 decode_216 decode_217 decode_218 decode_219 decode_220 decode_221 decode_222 decode_223 decode_224 decode_225 decode_226 decode_227 decode_228 decode_229 decode_230 decode_231 decode_232 decode_233 decode_234 decode_235 decode_236 decode_237 decode_238 decode_239 decode_240 decode_241 decode_242 decode_243 decode_244 decode_245 decode_246 decode_247 decode_248 decode_249 decode_250 decode_251 decode_252 decode_253 decode_254 decode_255 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : addr_7 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* OUTPUT: decode_65 
* OUTPUT: decode_66 
* OUTPUT: decode_67 
* OUTPUT: decode_68 
* OUTPUT: decode_69 
* OUTPUT: decode_70 
* OUTPUT: decode_71 
* OUTPUT: decode_72 
* OUTPUT: decode_73 
* OUTPUT: decode_74 
* OUTPUT: decode_75 
* OUTPUT: decode_76 
* OUTPUT: decode_77 
* OUTPUT: decode_78 
* OUTPUT: decode_79 
* OUTPUT: decode_80 
* OUTPUT: decode_81 
* OUTPUT: decode_82 
* OUTPUT: decode_83 
* OUTPUT: decode_84 
* OUTPUT: decode_85 
* OUTPUT: decode_86 
* OUTPUT: decode_87 
* OUTPUT: decode_88 
* OUTPUT: decode_89 
* OUTPUT: decode_90 
* OUTPUT: decode_91 
* OUTPUT: decode_92 
* OUTPUT: decode_93 
* OUTPUT: decode_94 
* OUTPUT: decode_95 
* OUTPUT: decode_96 
* OUTPUT: decode_97 
* OUTPUT: decode_98 
* OUTPUT: decode_99 
* OUTPUT: decode_100 
* OUTPUT: decode_101 
* OUTPUT: decode_102 
* OUTPUT: decode_103 
* OUTPUT: decode_104 
* OUTPUT: decode_105 
* OUTPUT: decode_106 
* OUTPUT: decode_107 
* OUTPUT: decode_108 
* OUTPUT: decode_109 
* OUTPUT: decode_110 
* OUTPUT: decode_111 
* OUTPUT: decode_112 
* OUTPUT: decode_113 
* OUTPUT: decode_114 
* OUTPUT: decode_115 
* OUTPUT: decode_116 
* OUTPUT: decode_117 
* OUTPUT: decode_118 
* OUTPUT: decode_119 
* OUTPUT: decode_120 
* OUTPUT: decode_121 
* OUTPUT: decode_122 
* OUTPUT: decode_123 
* OUTPUT: decode_124 
* OUTPUT: decode_125 
* OUTPUT: decode_126 
* OUTPUT: decode_127 
* OUTPUT: decode_128 
* OUTPUT: decode_129 
* OUTPUT: decode_130 
* OUTPUT: decode_131 
* OUTPUT: decode_132 
* OUTPUT: decode_133 
* OUTPUT: decode_134 
* OUTPUT: decode_135 
* OUTPUT: decode_136 
* OUTPUT: decode_137 
* OUTPUT: decode_138 
* OUTPUT: decode_139 
* OUTPUT: decode_140 
* OUTPUT: decode_141 
* OUTPUT: decode_142 
* OUTPUT: decode_143 
* OUTPUT: decode_144 
* OUTPUT: decode_145 
* OUTPUT: decode_146 
* OUTPUT: decode_147 
* OUTPUT: decode_148 
* OUTPUT: decode_149 
* OUTPUT: decode_150 
* OUTPUT: decode_151 
* OUTPUT: decode_152 
* OUTPUT: decode_153 
* OUTPUT: decode_154 
* OUTPUT: decode_155 
* OUTPUT: decode_156 
* OUTPUT: decode_157 
* OUTPUT: decode_158 
* OUTPUT: decode_159 
* OUTPUT: decode_160 
* OUTPUT: decode_161 
* OUTPUT: decode_162 
* OUTPUT: decode_163 
* OUTPUT: decode_164 
* OUTPUT: decode_165 
* OUTPUT: decode_166 
* OUTPUT: decode_167 
* OUTPUT: decode_168 
* OUTPUT: decode_169 
* OUTPUT: decode_170 
* OUTPUT: decode_171 
* OUTPUT: decode_172 
* OUTPUT: decode_173 
* OUTPUT: decode_174 
* OUTPUT: decode_175 
* OUTPUT: decode_176 
* OUTPUT: decode_177 
* OUTPUT: decode_178 
* OUTPUT: decode_179 
* OUTPUT: decode_180 
* OUTPUT: decode_181 
* OUTPUT: decode_182 
* OUTPUT: decode_183 
* OUTPUT: decode_184 
* OUTPUT: decode_185 
* OUTPUT: decode_186 
* OUTPUT: decode_187 
* OUTPUT: decode_188 
* OUTPUT: decode_189 
* OUTPUT: decode_190 
* OUTPUT: decode_191 
* OUTPUT: decode_192 
* OUTPUT: decode_193 
* OUTPUT: decode_194 
* OUTPUT: decode_195 
* OUTPUT: decode_196 
* OUTPUT: decode_197 
* OUTPUT: decode_198 
* OUTPUT: decode_199 
* OUTPUT: decode_200 
* OUTPUT: decode_201 
* OUTPUT: decode_202 
* OUTPUT: decode_203 
* OUTPUT: decode_204 
* OUTPUT: decode_205 
* OUTPUT: decode_206 
* OUTPUT: decode_207 
* OUTPUT: decode_208 
* OUTPUT: decode_209 
* OUTPUT: decode_210 
* OUTPUT: decode_211 
* OUTPUT: decode_212 
* OUTPUT: decode_213 
* OUTPUT: decode_214 
* OUTPUT: decode_215 
* OUTPUT: decode_216 
* OUTPUT: decode_217 
* OUTPUT: decode_218 
* OUTPUT: decode_219 
* OUTPUT: decode_220 
* OUTPUT: decode_221 
* OUTPUT: decode_222 
* OUTPUT: decode_223 
* OUTPUT: decode_224 
* OUTPUT: decode_225 
* OUTPUT: decode_226 
* OUTPUT: decode_227 
* OUTPUT: decode_228 
* OUTPUT: decode_229 
* OUTPUT: decode_230 
* OUTPUT: decode_231 
* OUTPUT: decode_232 
* OUTPUT: decode_233 
* OUTPUT: decode_234 
* OUTPUT: decode_235 
* OUTPUT: decode_236 
* OUTPUT: decode_237 
* OUTPUT: decode_238 
* OUTPUT: decode_239 
* OUTPUT: decode_240 
* OUTPUT: decode_241 
* OUTPUT: decode_242 
* OUTPUT: decode_243 
* OUTPUT: decode_244 
* OUTPUT: decode_245 
* OUTPUT: decode_246 
* OUTPUT: decode_247 
* OUTPUT: decode_248 
* OUTPUT: decode_249 
* OUTPUT: decode_250 
* OUTPUT: decode_251 
* OUTPUT: decode_252 
* OUTPUT: decode_253 
* OUTPUT: decode_254 
* OUTPUT: decode_255 
* POWER : vdd 
* GROUND: gnd 
Xpre_0 addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd hierarchical_predecode2x4_0
Xpre3x8_0 addr_2 addr_3 addr_4 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11 vdd gnd hierarchical_predecode3x8_0
Xpre3x8_1 addr_5 addr_6 addr_7 out_12 out_13 out_14 out_15 out_16 out_17 out_18 out_19 vdd gnd hierarchical_predecode3x8_0
XDEC_NAND_0 out_0 out_4 out_12 Z_0 vdd gnd pnand3_0
XDEC_NAND_32 out_0 out_4 out_13 Z_32 vdd gnd pnand3_0
XDEC_NAND_64 out_0 out_4 out_14 Z_64 vdd gnd pnand3_0
XDEC_NAND_96 out_0 out_4 out_15 Z_96 vdd gnd pnand3_0
XDEC_NAND_128 out_0 out_4 out_16 Z_128 vdd gnd pnand3_0
XDEC_NAND_160 out_0 out_4 out_17 Z_160 vdd gnd pnand3_0
XDEC_NAND_192 out_0 out_4 out_18 Z_192 vdd gnd pnand3_0
XDEC_NAND_224 out_0 out_4 out_19 Z_224 vdd gnd pnand3_0
XDEC_NAND_4 out_0 out_5 out_12 Z_4 vdd gnd pnand3_0
XDEC_NAND_36 out_0 out_5 out_13 Z_36 vdd gnd pnand3_0
XDEC_NAND_68 out_0 out_5 out_14 Z_68 vdd gnd pnand3_0
XDEC_NAND_100 out_0 out_5 out_15 Z_100 vdd gnd pnand3_0
XDEC_NAND_132 out_0 out_5 out_16 Z_132 vdd gnd pnand3_0
XDEC_NAND_164 out_0 out_5 out_17 Z_164 vdd gnd pnand3_0
XDEC_NAND_196 out_0 out_5 out_18 Z_196 vdd gnd pnand3_0
XDEC_NAND_228 out_0 out_5 out_19 Z_228 vdd gnd pnand3_0
XDEC_NAND_8 out_0 out_6 out_12 Z_8 vdd gnd pnand3_0
XDEC_NAND_40 out_0 out_6 out_13 Z_40 vdd gnd pnand3_0
XDEC_NAND_72 out_0 out_6 out_14 Z_72 vdd gnd pnand3_0
XDEC_NAND_104 out_0 out_6 out_15 Z_104 vdd gnd pnand3_0
XDEC_NAND_136 out_0 out_6 out_16 Z_136 vdd gnd pnand3_0
XDEC_NAND_168 out_0 out_6 out_17 Z_168 vdd gnd pnand3_0
XDEC_NAND_200 out_0 out_6 out_18 Z_200 vdd gnd pnand3_0
XDEC_NAND_232 out_0 out_6 out_19 Z_232 vdd gnd pnand3_0
XDEC_NAND_12 out_0 out_7 out_12 Z_12 vdd gnd pnand3_0
XDEC_NAND_44 out_0 out_7 out_13 Z_44 vdd gnd pnand3_0
XDEC_NAND_76 out_0 out_7 out_14 Z_76 vdd gnd pnand3_0
XDEC_NAND_108 out_0 out_7 out_15 Z_108 vdd gnd pnand3_0
XDEC_NAND_140 out_0 out_7 out_16 Z_140 vdd gnd pnand3_0
XDEC_NAND_172 out_0 out_7 out_17 Z_172 vdd gnd pnand3_0
XDEC_NAND_204 out_0 out_7 out_18 Z_204 vdd gnd pnand3_0
XDEC_NAND_236 out_0 out_7 out_19 Z_236 vdd gnd pnand3_0
XDEC_NAND_16 out_0 out_8 out_12 Z_16 vdd gnd pnand3_0
XDEC_NAND_48 out_0 out_8 out_13 Z_48 vdd gnd pnand3_0
XDEC_NAND_80 out_0 out_8 out_14 Z_80 vdd gnd pnand3_0
XDEC_NAND_112 out_0 out_8 out_15 Z_112 vdd gnd pnand3_0
XDEC_NAND_144 out_0 out_8 out_16 Z_144 vdd gnd pnand3_0
XDEC_NAND_176 out_0 out_8 out_17 Z_176 vdd gnd pnand3_0
XDEC_NAND_208 out_0 out_8 out_18 Z_208 vdd gnd pnand3_0
XDEC_NAND_240 out_0 out_8 out_19 Z_240 vdd gnd pnand3_0
XDEC_NAND_20 out_0 out_9 out_12 Z_20 vdd gnd pnand3_0
XDEC_NAND_52 out_0 out_9 out_13 Z_52 vdd gnd pnand3_0
XDEC_NAND_84 out_0 out_9 out_14 Z_84 vdd gnd pnand3_0
XDEC_NAND_116 out_0 out_9 out_15 Z_116 vdd gnd pnand3_0
XDEC_NAND_148 out_0 out_9 out_16 Z_148 vdd gnd pnand3_0
XDEC_NAND_180 out_0 out_9 out_17 Z_180 vdd gnd pnand3_0
XDEC_NAND_212 out_0 out_9 out_18 Z_212 vdd gnd pnand3_0
XDEC_NAND_244 out_0 out_9 out_19 Z_244 vdd gnd pnand3_0
XDEC_NAND_24 out_0 out_10 out_12 Z_24 vdd gnd pnand3_0
XDEC_NAND_56 out_0 out_10 out_13 Z_56 vdd gnd pnand3_0
XDEC_NAND_88 out_0 out_10 out_14 Z_88 vdd gnd pnand3_0
XDEC_NAND_120 out_0 out_10 out_15 Z_120 vdd gnd pnand3_0
XDEC_NAND_152 out_0 out_10 out_16 Z_152 vdd gnd pnand3_0
XDEC_NAND_184 out_0 out_10 out_17 Z_184 vdd gnd pnand3_0
XDEC_NAND_216 out_0 out_10 out_18 Z_216 vdd gnd pnand3_0
XDEC_NAND_248 out_0 out_10 out_19 Z_248 vdd gnd pnand3_0
XDEC_NAND_28 out_0 out_11 out_12 Z_28 vdd gnd pnand3_0
XDEC_NAND_60 out_0 out_11 out_13 Z_60 vdd gnd pnand3_0
XDEC_NAND_92 out_0 out_11 out_14 Z_92 vdd gnd pnand3_0
XDEC_NAND_124 out_0 out_11 out_15 Z_124 vdd gnd pnand3_0
XDEC_NAND_156 out_0 out_11 out_16 Z_156 vdd gnd pnand3_0
XDEC_NAND_188 out_0 out_11 out_17 Z_188 vdd gnd pnand3_0
XDEC_NAND_220 out_0 out_11 out_18 Z_220 vdd gnd pnand3_0
XDEC_NAND_252 out_0 out_11 out_19 Z_252 vdd gnd pnand3_0
XDEC_NAND_1 out_1 out_4 out_12 Z_1 vdd gnd pnand3_0
XDEC_NAND_33 out_1 out_4 out_13 Z_33 vdd gnd pnand3_0
XDEC_NAND_65 out_1 out_4 out_14 Z_65 vdd gnd pnand3_0
XDEC_NAND_97 out_1 out_4 out_15 Z_97 vdd gnd pnand3_0
XDEC_NAND_129 out_1 out_4 out_16 Z_129 vdd gnd pnand3_0
XDEC_NAND_161 out_1 out_4 out_17 Z_161 vdd gnd pnand3_0
XDEC_NAND_193 out_1 out_4 out_18 Z_193 vdd gnd pnand3_0
XDEC_NAND_225 out_1 out_4 out_19 Z_225 vdd gnd pnand3_0
XDEC_NAND_5 out_1 out_5 out_12 Z_5 vdd gnd pnand3_0
XDEC_NAND_37 out_1 out_5 out_13 Z_37 vdd gnd pnand3_0
XDEC_NAND_69 out_1 out_5 out_14 Z_69 vdd gnd pnand3_0
XDEC_NAND_101 out_1 out_5 out_15 Z_101 vdd gnd pnand3_0
XDEC_NAND_133 out_1 out_5 out_16 Z_133 vdd gnd pnand3_0
XDEC_NAND_165 out_1 out_5 out_17 Z_165 vdd gnd pnand3_0
XDEC_NAND_197 out_1 out_5 out_18 Z_197 vdd gnd pnand3_0
XDEC_NAND_229 out_1 out_5 out_19 Z_229 vdd gnd pnand3_0
XDEC_NAND_9 out_1 out_6 out_12 Z_9 vdd gnd pnand3_0
XDEC_NAND_41 out_1 out_6 out_13 Z_41 vdd gnd pnand3_0
XDEC_NAND_73 out_1 out_6 out_14 Z_73 vdd gnd pnand3_0
XDEC_NAND_105 out_1 out_6 out_15 Z_105 vdd gnd pnand3_0
XDEC_NAND_137 out_1 out_6 out_16 Z_137 vdd gnd pnand3_0
XDEC_NAND_169 out_1 out_6 out_17 Z_169 vdd gnd pnand3_0
XDEC_NAND_201 out_1 out_6 out_18 Z_201 vdd gnd pnand3_0
XDEC_NAND_233 out_1 out_6 out_19 Z_233 vdd gnd pnand3_0
XDEC_NAND_13 out_1 out_7 out_12 Z_13 vdd gnd pnand3_0
XDEC_NAND_45 out_1 out_7 out_13 Z_45 vdd gnd pnand3_0
XDEC_NAND_77 out_1 out_7 out_14 Z_77 vdd gnd pnand3_0
XDEC_NAND_109 out_1 out_7 out_15 Z_109 vdd gnd pnand3_0
XDEC_NAND_141 out_1 out_7 out_16 Z_141 vdd gnd pnand3_0
XDEC_NAND_173 out_1 out_7 out_17 Z_173 vdd gnd pnand3_0
XDEC_NAND_205 out_1 out_7 out_18 Z_205 vdd gnd pnand3_0
XDEC_NAND_237 out_1 out_7 out_19 Z_237 vdd gnd pnand3_0
XDEC_NAND_17 out_1 out_8 out_12 Z_17 vdd gnd pnand3_0
XDEC_NAND_49 out_1 out_8 out_13 Z_49 vdd gnd pnand3_0
XDEC_NAND_81 out_1 out_8 out_14 Z_81 vdd gnd pnand3_0
XDEC_NAND_113 out_1 out_8 out_15 Z_113 vdd gnd pnand3_0
XDEC_NAND_145 out_1 out_8 out_16 Z_145 vdd gnd pnand3_0
XDEC_NAND_177 out_1 out_8 out_17 Z_177 vdd gnd pnand3_0
XDEC_NAND_209 out_1 out_8 out_18 Z_209 vdd gnd pnand3_0
XDEC_NAND_241 out_1 out_8 out_19 Z_241 vdd gnd pnand3_0
XDEC_NAND_21 out_1 out_9 out_12 Z_21 vdd gnd pnand3_0
XDEC_NAND_53 out_1 out_9 out_13 Z_53 vdd gnd pnand3_0
XDEC_NAND_85 out_1 out_9 out_14 Z_85 vdd gnd pnand3_0
XDEC_NAND_117 out_1 out_9 out_15 Z_117 vdd gnd pnand3_0
XDEC_NAND_149 out_1 out_9 out_16 Z_149 vdd gnd pnand3_0
XDEC_NAND_181 out_1 out_9 out_17 Z_181 vdd gnd pnand3_0
XDEC_NAND_213 out_1 out_9 out_18 Z_213 vdd gnd pnand3_0
XDEC_NAND_245 out_1 out_9 out_19 Z_245 vdd gnd pnand3_0
XDEC_NAND_25 out_1 out_10 out_12 Z_25 vdd gnd pnand3_0
XDEC_NAND_57 out_1 out_10 out_13 Z_57 vdd gnd pnand3_0
XDEC_NAND_89 out_1 out_10 out_14 Z_89 vdd gnd pnand3_0
XDEC_NAND_121 out_1 out_10 out_15 Z_121 vdd gnd pnand3_0
XDEC_NAND_153 out_1 out_10 out_16 Z_153 vdd gnd pnand3_0
XDEC_NAND_185 out_1 out_10 out_17 Z_185 vdd gnd pnand3_0
XDEC_NAND_217 out_1 out_10 out_18 Z_217 vdd gnd pnand3_0
XDEC_NAND_249 out_1 out_10 out_19 Z_249 vdd gnd pnand3_0
XDEC_NAND_29 out_1 out_11 out_12 Z_29 vdd gnd pnand3_0
XDEC_NAND_61 out_1 out_11 out_13 Z_61 vdd gnd pnand3_0
XDEC_NAND_93 out_1 out_11 out_14 Z_93 vdd gnd pnand3_0
XDEC_NAND_125 out_1 out_11 out_15 Z_125 vdd gnd pnand3_0
XDEC_NAND_157 out_1 out_11 out_16 Z_157 vdd gnd pnand3_0
XDEC_NAND_189 out_1 out_11 out_17 Z_189 vdd gnd pnand3_0
XDEC_NAND_221 out_1 out_11 out_18 Z_221 vdd gnd pnand3_0
XDEC_NAND_253 out_1 out_11 out_19 Z_253 vdd gnd pnand3_0
XDEC_NAND_2 out_2 out_4 out_12 Z_2 vdd gnd pnand3_0
XDEC_NAND_34 out_2 out_4 out_13 Z_34 vdd gnd pnand3_0
XDEC_NAND_66 out_2 out_4 out_14 Z_66 vdd gnd pnand3_0
XDEC_NAND_98 out_2 out_4 out_15 Z_98 vdd gnd pnand3_0
XDEC_NAND_130 out_2 out_4 out_16 Z_130 vdd gnd pnand3_0
XDEC_NAND_162 out_2 out_4 out_17 Z_162 vdd gnd pnand3_0
XDEC_NAND_194 out_2 out_4 out_18 Z_194 vdd gnd pnand3_0
XDEC_NAND_226 out_2 out_4 out_19 Z_226 vdd gnd pnand3_0
XDEC_NAND_6 out_2 out_5 out_12 Z_6 vdd gnd pnand3_0
XDEC_NAND_38 out_2 out_5 out_13 Z_38 vdd gnd pnand3_0
XDEC_NAND_70 out_2 out_5 out_14 Z_70 vdd gnd pnand3_0
XDEC_NAND_102 out_2 out_5 out_15 Z_102 vdd gnd pnand3_0
XDEC_NAND_134 out_2 out_5 out_16 Z_134 vdd gnd pnand3_0
XDEC_NAND_166 out_2 out_5 out_17 Z_166 vdd gnd pnand3_0
XDEC_NAND_198 out_2 out_5 out_18 Z_198 vdd gnd pnand3_0
XDEC_NAND_230 out_2 out_5 out_19 Z_230 vdd gnd pnand3_0
XDEC_NAND_10 out_2 out_6 out_12 Z_10 vdd gnd pnand3_0
XDEC_NAND_42 out_2 out_6 out_13 Z_42 vdd gnd pnand3_0
XDEC_NAND_74 out_2 out_6 out_14 Z_74 vdd gnd pnand3_0
XDEC_NAND_106 out_2 out_6 out_15 Z_106 vdd gnd pnand3_0
XDEC_NAND_138 out_2 out_6 out_16 Z_138 vdd gnd pnand3_0
XDEC_NAND_170 out_2 out_6 out_17 Z_170 vdd gnd pnand3_0
XDEC_NAND_202 out_2 out_6 out_18 Z_202 vdd gnd pnand3_0
XDEC_NAND_234 out_2 out_6 out_19 Z_234 vdd gnd pnand3_0
XDEC_NAND_14 out_2 out_7 out_12 Z_14 vdd gnd pnand3_0
XDEC_NAND_46 out_2 out_7 out_13 Z_46 vdd gnd pnand3_0
XDEC_NAND_78 out_2 out_7 out_14 Z_78 vdd gnd pnand3_0
XDEC_NAND_110 out_2 out_7 out_15 Z_110 vdd gnd pnand3_0
XDEC_NAND_142 out_2 out_7 out_16 Z_142 vdd gnd pnand3_0
XDEC_NAND_174 out_2 out_7 out_17 Z_174 vdd gnd pnand3_0
XDEC_NAND_206 out_2 out_7 out_18 Z_206 vdd gnd pnand3_0
XDEC_NAND_238 out_2 out_7 out_19 Z_238 vdd gnd pnand3_0
XDEC_NAND_18 out_2 out_8 out_12 Z_18 vdd gnd pnand3_0
XDEC_NAND_50 out_2 out_8 out_13 Z_50 vdd gnd pnand3_0
XDEC_NAND_82 out_2 out_8 out_14 Z_82 vdd gnd pnand3_0
XDEC_NAND_114 out_2 out_8 out_15 Z_114 vdd gnd pnand3_0
XDEC_NAND_146 out_2 out_8 out_16 Z_146 vdd gnd pnand3_0
XDEC_NAND_178 out_2 out_8 out_17 Z_178 vdd gnd pnand3_0
XDEC_NAND_210 out_2 out_8 out_18 Z_210 vdd gnd pnand3_0
XDEC_NAND_242 out_2 out_8 out_19 Z_242 vdd gnd pnand3_0
XDEC_NAND_22 out_2 out_9 out_12 Z_22 vdd gnd pnand3_0
XDEC_NAND_54 out_2 out_9 out_13 Z_54 vdd gnd pnand3_0
XDEC_NAND_86 out_2 out_9 out_14 Z_86 vdd gnd pnand3_0
XDEC_NAND_118 out_2 out_9 out_15 Z_118 vdd gnd pnand3_0
XDEC_NAND_150 out_2 out_9 out_16 Z_150 vdd gnd pnand3_0
XDEC_NAND_182 out_2 out_9 out_17 Z_182 vdd gnd pnand3_0
XDEC_NAND_214 out_2 out_9 out_18 Z_214 vdd gnd pnand3_0
XDEC_NAND_246 out_2 out_9 out_19 Z_246 vdd gnd pnand3_0
XDEC_NAND_26 out_2 out_10 out_12 Z_26 vdd gnd pnand3_0
XDEC_NAND_58 out_2 out_10 out_13 Z_58 vdd gnd pnand3_0
XDEC_NAND_90 out_2 out_10 out_14 Z_90 vdd gnd pnand3_0
XDEC_NAND_122 out_2 out_10 out_15 Z_122 vdd gnd pnand3_0
XDEC_NAND_154 out_2 out_10 out_16 Z_154 vdd gnd pnand3_0
XDEC_NAND_186 out_2 out_10 out_17 Z_186 vdd gnd pnand3_0
XDEC_NAND_218 out_2 out_10 out_18 Z_218 vdd gnd pnand3_0
XDEC_NAND_250 out_2 out_10 out_19 Z_250 vdd gnd pnand3_0
XDEC_NAND_30 out_2 out_11 out_12 Z_30 vdd gnd pnand3_0
XDEC_NAND_62 out_2 out_11 out_13 Z_62 vdd gnd pnand3_0
XDEC_NAND_94 out_2 out_11 out_14 Z_94 vdd gnd pnand3_0
XDEC_NAND_126 out_2 out_11 out_15 Z_126 vdd gnd pnand3_0
XDEC_NAND_158 out_2 out_11 out_16 Z_158 vdd gnd pnand3_0
XDEC_NAND_190 out_2 out_11 out_17 Z_190 vdd gnd pnand3_0
XDEC_NAND_222 out_2 out_11 out_18 Z_222 vdd gnd pnand3_0
XDEC_NAND_254 out_2 out_11 out_19 Z_254 vdd gnd pnand3_0
XDEC_NAND_3 out_3 out_4 out_12 Z_3 vdd gnd pnand3_0
XDEC_NAND_35 out_3 out_4 out_13 Z_35 vdd gnd pnand3_0
XDEC_NAND_67 out_3 out_4 out_14 Z_67 vdd gnd pnand3_0
XDEC_NAND_99 out_3 out_4 out_15 Z_99 vdd gnd pnand3_0
XDEC_NAND_131 out_3 out_4 out_16 Z_131 vdd gnd pnand3_0
XDEC_NAND_163 out_3 out_4 out_17 Z_163 vdd gnd pnand3_0
XDEC_NAND_195 out_3 out_4 out_18 Z_195 vdd gnd pnand3_0
XDEC_NAND_227 out_3 out_4 out_19 Z_227 vdd gnd pnand3_0
XDEC_NAND_7 out_3 out_5 out_12 Z_7 vdd gnd pnand3_0
XDEC_NAND_39 out_3 out_5 out_13 Z_39 vdd gnd pnand3_0
XDEC_NAND_71 out_3 out_5 out_14 Z_71 vdd gnd pnand3_0
XDEC_NAND_103 out_3 out_5 out_15 Z_103 vdd gnd pnand3_0
XDEC_NAND_135 out_3 out_5 out_16 Z_135 vdd gnd pnand3_0
XDEC_NAND_167 out_3 out_5 out_17 Z_167 vdd gnd pnand3_0
XDEC_NAND_199 out_3 out_5 out_18 Z_199 vdd gnd pnand3_0
XDEC_NAND_231 out_3 out_5 out_19 Z_231 vdd gnd pnand3_0
XDEC_NAND_11 out_3 out_6 out_12 Z_11 vdd gnd pnand3_0
XDEC_NAND_43 out_3 out_6 out_13 Z_43 vdd gnd pnand3_0
XDEC_NAND_75 out_3 out_6 out_14 Z_75 vdd gnd pnand3_0
XDEC_NAND_107 out_3 out_6 out_15 Z_107 vdd gnd pnand3_0
XDEC_NAND_139 out_3 out_6 out_16 Z_139 vdd gnd pnand3_0
XDEC_NAND_171 out_3 out_6 out_17 Z_171 vdd gnd pnand3_0
XDEC_NAND_203 out_3 out_6 out_18 Z_203 vdd gnd pnand3_0
XDEC_NAND_235 out_3 out_6 out_19 Z_235 vdd gnd pnand3_0
XDEC_NAND_15 out_3 out_7 out_12 Z_15 vdd gnd pnand3_0
XDEC_NAND_47 out_3 out_7 out_13 Z_47 vdd gnd pnand3_0
XDEC_NAND_79 out_3 out_7 out_14 Z_79 vdd gnd pnand3_0
XDEC_NAND_111 out_3 out_7 out_15 Z_111 vdd gnd pnand3_0
XDEC_NAND_143 out_3 out_7 out_16 Z_143 vdd gnd pnand3_0
XDEC_NAND_175 out_3 out_7 out_17 Z_175 vdd gnd pnand3_0
XDEC_NAND_207 out_3 out_7 out_18 Z_207 vdd gnd pnand3_0
XDEC_NAND_239 out_3 out_7 out_19 Z_239 vdd gnd pnand3_0
XDEC_NAND_19 out_3 out_8 out_12 Z_19 vdd gnd pnand3_0
XDEC_NAND_51 out_3 out_8 out_13 Z_51 vdd gnd pnand3_0
XDEC_NAND_83 out_3 out_8 out_14 Z_83 vdd gnd pnand3_0
XDEC_NAND_115 out_3 out_8 out_15 Z_115 vdd gnd pnand3_0
XDEC_NAND_147 out_3 out_8 out_16 Z_147 vdd gnd pnand3_0
XDEC_NAND_179 out_3 out_8 out_17 Z_179 vdd gnd pnand3_0
XDEC_NAND_211 out_3 out_8 out_18 Z_211 vdd gnd pnand3_0
XDEC_NAND_243 out_3 out_8 out_19 Z_243 vdd gnd pnand3_0
XDEC_NAND_23 out_3 out_9 out_12 Z_23 vdd gnd pnand3_0
XDEC_NAND_55 out_3 out_9 out_13 Z_55 vdd gnd pnand3_0
XDEC_NAND_87 out_3 out_9 out_14 Z_87 vdd gnd pnand3_0
XDEC_NAND_119 out_3 out_9 out_15 Z_119 vdd gnd pnand3_0
XDEC_NAND_151 out_3 out_9 out_16 Z_151 vdd gnd pnand3_0
XDEC_NAND_183 out_3 out_9 out_17 Z_183 vdd gnd pnand3_0
XDEC_NAND_215 out_3 out_9 out_18 Z_215 vdd gnd pnand3_0
XDEC_NAND_247 out_3 out_9 out_19 Z_247 vdd gnd pnand3_0
XDEC_NAND_27 out_3 out_10 out_12 Z_27 vdd gnd pnand3_0
XDEC_NAND_59 out_3 out_10 out_13 Z_59 vdd gnd pnand3_0
XDEC_NAND_91 out_3 out_10 out_14 Z_91 vdd gnd pnand3_0
XDEC_NAND_123 out_3 out_10 out_15 Z_123 vdd gnd pnand3_0
XDEC_NAND_155 out_3 out_10 out_16 Z_155 vdd gnd pnand3_0
XDEC_NAND_187 out_3 out_10 out_17 Z_187 vdd gnd pnand3_0
XDEC_NAND_219 out_3 out_10 out_18 Z_219 vdd gnd pnand3_0
XDEC_NAND_251 out_3 out_10 out_19 Z_251 vdd gnd pnand3_0
XDEC_NAND_31 out_3 out_11 out_12 Z_31 vdd gnd pnand3_0
XDEC_NAND_63 out_3 out_11 out_13 Z_63 vdd gnd pnand3_0
XDEC_NAND_95 out_3 out_11 out_14 Z_95 vdd gnd pnand3_0
XDEC_NAND_127 out_3 out_11 out_15 Z_127 vdd gnd pnand3_0
XDEC_NAND_159 out_3 out_11 out_16 Z_159 vdd gnd pnand3_0
XDEC_NAND_191 out_3 out_11 out_17 Z_191 vdd gnd pnand3_0
XDEC_NAND_223 out_3 out_11 out_18 Z_223 vdd gnd pnand3_0
XDEC_NAND_255 out_3 out_11 out_19 Z_255 vdd gnd pnand3_0
XDEC_INV_0 Z_0 decode_0 vdd gnd pinv_0
XDEC_INV_1 Z_1 decode_1 vdd gnd pinv_0
XDEC_INV_2 Z_2 decode_2 vdd gnd pinv_0
XDEC_INV_3 Z_3 decode_3 vdd gnd pinv_0
XDEC_INV_4 Z_4 decode_4 vdd gnd pinv_0
XDEC_INV_5 Z_5 decode_5 vdd gnd pinv_0
XDEC_INV_6 Z_6 decode_6 vdd gnd pinv_0
XDEC_INV_7 Z_7 decode_7 vdd gnd pinv_0
XDEC_INV_8 Z_8 decode_8 vdd gnd pinv_0
XDEC_INV_9 Z_9 decode_9 vdd gnd pinv_0
XDEC_INV_10 Z_10 decode_10 vdd gnd pinv_0
XDEC_INV_11 Z_11 decode_11 vdd gnd pinv_0
XDEC_INV_12 Z_12 decode_12 vdd gnd pinv_0
XDEC_INV_13 Z_13 decode_13 vdd gnd pinv_0
XDEC_INV_14 Z_14 decode_14 vdd gnd pinv_0
XDEC_INV_15 Z_15 decode_15 vdd gnd pinv_0
XDEC_INV_16 Z_16 decode_16 vdd gnd pinv_0
XDEC_INV_17 Z_17 decode_17 vdd gnd pinv_0
XDEC_INV_18 Z_18 decode_18 vdd gnd pinv_0
XDEC_INV_19 Z_19 decode_19 vdd gnd pinv_0
XDEC_INV_20 Z_20 decode_20 vdd gnd pinv_0
XDEC_INV_21 Z_21 decode_21 vdd gnd pinv_0
XDEC_INV_22 Z_22 decode_22 vdd gnd pinv_0
XDEC_INV_23 Z_23 decode_23 vdd gnd pinv_0
XDEC_INV_24 Z_24 decode_24 vdd gnd pinv_0
XDEC_INV_25 Z_25 decode_25 vdd gnd pinv_0
XDEC_INV_26 Z_26 decode_26 vdd gnd pinv_0
XDEC_INV_27 Z_27 decode_27 vdd gnd pinv_0
XDEC_INV_28 Z_28 decode_28 vdd gnd pinv_0
XDEC_INV_29 Z_29 decode_29 vdd gnd pinv_0
XDEC_INV_30 Z_30 decode_30 vdd gnd pinv_0
XDEC_INV_31 Z_31 decode_31 vdd gnd pinv_0
XDEC_INV_32 Z_32 decode_32 vdd gnd pinv_0
XDEC_INV_33 Z_33 decode_33 vdd gnd pinv_0
XDEC_INV_34 Z_34 decode_34 vdd gnd pinv_0
XDEC_INV_35 Z_35 decode_35 vdd gnd pinv_0
XDEC_INV_36 Z_36 decode_36 vdd gnd pinv_0
XDEC_INV_37 Z_37 decode_37 vdd gnd pinv_0
XDEC_INV_38 Z_38 decode_38 vdd gnd pinv_0
XDEC_INV_39 Z_39 decode_39 vdd gnd pinv_0
XDEC_INV_40 Z_40 decode_40 vdd gnd pinv_0
XDEC_INV_41 Z_41 decode_41 vdd gnd pinv_0
XDEC_INV_42 Z_42 decode_42 vdd gnd pinv_0
XDEC_INV_43 Z_43 decode_43 vdd gnd pinv_0
XDEC_INV_44 Z_44 decode_44 vdd gnd pinv_0
XDEC_INV_45 Z_45 decode_45 vdd gnd pinv_0
XDEC_INV_46 Z_46 decode_46 vdd gnd pinv_0
XDEC_INV_47 Z_47 decode_47 vdd gnd pinv_0
XDEC_INV_48 Z_48 decode_48 vdd gnd pinv_0
XDEC_INV_49 Z_49 decode_49 vdd gnd pinv_0
XDEC_INV_50 Z_50 decode_50 vdd gnd pinv_0
XDEC_INV_51 Z_51 decode_51 vdd gnd pinv_0
XDEC_INV_52 Z_52 decode_52 vdd gnd pinv_0
XDEC_INV_53 Z_53 decode_53 vdd gnd pinv_0
XDEC_INV_54 Z_54 decode_54 vdd gnd pinv_0
XDEC_INV_55 Z_55 decode_55 vdd gnd pinv_0
XDEC_INV_56 Z_56 decode_56 vdd gnd pinv_0
XDEC_INV_57 Z_57 decode_57 vdd gnd pinv_0
XDEC_INV_58 Z_58 decode_58 vdd gnd pinv_0
XDEC_INV_59 Z_59 decode_59 vdd gnd pinv_0
XDEC_INV_60 Z_60 decode_60 vdd gnd pinv_0
XDEC_INV_61 Z_61 decode_61 vdd gnd pinv_0
XDEC_INV_62 Z_62 decode_62 vdd gnd pinv_0
XDEC_INV_63 Z_63 decode_63 vdd gnd pinv_0
XDEC_INV_64 Z_64 decode_64 vdd gnd pinv_0
XDEC_INV_65 Z_65 decode_65 vdd gnd pinv_0
XDEC_INV_66 Z_66 decode_66 vdd gnd pinv_0
XDEC_INV_67 Z_67 decode_67 vdd gnd pinv_0
XDEC_INV_68 Z_68 decode_68 vdd gnd pinv_0
XDEC_INV_69 Z_69 decode_69 vdd gnd pinv_0
XDEC_INV_70 Z_70 decode_70 vdd gnd pinv_0
XDEC_INV_71 Z_71 decode_71 vdd gnd pinv_0
XDEC_INV_72 Z_72 decode_72 vdd gnd pinv_0
XDEC_INV_73 Z_73 decode_73 vdd gnd pinv_0
XDEC_INV_74 Z_74 decode_74 vdd gnd pinv_0
XDEC_INV_75 Z_75 decode_75 vdd gnd pinv_0
XDEC_INV_76 Z_76 decode_76 vdd gnd pinv_0
XDEC_INV_77 Z_77 decode_77 vdd gnd pinv_0
XDEC_INV_78 Z_78 decode_78 vdd gnd pinv_0
XDEC_INV_79 Z_79 decode_79 vdd gnd pinv_0
XDEC_INV_80 Z_80 decode_80 vdd gnd pinv_0
XDEC_INV_81 Z_81 decode_81 vdd gnd pinv_0
XDEC_INV_82 Z_82 decode_82 vdd gnd pinv_0
XDEC_INV_83 Z_83 decode_83 vdd gnd pinv_0
XDEC_INV_84 Z_84 decode_84 vdd gnd pinv_0
XDEC_INV_85 Z_85 decode_85 vdd gnd pinv_0
XDEC_INV_86 Z_86 decode_86 vdd gnd pinv_0
XDEC_INV_87 Z_87 decode_87 vdd gnd pinv_0
XDEC_INV_88 Z_88 decode_88 vdd gnd pinv_0
XDEC_INV_89 Z_89 decode_89 vdd gnd pinv_0
XDEC_INV_90 Z_90 decode_90 vdd gnd pinv_0
XDEC_INV_91 Z_91 decode_91 vdd gnd pinv_0
XDEC_INV_92 Z_92 decode_92 vdd gnd pinv_0
XDEC_INV_93 Z_93 decode_93 vdd gnd pinv_0
XDEC_INV_94 Z_94 decode_94 vdd gnd pinv_0
XDEC_INV_95 Z_95 decode_95 vdd gnd pinv_0
XDEC_INV_96 Z_96 decode_96 vdd gnd pinv_0
XDEC_INV_97 Z_97 decode_97 vdd gnd pinv_0
XDEC_INV_98 Z_98 decode_98 vdd gnd pinv_0
XDEC_INV_99 Z_99 decode_99 vdd gnd pinv_0
XDEC_INV_100 Z_100 decode_100 vdd gnd pinv_0
XDEC_INV_101 Z_101 decode_101 vdd gnd pinv_0
XDEC_INV_102 Z_102 decode_102 vdd gnd pinv_0
XDEC_INV_103 Z_103 decode_103 vdd gnd pinv_0
XDEC_INV_104 Z_104 decode_104 vdd gnd pinv_0
XDEC_INV_105 Z_105 decode_105 vdd gnd pinv_0
XDEC_INV_106 Z_106 decode_106 vdd gnd pinv_0
XDEC_INV_107 Z_107 decode_107 vdd gnd pinv_0
XDEC_INV_108 Z_108 decode_108 vdd gnd pinv_0
XDEC_INV_109 Z_109 decode_109 vdd gnd pinv_0
XDEC_INV_110 Z_110 decode_110 vdd gnd pinv_0
XDEC_INV_111 Z_111 decode_111 vdd gnd pinv_0
XDEC_INV_112 Z_112 decode_112 vdd gnd pinv_0
XDEC_INV_113 Z_113 decode_113 vdd gnd pinv_0
XDEC_INV_114 Z_114 decode_114 vdd gnd pinv_0
XDEC_INV_115 Z_115 decode_115 vdd gnd pinv_0
XDEC_INV_116 Z_116 decode_116 vdd gnd pinv_0
XDEC_INV_117 Z_117 decode_117 vdd gnd pinv_0
XDEC_INV_118 Z_118 decode_118 vdd gnd pinv_0
XDEC_INV_119 Z_119 decode_119 vdd gnd pinv_0
XDEC_INV_120 Z_120 decode_120 vdd gnd pinv_0
XDEC_INV_121 Z_121 decode_121 vdd gnd pinv_0
XDEC_INV_122 Z_122 decode_122 vdd gnd pinv_0
XDEC_INV_123 Z_123 decode_123 vdd gnd pinv_0
XDEC_INV_124 Z_124 decode_124 vdd gnd pinv_0
XDEC_INV_125 Z_125 decode_125 vdd gnd pinv_0
XDEC_INV_126 Z_126 decode_126 vdd gnd pinv_0
XDEC_INV_127 Z_127 decode_127 vdd gnd pinv_0
XDEC_INV_128 Z_128 decode_128 vdd gnd pinv_0
XDEC_INV_129 Z_129 decode_129 vdd gnd pinv_0
XDEC_INV_130 Z_130 decode_130 vdd gnd pinv_0
XDEC_INV_131 Z_131 decode_131 vdd gnd pinv_0
XDEC_INV_132 Z_132 decode_132 vdd gnd pinv_0
XDEC_INV_133 Z_133 decode_133 vdd gnd pinv_0
XDEC_INV_134 Z_134 decode_134 vdd gnd pinv_0
XDEC_INV_135 Z_135 decode_135 vdd gnd pinv_0
XDEC_INV_136 Z_136 decode_136 vdd gnd pinv_0
XDEC_INV_137 Z_137 decode_137 vdd gnd pinv_0
XDEC_INV_138 Z_138 decode_138 vdd gnd pinv_0
XDEC_INV_139 Z_139 decode_139 vdd gnd pinv_0
XDEC_INV_140 Z_140 decode_140 vdd gnd pinv_0
XDEC_INV_141 Z_141 decode_141 vdd gnd pinv_0
XDEC_INV_142 Z_142 decode_142 vdd gnd pinv_0
XDEC_INV_143 Z_143 decode_143 vdd gnd pinv_0
XDEC_INV_144 Z_144 decode_144 vdd gnd pinv_0
XDEC_INV_145 Z_145 decode_145 vdd gnd pinv_0
XDEC_INV_146 Z_146 decode_146 vdd gnd pinv_0
XDEC_INV_147 Z_147 decode_147 vdd gnd pinv_0
XDEC_INV_148 Z_148 decode_148 vdd gnd pinv_0
XDEC_INV_149 Z_149 decode_149 vdd gnd pinv_0
XDEC_INV_150 Z_150 decode_150 vdd gnd pinv_0
XDEC_INV_151 Z_151 decode_151 vdd gnd pinv_0
XDEC_INV_152 Z_152 decode_152 vdd gnd pinv_0
XDEC_INV_153 Z_153 decode_153 vdd gnd pinv_0
XDEC_INV_154 Z_154 decode_154 vdd gnd pinv_0
XDEC_INV_155 Z_155 decode_155 vdd gnd pinv_0
XDEC_INV_156 Z_156 decode_156 vdd gnd pinv_0
XDEC_INV_157 Z_157 decode_157 vdd gnd pinv_0
XDEC_INV_158 Z_158 decode_158 vdd gnd pinv_0
XDEC_INV_159 Z_159 decode_159 vdd gnd pinv_0
XDEC_INV_160 Z_160 decode_160 vdd gnd pinv_0
XDEC_INV_161 Z_161 decode_161 vdd gnd pinv_0
XDEC_INV_162 Z_162 decode_162 vdd gnd pinv_0
XDEC_INV_163 Z_163 decode_163 vdd gnd pinv_0
XDEC_INV_164 Z_164 decode_164 vdd gnd pinv_0
XDEC_INV_165 Z_165 decode_165 vdd gnd pinv_0
XDEC_INV_166 Z_166 decode_166 vdd gnd pinv_0
XDEC_INV_167 Z_167 decode_167 vdd gnd pinv_0
XDEC_INV_168 Z_168 decode_168 vdd gnd pinv_0
XDEC_INV_169 Z_169 decode_169 vdd gnd pinv_0
XDEC_INV_170 Z_170 decode_170 vdd gnd pinv_0
XDEC_INV_171 Z_171 decode_171 vdd gnd pinv_0
XDEC_INV_172 Z_172 decode_172 vdd gnd pinv_0
XDEC_INV_173 Z_173 decode_173 vdd gnd pinv_0
XDEC_INV_174 Z_174 decode_174 vdd gnd pinv_0
XDEC_INV_175 Z_175 decode_175 vdd gnd pinv_0
XDEC_INV_176 Z_176 decode_176 vdd gnd pinv_0
XDEC_INV_177 Z_177 decode_177 vdd gnd pinv_0
XDEC_INV_178 Z_178 decode_178 vdd gnd pinv_0
XDEC_INV_179 Z_179 decode_179 vdd gnd pinv_0
XDEC_INV_180 Z_180 decode_180 vdd gnd pinv_0
XDEC_INV_181 Z_181 decode_181 vdd gnd pinv_0
XDEC_INV_182 Z_182 decode_182 vdd gnd pinv_0
XDEC_INV_183 Z_183 decode_183 vdd gnd pinv_0
XDEC_INV_184 Z_184 decode_184 vdd gnd pinv_0
XDEC_INV_185 Z_185 decode_185 vdd gnd pinv_0
XDEC_INV_186 Z_186 decode_186 vdd gnd pinv_0
XDEC_INV_187 Z_187 decode_187 vdd gnd pinv_0
XDEC_INV_188 Z_188 decode_188 vdd gnd pinv_0
XDEC_INV_189 Z_189 decode_189 vdd gnd pinv_0
XDEC_INV_190 Z_190 decode_190 vdd gnd pinv_0
XDEC_INV_191 Z_191 decode_191 vdd gnd pinv_0
XDEC_INV_192 Z_192 decode_192 vdd gnd pinv_0
XDEC_INV_193 Z_193 decode_193 vdd gnd pinv_0
XDEC_INV_194 Z_194 decode_194 vdd gnd pinv_0
XDEC_INV_195 Z_195 decode_195 vdd gnd pinv_0
XDEC_INV_196 Z_196 decode_196 vdd gnd pinv_0
XDEC_INV_197 Z_197 decode_197 vdd gnd pinv_0
XDEC_INV_198 Z_198 decode_198 vdd gnd pinv_0
XDEC_INV_199 Z_199 decode_199 vdd gnd pinv_0
XDEC_INV_200 Z_200 decode_200 vdd gnd pinv_0
XDEC_INV_201 Z_201 decode_201 vdd gnd pinv_0
XDEC_INV_202 Z_202 decode_202 vdd gnd pinv_0
XDEC_INV_203 Z_203 decode_203 vdd gnd pinv_0
XDEC_INV_204 Z_204 decode_204 vdd gnd pinv_0
XDEC_INV_205 Z_205 decode_205 vdd gnd pinv_0
XDEC_INV_206 Z_206 decode_206 vdd gnd pinv_0
XDEC_INV_207 Z_207 decode_207 vdd gnd pinv_0
XDEC_INV_208 Z_208 decode_208 vdd gnd pinv_0
XDEC_INV_209 Z_209 decode_209 vdd gnd pinv_0
XDEC_INV_210 Z_210 decode_210 vdd gnd pinv_0
XDEC_INV_211 Z_211 decode_211 vdd gnd pinv_0
XDEC_INV_212 Z_212 decode_212 vdd gnd pinv_0
XDEC_INV_213 Z_213 decode_213 vdd gnd pinv_0
XDEC_INV_214 Z_214 decode_214 vdd gnd pinv_0
XDEC_INV_215 Z_215 decode_215 vdd gnd pinv_0
XDEC_INV_216 Z_216 decode_216 vdd gnd pinv_0
XDEC_INV_217 Z_217 decode_217 vdd gnd pinv_0
XDEC_INV_218 Z_218 decode_218 vdd gnd pinv_0
XDEC_INV_219 Z_219 decode_219 vdd gnd pinv_0
XDEC_INV_220 Z_220 decode_220 vdd gnd pinv_0
XDEC_INV_221 Z_221 decode_221 vdd gnd pinv_0
XDEC_INV_222 Z_222 decode_222 vdd gnd pinv_0
XDEC_INV_223 Z_223 decode_223 vdd gnd pinv_0
XDEC_INV_224 Z_224 decode_224 vdd gnd pinv_0
XDEC_INV_225 Z_225 decode_225 vdd gnd pinv_0
XDEC_INV_226 Z_226 decode_226 vdd gnd pinv_0
XDEC_INV_227 Z_227 decode_227 vdd gnd pinv_0
XDEC_INV_228 Z_228 decode_228 vdd gnd pinv_0
XDEC_INV_229 Z_229 decode_229 vdd gnd pinv_0
XDEC_INV_230 Z_230 decode_230 vdd gnd pinv_0
XDEC_INV_231 Z_231 decode_231 vdd gnd pinv_0
XDEC_INV_232 Z_232 decode_232 vdd gnd pinv_0
XDEC_INV_233 Z_233 decode_233 vdd gnd pinv_0
XDEC_INV_234 Z_234 decode_234 vdd gnd pinv_0
XDEC_INV_235 Z_235 decode_235 vdd gnd pinv_0
XDEC_INV_236 Z_236 decode_236 vdd gnd pinv_0
XDEC_INV_237 Z_237 decode_237 vdd gnd pinv_0
XDEC_INV_238 Z_238 decode_238 vdd gnd pinv_0
XDEC_INV_239 Z_239 decode_239 vdd gnd pinv_0
XDEC_INV_240 Z_240 decode_240 vdd gnd pinv_0
XDEC_INV_241 Z_241 decode_241 vdd gnd pinv_0
XDEC_INV_242 Z_242 decode_242 vdd gnd pinv_0
XDEC_INV_243 Z_243 decode_243 vdd gnd pinv_0
XDEC_INV_244 Z_244 decode_244 vdd gnd pinv_0
XDEC_INV_245 Z_245 decode_245 vdd gnd pinv_0
XDEC_INV_246 Z_246 decode_246 vdd gnd pinv_0
XDEC_INV_247 Z_247 decode_247 vdd gnd pinv_0
XDEC_INV_248 Z_248 decode_248 vdd gnd pinv_0
XDEC_INV_249 Z_249 decode_249 vdd gnd pinv_0
XDEC_INV_250 Z_250 decode_250 vdd gnd pinv_0
XDEC_INV_251 Z_251 decode_251 vdd gnd pinv_0
XDEC_INV_252 Z_252 decode_252 vdd gnd pinv_0
XDEC_INV_253 Z_253 decode_253 vdd gnd pinv_0
XDEC_INV_254 Z_254 decode_254 vdd gnd pinv_0
XDEC_INV_255 Z_255 decode_255 vdd gnd pinv_0
.ENDS hierarchical_decoder_0

.SUBCKT pinv_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_1

* ptx M{0} {1} nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_2

* ptx M{0} {1} nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_3

* ptx M{0} {1} nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

.SUBCKT pinv_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_4

* ptx M{0} {1} nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

.SUBCKT pinv_5 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_5

.SUBCKT pdriver_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_1
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_1
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_1
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_2
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_3
Xbuf_inv6 Zb5_int Zb6_int vdd gnd pinv_4
Xbuf_inv7 Zb6_int Z vdd gnd pinv_5
.ENDS pdriver_0

.SUBCKT wordline_driver_0 in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67 in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78 in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89 in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100 in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110 in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120 in_121 in_122 in_123 in_124 in_125 in_126 in_127 in_128 in_129 in_130 in_131 in_132 in_133 in_134 in_135 in_136 in_137 in_138 in_139 in_140 in_141 in_142 in_143 in_144 in_145 in_146 in_147 in_148 in_149 in_150 in_151 in_152 in_153 in_154 in_155 in_156 in_157 in_158 in_159 in_160 in_161 in_162 in_163 in_164 in_165 in_166 in_167 in_168 in_169 in_170 in_171 in_172 in_173 in_174 in_175 in_176 in_177 in_178 in_179 in_180 in_181 in_182 in_183 in_184 in_185 in_186 in_187 in_188 in_189 in_190 in_191 in_192 in_193 in_194 in_195 in_196 in_197 in_198 in_199 in_200 in_201 in_202 in_203 in_204 in_205 in_206 in_207 in_208 in_209 in_210 in_211 in_212 in_213 in_214 in_215 in_216 in_217 in_218 in_219 in_220 in_221 in_222 in_223 in_224 in_225 in_226 in_227 in_228 in_229 in_230 in_231 in_232 in_233 in_234 in_235 in_236 in_237 in_238 in_239 in_240 in_241 in_242 in_243 in_244 in_245 in_246 in_247 in_248 in_249 in_250 in_251 in_252 in_253 in_254 in_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* INPUT : in_128 
* INPUT : in_129 
* INPUT : in_130 
* INPUT : in_131 
* INPUT : in_132 
* INPUT : in_133 
* INPUT : in_134 
* INPUT : in_135 
* INPUT : in_136 
* INPUT : in_137 
* INPUT : in_138 
* INPUT : in_139 
* INPUT : in_140 
* INPUT : in_141 
* INPUT : in_142 
* INPUT : in_143 
* INPUT : in_144 
* INPUT : in_145 
* INPUT : in_146 
* INPUT : in_147 
* INPUT : in_148 
* INPUT : in_149 
* INPUT : in_150 
* INPUT : in_151 
* INPUT : in_152 
* INPUT : in_153 
* INPUT : in_154 
* INPUT : in_155 
* INPUT : in_156 
* INPUT : in_157 
* INPUT : in_158 
* INPUT : in_159 
* INPUT : in_160 
* INPUT : in_161 
* INPUT : in_162 
* INPUT : in_163 
* INPUT : in_164 
* INPUT : in_165 
* INPUT : in_166 
* INPUT : in_167 
* INPUT : in_168 
* INPUT : in_169 
* INPUT : in_170 
* INPUT : in_171 
* INPUT : in_172 
* INPUT : in_173 
* INPUT : in_174 
* INPUT : in_175 
* INPUT : in_176 
* INPUT : in_177 
* INPUT : in_178 
* INPUT : in_179 
* INPUT : in_180 
* INPUT : in_181 
* INPUT : in_182 
* INPUT : in_183 
* INPUT : in_184 
* INPUT : in_185 
* INPUT : in_186 
* INPUT : in_187 
* INPUT : in_188 
* INPUT : in_189 
* INPUT : in_190 
* INPUT : in_191 
* INPUT : in_192 
* INPUT : in_193 
* INPUT : in_194 
* INPUT : in_195 
* INPUT : in_196 
* INPUT : in_197 
* INPUT : in_198 
* INPUT : in_199 
* INPUT : in_200 
* INPUT : in_201 
* INPUT : in_202 
* INPUT : in_203 
* INPUT : in_204 
* INPUT : in_205 
* INPUT : in_206 
* INPUT : in_207 
* INPUT : in_208 
* INPUT : in_209 
* INPUT : in_210 
* INPUT : in_211 
* INPUT : in_212 
* INPUT : in_213 
* INPUT : in_214 
* INPUT : in_215 
* INPUT : in_216 
* INPUT : in_217 
* INPUT : in_218 
* INPUT : in_219 
* INPUT : in_220 
* INPUT : in_221 
* INPUT : in_222 
* INPUT : in_223 
* INPUT : in_224 
* INPUT : in_225 
* INPUT : in_226 
* INPUT : in_227 
* INPUT : in_228 
* INPUT : in_229 
* INPUT : in_230 
* INPUT : in_231 
* INPUT : in_232 
* INPUT : in_233 
* INPUT : in_234 
* INPUT : in_235 
* INPUT : in_236 
* INPUT : in_237 
* INPUT : in_238 
* INPUT : in_239 
* INPUT : in_240 
* INPUT : in_241 
* INPUT : in_242 
* INPUT : in_243 
* INPUT : in_244 
* INPUT : in_245 
* INPUT : in_246 
* INPUT : in_247 
* INPUT : in_248 
* INPUT : in_249 
* INPUT : in_250 
* INPUT : in_251 
* INPUT : in_252 
* INPUT : in_253 
* INPUT : in_254 
* INPUT : in_255 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* OUTPUT: wl_128 
* OUTPUT: wl_129 
* OUTPUT: wl_130 
* OUTPUT: wl_131 
* OUTPUT: wl_132 
* OUTPUT: wl_133 
* OUTPUT: wl_134 
* OUTPUT: wl_135 
* OUTPUT: wl_136 
* OUTPUT: wl_137 
* OUTPUT: wl_138 
* OUTPUT: wl_139 
* OUTPUT: wl_140 
* OUTPUT: wl_141 
* OUTPUT: wl_142 
* OUTPUT: wl_143 
* OUTPUT: wl_144 
* OUTPUT: wl_145 
* OUTPUT: wl_146 
* OUTPUT: wl_147 
* OUTPUT: wl_148 
* OUTPUT: wl_149 
* OUTPUT: wl_150 
* OUTPUT: wl_151 
* OUTPUT: wl_152 
* OUTPUT: wl_153 
* OUTPUT: wl_154 
* OUTPUT: wl_155 
* OUTPUT: wl_156 
* OUTPUT: wl_157 
* OUTPUT: wl_158 
* OUTPUT: wl_159 
* OUTPUT: wl_160 
* OUTPUT: wl_161 
* OUTPUT: wl_162 
* OUTPUT: wl_163 
* OUTPUT: wl_164 
* OUTPUT: wl_165 
* OUTPUT: wl_166 
* OUTPUT: wl_167 
* OUTPUT: wl_168 
* OUTPUT: wl_169 
* OUTPUT: wl_170 
* OUTPUT: wl_171 
* OUTPUT: wl_172 
* OUTPUT: wl_173 
* OUTPUT: wl_174 
* OUTPUT: wl_175 
* OUTPUT: wl_176 
* OUTPUT: wl_177 
* OUTPUT: wl_178 
* OUTPUT: wl_179 
* OUTPUT: wl_180 
* OUTPUT: wl_181 
* OUTPUT: wl_182 
* OUTPUT: wl_183 
* OUTPUT: wl_184 
* OUTPUT: wl_185 
* OUTPUT: wl_186 
* OUTPUT: wl_187 
* OUTPUT: wl_188 
* OUTPUT: wl_189 
* OUTPUT: wl_190 
* OUTPUT: wl_191 
* OUTPUT: wl_192 
* OUTPUT: wl_193 
* OUTPUT: wl_194 
* OUTPUT: wl_195 
* OUTPUT: wl_196 
* OUTPUT: wl_197 
* OUTPUT: wl_198 
* OUTPUT: wl_199 
* OUTPUT: wl_200 
* OUTPUT: wl_201 
* OUTPUT: wl_202 
* OUTPUT: wl_203 
* OUTPUT: wl_204 
* OUTPUT: wl_205 
* OUTPUT: wl_206 
* OUTPUT: wl_207 
* OUTPUT: wl_208 
* OUTPUT: wl_209 
* OUTPUT: wl_210 
* OUTPUT: wl_211 
* OUTPUT: wl_212 
* OUTPUT: wl_213 
* OUTPUT: wl_214 
* OUTPUT: wl_215 
* OUTPUT: wl_216 
* OUTPUT: wl_217 
* OUTPUT: wl_218 
* OUTPUT: wl_219 
* OUTPUT: wl_220 
* OUTPUT: wl_221 
* OUTPUT: wl_222 
* OUTPUT: wl_223 
* OUTPUT: wl_224 
* OUTPUT: wl_225 
* OUTPUT: wl_226 
* OUTPUT: wl_227 
* OUTPUT: wl_228 
* OUTPUT: wl_229 
* OUTPUT: wl_230 
* OUTPUT: wl_231 
* OUTPUT: wl_232 
* OUTPUT: wl_233 
* OUTPUT: wl_234 
* OUTPUT: wl_235 
* OUTPUT: wl_236 
* OUTPUT: wl_237 
* OUTPUT: wl_238 
* OUTPUT: wl_239 
* OUTPUT: wl_240 
* OUTPUT: wl_241 
* OUTPUT: wl_242 
* OUTPUT: wl_243 
* OUTPUT: wl_244 
* OUTPUT: wl_245 
* OUTPUT: wl_246 
* OUTPUT: wl_247 
* OUTPUT: wl_248 
* OUTPUT: wl_249 
* OUTPUT: wl_250 
* OUTPUT: wl_251 
* OUTPUT: wl_252 
* OUTPUT: wl_253 
* OUTPUT: wl_254 
* OUTPUT: wl_255 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 256 cols: 256
Xwl_driver_nand0 en in_0 wl_bar_0 vdd gnd pnand2_0
Xwl_driver_inv0 wl_bar_0 wl_0 vdd gnd pdriver_0
Xwl_driver_nand1 en in_1 wl_bar_1 vdd gnd pnand2_0
Xwl_driver_inv1 wl_bar_1 wl_1 vdd gnd pdriver_0
Xwl_driver_nand2 en in_2 wl_bar_2 vdd gnd pnand2_0
Xwl_driver_inv2 wl_bar_2 wl_2 vdd gnd pdriver_0
Xwl_driver_nand3 en in_3 wl_bar_3 vdd gnd pnand2_0
Xwl_driver_inv3 wl_bar_3 wl_3 vdd gnd pdriver_0
Xwl_driver_nand4 en in_4 wl_bar_4 vdd gnd pnand2_0
Xwl_driver_inv4 wl_bar_4 wl_4 vdd gnd pdriver_0
Xwl_driver_nand5 en in_5 wl_bar_5 vdd gnd pnand2_0
Xwl_driver_inv5 wl_bar_5 wl_5 vdd gnd pdriver_0
Xwl_driver_nand6 en in_6 wl_bar_6 vdd gnd pnand2_0
Xwl_driver_inv6 wl_bar_6 wl_6 vdd gnd pdriver_0
Xwl_driver_nand7 en in_7 wl_bar_7 vdd gnd pnand2_0
Xwl_driver_inv7 wl_bar_7 wl_7 vdd gnd pdriver_0
Xwl_driver_nand8 en in_8 wl_bar_8 vdd gnd pnand2_0
Xwl_driver_inv8 wl_bar_8 wl_8 vdd gnd pdriver_0
Xwl_driver_nand9 en in_9 wl_bar_9 vdd gnd pnand2_0
Xwl_driver_inv9 wl_bar_9 wl_9 vdd gnd pdriver_0
Xwl_driver_nand10 en in_10 wl_bar_10 vdd gnd pnand2_0
Xwl_driver_inv10 wl_bar_10 wl_10 vdd gnd pdriver_0
Xwl_driver_nand11 en in_11 wl_bar_11 vdd gnd pnand2_0
Xwl_driver_inv11 wl_bar_11 wl_11 vdd gnd pdriver_0
Xwl_driver_nand12 en in_12 wl_bar_12 vdd gnd pnand2_0
Xwl_driver_inv12 wl_bar_12 wl_12 vdd gnd pdriver_0
Xwl_driver_nand13 en in_13 wl_bar_13 vdd gnd pnand2_0
Xwl_driver_inv13 wl_bar_13 wl_13 vdd gnd pdriver_0
Xwl_driver_nand14 en in_14 wl_bar_14 vdd gnd pnand2_0
Xwl_driver_inv14 wl_bar_14 wl_14 vdd gnd pdriver_0
Xwl_driver_nand15 en in_15 wl_bar_15 vdd gnd pnand2_0
Xwl_driver_inv15 wl_bar_15 wl_15 vdd gnd pdriver_0
Xwl_driver_nand16 en in_16 wl_bar_16 vdd gnd pnand2_0
Xwl_driver_inv16 wl_bar_16 wl_16 vdd gnd pdriver_0
Xwl_driver_nand17 en in_17 wl_bar_17 vdd gnd pnand2_0
Xwl_driver_inv17 wl_bar_17 wl_17 vdd gnd pdriver_0
Xwl_driver_nand18 en in_18 wl_bar_18 vdd gnd pnand2_0
Xwl_driver_inv18 wl_bar_18 wl_18 vdd gnd pdriver_0
Xwl_driver_nand19 en in_19 wl_bar_19 vdd gnd pnand2_0
Xwl_driver_inv19 wl_bar_19 wl_19 vdd gnd pdriver_0
Xwl_driver_nand20 en in_20 wl_bar_20 vdd gnd pnand2_0
Xwl_driver_inv20 wl_bar_20 wl_20 vdd gnd pdriver_0
Xwl_driver_nand21 en in_21 wl_bar_21 vdd gnd pnand2_0
Xwl_driver_inv21 wl_bar_21 wl_21 vdd gnd pdriver_0
Xwl_driver_nand22 en in_22 wl_bar_22 vdd gnd pnand2_0
Xwl_driver_inv22 wl_bar_22 wl_22 vdd gnd pdriver_0
Xwl_driver_nand23 en in_23 wl_bar_23 vdd gnd pnand2_0
Xwl_driver_inv23 wl_bar_23 wl_23 vdd gnd pdriver_0
Xwl_driver_nand24 en in_24 wl_bar_24 vdd gnd pnand2_0
Xwl_driver_inv24 wl_bar_24 wl_24 vdd gnd pdriver_0
Xwl_driver_nand25 en in_25 wl_bar_25 vdd gnd pnand2_0
Xwl_driver_inv25 wl_bar_25 wl_25 vdd gnd pdriver_0
Xwl_driver_nand26 en in_26 wl_bar_26 vdd gnd pnand2_0
Xwl_driver_inv26 wl_bar_26 wl_26 vdd gnd pdriver_0
Xwl_driver_nand27 en in_27 wl_bar_27 vdd gnd pnand2_0
Xwl_driver_inv27 wl_bar_27 wl_27 vdd gnd pdriver_0
Xwl_driver_nand28 en in_28 wl_bar_28 vdd gnd pnand2_0
Xwl_driver_inv28 wl_bar_28 wl_28 vdd gnd pdriver_0
Xwl_driver_nand29 en in_29 wl_bar_29 vdd gnd pnand2_0
Xwl_driver_inv29 wl_bar_29 wl_29 vdd gnd pdriver_0
Xwl_driver_nand30 en in_30 wl_bar_30 vdd gnd pnand2_0
Xwl_driver_inv30 wl_bar_30 wl_30 vdd gnd pdriver_0
Xwl_driver_nand31 en in_31 wl_bar_31 vdd gnd pnand2_0
Xwl_driver_inv31 wl_bar_31 wl_31 vdd gnd pdriver_0
Xwl_driver_nand32 en in_32 wl_bar_32 vdd gnd pnand2_0
Xwl_driver_inv32 wl_bar_32 wl_32 vdd gnd pdriver_0
Xwl_driver_nand33 en in_33 wl_bar_33 vdd gnd pnand2_0
Xwl_driver_inv33 wl_bar_33 wl_33 vdd gnd pdriver_0
Xwl_driver_nand34 en in_34 wl_bar_34 vdd gnd pnand2_0
Xwl_driver_inv34 wl_bar_34 wl_34 vdd gnd pdriver_0
Xwl_driver_nand35 en in_35 wl_bar_35 vdd gnd pnand2_0
Xwl_driver_inv35 wl_bar_35 wl_35 vdd gnd pdriver_0
Xwl_driver_nand36 en in_36 wl_bar_36 vdd gnd pnand2_0
Xwl_driver_inv36 wl_bar_36 wl_36 vdd gnd pdriver_0
Xwl_driver_nand37 en in_37 wl_bar_37 vdd gnd pnand2_0
Xwl_driver_inv37 wl_bar_37 wl_37 vdd gnd pdriver_0
Xwl_driver_nand38 en in_38 wl_bar_38 vdd gnd pnand2_0
Xwl_driver_inv38 wl_bar_38 wl_38 vdd gnd pdriver_0
Xwl_driver_nand39 en in_39 wl_bar_39 vdd gnd pnand2_0
Xwl_driver_inv39 wl_bar_39 wl_39 vdd gnd pdriver_0
Xwl_driver_nand40 en in_40 wl_bar_40 vdd gnd pnand2_0
Xwl_driver_inv40 wl_bar_40 wl_40 vdd gnd pdriver_0
Xwl_driver_nand41 en in_41 wl_bar_41 vdd gnd pnand2_0
Xwl_driver_inv41 wl_bar_41 wl_41 vdd gnd pdriver_0
Xwl_driver_nand42 en in_42 wl_bar_42 vdd gnd pnand2_0
Xwl_driver_inv42 wl_bar_42 wl_42 vdd gnd pdriver_0
Xwl_driver_nand43 en in_43 wl_bar_43 vdd gnd pnand2_0
Xwl_driver_inv43 wl_bar_43 wl_43 vdd gnd pdriver_0
Xwl_driver_nand44 en in_44 wl_bar_44 vdd gnd pnand2_0
Xwl_driver_inv44 wl_bar_44 wl_44 vdd gnd pdriver_0
Xwl_driver_nand45 en in_45 wl_bar_45 vdd gnd pnand2_0
Xwl_driver_inv45 wl_bar_45 wl_45 vdd gnd pdriver_0
Xwl_driver_nand46 en in_46 wl_bar_46 vdd gnd pnand2_0
Xwl_driver_inv46 wl_bar_46 wl_46 vdd gnd pdriver_0
Xwl_driver_nand47 en in_47 wl_bar_47 vdd gnd pnand2_0
Xwl_driver_inv47 wl_bar_47 wl_47 vdd gnd pdriver_0
Xwl_driver_nand48 en in_48 wl_bar_48 vdd gnd pnand2_0
Xwl_driver_inv48 wl_bar_48 wl_48 vdd gnd pdriver_0
Xwl_driver_nand49 en in_49 wl_bar_49 vdd gnd pnand2_0
Xwl_driver_inv49 wl_bar_49 wl_49 vdd gnd pdriver_0
Xwl_driver_nand50 en in_50 wl_bar_50 vdd gnd pnand2_0
Xwl_driver_inv50 wl_bar_50 wl_50 vdd gnd pdriver_0
Xwl_driver_nand51 en in_51 wl_bar_51 vdd gnd pnand2_0
Xwl_driver_inv51 wl_bar_51 wl_51 vdd gnd pdriver_0
Xwl_driver_nand52 en in_52 wl_bar_52 vdd gnd pnand2_0
Xwl_driver_inv52 wl_bar_52 wl_52 vdd gnd pdriver_0
Xwl_driver_nand53 en in_53 wl_bar_53 vdd gnd pnand2_0
Xwl_driver_inv53 wl_bar_53 wl_53 vdd gnd pdriver_0
Xwl_driver_nand54 en in_54 wl_bar_54 vdd gnd pnand2_0
Xwl_driver_inv54 wl_bar_54 wl_54 vdd gnd pdriver_0
Xwl_driver_nand55 en in_55 wl_bar_55 vdd gnd pnand2_0
Xwl_driver_inv55 wl_bar_55 wl_55 vdd gnd pdriver_0
Xwl_driver_nand56 en in_56 wl_bar_56 vdd gnd pnand2_0
Xwl_driver_inv56 wl_bar_56 wl_56 vdd gnd pdriver_0
Xwl_driver_nand57 en in_57 wl_bar_57 vdd gnd pnand2_0
Xwl_driver_inv57 wl_bar_57 wl_57 vdd gnd pdriver_0
Xwl_driver_nand58 en in_58 wl_bar_58 vdd gnd pnand2_0
Xwl_driver_inv58 wl_bar_58 wl_58 vdd gnd pdriver_0
Xwl_driver_nand59 en in_59 wl_bar_59 vdd gnd pnand2_0
Xwl_driver_inv59 wl_bar_59 wl_59 vdd gnd pdriver_0
Xwl_driver_nand60 en in_60 wl_bar_60 vdd gnd pnand2_0
Xwl_driver_inv60 wl_bar_60 wl_60 vdd gnd pdriver_0
Xwl_driver_nand61 en in_61 wl_bar_61 vdd gnd pnand2_0
Xwl_driver_inv61 wl_bar_61 wl_61 vdd gnd pdriver_0
Xwl_driver_nand62 en in_62 wl_bar_62 vdd gnd pnand2_0
Xwl_driver_inv62 wl_bar_62 wl_62 vdd gnd pdriver_0
Xwl_driver_nand63 en in_63 wl_bar_63 vdd gnd pnand2_0
Xwl_driver_inv63 wl_bar_63 wl_63 vdd gnd pdriver_0
Xwl_driver_nand64 en in_64 wl_bar_64 vdd gnd pnand2_0
Xwl_driver_inv64 wl_bar_64 wl_64 vdd gnd pdriver_0
Xwl_driver_nand65 en in_65 wl_bar_65 vdd gnd pnand2_0
Xwl_driver_inv65 wl_bar_65 wl_65 vdd gnd pdriver_0
Xwl_driver_nand66 en in_66 wl_bar_66 vdd gnd pnand2_0
Xwl_driver_inv66 wl_bar_66 wl_66 vdd gnd pdriver_0
Xwl_driver_nand67 en in_67 wl_bar_67 vdd gnd pnand2_0
Xwl_driver_inv67 wl_bar_67 wl_67 vdd gnd pdriver_0
Xwl_driver_nand68 en in_68 wl_bar_68 vdd gnd pnand2_0
Xwl_driver_inv68 wl_bar_68 wl_68 vdd gnd pdriver_0
Xwl_driver_nand69 en in_69 wl_bar_69 vdd gnd pnand2_0
Xwl_driver_inv69 wl_bar_69 wl_69 vdd gnd pdriver_0
Xwl_driver_nand70 en in_70 wl_bar_70 vdd gnd pnand2_0
Xwl_driver_inv70 wl_bar_70 wl_70 vdd gnd pdriver_0
Xwl_driver_nand71 en in_71 wl_bar_71 vdd gnd pnand2_0
Xwl_driver_inv71 wl_bar_71 wl_71 vdd gnd pdriver_0
Xwl_driver_nand72 en in_72 wl_bar_72 vdd gnd pnand2_0
Xwl_driver_inv72 wl_bar_72 wl_72 vdd gnd pdriver_0
Xwl_driver_nand73 en in_73 wl_bar_73 vdd gnd pnand2_0
Xwl_driver_inv73 wl_bar_73 wl_73 vdd gnd pdriver_0
Xwl_driver_nand74 en in_74 wl_bar_74 vdd gnd pnand2_0
Xwl_driver_inv74 wl_bar_74 wl_74 vdd gnd pdriver_0
Xwl_driver_nand75 en in_75 wl_bar_75 vdd gnd pnand2_0
Xwl_driver_inv75 wl_bar_75 wl_75 vdd gnd pdriver_0
Xwl_driver_nand76 en in_76 wl_bar_76 vdd gnd pnand2_0
Xwl_driver_inv76 wl_bar_76 wl_76 vdd gnd pdriver_0
Xwl_driver_nand77 en in_77 wl_bar_77 vdd gnd pnand2_0
Xwl_driver_inv77 wl_bar_77 wl_77 vdd gnd pdriver_0
Xwl_driver_nand78 en in_78 wl_bar_78 vdd gnd pnand2_0
Xwl_driver_inv78 wl_bar_78 wl_78 vdd gnd pdriver_0
Xwl_driver_nand79 en in_79 wl_bar_79 vdd gnd pnand2_0
Xwl_driver_inv79 wl_bar_79 wl_79 vdd gnd pdriver_0
Xwl_driver_nand80 en in_80 wl_bar_80 vdd gnd pnand2_0
Xwl_driver_inv80 wl_bar_80 wl_80 vdd gnd pdriver_0
Xwl_driver_nand81 en in_81 wl_bar_81 vdd gnd pnand2_0
Xwl_driver_inv81 wl_bar_81 wl_81 vdd gnd pdriver_0
Xwl_driver_nand82 en in_82 wl_bar_82 vdd gnd pnand2_0
Xwl_driver_inv82 wl_bar_82 wl_82 vdd gnd pdriver_0
Xwl_driver_nand83 en in_83 wl_bar_83 vdd gnd pnand2_0
Xwl_driver_inv83 wl_bar_83 wl_83 vdd gnd pdriver_0
Xwl_driver_nand84 en in_84 wl_bar_84 vdd gnd pnand2_0
Xwl_driver_inv84 wl_bar_84 wl_84 vdd gnd pdriver_0
Xwl_driver_nand85 en in_85 wl_bar_85 vdd gnd pnand2_0
Xwl_driver_inv85 wl_bar_85 wl_85 vdd gnd pdriver_0
Xwl_driver_nand86 en in_86 wl_bar_86 vdd gnd pnand2_0
Xwl_driver_inv86 wl_bar_86 wl_86 vdd gnd pdriver_0
Xwl_driver_nand87 en in_87 wl_bar_87 vdd gnd pnand2_0
Xwl_driver_inv87 wl_bar_87 wl_87 vdd gnd pdriver_0
Xwl_driver_nand88 en in_88 wl_bar_88 vdd gnd pnand2_0
Xwl_driver_inv88 wl_bar_88 wl_88 vdd gnd pdriver_0
Xwl_driver_nand89 en in_89 wl_bar_89 vdd gnd pnand2_0
Xwl_driver_inv89 wl_bar_89 wl_89 vdd gnd pdriver_0
Xwl_driver_nand90 en in_90 wl_bar_90 vdd gnd pnand2_0
Xwl_driver_inv90 wl_bar_90 wl_90 vdd gnd pdriver_0
Xwl_driver_nand91 en in_91 wl_bar_91 vdd gnd pnand2_0
Xwl_driver_inv91 wl_bar_91 wl_91 vdd gnd pdriver_0
Xwl_driver_nand92 en in_92 wl_bar_92 vdd gnd pnand2_0
Xwl_driver_inv92 wl_bar_92 wl_92 vdd gnd pdriver_0
Xwl_driver_nand93 en in_93 wl_bar_93 vdd gnd pnand2_0
Xwl_driver_inv93 wl_bar_93 wl_93 vdd gnd pdriver_0
Xwl_driver_nand94 en in_94 wl_bar_94 vdd gnd pnand2_0
Xwl_driver_inv94 wl_bar_94 wl_94 vdd gnd pdriver_0
Xwl_driver_nand95 en in_95 wl_bar_95 vdd gnd pnand2_0
Xwl_driver_inv95 wl_bar_95 wl_95 vdd gnd pdriver_0
Xwl_driver_nand96 en in_96 wl_bar_96 vdd gnd pnand2_0
Xwl_driver_inv96 wl_bar_96 wl_96 vdd gnd pdriver_0
Xwl_driver_nand97 en in_97 wl_bar_97 vdd gnd pnand2_0
Xwl_driver_inv97 wl_bar_97 wl_97 vdd gnd pdriver_0
Xwl_driver_nand98 en in_98 wl_bar_98 vdd gnd pnand2_0
Xwl_driver_inv98 wl_bar_98 wl_98 vdd gnd pdriver_0
Xwl_driver_nand99 en in_99 wl_bar_99 vdd gnd pnand2_0
Xwl_driver_inv99 wl_bar_99 wl_99 vdd gnd pdriver_0
Xwl_driver_nand100 en in_100 wl_bar_100 vdd gnd pnand2_0
Xwl_driver_inv100 wl_bar_100 wl_100 vdd gnd pdriver_0
Xwl_driver_nand101 en in_101 wl_bar_101 vdd gnd pnand2_0
Xwl_driver_inv101 wl_bar_101 wl_101 vdd gnd pdriver_0
Xwl_driver_nand102 en in_102 wl_bar_102 vdd gnd pnand2_0
Xwl_driver_inv102 wl_bar_102 wl_102 vdd gnd pdriver_0
Xwl_driver_nand103 en in_103 wl_bar_103 vdd gnd pnand2_0
Xwl_driver_inv103 wl_bar_103 wl_103 vdd gnd pdriver_0
Xwl_driver_nand104 en in_104 wl_bar_104 vdd gnd pnand2_0
Xwl_driver_inv104 wl_bar_104 wl_104 vdd gnd pdriver_0
Xwl_driver_nand105 en in_105 wl_bar_105 vdd gnd pnand2_0
Xwl_driver_inv105 wl_bar_105 wl_105 vdd gnd pdriver_0
Xwl_driver_nand106 en in_106 wl_bar_106 vdd gnd pnand2_0
Xwl_driver_inv106 wl_bar_106 wl_106 vdd gnd pdriver_0
Xwl_driver_nand107 en in_107 wl_bar_107 vdd gnd pnand2_0
Xwl_driver_inv107 wl_bar_107 wl_107 vdd gnd pdriver_0
Xwl_driver_nand108 en in_108 wl_bar_108 vdd gnd pnand2_0
Xwl_driver_inv108 wl_bar_108 wl_108 vdd gnd pdriver_0
Xwl_driver_nand109 en in_109 wl_bar_109 vdd gnd pnand2_0
Xwl_driver_inv109 wl_bar_109 wl_109 vdd gnd pdriver_0
Xwl_driver_nand110 en in_110 wl_bar_110 vdd gnd pnand2_0
Xwl_driver_inv110 wl_bar_110 wl_110 vdd gnd pdriver_0
Xwl_driver_nand111 en in_111 wl_bar_111 vdd gnd pnand2_0
Xwl_driver_inv111 wl_bar_111 wl_111 vdd gnd pdriver_0
Xwl_driver_nand112 en in_112 wl_bar_112 vdd gnd pnand2_0
Xwl_driver_inv112 wl_bar_112 wl_112 vdd gnd pdriver_0
Xwl_driver_nand113 en in_113 wl_bar_113 vdd gnd pnand2_0
Xwl_driver_inv113 wl_bar_113 wl_113 vdd gnd pdriver_0
Xwl_driver_nand114 en in_114 wl_bar_114 vdd gnd pnand2_0
Xwl_driver_inv114 wl_bar_114 wl_114 vdd gnd pdriver_0
Xwl_driver_nand115 en in_115 wl_bar_115 vdd gnd pnand2_0
Xwl_driver_inv115 wl_bar_115 wl_115 vdd gnd pdriver_0
Xwl_driver_nand116 en in_116 wl_bar_116 vdd gnd pnand2_0
Xwl_driver_inv116 wl_bar_116 wl_116 vdd gnd pdriver_0
Xwl_driver_nand117 en in_117 wl_bar_117 vdd gnd pnand2_0
Xwl_driver_inv117 wl_bar_117 wl_117 vdd gnd pdriver_0
Xwl_driver_nand118 en in_118 wl_bar_118 vdd gnd pnand2_0
Xwl_driver_inv118 wl_bar_118 wl_118 vdd gnd pdriver_0
Xwl_driver_nand119 en in_119 wl_bar_119 vdd gnd pnand2_0
Xwl_driver_inv119 wl_bar_119 wl_119 vdd gnd pdriver_0
Xwl_driver_nand120 en in_120 wl_bar_120 vdd gnd pnand2_0
Xwl_driver_inv120 wl_bar_120 wl_120 vdd gnd pdriver_0
Xwl_driver_nand121 en in_121 wl_bar_121 vdd gnd pnand2_0
Xwl_driver_inv121 wl_bar_121 wl_121 vdd gnd pdriver_0
Xwl_driver_nand122 en in_122 wl_bar_122 vdd gnd pnand2_0
Xwl_driver_inv122 wl_bar_122 wl_122 vdd gnd pdriver_0
Xwl_driver_nand123 en in_123 wl_bar_123 vdd gnd pnand2_0
Xwl_driver_inv123 wl_bar_123 wl_123 vdd gnd pdriver_0
Xwl_driver_nand124 en in_124 wl_bar_124 vdd gnd pnand2_0
Xwl_driver_inv124 wl_bar_124 wl_124 vdd gnd pdriver_0
Xwl_driver_nand125 en in_125 wl_bar_125 vdd gnd pnand2_0
Xwl_driver_inv125 wl_bar_125 wl_125 vdd gnd pdriver_0
Xwl_driver_nand126 en in_126 wl_bar_126 vdd gnd pnand2_0
Xwl_driver_inv126 wl_bar_126 wl_126 vdd gnd pdriver_0
Xwl_driver_nand127 en in_127 wl_bar_127 vdd gnd pnand2_0
Xwl_driver_inv127 wl_bar_127 wl_127 vdd gnd pdriver_0
Xwl_driver_nand128 en in_128 wl_bar_128 vdd gnd pnand2_0
Xwl_driver_inv128 wl_bar_128 wl_128 vdd gnd pdriver_0
Xwl_driver_nand129 en in_129 wl_bar_129 vdd gnd pnand2_0
Xwl_driver_inv129 wl_bar_129 wl_129 vdd gnd pdriver_0
Xwl_driver_nand130 en in_130 wl_bar_130 vdd gnd pnand2_0
Xwl_driver_inv130 wl_bar_130 wl_130 vdd gnd pdriver_0
Xwl_driver_nand131 en in_131 wl_bar_131 vdd gnd pnand2_0
Xwl_driver_inv131 wl_bar_131 wl_131 vdd gnd pdriver_0
Xwl_driver_nand132 en in_132 wl_bar_132 vdd gnd pnand2_0
Xwl_driver_inv132 wl_bar_132 wl_132 vdd gnd pdriver_0
Xwl_driver_nand133 en in_133 wl_bar_133 vdd gnd pnand2_0
Xwl_driver_inv133 wl_bar_133 wl_133 vdd gnd pdriver_0
Xwl_driver_nand134 en in_134 wl_bar_134 vdd gnd pnand2_0
Xwl_driver_inv134 wl_bar_134 wl_134 vdd gnd pdriver_0
Xwl_driver_nand135 en in_135 wl_bar_135 vdd gnd pnand2_0
Xwl_driver_inv135 wl_bar_135 wl_135 vdd gnd pdriver_0
Xwl_driver_nand136 en in_136 wl_bar_136 vdd gnd pnand2_0
Xwl_driver_inv136 wl_bar_136 wl_136 vdd gnd pdriver_0
Xwl_driver_nand137 en in_137 wl_bar_137 vdd gnd pnand2_0
Xwl_driver_inv137 wl_bar_137 wl_137 vdd gnd pdriver_0
Xwl_driver_nand138 en in_138 wl_bar_138 vdd gnd pnand2_0
Xwl_driver_inv138 wl_bar_138 wl_138 vdd gnd pdriver_0
Xwl_driver_nand139 en in_139 wl_bar_139 vdd gnd pnand2_0
Xwl_driver_inv139 wl_bar_139 wl_139 vdd gnd pdriver_0
Xwl_driver_nand140 en in_140 wl_bar_140 vdd gnd pnand2_0
Xwl_driver_inv140 wl_bar_140 wl_140 vdd gnd pdriver_0
Xwl_driver_nand141 en in_141 wl_bar_141 vdd gnd pnand2_0
Xwl_driver_inv141 wl_bar_141 wl_141 vdd gnd pdriver_0
Xwl_driver_nand142 en in_142 wl_bar_142 vdd gnd pnand2_0
Xwl_driver_inv142 wl_bar_142 wl_142 vdd gnd pdriver_0
Xwl_driver_nand143 en in_143 wl_bar_143 vdd gnd pnand2_0
Xwl_driver_inv143 wl_bar_143 wl_143 vdd gnd pdriver_0
Xwl_driver_nand144 en in_144 wl_bar_144 vdd gnd pnand2_0
Xwl_driver_inv144 wl_bar_144 wl_144 vdd gnd pdriver_0
Xwl_driver_nand145 en in_145 wl_bar_145 vdd gnd pnand2_0
Xwl_driver_inv145 wl_bar_145 wl_145 vdd gnd pdriver_0
Xwl_driver_nand146 en in_146 wl_bar_146 vdd gnd pnand2_0
Xwl_driver_inv146 wl_bar_146 wl_146 vdd gnd pdriver_0
Xwl_driver_nand147 en in_147 wl_bar_147 vdd gnd pnand2_0
Xwl_driver_inv147 wl_bar_147 wl_147 vdd gnd pdriver_0
Xwl_driver_nand148 en in_148 wl_bar_148 vdd gnd pnand2_0
Xwl_driver_inv148 wl_bar_148 wl_148 vdd gnd pdriver_0
Xwl_driver_nand149 en in_149 wl_bar_149 vdd gnd pnand2_0
Xwl_driver_inv149 wl_bar_149 wl_149 vdd gnd pdriver_0
Xwl_driver_nand150 en in_150 wl_bar_150 vdd gnd pnand2_0
Xwl_driver_inv150 wl_bar_150 wl_150 vdd gnd pdriver_0
Xwl_driver_nand151 en in_151 wl_bar_151 vdd gnd pnand2_0
Xwl_driver_inv151 wl_bar_151 wl_151 vdd gnd pdriver_0
Xwl_driver_nand152 en in_152 wl_bar_152 vdd gnd pnand2_0
Xwl_driver_inv152 wl_bar_152 wl_152 vdd gnd pdriver_0
Xwl_driver_nand153 en in_153 wl_bar_153 vdd gnd pnand2_0
Xwl_driver_inv153 wl_bar_153 wl_153 vdd gnd pdriver_0
Xwl_driver_nand154 en in_154 wl_bar_154 vdd gnd pnand2_0
Xwl_driver_inv154 wl_bar_154 wl_154 vdd gnd pdriver_0
Xwl_driver_nand155 en in_155 wl_bar_155 vdd gnd pnand2_0
Xwl_driver_inv155 wl_bar_155 wl_155 vdd gnd pdriver_0
Xwl_driver_nand156 en in_156 wl_bar_156 vdd gnd pnand2_0
Xwl_driver_inv156 wl_bar_156 wl_156 vdd gnd pdriver_0
Xwl_driver_nand157 en in_157 wl_bar_157 vdd gnd pnand2_0
Xwl_driver_inv157 wl_bar_157 wl_157 vdd gnd pdriver_0
Xwl_driver_nand158 en in_158 wl_bar_158 vdd gnd pnand2_0
Xwl_driver_inv158 wl_bar_158 wl_158 vdd gnd pdriver_0
Xwl_driver_nand159 en in_159 wl_bar_159 vdd gnd pnand2_0
Xwl_driver_inv159 wl_bar_159 wl_159 vdd gnd pdriver_0
Xwl_driver_nand160 en in_160 wl_bar_160 vdd gnd pnand2_0
Xwl_driver_inv160 wl_bar_160 wl_160 vdd gnd pdriver_0
Xwl_driver_nand161 en in_161 wl_bar_161 vdd gnd pnand2_0
Xwl_driver_inv161 wl_bar_161 wl_161 vdd gnd pdriver_0
Xwl_driver_nand162 en in_162 wl_bar_162 vdd gnd pnand2_0
Xwl_driver_inv162 wl_bar_162 wl_162 vdd gnd pdriver_0
Xwl_driver_nand163 en in_163 wl_bar_163 vdd gnd pnand2_0
Xwl_driver_inv163 wl_bar_163 wl_163 vdd gnd pdriver_0
Xwl_driver_nand164 en in_164 wl_bar_164 vdd gnd pnand2_0
Xwl_driver_inv164 wl_bar_164 wl_164 vdd gnd pdriver_0
Xwl_driver_nand165 en in_165 wl_bar_165 vdd gnd pnand2_0
Xwl_driver_inv165 wl_bar_165 wl_165 vdd gnd pdriver_0
Xwl_driver_nand166 en in_166 wl_bar_166 vdd gnd pnand2_0
Xwl_driver_inv166 wl_bar_166 wl_166 vdd gnd pdriver_0
Xwl_driver_nand167 en in_167 wl_bar_167 vdd gnd pnand2_0
Xwl_driver_inv167 wl_bar_167 wl_167 vdd gnd pdriver_0
Xwl_driver_nand168 en in_168 wl_bar_168 vdd gnd pnand2_0
Xwl_driver_inv168 wl_bar_168 wl_168 vdd gnd pdriver_0
Xwl_driver_nand169 en in_169 wl_bar_169 vdd gnd pnand2_0
Xwl_driver_inv169 wl_bar_169 wl_169 vdd gnd pdriver_0
Xwl_driver_nand170 en in_170 wl_bar_170 vdd gnd pnand2_0
Xwl_driver_inv170 wl_bar_170 wl_170 vdd gnd pdriver_0
Xwl_driver_nand171 en in_171 wl_bar_171 vdd gnd pnand2_0
Xwl_driver_inv171 wl_bar_171 wl_171 vdd gnd pdriver_0
Xwl_driver_nand172 en in_172 wl_bar_172 vdd gnd pnand2_0
Xwl_driver_inv172 wl_bar_172 wl_172 vdd gnd pdriver_0
Xwl_driver_nand173 en in_173 wl_bar_173 vdd gnd pnand2_0
Xwl_driver_inv173 wl_bar_173 wl_173 vdd gnd pdriver_0
Xwl_driver_nand174 en in_174 wl_bar_174 vdd gnd pnand2_0
Xwl_driver_inv174 wl_bar_174 wl_174 vdd gnd pdriver_0
Xwl_driver_nand175 en in_175 wl_bar_175 vdd gnd pnand2_0
Xwl_driver_inv175 wl_bar_175 wl_175 vdd gnd pdriver_0
Xwl_driver_nand176 en in_176 wl_bar_176 vdd gnd pnand2_0
Xwl_driver_inv176 wl_bar_176 wl_176 vdd gnd pdriver_0
Xwl_driver_nand177 en in_177 wl_bar_177 vdd gnd pnand2_0
Xwl_driver_inv177 wl_bar_177 wl_177 vdd gnd pdriver_0
Xwl_driver_nand178 en in_178 wl_bar_178 vdd gnd pnand2_0
Xwl_driver_inv178 wl_bar_178 wl_178 vdd gnd pdriver_0
Xwl_driver_nand179 en in_179 wl_bar_179 vdd gnd pnand2_0
Xwl_driver_inv179 wl_bar_179 wl_179 vdd gnd pdriver_0
Xwl_driver_nand180 en in_180 wl_bar_180 vdd gnd pnand2_0
Xwl_driver_inv180 wl_bar_180 wl_180 vdd gnd pdriver_0
Xwl_driver_nand181 en in_181 wl_bar_181 vdd gnd pnand2_0
Xwl_driver_inv181 wl_bar_181 wl_181 vdd gnd pdriver_0
Xwl_driver_nand182 en in_182 wl_bar_182 vdd gnd pnand2_0
Xwl_driver_inv182 wl_bar_182 wl_182 vdd gnd pdriver_0
Xwl_driver_nand183 en in_183 wl_bar_183 vdd gnd pnand2_0
Xwl_driver_inv183 wl_bar_183 wl_183 vdd gnd pdriver_0
Xwl_driver_nand184 en in_184 wl_bar_184 vdd gnd pnand2_0
Xwl_driver_inv184 wl_bar_184 wl_184 vdd gnd pdriver_0
Xwl_driver_nand185 en in_185 wl_bar_185 vdd gnd pnand2_0
Xwl_driver_inv185 wl_bar_185 wl_185 vdd gnd pdriver_0
Xwl_driver_nand186 en in_186 wl_bar_186 vdd gnd pnand2_0
Xwl_driver_inv186 wl_bar_186 wl_186 vdd gnd pdriver_0
Xwl_driver_nand187 en in_187 wl_bar_187 vdd gnd pnand2_0
Xwl_driver_inv187 wl_bar_187 wl_187 vdd gnd pdriver_0
Xwl_driver_nand188 en in_188 wl_bar_188 vdd gnd pnand2_0
Xwl_driver_inv188 wl_bar_188 wl_188 vdd gnd pdriver_0
Xwl_driver_nand189 en in_189 wl_bar_189 vdd gnd pnand2_0
Xwl_driver_inv189 wl_bar_189 wl_189 vdd gnd pdriver_0
Xwl_driver_nand190 en in_190 wl_bar_190 vdd gnd pnand2_0
Xwl_driver_inv190 wl_bar_190 wl_190 vdd gnd pdriver_0
Xwl_driver_nand191 en in_191 wl_bar_191 vdd gnd pnand2_0
Xwl_driver_inv191 wl_bar_191 wl_191 vdd gnd pdriver_0
Xwl_driver_nand192 en in_192 wl_bar_192 vdd gnd pnand2_0
Xwl_driver_inv192 wl_bar_192 wl_192 vdd gnd pdriver_0
Xwl_driver_nand193 en in_193 wl_bar_193 vdd gnd pnand2_0
Xwl_driver_inv193 wl_bar_193 wl_193 vdd gnd pdriver_0
Xwl_driver_nand194 en in_194 wl_bar_194 vdd gnd pnand2_0
Xwl_driver_inv194 wl_bar_194 wl_194 vdd gnd pdriver_0
Xwl_driver_nand195 en in_195 wl_bar_195 vdd gnd pnand2_0
Xwl_driver_inv195 wl_bar_195 wl_195 vdd gnd pdriver_0
Xwl_driver_nand196 en in_196 wl_bar_196 vdd gnd pnand2_0
Xwl_driver_inv196 wl_bar_196 wl_196 vdd gnd pdriver_0
Xwl_driver_nand197 en in_197 wl_bar_197 vdd gnd pnand2_0
Xwl_driver_inv197 wl_bar_197 wl_197 vdd gnd pdriver_0
Xwl_driver_nand198 en in_198 wl_bar_198 vdd gnd pnand2_0
Xwl_driver_inv198 wl_bar_198 wl_198 vdd gnd pdriver_0
Xwl_driver_nand199 en in_199 wl_bar_199 vdd gnd pnand2_0
Xwl_driver_inv199 wl_bar_199 wl_199 vdd gnd pdriver_0
Xwl_driver_nand200 en in_200 wl_bar_200 vdd gnd pnand2_0
Xwl_driver_inv200 wl_bar_200 wl_200 vdd gnd pdriver_0
Xwl_driver_nand201 en in_201 wl_bar_201 vdd gnd pnand2_0
Xwl_driver_inv201 wl_bar_201 wl_201 vdd gnd pdriver_0
Xwl_driver_nand202 en in_202 wl_bar_202 vdd gnd pnand2_0
Xwl_driver_inv202 wl_bar_202 wl_202 vdd gnd pdriver_0
Xwl_driver_nand203 en in_203 wl_bar_203 vdd gnd pnand2_0
Xwl_driver_inv203 wl_bar_203 wl_203 vdd gnd pdriver_0
Xwl_driver_nand204 en in_204 wl_bar_204 vdd gnd pnand2_0
Xwl_driver_inv204 wl_bar_204 wl_204 vdd gnd pdriver_0
Xwl_driver_nand205 en in_205 wl_bar_205 vdd gnd pnand2_0
Xwl_driver_inv205 wl_bar_205 wl_205 vdd gnd pdriver_0
Xwl_driver_nand206 en in_206 wl_bar_206 vdd gnd pnand2_0
Xwl_driver_inv206 wl_bar_206 wl_206 vdd gnd pdriver_0
Xwl_driver_nand207 en in_207 wl_bar_207 vdd gnd pnand2_0
Xwl_driver_inv207 wl_bar_207 wl_207 vdd gnd pdriver_0
Xwl_driver_nand208 en in_208 wl_bar_208 vdd gnd pnand2_0
Xwl_driver_inv208 wl_bar_208 wl_208 vdd gnd pdriver_0
Xwl_driver_nand209 en in_209 wl_bar_209 vdd gnd pnand2_0
Xwl_driver_inv209 wl_bar_209 wl_209 vdd gnd pdriver_0
Xwl_driver_nand210 en in_210 wl_bar_210 vdd gnd pnand2_0
Xwl_driver_inv210 wl_bar_210 wl_210 vdd gnd pdriver_0
Xwl_driver_nand211 en in_211 wl_bar_211 vdd gnd pnand2_0
Xwl_driver_inv211 wl_bar_211 wl_211 vdd gnd pdriver_0
Xwl_driver_nand212 en in_212 wl_bar_212 vdd gnd pnand2_0
Xwl_driver_inv212 wl_bar_212 wl_212 vdd gnd pdriver_0
Xwl_driver_nand213 en in_213 wl_bar_213 vdd gnd pnand2_0
Xwl_driver_inv213 wl_bar_213 wl_213 vdd gnd pdriver_0
Xwl_driver_nand214 en in_214 wl_bar_214 vdd gnd pnand2_0
Xwl_driver_inv214 wl_bar_214 wl_214 vdd gnd pdriver_0
Xwl_driver_nand215 en in_215 wl_bar_215 vdd gnd pnand2_0
Xwl_driver_inv215 wl_bar_215 wl_215 vdd gnd pdriver_0
Xwl_driver_nand216 en in_216 wl_bar_216 vdd gnd pnand2_0
Xwl_driver_inv216 wl_bar_216 wl_216 vdd gnd pdriver_0
Xwl_driver_nand217 en in_217 wl_bar_217 vdd gnd pnand2_0
Xwl_driver_inv217 wl_bar_217 wl_217 vdd gnd pdriver_0
Xwl_driver_nand218 en in_218 wl_bar_218 vdd gnd pnand2_0
Xwl_driver_inv218 wl_bar_218 wl_218 vdd gnd pdriver_0
Xwl_driver_nand219 en in_219 wl_bar_219 vdd gnd pnand2_0
Xwl_driver_inv219 wl_bar_219 wl_219 vdd gnd pdriver_0
Xwl_driver_nand220 en in_220 wl_bar_220 vdd gnd pnand2_0
Xwl_driver_inv220 wl_bar_220 wl_220 vdd gnd pdriver_0
Xwl_driver_nand221 en in_221 wl_bar_221 vdd gnd pnand2_0
Xwl_driver_inv221 wl_bar_221 wl_221 vdd gnd pdriver_0
Xwl_driver_nand222 en in_222 wl_bar_222 vdd gnd pnand2_0
Xwl_driver_inv222 wl_bar_222 wl_222 vdd gnd pdriver_0
Xwl_driver_nand223 en in_223 wl_bar_223 vdd gnd pnand2_0
Xwl_driver_inv223 wl_bar_223 wl_223 vdd gnd pdriver_0
Xwl_driver_nand224 en in_224 wl_bar_224 vdd gnd pnand2_0
Xwl_driver_inv224 wl_bar_224 wl_224 vdd gnd pdriver_0
Xwl_driver_nand225 en in_225 wl_bar_225 vdd gnd pnand2_0
Xwl_driver_inv225 wl_bar_225 wl_225 vdd gnd pdriver_0
Xwl_driver_nand226 en in_226 wl_bar_226 vdd gnd pnand2_0
Xwl_driver_inv226 wl_bar_226 wl_226 vdd gnd pdriver_0
Xwl_driver_nand227 en in_227 wl_bar_227 vdd gnd pnand2_0
Xwl_driver_inv227 wl_bar_227 wl_227 vdd gnd pdriver_0
Xwl_driver_nand228 en in_228 wl_bar_228 vdd gnd pnand2_0
Xwl_driver_inv228 wl_bar_228 wl_228 vdd gnd pdriver_0
Xwl_driver_nand229 en in_229 wl_bar_229 vdd gnd pnand2_0
Xwl_driver_inv229 wl_bar_229 wl_229 vdd gnd pdriver_0
Xwl_driver_nand230 en in_230 wl_bar_230 vdd gnd pnand2_0
Xwl_driver_inv230 wl_bar_230 wl_230 vdd gnd pdriver_0
Xwl_driver_nand231 en in_231 wl_bar_231 vdd gnd pnand2_0
Xwl_driver_inv231 wl_bar_231 wl_231 vdd gnd pdriver_0
Xwl_driver_nand232 en in_232 wl_bar_232 vdd gnd pnand2_0
Xwl_driver_inv232 wl_bar_232 wl_232 vdd gnd pdriver_0
Xwl_driver_nand233 en in_233 wl_bar_233 vdd gnd pnand2_0
Xwl_driver_inv233 wl_bar_233 wl_233 vdd gnd pdriver_0
Xwl_driver_nand234 en in_234 wl_bar_234 vdd gnd pnand2_0
Xwl_driver_inv234 wl_bar_234 wl_234 vdd gnd pdriver_0
Xwl_driver_nand235 en in_235 wl_bar_235 vdd gnd pnand2_0
Xwl_driver_inv235 wl_bar_235 wl_235 vdd gnd pdriver_0
Xwl_driver_nand236 en in_236 wl_bar_236 vdd gnd pnand2_0
Xwl_driver_inv236 wl_bar_236 wl_236 vdd gnd pdriver_0
Xwl_driver_nand237 en in_237 wl_bar_237 vdd gnd pnand2_0
Xwl_driver_inv237 wl_bar_237 wl_237 vdd gnd pdriver_0
Xwl_driver_nand238 en in_238 wl_bar_238 vdd gnd pnand2_0
Xwl_driver_inv238 wl_bar_238 wl_238 vdd gnd pdriver_0
Xwl_driver_nand239 en in_239 wl_bar_239 vdd gnd pnand2_0
Xwl_driver_inv239 wl_bar_239 wl_239 vdd gnd pdriver_0
Xwl_driver_nand240 en in_240 wl_bar_240 vdd gnd pnand2_0
Xwl_driver_inv240 wl_bar_240 wl_240 vdd gnd pdriver_0
Xwl_driver_nand241 en in_241 wl_bar_241 vdd gnd pnand2_0
Xwl_driver_inv241 wl_bar_241 wl_241 vdd gnd pdriver_0
Xwl_driver_nand242 en in_242 wl_bar_242 vdd gnd pnand2_0
Xwl_driver_inv242 wl_bar_242 wl_242 vdd gnd pdriver_0
Xwl_driver_nand243 en in_243 wl_bar_243 vdd gnd pnand2_0
Xwl_driver_inv243 wl_bar_243 wl_243 vdd gnd pdriver_0
Xwl_driver_nand244 en in_244 wl_bar_244 vdd gnd pnand2_0
Xwl_driver_inv244 wl_bar_244 wl_244 vdd gnd pdriver_0
Xwl_driver_nand245 en in_245 wl_bar_245 vdd gnd pnand2_0
Xwl_driver_inv245 wl_bar_245 wl_245 vdd gnd pdriver_0
Xwl_driver_nand246 en in_246 wl_bar_246 vdd gnd pnand2_0
Xwl_driver_inv246 wl_bar_246 wl_246 vdd gnd pdriver_0
Xwl_driver_nand247 en in_247 wl_bar_247 vdd gnd pnand2_0
Xwl_driver_inv247 wl_bar_247 wl_247 vdd gnd pdriver_0
Xwl_driver_nand248 en in_248 wl_bar_248 vdd gnd pnand2_0
Xwl_driver_inv248 wl_bar_248 wl_248 vdd gnd pdriver_0
Xwl_driver_nand249 en in_249 wl_bar_249 vdd gnd pnand2_0
Xwl_driver_inv249 wl_bar_249 wl_249 vdd gnd pdriver_0
Xwl_driver_nand250 en in_250 wl_bar_250 vdd gnd pnand2_0
Xwl_driver_inv250 wl_bar_250 wl_250 vdd gnd pdriver_0
Xwl_driver_nand251 en in_251 wl_bar_251 vdd gnd pnand2_0
Xwl_driver_inv251 wl_bar_251 wl_251 vdd gnd pdriver_0
Xwl_driver_nand252 en in_252 wl_bar_252 vdd gnd pnand2_0
Xwl_driver_inv252 wl_bar_252 wl_252 vdd gnd pdriver_0
Xwl_driver_nand253 en in_253 wl_bar_253 vdd gnd pnand2_0
Xwl_driver_inv253 wl_bar_253 wl_253 vdd gnd pdriver_0
Xwl_driver_nand254 en in_254 wl_bar_254 vdd gnd pnand2_0
Xwl_driver_inv254 wl_bar_254 wl_254 vdd gnd pdriver_0
Xwl_driver_nand255 en in_255 wl_bar_255 vdd gnd pnand2_0
Xwl_driver_inv255 wl_bar_255 wl_255 vdd gnd pdriver_0
.ENDS wordline_driver_0

.SUBCKT port_address_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : addr_7 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* OUTPUT: wl_128 
* OUTPUT: wl_129 
* OUTPUT: wl_130 
* OUTPUT: wl_131 
* OUTPUT: wl_132 
* OUTPUT: wl_133 
* OUTPUT: wl_134 
* OUTPUT: wl_135 
* OUTPUT: wl_136 
* OUTPUT: wl_137 
* OUTPUT: wl_138 
* OUTPUT: wl_139 
* OUTPUT: wl_140 
* OUTPUT: wl_141 
* OUTPUT: wl_142 
* OUTPUT: wl_143 
* OUTPUT: wl_144 
* OUTPUT: wl_145 
* OUTPUT: wl_146 
* OUTPUT: wl_147 
* OUTPUT: wl_148 
* OUTPUT: wl_149 
* OUTPUT: wl_150 
* OUTPUT: wl_151 
* OUTPUT: wl_152 
* OUTPUT: wl_153 
* OUTPUT: wl_154 
* OUTPUT: wl_155 
* OUTPUT: wl_156 
* OUTPUT: wl_157 
* OUTPUT: wl_158 
* OUTPUT: wl_159 
* OUTPUT: wl_160 
* OUTPUT: wl_161 
* OUTPUT: wl_162 
* OUTPUT: wl_163 
* OUTPUT: wl_164 
* OUTPUT: wl_165 
* OUTPUT: wl_166 
* OUTPUT: wl_167 
* OUTPUT: wl_168 
* OUTPUT: wl_169 
* OUTPUT: wl_170 
* OUTPUT: wl_171 
* OUTPUT: wl_172 
* OUTPUT: wl_173 
* OUTPUT: wl_174 
* OUTPUT: wl_175 
* OUTPUT: wl_176 
* OUTPUT: wl_177 
* OUTPUT: wl_178 
* OUTPUT: wl_179 
* OUTPUT: wl_180 
* OUTPUT: wl_181 
* OUTPUT: wl_182 
* OUTPUT: wl_183 
* OUTPUT: wl_184 
* OUTPUT: wl_185 
* OUTPUT: wl_186 
* OUTPUT: wl_187 
* OUTPUT: wl_188 
* OUTPUT: wl_189 
* OUTPUT: wl_190 
* OUTPUT: wl_191 
* OUTPUT: wl_192 
* OUTPUT: wl_193 
* OUTPUT: wl_194 
* OUTPUT: wl_195 
* OUTPUT: wl_196 
* OUTPUT: wl_197 
* OUTPUT: wl_198 
* OUTPUT: wl_199 
* OUTPUT: wl_200 
* OUTPUT: wl_201 
* OUTPUT: wl_202 
* OUTPUT: wl_203 
* OUTPUT: wl_204 
* OUTPUT: wl_205 
* OUTPUT: wl_206 
* OUTPUT: wl_207 
* OUTPUT: wl_208 
* OUTPUT: wl_209 
* OUTPUT: wl_210 
* OUTPUT: wl_211 
* OUTPUT: wl_212 
* OUTPUT: wl_213 
* OUTPUT: wl_214 
* OUTPUT: wl_215 
* OUTPUT: wl_216 
* OUTPUT: wl_217 
* OUTPUT: wl_218 
* OUTPUT: wl_219 
* OUTPUT: wl_220 
* OUTPUT: wl_221 
* OUTPUT: wl_222 
* OUTPUT: wl_223 
* OUTPUT: wl_224 
* OUTPUT: wl_225 
* OUTPUT: wl_226 
* OUTPUT: wl_227 
* OUTPUT: wl_228 
* OUTPUT: wl_229 
* OUTPUT: wl_230 
* OUTPUT: wl_231 
* OUTPUT: wl_232 
* OUTPUT: wl_233 
* OUTPUT: wl_234 
* OUTPUT: wl_235 
* OUTPUT: wl_236 
* OUTPUT: wl_237 
* OUTPUT: wl_238 
* OUTPUT: wl_239 
* OUTPUT: wl_240 
* OUTPUT: wl_241 
* OUTPUT: wl_242 
* OUTPUT: wl_243 
* OUTPUT: wl_244 
* OUTPUT: wl_245 
* OUTPUT: wl_246 
* OUTPUT: wl_247 
* OUTPUT: wl_248 
* OUTPUT: wl_249 
* OUTPUT: wl_250 
* OUTPUT: wl_251 
* OUTPUT: wl_252 
* OUTPUT: wl_253 
* OUTPUT: wl_254 
* OUTPUT: wl_255 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 dec_out_128 dec_out_129 dec_out_130 dec_out_131 dec_out_132 dec_out_133 dec_out_134 dec_out_135 dec_out_136 dec_out_137 dec_out_138 dec_out_139 dec_out_140 dec_out_141 dec_out_142 dec_out_143 dec_out_144 dec_out_145 dec_out_146 dec_out_147 dec_out_148 dec_out_149 dec_out_150 dec_out_151 dec_out_152 dec_out_153 dec_out_154 dec_out_155 dec_out_156 dec_out_157 dec_out_158 dec_out_159 dec_out_160 dec_out_161 dec_out_162 dec_out_163 dec_out_164 dec_out_165 dec_out_166 dec_out_167 dec_out_168 dec_out_169 dec_out_170 dec_out_171 dec_out_172 dec_out_173 dec_out_174 dec_out_175 dec_out_176 dec_out_177 dec_out_178 dec_out_179 dec_out_180 dec_out_181 dec_out_182 dec_out_183 dec_out_184 dec_out_185 dec_out_186 dec_out_187 dec_out_188 dec_out_189 dec_out_190 dec_out_191 dec_out_192 dec_out_193 dec_out_194 dec_out_195 dec_out_196 dec_out_197 dec_out_198 dec_out_199 dec_out_200 dec_out_201 dec_out_202 dec_out_203 dec_out_204 dec_out_205 dec_out_206 dec_out_207 dec_out_208 dec_out_209 dec_out_210 dec_out_211 dec_out_212 dec_out_213 dec_out_214 dec_out_215 dec_out_216 dec_out_217 dec_out_218 dec_out_219 dec_out_220 dec_out_221 dec_out_222 dec_out_223 dec_out_224 dec_out_225 dec_out_226 dec_out_227 dec_out_228 dec_out_229 dec_out_230 dec_out_231 dec_out_232 dec_out_233 dec_out_234 dec_out_235 dec_out_236 dec_out_237 dec_out_238 dec_out_239 dec_out_240 dec_out_241 dec_out_242 dec_out_243 dec_out_244 dec_out_245 dec_out_246 dec_out_247 dec_out_248 dec_out_249 dec_out_250 dec_out_251 dec_out_252 dec_out_253 dec_out_254 dec_out_255 vdd gnd hierarchical_decoder_0
Xwordline_driver dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 dec_out_128 dec_out_129 dec_out_130 dec_out_131 dec_out_132 dec_out_133 dec_out_134 dec_out_135 dec_out_136 dec_out_137 dec_out_138 dec_out_139 dec_out_140 dec_out_141 dec_out_142 dec_out_143 dec_out_144 dec_out_145 dec_out_146 dec_out_147 dec_out_148 dec_out_149 dec_out_150 dec_out_151 dec_out_152 dec_out_153 dec_out_154 dec_out_155 dec_out_156 dec_out_157 dec_out_158 dec_out_159 dec_out_160 dec_out_161 dec_out_162 dec_out_163 dec_out_164 dec_out_165 dec_out_166 dec_out_167 dec_out_168 dec_out_169 dec_out_170 dec_out_171 dec_out_172 dec_out_173 dec_out_174 dec_out_175 dec_out_176 dec_out_177 dec_out_178 dec_out_179 dec_out_180 dec_out_181 dec_out_182 dec_out_183 dec_out_184 dec_out_185 dec_out_186 dec_out_187 dec_out_188 dec_out_189 dec_out_190 dec_out_191 dec_out_192 dec_out_193 dec_out_194 dec_out_195 dec_out_196 dec_out_197 dec_out_198 dec_out_199 dec_out_200 dec_out_201 dec_out_202 dec_out_203 dec_out_204 dec_out_205 dec_out_206 dec_out_207 dec_out_208 dec_out_209 dec_out_210 dec_out_211 dec_out_212 dec_out_213 dec_out_214 dec_out_215 dec_out_216 dec_out_217 dec_out_218 dec_out_219 dec_out_220 dec_out_221 dec_out_222 dec_out_223 dec_out_224 dec_out_225 dec_out_226 dec_out_227 dec_out_228 dec_out_229 dec_out_230 dec_out_231 dec_out_232 dec_out_233 dec_out_234 dec_out_235 dec_out_236 dec_out_237 dec_out_238 dec_out_239 dec_out_240 dec_out_241 dec_out_242 dec_out_243 dec_out_244 dec_out_245 dec_out_246 dec_out_247 dec_out_248 dec_out_249 dec_out_250 dec_out_251 dec_out_252 dec_out_253 dec_out_254 dec_out_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 wl_en vdd gnd wordline_driver_0
.ENDS port_address_0

.SUBCKT cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* INPUT : wl_131 
* INPUT : wl_132 
* INPUT : wl_133 
* INPUT : wl_134 
* INPUT : wl_135 
* INPUT : wl_136 
* INPUT : wl_137 
* INPUT : wl_138 
* INPUT : wl_139 
* INPUT : wl_140 
* INPUT : wl_141 
* INPUT : wl_142 
* INPUT : wl_143 
* INPUT : wl_144 
* INPUT : wl_145 
* INPUT : wl_146 
* INPUT : wl_147 
* INPUT : wl_148 
* INPUT : wl_149 
* INPUT : wl_150 
* INPUT : wl_151 
* INPUT : wl_152 
* INPUT : wl_153 
* INPUT : wl_154 
* INPUT : wl_155 
* INPUT : wl_156 
* INPUT : wl_157 
* INPUT : wl_158 
* INPUT : wl_159 
* INPUT : wl_160 
* INPUT : wl_161 
* INPUT : wl_162 
* INPUT : wl_163 
* INPUT : wl_164 
* INPUT : wl_165 
* INPUT : wl_166 
* INPUT : wl_167 
* INPUT : wl_168 
* INPUT : wl_169 
* INPUT : wl_170 
* INPUT : wl_171 
* INPUT : wl_172 
* INPUT : wl_173 
* INPUT : wl_174 
* INPUT : wl_175 
* INPUT : wl_176 
* INPUT : wl_177 
* INPUT : wl_178 
* INPUT : wl_179 
* INPUT : wl_180 
* INPUT : wl_181 
* INPUT : wl_182 
* INPUT : wl_183 
* INPUT : wl_184 
* INPUT : wl_185 
* INPUT : wl_186 
* INPUT : wl_187 
* INPUT : wl_188 
* INPUT : wl_189 
* INPUT : wl_190 
* INPUT : wl_191 
* INPUT : wl_192 
* INPUT : wl_193 
* INPUT : wl_194 
* INPUT : wl_195 
* INPUT : wl_196 
* INPUT : wl_197 
* INPUT : wl_198 
* INPUT : wl_199 
* INPUT : wl_200 
* INPUT : wl_201 
* INPUT : wl_202 
* INPUT : wl_203 
* INPUT : wl_204 
* INPUT : wl_205 
* INPUT : wl_206 
* INPUT : wl_207 
* INPUT : wl_208 
* INPUT : wl_209 
* INPUT : wl_210 
* INPUT : wl_211 
* INPUT : wl_212 
* INPUT : wl_213 
* INPUT : wl_214 
* INPUT : wl_215 
* INPUT : wl_216 
* INPUT : wl_217 
* INPUT : wl_218 
* INPUT : wl_219 
* INPUT : wl_220 
* INPUT : wl_221 
* INPUT : wl_222 
* INPUT : wl_223 
* INPUT : wl_224 
* INPUT : wl_225 
* INPUT : wl_226 
* INPUT : wl_227 
* INPUT : wl_228 
* INPUT : wl_229 
* INPUT : wl_230 
* INPUT : wl_231 
* INPUT : wl_232 
* INPUT : wl_233 
* INPUT : wl_234 
* INPUT : wl_235 
* INPUT : wl_236 
* INPUT : wl_237 
* INPUT : wl_238 
* INPUT : wl_239 
* INPUT : wl_240 
* INPUT : wl_241 
* INPUT : wl_242 
* INPUT : wl_243 
* INPUT : wl_244 
* INPUT : wl_245 
* INPUT : wl_246 
* INPUT : wl_247 
* INPUT : wl_248 
* INPUT : wl_249 
* INPUT : wl_250 
* INPUT : wl_251 
* INPUT : wl_252 
* INPUT : wl_253 
* INPUT : wl_254 
* INPUT : wl_255 
* POWER : vdd 
* GROUND: gnd 
* rows: 256 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd cell_6t
Xbit_r128_c0 bl_0 br_0 wl_128 vdd gnd cell_6t
Xbit_r129_c0 bl_0 br_0 wl_129 vdd gnd cell_6t
Xbit_r130_c0 bl_0 br_0 wl_130 vdd gnd cell_6t
Xbit_r131_c0 bl_0 br_0 wl_131 vdd gnd cell_6t
Xbit_r132_c0 bl_0 br_0 wl_132 vdd gnd cell_6t
Xbit_r133_c0 bl_0 br_0 wl_133 vdd gnd cell_6t
Xbit_r134_c0 bl_0 br_0 wl_134 vdd gnd cell_6t
Xbit_r135_c0 bl_0 br_0 wl_135 vdd gnd cell_6t
Xbit_r136_c0 bl_0 br_0 wl_136 vdd gnd cell_6t
Xbit_r137_c0 bl_0 br_0 wl_137 vdd gnd cell_6t
Xbit_r138_c0 bl_0 br_0 wl_138 vdd gnd cell_6t
Xbit_r139_c0 bl_0 br_0 wl_139 vdd gnd cell_6t
Xbit_r140_c0 bl_0 br_0 wl_140 vdd gnd cell_6t
Xbit_r141_c0 bl_0 br_0 wl_141 vdd gnd cell_6t
Xbit_r142_c0 bl_0 br_0 wl_142 vdd gnd cell_6t
Xbit_r143_c0 bl_0 br_0 wl_143 vdd gnd cell_6t
Xbit_r144_c0 bl_0 br_0 wl_144 vdd gnd cell_6t
Xbit_r145_c0 bl_0 br_0 wl_145 vdd gnd cell_6t
Xbit_r146_c0 bl_0 br_0 wl_146 vdd gnd cell_6t
Xbit_r147_c0 bl_0 br_0 wl_147 vdd gnd cell_6t
Xbit_r148_c0 bl_0 br_0 wl_148 vdd gnd cell_6t
Xbit_r149_c0 bl_0 br_0 wl_149 vdd gnd cell_6t
Xbit_r150_c0 bl_0 br_0 wl_150 vdd gnd cell_6t
Xbit_r151_c0 bl_0 br_0 wl_151 vdd gnd cell_6t
Xbit_r152_c0 bl_0 br_0 wl_152 vdd gnd cell_6t
Xbit_r153_c0 bl_0 br_0 wl_153 vdd gnd cell_6t
Xbit_r154_c0 bl_0 br_0 wl_154 vdd gnd cell_6t
Xbit_r155_c0 bl_0 br_0 wl_155 vdd gnd cell_6t
Xbit_r156_c0 bl_0 br_0 wl_156 vdd gnd cell_6t
Xbit_r157_c0 bl_0 br_0 wl_157 vdd gnd cell_6t
Xbit_r158_c0 bl_0 br_0 wl_158 vdd gnd cell_6t
Xbit_r159_c0 bl_0 br_0 wl_159 vdd gnd cell_6t
Xbit_r160_c0 bl_0 br_0 wl_160 vdd gnd cell_6t
Xbit_r161_c0 bl_0 br_0 wl_161 vdd gnd cell_6t
Xbit_r162_c0 bl_0 br_0 wl_162 vdd gnd cell_6t
Xbit_r163_c0 bl_0 br_0 wl_163 vdd gnd cell_6t
Xbit_r164_c0 bl_0 br_0 wl_164 vdd gnd cell_6t
Xbit_r165_c0 bl_0 br_0 wl_165 vdd gnd cell_6t
Xbit_r166_c0 bl_0 br_0 wl_166 vdd gnd cell_6t
Xbit_r167_c0 bl_0 br_0 wl_167 vdd gnd cell_6t
Xbit_r168_c0 bl_0 br_0 wl_168 vdd gnd cell_6t
Xbit_r169_c0 bl_0 br_0 wl_169 vdd gnd cell_6t
Xbit_r170_c0 bl_0 br_0 wl_170 vdd gnd cell_6t
Xbit_r171_c0 bl_0 br_0 wl_171 vdd gnd cell_6t
Xbit_r172_c0 bl_0 br_0 wl_172 vdd gnd cell_6t
Xbit_r173_c0 bl_0 br_0 wl_173 vdd gnd cell_6t
Xbit_r174_c0 bl_0 br_0 wl_174 vdd gnd cell_6t
Xbit_r175_c0 bl_0 br_0 wl_175 vdd gnd cell_6t
Xbit_r176_c0 bl_0 br_0 wl_176 vdd gnd cell_6t
Xbit_r177_c0 bl_0 br_0 wl_177 vdd gnd cell_6t
Xbit_r178_c0 bl_0 br_0 wl_178 vdd gnd cell_6t
Xbit_r179_c0 bl_0 br_0 wl_179 vdd gnd cell_6t
Xbit_r180_c0 bl_0 br_0 wl_180 vdd gnd cell_6t
Xbit_r181_c0 bl_0 br_0 wl_181 vdd gnd cell_6t
Xbit_r182_c0 bl_0 br_0 wl_182 vdd gnd cell_6t
Xbit_r183_c0 bl_0 br_0 wl_183 vdd gnd cell_6t
Xbit_r184_c0 bl_0 br_0 wl_184 vdd gnd cell_6t
Xbit_r185_c0 bl_0 br_0 wl_185 vdd gnd cell_6t
Xbit_r186_c0 bl_0 br_0 wl_186 vdd gnd cell_6t
Xbit_r187_c0 bl_0 br_0 wl_187 vdd gnd cell_6t
Xbit_r188_c0 bl_0 br_0 wl_188 vdd gnd cell_6t
Xbit_r189_c0 bl_0 br_0 wl_189 vdd gnd cell_6t
Xbit_r190_c0 bl_0 br_0 wl_190 vdd gnd cell_6t
Xbit_r191_c0 bl_0 br_0 wl_191 vdd gnd cell_6t
Xbit_r192_c0 bl_0 br_0 wl_192 vdd gnd cell_6t
Xbit_r193_c0 bl_0 br_0 wl_193 vdd gnd cell_6t
Xbit_r194_c0 bl_0 br_0 wl_194 vdd gnd cell_6t
Xbit_r195_c0 bl_0 br_0 wl_195 vdd gnd cell_6t
Xbit_r196_c0 bl_0 br_0 wl_196 vdd gnd cell_6t
Xbit_r197_c0 bl_0 br_0 wl_197 vdd gnd cell_6t
Xbit_r198_c0 bl_0 br_0 wl_198 vdd gnd cell_6t
Xbit_r199_c0 bl_0 br_0 wl_199 vdd gnd cell_6t
Xbit_r200_c0 bl_0 br_0 wl_200 vdd gnd cell_6t
Xbit_r201_c0 bl_0 br_0 wl_201 vdd gnd cell_6t
Xbit_r202_c0 bl_0 br_0 wl_202 vdd gnd cell_6t
Xbit_r203_c0 bl_0 br_0 wl_203 vdd gnd cell_6t
Xbit_r204_c0 bl_0 br_0 wl_204 vdd gnd cell_6t
Xbit_r205_c0 bl_0 br_0 wl_205 vdd gnd cell_6t
Xbit_r206_c0 bl_0 br_0 wl_206 vdd gnd cell_6t
Xbit_r207_c0 bl_0 br_0 wl_207 vdd gnd cell_6t
Xbit_r208_c0 bl_0 br_0 wl_208 vdd gnd cell_6t
Xbit_r209_c0 bl_0 br_0 wl_209 vdd gnd cell_6t
Xbit_r210_c0 bl_0 br_0 wl_210 vdd gnd cell_6t
Xbit_r211_c0 bl_0 br_0 wl_211 vdd gnd cell_6t
Xbit_r212_c0 bl_0 br_0 wl_212 vdd gnd cell_6t
Xbit_r213_c0 bl_0 br_0 wl_213 vdd gnd cell_6t
Xbit_r214_c0 bl_0 br_0 wl_214 vdd gnd cell_6t
Xbit_r215_c0 bl_0 br_0 wl_215 vdd gnd cell_6t
Xbit_r216_c0 bl_0 br_0 wl_216 vdd gnd cell_6t
Xbit_r217_c0 bl_0 br_0 wl_217 vdd gnd cell_6t
Xbit_r218_c0 bl_0 br_0 wl_218 vdd gnd cell_6t
Xbit_r219_c0 bl_0 br_0 wl_219 vdd gnd cell_6t
Xbit_r220_c0 bl_0 br_0 wl_220 vdd gnd cell_6t
Xbit_r221_c0 bl_0 br_0 wl_221 vdd gnd cell_6t
Xbit_r222_c0 bl_0 br_0 wl_222 vdd gnd cell_6t
Xbit_r223_c0 bl_0 br_0 wl_223 vdd gnd cell_6t
Xbit_r224_c0 bl_0 br_0 wl_224 vdd gnd cell_6t
Xbit_r225_c0 bl_0 br_0 wl_225 vdd gnd cell_6t
Xbit_r226_c0 bl_0 br_0 wl_226 vdd gnd cell_6t
Xbit_r227_c0 bl_0 br_0 wl_227 vdd gnd cell_6t
Xbit_r228_c0 bl_0 br_0 wl_228 vdd gnd cell_6t
Xbit_r229_c0 bl_0 br_0 wl_229 vdd gnd cell_6t
Xbit_r230_c0 bl_0 br_0 wl_230 vdd gnd cell_6t
Xbit_r231_c0 bl_0 br_0 wl_231 vdd gnd cell_6t
Xbit_r232_c0 bl_0 br_0 wl_232 vdd gnd cell_6t
Xbit_r233_c0 bl_0 br_0 wl_233 vdd gnd cell_6t
Xbit_r234_c0 bl_0 br_0 wl_234 vdd gnd cell_6t
Xbit_r235_c0 bl_0 br_0 wl_235 vdd gnd cell_6t
Xbit_r236_c0 bl_0 br_0 wl_236 vdd gnd cell_6t
Xbit_r237_c0 bl_0 br_0 wl_237 vdd gnd cell_6t
Xbit_r238_c0 bl_0 br_0 wl_238 vdd gnd cell_6t
Xbit_r239_c0 bl_0 br_0 wl_239 vdd gnd cell_6t
Xbit_r240_c0 bl_0 br_0 wl_240 vdd gnd cell_6t
Xbit_r241_c0 bl_0 br_0 wl_241 vdd gnd cell_6t
Xbit_r242_c0 bl_0 br_0 wl_242 vdd gnd cell_6t
Xbit_r243_c0 bl_0 br_0 wl_243 vdd gnd cell_6t
Xbit_r244_c0 bl_0 br_0 wl_244 vdd gnd cell_6t
Xbit_r245_c0 bl_0 br_0 wl_245 vdd gnd cell_6t
Xbit_r246_c0 bl_0 br_0 wl_246 vdd gnd cell_6t
Xbit_r247_c0 bl_0 br_0 wl_247 vdd gnd cell_6t
Xbit_r248_c0 bl_0 br_0 wl_248 vdd gnd cell_6t
Xbit_r249_c0 bl_0 br_0 wl_249 vdd gnd cell_6t
Xbit_r250_c0 bl_0 br_0 wl_250 vdd gnd cell_6t
Xbit_r251_c0 bl_0 br_0 wl_251 vdd gnd cell_6t
Xbit_r252_c0 bl_0 br_0 wl_252 vdd gnd cell_6t
Xbit_r253_c0 bl_0 br_0 wl_253 vdd gnd cell_6t
Xbit_r254_c0 bl_0 br_0 wl_254 vdd gnd cell_6t
Xbit_r255_c0 bl_0 br_0 wl_255 vdd gnd cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd cell_6t
Xbit_r1_c1 bl_1 br_1 wl_1 vdd gnd cell_6t
Xbit_r2_c1 bl_1 br_1 wl_2 vdd gnd cell_6t
Xbit_r3_c1 bl_1 br_1 wl_3 vdd gnd cell_6t
Xbit_r4_c1 bl_1 br_1 wl_4 vdd gnd cell_6t
Xbit_r5_c1 bl_1 br_1 wl_5 vdd gnd cell_6t
Xbit_r6_c1 bl_1 br_1 wl_6 vdd gnd cell_6t
Xbit_r7_c1 bl_1 br_1 wl_7 vdd gnd cell_6t
Xbit_r8_c1 bl_1 br_1 wl_8 vdd gnd cell_6t
Xbit_r9_c1 bl_1 br_1 wl_9 vdd gnd cell_6t
Xbit_r10_c1 bl_1 br_1 wl_10 vdd gnd cell_6t
Xbit_r11_c1 bl_1 br_1 wl_11 vdd gnd cell_6t
Xbit_r12_c1 bl_1 br_1 wl_12 vdd gnd cell_6t
Xbit_r13_c1 bl_1 br_1 wl_13 vdd gnd cell_6t
Xbit_r14_c1 bl_1 br_1 wl_14 vdd gnd cell_6t
Xbit_r15_c1 bl_1 br_1 wl_15 vdd gnd cell_6t
Xbit_r16_c1 bl_1 br_1 wl_16 vdd gnd cell_6t
Xbit_r17_c1 bl_1 br_1 wl_17 vdd gnd cell_6t
Xbit_r18_c1 bl_1 br_1 wl_18 vdd gnd cell_6t
Xbit_r19_c1 bl_1 br_1 wl_19 vdd gnd cell_6t
Xbit_r20_c1 bl_1 br_1 wl_20 vdd gnd cell_6t
Xbit_r21_c1 bl_1 br_1 wl_21 vdd gnd cell_6t
Xbit_r22_c1 bl_1 br_1 wl_22 vdd gnd cell_6t
Xbit_r23_c1 bl_1 br_1 wl_23 vdd gnd cell_6t
Xbit_r24_c1 bl_1 br_1 wl_24 vdd gnd cell_6t
Xbit_r25_c1 bl_1 br_1 wl_25 vdd gnd cell_6t
Xbit_r26_c1 bl_1 br_1 wl_26 vdd gnd cell_6t
Xbit_r27_c1 bl_1 br_1 wl_27 vdd gnd cell_6t
Xbit_r28_c1 bl_1 br_1 wl_28 vdd gnd cell_6t
Xbit_r29_c1 bl_1 br_1 wl_29 vdd gnd cell_6t
Xbit_r30_c1 bl_1 br_1 wl_30 vdd gnd cell_6t
Xbit_r31_c1 bl_1 br_1 wl_31 vdd gnd cell_6t
Xbit_r32_c1 bl_1 br_1 wl_32 vdd gnd cell_6t
Xbit_r33_c1 bl_1 br_1 wl_33 vdd gnd cell_6t
Xbit_r34_c1 bl_1 br_1 wl_34 vdd gnd cell_6t
Xbit_r35_c1 bl_1 br_1 wl_35 vdd gnd cell_6t
Xbit_r36_c1 bl_1 br_1 wl_36 vdd gnd cell_6t
Xbit_r37_c1 bl_1 br_1 wl_37 vdd gnd cell_6t
Xbit_r38_c1 bl_1 br_1 wl_38 vdd gnd cell_6t
Xbit_r39_c1 bl_1 br_1 wl_39 vdd gnd cell_6t
Xbit_r40_c1 bl_1 br_1 wl_40 vdd gnd cell_6t
Xbit_r41_c1 bl_1 br_1 wl_41 vdd gnd cell_6t
Xbit_r42_c1 bl_1 br_1 wl_42 vdd gnd cell_6t
Xbit_r43_c1 bl_1 br_1 wl_43 vdd gnd cell_6t
Xbit_r44_c1 bl_1 br_1 wl_44 vdd gnd cell_6t
Xbit_r45_c1 bl_1 br_1 wl_45 vdd gnd cell_6t
Xbit_r46_c1 bl_1 br_1 wl_46 vdd gnd cell_6t
Xbit_r47_c1 bl_1 br_1 wl_47 vdd gnd cell_6t
Xbit_r48_c1 bl_1 br_1 wl_48 vdd gnd cell_6t
Xbit_r49_c1 bl_1 br_1 wl_49 vdd gnd cell_6t
Xbit_r50_c1 bl_1 br_1 wl_50 vdd gnd cell_6t
Xbit_r51_c1 bl_1 br_1 wl_51 vdd gnd cell_6t
Xbit_r52_c1 bl_1 br_1 wl_52 vdd gnd cell_6t
Xbit_r53_c1 bl_1 br_1 wl_53 vdd gnd cell_6t
Xbit_r54_c1 bl_1 br_1 wl_54 vdd gnd cell_6t
Xbit_r55_c1 bl_1 br_1 wl_55 vdd gnd cell_6t
Xbit_r56_c1 bl_1 br_1 wl_56 vdd gnd cell_6t
Xbit_r57_c1 bl_1 br_1 wl_57 vdd gnd cell_6t
Xbit_r58_c1 bl_1 br_1 wl_58 vdd gnd cell_6t
Xbit_r59_c1 bl_1 br_1 wl_59 vdd gnd cell_6t
Xbit_r60_c1 bl_1 br_1 wl_60 vdd gnd cell_6t
Xbit_r61_c1 bl_1 br_1 wl_61 vdd gnd cell_6t
Xbit_r62_c1 bl_1 br_1 wl_62 vdd gnd cell_6t
Xbit_r63_c1 bl_1 br_1 wl_63 vdd gnd cell_6t
Xbit_r64_c1 bl_1 br_1 wl_64 vdd gnd cell_6t
Xbit_r65_c1 bl_1 br_1 wl_65 vdd gnd cell_6t
Xbit_r66_c1 bl_1 br_1 wl_66 vdd gnd cell_6t
Xbit_r67_c1 bl_1 br_1 wl_67 vdd gnd cell_6t
Xbit_r68_c1 bl_1 br_1 wl_68 vdd gnd cell_6t
Xbit_r69_c1 bl_1 br_1 wl_69 vdd gnd cell_6t
Xbit_r70_c1 bl_1 br_1 wl_70 vdd gnd cell_6t
Xbit_r71_c1 bl_1 br_1 wl_71 vdd gnd cell_6t
Xbit_r72_c1 bl_1 br_1 wl_72 vdd gnd cell_6t
Xbit_r73_c1 bl_1 br_1 wl_73 vdd gnd cell_6t
Xbit_r74_c1 bl_1 br_1 wl_74 vdd gnd cell_6t
Xbit_r75_c1 bl_1 br_1 wl_75 vdd gnd cell_6t
Xbit_r76_c1 bl_1 br_1 wl_76 vdd gnd cell_6t
Xbit_r77_c1 bl_1 br_1 wl_77 vdd gnd cell_6t
Xbit_r78_c1 bl_1 br_1 wl_78 vdd gnd cell_6t
Xbit_r79_c1 bl_1 br_1 wl_79 vdd gnd cell_6t
Xbit_r80_c1 bl_1 br_1 wl_80 vdd gnd cell_6t
Xbit_r81_c1 bl_1 br_1 wl_81 vdd gnd cell_6t
Xbit_r82_c1 bl_1 br_1 wl_82 vdd gnd cell_6t
Xbit_r83_c1 bl_1 br_1 wl_83 vdd gnd cell_6t
Xbit_r84_c1 bl_1 br_1 wl_84 vdd gnd cell_6t
Xbit_r85_c1 bl_1 br_1 wl_85 vdd gnd cell_6t
Xbit_r86_c1 bl_1 br_1 wl_86 vdd gnd cell_6t
Xbit_r87_c1 bl_1 br_1 wl_87 vdd gnd cell_6t
Xbit_r88_c1 bl_1 br_1 wl_88 vdd gnd cell_6t
Xbit_r89_c1 bl_1 br_1 wl_89 vdd gnd cell_6t
Xbit_r90_c1 bl_1 br_1 wl_90 vdd gnd cell_6t
Xbit_r91_c1 bl_1 br_1 wl_91 vdd gnd cell_6t
Xbit_r92_c1 bl_1 br_1 wl_92 vdd gnd cell_6t
Xbit_r93_c1 bl_1 br_1 wl_93 vdd gnd cell_6t
Xbit_r94_c1 bl_1 br_1 wl_94 vdd gnd cell_6t
Xbit_r95_c1 bl_1 br_1 wl_95 vdd gnd cell_6t
Xbit_r96_c1 bl_1 br_1 wl_96 vdd gnd cell_6t
Xbit_r97_c1 bl_1 br_1 wl_97 vdd gnd cell_6t
Xbit_r98_c1 bl_1 br_1 wl_98 vdd gnd cell_6t
Xbit_r99_c1 bl_1 br_1 wl_99 vdd gnd cell_6t
Xbit_r100_c1 bl_1 br_1 wl_100 vdd gnd cell_6t
Xbit_r101_c1 bl_1 br_1 wl_101 vdd gnd cell_6t
Xbit_r102_c1 bl_1 br_1 wl_102 vdd gnd cell_6t
Xbit_r103_c1 bl_1 br_1 wl_103 vdd gnd cell_6t
Xbit_r104_c1 bl_1 br_1 wl_104 vdd gnd cell_6t
Xbit_r105_c1 bl_1 br_1 wl_105 vdd gnd cell_6t
Xbit_r106_c1 bl_1 br_1 wl_106 vdd gnd cell_6t
Xbit_r107_c1 bl_1 br_1 wl_107 vdd gnd cell_6t
Xbit_r108_c1 bl_1 br_1 wl_108 vdd gnd cell_6t
Xbit_r109_c1 bl_1 br_1 wl_109 vdd gnd cell_6t
Xbit_r110_c1 bl_1 br_1 wl_110 vdd gnd cell_6t
Xbit_r111_c1 bl_1 br_1 wl_111 vdd gnd cell_6t
Xbit_r112_c1 bl_1 br_1 wl_112 vdd gnd cell_6t
Xbit_r113_c1 bl_1 br_1 wl_113 vdd gnd cell_6t
Xbit_r114_c1 bl_1 br_1 wl_114 vdd gnd cell_6t
Xbit_r115_c1 bl_1 br_1 wl_115 vdd gnd cell_6t
Xbit_r116_c1 bl_1 br_1 wl_116 vdd gnd cell_6t
Xbit_r117_c1 bl_1 br_1 wl_117 vdd gnd cell_6t
Xbit_r118_c1 bl_1 br_1 wl_118 vdd gnd cell_6t
Xbit_r119_c1 bl_1 br_1 wl_119 vdd gnd cell_6t
Xbit_r120_c1 bl_1 br_1 wl_120 vdd gnd cell_6t
Xbit_r121_c1 bl_1 br_1 wl_121 vdd gnd cell_6t
Xbit_r122_c1 bl_1 br_1 wl_122 vdd gnd cell_6t
Xbit_r123_c1 bl_1 br_1 wl_123 vdd gnd cell_6t
Xbit_r124_c1 bl_1 br_1 wl_124 vdd gnd cell_6t
Xbit_r125_c1 bl_1 br_1 wl_125 vdd gnd cell_6t
Xbit_r126_c1 bl_1 br_1 wl_126 vdd gnd cell_6t
Xbit_r127_c1 bl_1 br_1 wl_127 vdd gnd cell_6t
Xbit_r128_c1 bl_1 br_1 wl_128 vdd gnd cell_6t
Xbit_r129_c1 bl_1 br_1 wl_129 vdd gnd cell_6t
Xbit_r130_c1 bl_1 br_1 wl_130 vdd gnd cell_6t
Xbit_r131_c1 bl_1 br_1 wl_131 vdd gnd cell_6t
Xbit_r132_c1 bl_1 br_1 wl_132 vdd gnd cell_6t
Xbit_r133_c1 bl_1 br_1 wl_133 vdd gnd cell_6t
Xbit_r134_c1 bl_1 br_1 wl_134 vdd gnd cell_6t
Xbit_r135_c1 bl_1 br_1 wl_135 vdd gnd cell_6t
Xbit_r136_c1 bl_1 br_1 wl_136 vdd gnd cell_6t
Xbit_r137_c1 bl_1 br_1 wl_137 vdd gnd cell_6t
Xbit_r138_c1 bl_1 br_1 wl_138 vdd gnd cell_6t
Xbit_r139_c1 bl_1 br_1 wl_139 vdd gnd cell_6t
Xbit_r140_c1 bl_1 br_1 wl_140 vdd gnd cell_6t
Xbit_r141_c1 bl_1 br_1 wl_141 vdd gnd cell_6t
Xbit_r142_c1 bl_1 br_1 wl_142 vdd gnd cell_6t
Xbit_r143_c1 bl_1 br_1 wl_143 vdd gnd cell_6t
Xbit_r144_c1 bl_1 br_1 wl_144 vdd gnd cell_6t
Xbit_r145_c1 bl_1 br_1 wl_145 vdd gnd cell_6t
Xbit_r146_c1 bl_1 br_1 wl_146 vdd gnd cell_6t
Xbit_r147_c1 bl_1 br_1 wl_147 vdd gnd cell_6t
Xbit_r148_c1 bl_1 br_1 wl_148 vdd gnd cell_6t
Xbit_r149_c1 bl_1 br_1 wl_149 vdd gnd cell_6t
Xbit_r150_c1 bl_1 br_1 wl_150 vdd gnd cell_6t
Xbit_r151_c1 bl_1 br_1 wl_151 vdd gnd cell_6t
Xbit_r152_c1 bl_1 br_1 wl_152 vdd gnd cell_6t
Xbit_r153_c1 bl_1 br_1 wl_153 vdd gnd cell_6t
Xbit_r154_c1 bl_1 br_1 wl_154 vdd gnd cell_6t
Xbit_r155_c1 bl_1 br_1 wl_155 vdd gnd cell_6t
Xbit_r156_c1 bl_1 br_1 wl_156 vdd gnd cell_6t
Xbit_r157_c1 bl_1 br_1 wl_157 vdd gnd cell_6t
Xbit_r158_c1 bl_1 br_1 wl_158 vdd gnd cell_6t
Xbit_r159_c1 bl_1 br_1 wl_159 vdd gnd cell_6t
Xbit_r160_c1 bl_1 br_1 wl_160 vdd gnd cell_6t
Xbit_r161_c1 bl_1 br_1 wl_161 vdd gnd cell_6t
Xbit_r162_c1 bl_1 br_1 wl_162 vdd gnd cell_6t
Xbit_r163_c1 bl_1 br_1 wl_163 vdd gnd cell_6t
Xbit_r164_c1 bl_1 br_1 wl_164 vdd gnd cell_6t
Xbit_r165_c1 bl_1 br_1 wl_165 vdd gnd cell_6t
Xbit_r166_c1 bl_1 br_1 wl_166 vdd gnd cell_6t
Xbit_r167_c1 bl_1 br_1 wl_167 vdd gnd cell_6t
Xbit_r168_c1 bl_1 br_1 wl_168 vdd gnd cell_6t
Xbit_r169_c1 bl_1 br_1 wl_169 vdd gnd cell_6t
Xbit_r170_c1 bl_1 br_1 wl_170 vdd gnd cell_6t
Xbit_r171_c1 bl_1 br_1 wl_171 vdd gnd cell_6t
Xbit_r172_c1 bl_1 br_1 wl_172 vdd gnd cell_6t
Xbit_r173_c1 bl_1 br_1 wl_173 vdd gnd cell_6t
Xbit_r174_c1 bl_1 br_1 wl_174 vdd gnd cell_6t
Xbit_r175_c1 bl_1 br_1 wl_175 vdd gnd cell_6t
Xbit_r176_c1 bl_1 br_1 wl_176 vdd gnd cell_6t
Xbit_r177_c1 bl_1 br_1 wl_177 vdd gnd cell_6t
Xbit_r178_c1 bl_1 br_1 wl_178 vdd gnd cell_6t
Xbit_r179_c1 bl_1 br_1 wl_179 vdd gnd cell_6t
Xbit_r180_c1 bl_1 br_1 wl_180 vdd gnd cell_6t
Xbit_r181_c1 bl_1 br_1 wl_181 vdd gnd cell_6t
Xbit_r182_c1 bl_1 br_1 wl_182 vdd gnd cell_6t
Xbit_r183_c1 bl_1 br_1 wl_183 vdd gnd cell_6t
Xbit_r184_c1 bl_1 br_1 wl_184 vdd gnd cell_6t
Xbit_r185_c1 bl_1 br_1 wl_185 vdd gnd cell_6t
Xbit_r186_c1 bl_1 br_1 wl_186 vdd gnd cell_6t
Xbit_r187_c1 bl_1 br_1 wl_187 vdd gnd cell_6t
Xbit_r188_c1 bl_1 br_1 wl_188 vdd gnd cell_6t
Xbit_r189_c1 bl_1 br_1 wl_189 vdd gnd cell_6t
Xbit_r190_c1 bl_1 br_1 wl_190 vdd gnd cell_6t
Xbit_r191_c1 bl_1 br_1 wl_191 vdd gnd cell_6t
Xbit_r192_c1 bl_1 br_1 wl_192 vdd gnd cell_6t
Xbit_r193_c1 bl_1 br_1 wl_193 vdd gnd cell_6t
Xbit_r194_c1 bl_1 br_1 wl_194 vdd gnd cell_6t
Xbit_r195_c1 bl_1 br_1 wl_195 vdd gnd cell_6t
Xbit_r196_c1 bl_1 br_1 wl_196 vdd gnd cell_6t
Xbit_r197_c1 bl_1 br_1 wl_197 vdd gnd cell_6t
Xbit_r198_c1 bl_1 br_1 wl_198 vdd gnd cell_6t
Xbit_r199_c1 bl_1 br_1 wl_199 vdd gnd cell_6t
Xbit_r200_c1 bl_1 br_1 wl_200 vdd gnd cell_6t
Xbit_r201_c1 bl_1 br_1 wl_201 vdd gnd cell_6t
Xbit_r202_c1 bl_1 br_1 wl_202 vdd gnd cell_6t
Xbit_r203_c1 bl_1 br_1 wl_203 vdd gnd cell_6t
Xbit_r204_c1 bl_1 br_1 wl_204 vdd gnd cell_6t
Xbit_r205_c1 bl_1 br_1 wl_205 vdd gnd cell_6t
Xbit_r206_c1 bl_1 br_1 wl_206 vdd gnd cell_6t
Xbit_r207_c1 bl_1 br_1 wl_207 vdd gnd cell_6t
Xbit_r208_c1 bl_1 br_1 wl_208 vdd gnd cell_6t
Xbit_r209_c1 bl_1 br_1 wl_209 vdd gnd cell_6t
Xbit_r210_c1 bl_1 br_1 wl_210 vdd gnd cell_6t
Xbit_r211_c1 bl_1 br_1 wl_211 vdd gnd cell_6t
Xbit_r212_c1 bl_1 br_1 wl_212 vdd gnd cell_6t
Xbit_r213_c1 bl_1 br_1 wl_213 vdd gnd cell_6t
Xbit_r214_c1 bl_1 br_1 wl_214 vdd gnd cell_6t
Xbit_r215_c1 bl_1 br_1 wl_215 vdd gnd cell_6t
Xbit_r216_c1 bl_1 br_1 wl_216 vdd gnd cell_6t
Xbit_r217_c1 bl_1 br_1 wl_217 vdd gnd cell_6t
Xbit_r218_c1 bl_1 br_1 wl_218 vdd gnd cell_6t
Xbit_r219_c1 bl_1 br_1 wl_219 vdd gnd cell_6t
Xbit_r220_c1 bl_1 br_1 wl_220 vdd gnd cell_6t
Xbit_r221_c1 bl_1 br_1 wl_221 vdd gnd cell_6t
Xbit_r222_c1 bl_1 br_1 wl_222 vdd gnd cell_6t
Xbit_r223_c1 bl_1 br_1 wl_223 vdd gnd cell_6t
Xbit_r224_c1 bl_1 br_1 wl_224 vdd gnd cell_6t
Xbit_r225_c1 bl_1 br_1 wl_225 vdd gnd cell_6t
Xbit_r226_c1 bl_1 br_1 wl_226 vdd gnd cell_6t
Xbit_r227_c1 bl_1 br_1 wl_227 vdd gnd cell_6t
Xbit_r228_c1 bl_1 br_1 wl_228 vdd gnd cell_6t
Xbit_r229_c1 bl_1 br_1 wl_229 vdd gnd cell_6t
Xbit_r230_c1 bl_1 br_1 wl_230 vdd gnd cell_6t
Xbit_r231_c1 bl_1 br_1 wl_231 vdd gnd cell_6t
Xbit_r232_c1 bl_1 br_1 wl_232 vdd gnd cell_6t
Xbit_r233_c1 bl_1 br_1 wl_233 vdd gnd cell_6t
Xbit_r234_c1 bl_1 br_1 wl_234 vdd gnd cell_6t
Xbit_r235_c1 bl_1 br_1 wl_235 vdd gnd cell_6t
Xbit_r236_c1 bl_1 br_1 wl_236 vdd gnd cell_6t
Xbit_r237_c1 bl_1 br_1 wl_237 vdd gnd cell_6t
Xbit_r238_c1 bl_1 br_1 wl_238 vdd gnd cell_6t
Xbit_r239_c1 bl_1 br_1 wl_239 vdd gnd cell_6t
Xbit_r240_c1 bl_1 br_1 wl_240 vdd gnd cell_6t
Xbit_r241_c1 bl_1 br_1 wl_241 vdd gnd cell_6t
Xbit_r242_c1 bl_1 br_1 wl_242 vdd gnd cell_6t
Xbit_r243_c1 bl_1 br_1 wl_243 vdd gnd cell_6t
Xbit_r244_c1 bl_1 br_1 wl_244 vdd gnd cell_6t
Xbit_r245_c1 bl_1 br_1 wl_245 vdd gnd cell_6t
Xbit_r246_c1 bl_1 br_1 wl_246 vdd gnd cell_6t
Xbit_r247_c1 bl_1 br_1 wl_247 vdd gnd cell_6t
Xbit_r248_c1 bl_1 br_1 wl_248 vdd gnd cell_6t
Xbit_r249_c1 bl_1 br_1 wl_249 vdd gnd cell_6t
Xbit_r250_c1 bl_1 br_1 wl_250 vdd gnd cell_6t
Xbit_r251_c1 bl_1 br_1 wl_251 vdd gnd cell_6t
Xbit_r252_c1 bl_1 br_1 wl_252 vdd gnd cell_6t
Xbit_r253_c1 bl_1 br_1 wl_253 vdd gnd cell_6t
Xbit_r254_c1 bl_1 br_1 wl_254 vdd gnd cell_6t
Xbit_r255_c1 bl_1 br_1 wl_255 vdd gnd cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd cell_6t
Xbit_r1_c2 bl_2 br_2 wl_1 vdd gnd cell_6t
Xbit_r2_c2 bl_2 br_2 wl_2 vdd gnd cell_6t
Xbit_r3_c2 bl_2 br_2 wl_3 vdd gnd cell_6t
Xbit_r4_c2 bl_2 br_2 wl_4 vdd gnd cell_6t
Xbit_r5_c2 bl_2 br_2 wl_5 vdd gnd cell_6t
Xbit_r6_c2 bl_2 br_2 wl_6 vdd gnd cell_6t
Xbit_r7_c2 bl_2 br_2 wl_7 vdd gnd cell_6t
Xbit_r8_c2 bl_2 br_2 wl_8 vdd gnd cell_6t
Xbit_r9_c2 bl_2 br_2 wl_9 vdd gnd cell_6t
Xbit_r10_c2 bl_2 br_2 wl_10 vdd gnd cell_6t
Xbit_r11_c2 bl_2 br_2 wl_11 vdd gnd cell_6t
Xbit_r12_c2 bl_2 br_2 wl_12 vdd gnd cell_6t
Xbit_r13_c2 bl_2 br_2 wl_13 vdd gnd cell_6t
Xbit_r14_c2 bl_2 br_2 wl_14 vdd gnd cell_6t
Xbit_r15_c2 bl_2 br_2 wl_15 vdd gnd cell_6t
Xbit_r16_c2 bl_2 br_2 wl_16 vdd gnd cell_6t
Xbit_r17_c2 bl_2 br_2 wl_17 vdd gnd cell_6t
Xbit_r18_c2 bl_2 br_2 wl_18 vdd gnd cell_6t
Xbit_r19_c2 bl_2 br_2 wl_19 vdd gnd cell_6t
Xbit_r20_c2 bl_2 br_2 wl_20 vdd gnd cell_6t
Xbit_r21_c2 bl_2 br_2 wl_21 vdd gnd cell_6t
Xbit_r22_c2 bl_2 br_2 wl_22 vdd gnd cell_6t
Xbit_r23_c2 bl_2 br_2 wl_23 vdd gnd cell_6t
Xbit_r24_c2 bl_2 br_2 wl_24 vdd gnd cell_6t
Xbit_r25_c2 bl_2 br_2 wl_25 vdd gnd cell_6t
Xbit_r26_c2 bl_2 br_2 wl_26 vdd gnd cell_6t
Xbit_r27_c2 bl_2 br_2 wl_27 vdd gnd cell_6t
Xbit_r28_c2 bl_2 br_2 wl_28 vdd gnd cell_6t
Xbit_r29_c2 bl_2 br_2 wl_29 vdd gnd cell_6t
Xbit_r30_c2 bl_2 br_2 wl_30 vdd gnd cell_6t
Xbit_r31_c2 bl_2 br_2 wl_31 vdd gnd cell_6t
Xbit_r32_c2 bl_2 br_2 wl_32 vdd gnd cell_6t
Xbit_r33_c2 bl_2 br_2 wl_33 vdd gnd cell_6t
Xbit_r34_c2 bl_2 br_2 wl_34 vdd gnd cell_6t
Xbit_r35_c2 bl_2 br_2 wl_35 vdd gnd cell_6t
Xbit_r36_c2 bl_2 br_2 wl_36 vdd gnd cell_6t
Xbit_r37_c2 bl_2 br_2 wl_37 vdd gnd cell_6t
Xbit_r38_c2 bl_2 br_2 wl_38 vdd gnd cell_6t
Xbit_r39_c2 bl_2 br_2 wl_39 vdd gnd cell_6t
Xbit_r40_c2 bl_2 br_2 wl_40 vdd gnd cell_6t
Xbit_r41_c2 bl_2 br_2 wl_41 vdd gnd cell_6t
Xbit_r42_c2 bl_2 br_2 wl_42 vdd gnd cell_6t
Xbit_r43_c2 bl_2 br_2 wl_43 vdd gnd cell_6t
Xbit_r44_c2 bl_2 br_2 wl_44 vdd gnd cell_6t
Xbit_r45_c2 bl_2 br_2 wl_45 vdd gnd cell_6t
Xbit_r46_c2 bl_2 br_2 wl_46 vdd gnd cell_6t
Xbit_r47_c2 bl_2 br_2 wl_47 vdd gnd cell_6t
Xbit_r48_c2 bl_2 br_2 wl_48 vdd gnd cell_6t
Xbit_r49_c2 bl_2 br_2 wl_49 vdd gnd cell_6t
Xbit_r50_c2 bl_2 br_2 wl_50 vdd gnd cell_6t
Xbit_r51_c2 bl_2 br_2 wl_51 vdd gnd cell_6t
Xbit_r52_c2 bl_2 br_2 wl_52 vdd gnd cell_6t
Xbit_r53_c2 bl_2 br_2 wl_53 vdd gnd cell_6t
Xbit_r54_c2 bl_2 br_2 wl_54 vdd gnd cell_6t
Xbit_r55_c2 bl_2 br_2 wl_55 vdd gnd cell_6t
Xbit_r56_c2 bl_2 br_2 wl_56 vdd gnd cell_6t
Xbit_r57_c2 bl_2 br_2 wl_57 vdd gnd cell_6t
Xbit_r58_c2 bl_2 br_2 wl_58 vdd gnd cell_6t
Xbit_r59_c2 bl_2 br_2 wl_59 vdd gnd cell_6t
Xbit_r60_c2 bl_2 br_2 wl_60 vdd gnd cell_6t
Xbit_r61_c2 bl_2 br_2 wl_61 vdd gnd cell_6t
Xbit_r62_c2 bl_2 br_2 wl_62 vdd gnd cell_6t
Xbit_r63_c2 bl_2 br_2 wl_63 vdd gnd cell_6t
Xbit_r64_c2 bl_2 br_2 wl_64 vdd gnd cell_6t
Xbit_r65_c2 bl_2 br_2 wl_65 vdd gnd cell_6t
Xbit_r66_c2 bl_2 br_2 wl_66 vdd gnd cell_6t
Xbit_r67_c2 bl_2 br_2 wl_67 vdd gnd cell_6t
Xbit_r68_c2 bl_2 br_2 wl_68 vdd gnd cell_6t
Xbit_r69_c2 bl_2 br_2 wl_69 vdd gnd cell_6t
Xbit_r70_c2 bl_2 br_2 wl_70 vdd gnd cell_6t
Xbit_r71_c2 bl_2 br_2 wl_71 vdd gnd cell_6t
Xbit_r72_c2 bl_2 br_2 wl_72 vdd gnd cell_6t
Xbit_r73_c2 bl_2 br_2 wl_73 vdd gnd cell_6t
Xbit_r74_c2 bl_2 br_2 wl_74 vdd gnd cell_6t
Xbit_r75_c2 bl_2 br_2 wl_75 vdd gnd cell_6t
Xbit_r76_c2 bl_2 br_2 wl_76 vdd gnd cell_6t
Xbit_r77_c2 bl_2 br_2 wl_77 vdd gnd cell_6t
Xbit_r78_c2 bl_2 br_2 wl_78 vdd gnd cell_6t
Xbit_r79_c2 bl_2 br_2 wl_79 vdd gnd cell_6t
Xbit_r80_c2 bl_2 br_2 wl_80 vdd gnd cell_6t
Xbit_r81_c2 bl_2 br_2 wl_81 vdd gnd cell_6t
Xbit_r82_c2 bl_2 br_2 wl_82 vdd gnd cell_6t
Xbit_r83_c2 bl_2 br_2 wl_83 vdd gnd cell_6t
Xbit_r84_c2 bl_2 br_2 wl_84 vdd gnd cell_6t
Xbit_r85_c2 bl_2 br_2 wl_85 vdd gnd cell_6t
Xbit_r86_c2 bl_2 br_2 wl_86 vdd gnd cell_6t
Xbit_r87_c2 bl_2 br_2 wl_87 vdd gnd cell_6t
Xbit_r88_c2 bl_2 br_2 wl_88 vdd gnd cell_6t
Xbit_r89_c2 bl_2 br_2 wl_89 vdd gnd cell_6t
Xbit_r90_c2 bl_2 br_2 wl_90 vdd gnd cell_6t
Xbit_r91_c2 bl_2 br_2 wl_91 vdd gnd cell_6t
Xbit_r92_c2 bl_2 br_2 wl_92 vdd gnd cell_6t
Xbit_r93_c2 bl_2 br_2 wl_93 vdd gnd cell_6t
Xbit_r94_c2 bl_2 br_2 wl_94 vdd gnd cell_6t
Xbit_r95_c2 bl_2 br_2 wl_95 vdd gnd cell_6t
Xbit_r96_c2 bl_2 br_2 wl_96 vdd gnd cell_6t
Xbit_r97_c2 bl_2 br_2 wl_97 vdd gnd cell_6t
Xbit_r98_c2 bl_2 br_2 wl_98 vdd gnd cell_6t
Xbit_r99_c2 bl_2 br_2 wl_99 vdd gnd cell_6t
Xbit_r100_c2 bl_2 br_2 wl_100 vdd gnd cell_6t
Xbit_r101_c2 bl_2 br_2 wl_101 vdd gnd cell_6t
Xbit_r102_c2 bl_2 br_2 wl_102 vdd gnd cell_6t
Xbit_r103_c2 bl_2 br_2 wl_103 vdd gnd cell_6t
Xbit_r104_c2 bl_2 br_2 wl_104 vdd gnd cell_6t
Xbit_r105_c2 bl_2 br_2 wl_105 vdd gnd cell_6t
Xbit_r106_c2 bl_2 br_2 wl_106 vdd gnd cell_6t
Xbit_r107_c2 bl_2 br_2 wl_107 vdd gnd cell_6t
Xbit_r108_c2 bl_2 br_2 wl_108 vdd gnd cell_6t
Xbit_r109_c2 bl_2 br_2 wl_109 vdd gnd cell_6t
Xbit_r110_c2 bl_2 br_2 wl_110 vdd gnd cell_6t
Xbit_r111_c2 bl_2 br_2 wl_111 vdd gnd cell_6t
Xbit_r112_c2 bl_2 br_2 wl_112 vdd gnd cell_6t
Xbit_r113_c2 bl_2 br_2 wl_113 vdd gnd cell_6t
Xbit_r114_c2 bl_2 br_2 wl_114 vdd gnd cell_6t
Xbit_r115_c2 bl_2 br_2 wl_115 vdd gnd cell_6t
Xbit_r116_c2 bl_2 br_2 wl_116 vdd gnd cell_6t
Xbit_r117_c2 bl_2 br_2 wl_117 vdd gnd cell_6t
Xbit_r118_c2 bl_2 br_2 wl_118 vdd gnd cell_6t
Xbit_r119_c2 bl_2 br_2 wl_119 vdd gnd cell_6t
Xbit_r120_c2 bl_2 br_2 wl_120 vdd gnd cell_6t
Xbit_r121_c2 bl_2 br_2 wl_121 vdd gnd cell_6t
Xbit_r122_c2 bl_2 br_2 wl_122 vdd gnd cell_6t
Xbit_r123_c2 bl_2 br_2 wl_123 vdd gnd cell_6t
Xbit_r124_c2 bl_2 br_2 wl_124 vdd gnd cell_6t
Xbit_r125_c2 bl_2 br_2 wl_125 vdd gnd cell_6t
Xbit_r126_c2 bl_2 br_2 wl_126 vdd gnd cell_6t
Xbit_r127_c2 bl_2 br_2 wl_127 vdd gnd cell_6t
Xbit_r128_c2 bl_2 br_2 wl_128 vdd gnd cell_6t
Xbit_r129_c2 bl_2 br_2 wl_129 vdd gnd cell_6t
Xbit_r130_c2 bl_2 br_2 wl_130 vdd gnd cell_6t
Xbit_r131_c2 bl_2 br_2 wl_131 vdd gnd cell_6t
Xbit_r132_c2 bl_2 br_2 wl_132 vdd gnd cell_6t
Xbit_r133_c2 bl_2 br_2 wl_133 vdd gnd cell_6t
Xbit_r134_c2 bl_2 br_2 wl_134 vdd gnd cell_6t
Xbit_r135_c2 bl_2 br_2 wl_135 vdd gnd cell_6t
Xbit_r136_c2 bl_2 br_2 wl_136 vdd gnd cell_6t
Xbit_r137_c2 bl_2 br_2 wl_137 vdd gnd cell_6t
Xbit_r138_c2 bl_2 br_2 wl_138 vdd gnd cell_6t
Xbit_r139_c2 bl_2 br_2 wl_139 vdd gnd cell_6t
Xbit_r140_c2 bl_2 br_2 wl_140 vdd gnd cell_6t
Xbit_r141_c2 bl_2 br_2 wl_141 vdd gnd cell_6t
Xbit_r142_c2 bl_2 br_2 wl_142 vdd gnd cell_6t
Xbit_r143_c2 bl_2 br_2 wl_143 vdd gnd cell_6t
Xbit_r144_c2 bl_2 br_2 wl_144 vdd gnd cell_6t
Xbit_r145_c2 bl_2 br_2 wl_145 vdd gnd cell_6t
Xbit_r146_c2 bl_2 br_2 wl_146 vdd gnd cell_6t
Xbit_r147_c2 bl_2 br_2 wl_147 vdd gnd cell_6t
Xbit_r148_c2 bl_2 br_2 wl_148 vdd gnd cell_6t
Xbit_r149_c2 bl_2 br_2 wl_149 vdd gnd cell_6t
Xbit_r150_c2 bl_2 br_2 wl_150 vdd gnd cell_6t
Xbit_r151_c2 bl_2 br_2 wl_151 vdd gnd cell_6t
Xbit_r152_c2 bl_2 br_2 wl_152 vdd gnd cell_6t
Xbit_r153_c2 bl_2 br_2 wl_153 vdd gnd cell_6t
Xbit_r154_c2 bl_2 br_2 wl_154 vdd gnd cell_6t
Xbit_r155_c2 bl_2 br_2 wl_155 vdd gnd cell_6t
Xbit_r156_c2 bl_2 br_2 wl_156 vdd gnd cell_6t
Xbit_r157_c2 bl_2 br_2 wl_157 vdd gnd cell_6t
Xbit_r158_c2 bl_2 br_2 wl_158 vdd gnd cell_6t
Xbit_r159_c2 bl_2 br_2 wl_159 vdd gnd cell_6t
Xbit_r160_c2 bl_2 br_2 wl_160 vdd gnd cell_6t
Xbit_r161_c2 bl_2 br_2 wl_161 vdd gnd cell_6t
Xbit_r162_c2 bl_2 br_2 wl_162 vdd gnd cell_6t
Xbit_r163_c2 bl_2 br_2 wl_163 vdd gnd cell_6t
Xbit_r164_c2 bl_2 br_2 wl_164 vdd gnd cell_6t
Xbit_r165_c2 bl_2 br_2 wl_165 vdd gnd cell_6t
Xbit_r166_c2 bl_2 br_2 wl_166 vdd gnd cell_6t
Xbit_r167_c2 bl_2 br_2 wl_167 vdd gnd cell_6t
Xbit_r168_c2 bl_2 br_2 wl_168 vdd gnd cell_6t
Xbit_r169_c2 bl_2 br_2 wl_169 vdd gnd cell_6t
Xbit_r170_c2 bl_2 br_2 wl_170 vdd gnd cell_6t
Xbit_r171_c2 bl_2 br_2 wl_171 vdd gnd cell_6t
Xbit_r172_c2 bl_2 br_2 wl_172 vdd gnd cell_6t
Xbit_r173_c2 bl_2 br_2 wl_173 vdd gnd cell_6t
Xbit_r174_c2 bl_2 br_2 wl_174 vdd gnd cell_6t
Xbit_r175_c2 bl_2 br_2 wl_175 vdd gnd cell_6t
Xbit_r176_c2 bl_2 br_2 wl_176 vdd gnd cell_6t
Xbit_r177_c2 bl_2 br_2 wl_177 vdd gnd cell_6t
Xbit_r178_c2 bl_2 br_2 wl_178 vdd gnd cell_6t
Xbit_r179_c2 bl_2 br_2 wl_179 vdd gnd cell_6t
Xbit_r180_c2 bl_2 br_2 wl_180 vdd gnd cell_6t
Xbit_r181_c2 bl_2 br_2 wl_181 vdd gnd cell_6t
Xbit_r182_c2 bl_2 br_2 wl_182 vdd gnd cell_6t
Xbit_r183_c2 bl_2 br_2 wl_183 vdd gnd cell_6t
Xbit_r184_c2 bl_2 br_2 wl_184 vdd gnd cell_6t
Xbit_r185_c2 bl_2 br_2 wl_185 vdd gnd cell_6t
Xbit_r186_c2 bl_2 br_2 wl_186 vdd gnd cell_6t
Xbit_r187_c2 bl_2 br_2 wl_187 vdd gnd cell_6t
Xbit_r188_c2 bl_2 br_2 wl_188 vdd gnd cell_6t
Xbit_r189_c2 bl_2 br_2 wl_189 vdd gnd cell_6t
Xbit_r190_c2 bl_2 br_2 wl_190 vdd gnd cell_6t
Xbit_r191_c2 bl_2 br_2 wl_191 vdd gnd cell_6t
Xbit_r192_c2 bl_2 br_2 wl_192 vdd gnd cell_6t
Xbit_r193_c2 bl_2 br_2 wl_193 vdd gnd cell_6t
Xbit_r194_c2 bl_2 br_2 wl_194 vdd gnd cell_6t
Xbit_r195_c2 bl_2 br_2 wl_195 vdd gnd cell_6t
Xbit_r196_c2 bl_2 br_2 wl_196 vdd gnd cell_6t
Xbit_r197_c2 bl_2 br_2 wl_197 vdd gnd cell_6t
Xbit_r198_c2 bl_2 br_2 wl_198 vdd gnd cell_6t
Xbit_r199_c2 bl_2 br_2 wl_199 vdd gnd cell_6t
Xbit_r200_c2 bl_2 br_2 wl_200 vdd gnd cell_6t
Xbit_r201_c2 bl_2 br_2 wl_201 vdd gnd cell_6t
Xbit_r202_c2 bl_2 br_2 wl_202 vdd gnd cell_6t
Xbit_r203_c2 bl_2 br_2 wl_203 vdd gnd cell_6t
Xbit_r204_c2 bl_2 br_2 wl_204 vdd gnd cell_6t
Xbit_r205_c2 bl_2 br_2 wl_205 vdd gnd cell_6t
Xbit_r206_c2 bl_2 br_2 wl_206 vdd gnd cell_6t
Xbit_r207_c2 bl_2 br_2 wl_207 vdd gnd cell_6t
Xbit_r208_c2 bl_2 br_2 wl_208 vdd gnd cell_6t
Xbit_r209_c2 bl_2 br_2 wl_209 vdd gnd cell_6t
Xbit_r210_c2 bl_2 br_2 wl_210 vdd gnd cell_6t
Xbit_r211_c2 bl_2 br_2 wl_211 vdd gnd cell_6t
Xbit_r212_c2 bl_2 br_2 wl_212 vdd gnd cell_6t
Xbit_r213_c2 bl_2 br_2 wl_213 vdd gnd cell_6t
Xbit_r214_c2 bl_2 br_2 wl_214 vdd gnd cell_6t
Xbit_r215_c2 bl_2 br_2 wl_215 vdd gnd cell_6t
Xbit_r216_c2 bl_2 br_2 wl_216 vdd gnd cell_6t
Xbit_r217_c2 bl_2 br_2 wl_217 vdd gnd cell_6t
Xbit_r218_c2 bl_2 br_2 wl_218 vdd gnd cell_6t
Xbit_r219_c2 bl_2 br_2 wl_219 vdd gnd cell_6t
Xbit_r220_c2 bl_2 br_2 wl_220 vdd gnd cell_6t
Xbit_r221_c2 bl_2 br_2 wl_221 vdd gnd cell_6t
Xbit_r222_c2 bl_2 br_2 wl_222 vdd gnd cell_6t
Xbit_r223_c2 bl_2 br_2 wl_223 vdd gnd cell_6t
Xbit_r224_c2 bl_2 br_2 wl_224 vdd gnd cell_6t
Xbit_r225_c2 bl_2 br_2 wl_225 vdd gnd cell_6t
Xbit_r226_c2 bl_2 br_2 wl_226 vdd gnd cell_6t
Xbit_r227_c2 bl_2 br_2 wl_227 vdd gnd cell_6t
Xbit_r228_c2 bl_2 br_2 wl_228 vdd gnd cell_6t
Xbit_r229_c2 bl_2 br_2 wl_229 vdd gnd cell_6t
Xbit_r230_c2 bl_2 br_2 wl_230 vdd gnd cell_6t
Xbit_r231_c2 bl_2 br_2 wl_231 vdd gnd cell_6t
Xbit_r232_c2 bl_2 br_2 wl_232 vdd gnd cell_6t
Xbit_r233_c2 bl_2 br_2 wl_233 vdd gnd cell_6t
Xbit_r234_c2 bl_2 br_2 wl_234 vdd gnd cell_6t
Xbit_r235_c2 bl_2 br_2 wl_235 vdd gnd cell_6t
Xbit_r236_c2 bl_2 br_2 wl_236 vdd gnd cell_6t
Xbit_r237_c2 bl_2 br_2 wl_237 vdd gnd cell_6t
Xbit_r238_c2 bl_2 br_2 wl_238 vdd gnd cell_6t
Xbit_r239_c2 bl_2 br_2 wl_239 vdd gnd cell_6t
Xbit_r240_c2 bl_2 br_2 wl_240 vdd gnd cell_6t
Xbit_r241_c2 bl_2 br_2 wl_241 vdd gnd cell_6t
Xbit_r242_c2 bl_2 br_2 wl_242 vdd gnd cell_6t
Xbit_r243_c2 bl_2 br_2 wl_243 vdd gnd cell_6t
Xbit_r244_c2 bl_2 br_2 wl_244 vdd gnd cell_6t
Xbit_r245_c2 bl_2 br_2 wl_245 vdd gnd cell_6t
Xbit_r246_c2 bl_2 br_2 wl_246 vdd gnd cell_6t
Xbit_r247_c2 bl_2 br_2 wl_247 vdd gnd cell_6t
Xbit_r248_c2 bl_2 br_2 wl_248 vdd gnd cell_6t
Xbit_r249_c2 bl_2 br_2 wl_249 vdd gnd cell_6t
Xbit_r250_c2 bl_2 br_2 wl_250 vdd gnd cell_6t
Xbit_r251_c2 bl_2 br_2 wl_251 vdd gnd cell_6t
Xbit_r252_c2 bl_2 br_2 wl_252 vdd gnd cell_6t
Xbit_r253_c2 bl_2 br_2 wl_253 vdd gnd cell_6t
Xbit_r254_c2 bl_2 br_2 wl_254 vdd gnd cell_6t
Xbit_r255_c2 bl_2 br_2 wl_255 vdd gnd cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd cell_6t
Xbit_r1_c3 bl_3 br_3 wl_1 vdd gnd cell_6t
Xbit_r2_c3 bl_3 br_3 wl_2 vdd gnd cell_6t
Xbit_r3_c3 bl_3 br_3 wl_3 vdd gnd cell_6t
Xbit_r4_c3 bl_3 br_3 wl_4 vdd gnd cell_6t
Xbit_r5_c3 bl_3 br_3 wl_5 vdd gnd cell_6t
Xbit_r6_c3 bl_3 br_3 wl_6 vdd gnd cell_6t
Xbit_r7_c3 bl_3 br_3 wl_7 vdd gnd cell_6t
Xbit_r8_c3 bl_3 br_3 wl_8 vdd gnd cell_6t
Xbit_r9_c3 bl_3 br_3 wl_9 vdd gnd cell_6t
Xbit_r10_c3 bl_3 br_3 wl_10 vdd gnd cell_6t
Xbit_r11_c3 bl_3 br_3 wl_11 vdd gnd cell_6t
Xbit_r12_c3 bl_3 br_3 wl_12 vdd gnd cell_6t
Xbit_r13_c3 bl_3 br_3 wl_13 vdd gnd cell_6t
Xbit_r14_c3 bl_3 br_3 wl_14 vdd gnd cell_6t
Xbit_r15_c3 bl_3 br_3 wl_15 vdd gnd cell_6t
Xbit_r16_c3 bl_3 br_3 wl_16 vdd gnd cell_6t
Xbit_r17_c3 bl_3 br_3 wl_17 vdd gnd cell_6t
Xbit_r18_c3 bl_3 br_3 wl_18 vdd gnd cell_6t
Xbit_r19_c3 bl_3 br_3 wl_19 vdd gnd cell_6t
Xbit_r20_c3 bl_3 br_3 wl_20 vdd gnd cell_6t
Xbit_r21_c3 bl_3 br_3 wl_21 vdd gnd cell_6t
Xbit_r22_c3 bl_3 br_3 wl_22 vdd gnd cell_6t
Xbit_r23_c3 bl_3 br_3 wl_23 vdd gnd cell_6t
Xbit_r24_c3 bl_3 br_3 wl_24 vdd gnd cell_6t
Xbit_r25_c3 bl_3 br_3 wl_25 vdd gnd cell_6t
Xbit_r26_c3 bl_3 br_3 wl_26 vdd gnd cell_6t
Xbit_r27_c3 bl_3 br_3 wl_27 vdd gnd cell_6t
Xbit_r28_c3 bl_3 br_3 wl_28 vdd gnd cell_6t
Xbit_r29_c3 bl_3 br_3 wl_29 vdd gnd cell_6t
Xbit_r30_c3 bl_3 br_3 wl_30 vdd gnd cell_6t
Xbit_r31_c3 bl_3 br_3 wl_31 vdd gnd cell_6t
Xbit_r32_c3 bl_3 br_3 wl_32 vdd gnd cell_6t
Xbit_r33_c3 bl_3 br_3 wl_33 vdd gnd cell_6t
Xbit_r34_c3 bl_3 br_3 wl_34 vdd gnd cell_6t
Xbit_r35_c3 bl_3 br_3 wl_35 vdd gnd cell_6t
Xbit_r36_c3 bl_3 br_3 wl_36 vdd gnd cell_6t
Xbit_r37_c3 bl_3 br_3 wl_37 vdd gnd cell_6t
Xbit_r38_c3 bl_3 br_3 wl_38 vdd gnd cell_6t
Xbit_r39_c3 bl_3 br_3 wl_39 vdd gnd cell_6t
Xbit_r40_c3 bl_3 br_3 wl_40 vdd gnd cell_6t
Xbit_r41_c3 bl_3 br_3 wl_41 vdd gnd cell_6t
Xbit_r42_c3 bl_3 br_3 wl_42 vdd gnd cell_6t
Xbit_r43_c3 bl_3 br_3 wl_43 vdd gnd cell_6t
Xbit_r44_c3 bl_3 br_3 wl_44 vdd gnd cell_6t
Xbit_r45_c3 bl_3 br_3 wl_45 vdd gnd cell_6t
Xbit_r46_c3 bl_3 br_3 wl_46 vdd gnd cell_6t
Xbit_r47_c3 bl_3 br_3 wl_47 vdd gnd cell_6t
Xbit_r48_c3 bl_3 br_3 wl_48 vdd gnd cell_6t
Xbit_r49_c3 bl_3 br_3 wl_49 vdd gnd cell_6t
Xbit_r50_c3 bl_3 br_3 wl_50 vdd gnd cell_6t
Xbit_r51_c3 bl_3 br_3 wl_51 vdd gnd cell_6t
Xbit_r52_c3 bl_3 br_3 wl_52 vdd gnd cell_6t
Xbit_r53_c3 bl_3 br_3 wl_53 vdd gnd cell_6t
Xbit_r54_c3 bl_3 br_3 wl_54 vdd gnd cell_6t
Xbit_r55_c3 bl_3 br_3 wl_55 vdd gnd cell_6t
Xbit_r56_c3 bl_3 br_3 wl_56 vdd gnd cell_6t
Xbit_r57_c3 bl_3 br_3 wl_57 vdd gnd cell_6t
Xbit_r58_c3 bl_3 br_3 wl_58 vdd gnd cell_6t
Xbit_r59_c3 bl_3 br_3 wl_59 vdd gnd cell_6t
Xbit_r60_c3 bl_3 br_3 wl_60 vdd gnd cell_6t
Xbit_r61_c3 bl_3 br_3 wl_61 vdd gnd cell_6t
Xbit_r62_c3 bl_3 br_3 wl_62 vdd gnd cell_6t
Xbit_r63_c3 bl_3 br_3 wl_63 vdd gnd cell_6t
Xbit_r64_c3 bl_3 br_3 wl_64 vdd gnd cell_6t
Xbit_r65_c3 bl_3 br_3 wl_65 vdd gnd cell_6t
Xbit_r66_c3 bl_3 br_3 wl_66 vdd gnd cell_6t
Xbit_r67_c3 bl_3 br_3 wl_67 vdd gnd cell_6t
Xbit_r68_c3 bl_3 br_3 wl_68 vdd gnd cell_6t
Xbit_r69_c3 bl_3 br_3 wl_69 vdd gnd cell_6t
Xbit_r70_c3 bl_3 br_3 wl_70 vdd gnd cell_6t
Xbit_r71_c3 bl_3 br_3 wl_71 vdd gnd cell_6t
Xbit_r72_c3 bl_3 br_3 wl_72 vdd gnd cell_6t
Xbit_r73_c3 bl_3 br_3 wl_73 vdd gnd cell_6t
Xbit_r74_c3 bl_3 br_3 wl_74 vdd gnd cell_6t
Xbit_r75_c3 bl_3 br_3 wl_75 vdd gnd cell_6t
Xbit_r76_c3 bl_3 br_3 wl_76 vdd gnd cell_6t
Xbit_r77_c3 bl_3 br_3 wl_77 vdd gnd cell_6t
Xbit_r78_c3 bl_3 br_3 wl_78 vdd gnd cell_6t
Xbit_r79_c3 bl_3 br_3 wl_79 vdd gnd cell_6t
Xbit_r80_c3 bl_3 br_3 wl_80 vdd gnd cell_6t
Xbit_r81_c3 bl_3 br_3 wl_81 vdd gnd cell_6t
Xbit_r82_c3 bl_3 br_3 wl_82 vdd gnd cell_6t
Xbit_r83_c3 bl_3 br_3 wl_83 vdd gnd cell_6t
Xbit_r84_c3 bl_3 br_3 wl_84 vdd gnd cell_6t
Xbit_r85_c3 bl_3 br_3 wl_85 vdd gnd cell_6t
Xbit_r86_c3 bl_3 br_3 wl_86 vdd gnd cell_6t
Xbit_r87_c3 bl_3 br_3 wl_87 vdd gnd cell_6t
Xbit_r88_c3 bl_3 br_3 wl_88 vdd gnd cell_6t
Xbit_r89_c3 bl_3 br_3 wl_89 vdd gnd cell_6t
Xbit_r90_c3 bl_3 br_3 wl_90 vdd gnd cell_6t
Xbit_r91_c3 bl_3 br_3 wl_91 vdd gnd cell_6t
Xbit_r92_c3 bl_3 br_3 wl_92 vdd gnd cell_6t
Xbit_r93_c3 bl_3 br_3 wl_93 vdd gnd cell_6t
Xbit_r94_c3 bl_3 br_3 wl_94 vdd gnd cell_6t
Xbit_r95_c3 bl_3 br_3 wl_95 vdd gnd cell_6t
Xbit_r96_c3 bl_3 br_3 wl_96 vdd gnd cell_6t
Xbit_r97_c3 bl_3 br_3 wl_97 vdd gnd cell_6t
Xbit_r98_c3 bl_3 br_3 wl_98 vdd gnd cell_6t
Xbit_r99_c3 bl_3 br_3 wl_99 vdd gnd cell_6t
Xbit_r100_c3 bl_3 br_3 wl_100 vdd gnd cell_6t
Xbit_r101_c3 bl_3 br_3 wl_101 vdd gnd cell_6t
Xbit_r102_c3 bl_3 br_3 wl_102 vdd gnd cell_6t
Xbit_r103_c3 bl_3 br_3 wl_103 vdd gnd cell_6t
Xbit_r104_c3 bl_3 br_3 wl_104 vdd gnd cell_6t
Xbit_r105_c3 bl_3 br_3 wl_105 vdd gnd cell_6t
Xbit_r106_c3 bl_3 br_3 wl_106 vdd gnd cell_6t
Xbit_r107_c3 bl_3 br_3 wl_107 vdd gnd cell_6t
Xbit_r108_c3 bl_3 br_3 wl_108 vdd gnd cell_6t
Xbit_r109_c3 bl_3 br_3 wl_109 vdd gnd cell_6t
Xbit_r110_c3 bl_3 br_3 wl_110 vdd gnd cell_6t
Xbit_r111_c3 bl_3 br_3 wl_111 vdd gnd cell_6t
Xbit_r112_c3 bl_3 br_3 wl_112 vdd gnd cell_6t
Xbit_r113_c3 bl_3 br_3 wl_113 vdd gnd cell_6t
Xbit_r114_c3 bl_3 br_3 wl_114 vdd gnd cell_6t
Xbit_r115_c3 bl_3 br_3 wl_115 vdd gnd cell_6t
Xbit_r116_c3 bl_3 br_3 wl_116 vdd gnd cell_6t
Xbit_r117_c3 bl_3 br_3 wl_117 vdd gnd cell_6t
Xbit_r118_c3 bl_3 br_3 wl_118 vdd gnd cell_6t
Xbit_r119_c3 bl_3 br_3 wl_119 vdd gnd cell_6t
Xbit_r120_c3 bl_3 br_3 wl_120 vdd gnd cell_6t
Xbit_r121_c3 bl_3 br_3 wl_121 vdd gnd cell_6t
Xbit_r122_c3 bl_3 br_3 wl_122 vdd gnd cell_6t
Xbit_r123_c3 bl_3 br_3 wl_123 vdd gnd cell_6t
Xbit_r124_c3 bl_3 br_3 wl_124 vdd gnd cell_6t
Xbit_r125_c3 bl_3 br_3 wl_125 vdd gnd cell_6t
Xbit_r126_c3 bl_3 br_3 wl_126 vdd gnd cell_6t
Xbit_r127_c3 bl_3 br_3 wl_127 vdd gnd cell_6t
Xbit_r128_c3 bl_3 br_3 wl_128 vdd gnd cell_6t
Xbit_r129_c3 bl_3 br_3 wl_129 vdd gnd cell_6t
Xbit_r130_c3 bl_3 br_3 wl_130 vdd gnd cell_6t
Xbit_r131_c3 bl_3 br_3 wl_131 vdd gnd cell_6t
Xbit_r132_c3 bl_3 br_3 wl_132 vdd gnd cell_6t
Xbit_r133_c3 bl_3 br_3 wl_133 vdd gnd cell_6t
Xbit_r134_c3 bl_3 br_3 wl_134 vdd gnd cell_6t
Xbit_r135_c3 bl_3 br_3 wl_135 vdd gnd cell_6t
Xbit_r136_c3 bl_3 br_3 wl_136 vdd gnd cell_6t
Xbit_r137_c3 bl_3 br_3 wl_137 vdd gnd cell_6t
Xbit_r138_c3 bl_3 br_3 wl_138 vdd gnd cell_6t
Xbit_r139_c3 bl_3 br_3 wl_139 vdd gnd cell_6t
Xbit_r140_c3 bl_3 br_3 wl_140 vdd gnd cell_6t
Xbit_r141_c3 bl_3 br_3 wl_141 vdd gnd cell_6t
Xbit_r142_c3 bl_3 br_3 wl_142 vdd gnd cell_6t
Xbit_r143_c3 bl_3 br_3 wl_143 vdd gnd cell_6t
Xbit_r144_c3 bl_3 br_3 wl_144 vdd gnd cell_6t
Xbit_r145_c3 bl_3 br_3 wl_145 vdd gnd cell_6t
Xbit_r146_c3 bl_3 br_3 wl_146 vdd gnd cell_6t
Xbit_r147_c3 bl_3 br_3 wl_147 vdd gnd cell_6t
Xbit_r148_c3 bl_3 br_3 wl_148 vdd gnd cell_6t
Xbit_r149_c3 bl_3 br_3 wl_149 vdd gnd cell_6t
Xbit_r150_c3 bl_3 br_3 wl_150 vdd gnd cell_6t
Xbit_r151_c3 bl_3 br_3 wl_151 vdd gnd cell_6t
Xbit_r152_c3 bl_3 br_3 wl_152 vdd gnd cell_6t
Xbit_r153_c3 bl_3 br_3 wl_153 vdd gnd cell_6t
Xbit_r154_c3 bl_3 br_3 wl_154 vdd gnd cell_6t
Xbit_r155_c3 bl_3 br_3 wl_155 vdd gnd cell_6t
Xbit_r156_c3 bl_3 br_3 wl_156 vdd gnd cell_6t
Xbit_r157_c3 bl_3 br_3 wl_157 vdd gnd cell_6t
Xbit_r158_c3 bl_3 br_3 wl_158 vdd gnd cell_6t
Xbit_r159_c3 bl_3 br_3 wl_159 vdd gnd cell_6t
Xbit_r160_c3 bl_3 br_3 wl_160 vdd gnd cell_6t
Xbit_r161_c3 bl_3 br_3 wl_161 vdd gnd cell_6t
Xbit_r162_c3 bl_3 br_3 wl_162 vdd gnd cell_6t
Xbit_r163_c3 bl_3 br_3 wl_163 vdd gnd cell_6t
Xbit_r164_c3 bl_3 br_3 wl_164 vdd gnd cell_6t
Xbit_r165_c3 bl_3 br_3 wl_165 vdd gnd cell_6t
Xbit_r166_c3 bl_3 br_3 wl_166 vdd gnd cell_6t
Xbit_r167_c3 bl_3 br_3 wl_167 vdd gnd cell_6t
Xbit_r168_c3 bl_3 br_3 wl_168 vdd gnd cell_6t
Xbit_r169_c3 bl_3 br_3 wl_169 vdd gnd cell_6t
Xbit_r170_c3 bl_3 br_3 wl_170 vdd gnd cell_6t
Xbit_r171_c3 bl_3 br_3 wl_171 vdd gnd cell_6t
Xbit_r172_c3 bl_3 br_3 wl_172 vdd gnd cell_6t
Xbit_r173_c3 bl_3 br_3 wl_173 vdd gnd cell_6t
Xbit_r174_c3 bl_3 br_3 wl_174 vdd gnd cell_6t
Xbit_r175_c3 bl_3 br_3 wl_175 vdd gnd cell_6t
Xbit_r176_c3 bl_3 br_3 wl_176 vdd gnd cell_6t
Xbit_r177_c3 bl_3 br_3 wl_177 vdd gnd cell_6t
Xbit_r178_c3 bl_3 br_3 wl_178 vdd gnd cell_6t
Xbit_r179_c3 bl_3 br_3 wl_179 vdd gnd cell_6t
Xbit_r180_c3 bl_3 br_3 wl_180 vdd gnd cell_6t
Xbit_r181_c3 bl_3 br_3 wl_181 vdd gnd cell_6t
Xbit_r182_c3 bl_3 br_3 wl_182 vdd gnd cell_6t
Xbit_r183_c3 bl_3 br_3 wl_183 vdd gnd cell_6t
Xbit_r184_c3 bl_3 br_3 wl_184 vdd gnd cell_6t
Xbit_r185_c3 bl_3 br_3 wl_185 vdd gnd cell_6t
Xbit_r186_c3 bl_3 br_3 wl_186 vdd gnd cell_6t
Xbit_r187_c3 bl_3 br_3 wl_187 vdd gnd cell_6t
Xbit_r188_c3 bl_3 br_3 wl_188 vdd gnd cell_6t
Xbit_r189_c3 bl_3 br_3 wl_189 vdd gnd cell_6t
Xbit_r190_c3 bl_3 br_3 wl_190 vdd gnd cell_6t
Xbit_r191_c3 bl_3 br_3 wl_191 vdd gnd cell_6t
Xbit_r192_c3 bl_3 br_3 wl_192 vdd gnd cell_6t
Xbit_r193_c3 bl_3 br_3 wl_193 vdd gnd cell_6t
Xbit_r194_c3 bl_3 br_3 wl_194 vdd gnd cell_6t
Xbit_r195_c3 bl_3 br_3 wl_195 vdd gnd cell_6t
Xbit_r196_c3 bl_3 br_3 wl_196 vdd gnd cell_6t
Xbit_r197_c3 bl_3 br_3 wl_197 vdd gnd cell_6t
Xbit_r198_c3 bl_3 br_3 wl_198 vdd gnd cell_6t
Xbit_r199_c3 bl_3 br_3 wl_199 vdd gnd cell_6t
Xbit_r200_c3 bl_3 br_3 wl_200 vdd gnd cell_6t
Xbit_r201_c3 bl_3 br_3 wl_201 vdd gnd cell_6t
Xbit_r202_c3 bl_3 br_3 wl_202 vdd gnd cell_6t
Xbit_r203_c3 bl_3 br_3 wl_203 vdd gnd cell_6t
Xbit_r204_c3 bl_3 br_3 wl_204 vdd gnd cell_6t
Xbit_r205_c3 bl_3 br_3 wl_205 vdd gnd cell_6t
Xbit_r206_c3 bl_3 br_3 wl_206 vdd gnd cell_6t
Xbit_r207_c3 bl_3 br_3 wl_207 vdd gnd cell_6t
Xbit_r208_c3 bl_3 br_3 wl_208 vdd gnd cell_6t
Xbit_r209_c3 bl_3 br_3 wl_209 vdd gnd cell_6t
Xbit_r210_c3 bl_3 br_3 wl_210 vdd gnd cell_6t
Xbit_r211_c3 bl_3 br_3 wl_211 vdd gnd cell_6t
Xbit_r212_c3 bl_3 br_3 wl_212 vdd gnd cell_6t
Xbit_r213_c3 bl_3 br_3 wl_213 vdd gnd cell_6t
Xbit_r214_c3 bl_3 br_3 wl_214 vdd gnd cell_6t
Xbit_r215_c3 bl_3 br_3 wl_215 vdd gnd cell_6t
Xbit_r216_c3 bl_3 br_3 wl_216 vdd gnd cell_6t
Xbit_r217_c3 bl_3 br_3 wl_217 vdd gnd cell_6t
Xbit_r218_c3 bl_3 br_3 wl_218 vdd gnd cell_6t
Xbit_r219_c3 bl_3 br_3 wl_219 vdd gnd cell_6t
Xbit_r220_c3 bl_3 br_3 wl_220 vdd gnd cell_6t
Xbit_r221_c3 bl_3 br_3 wl_221 vdd gnd cell_6t
Xbit_r222_c3 bl_3 br_3 wl_222 vdd gnd cell_6t
Xbit_r223_c3 bl_3 br_3 wl_223 vdd gnd cell_6t
Xbit_r224_c3 bl_3 br_3 wl_224 vdd gnd cell_6t
Xbit_r225_c3 bl_3 br_3 wl_225 vdd gnd cell_6t
Xbit_r226_c3 bl_3 br_3 wl_226 vdd gnd cell_6t
Xbit_r227_c3 bl_3 br_3 wl_227 vdd gnd cell_6t
Xbit_r228_c3 bl_3 br_3 wl_228 vdd gnd cell_6t
Xbit_r229_c3 bl_3 br_3 wl_229 vdd gnd cell_6t
Xbit_r230_c3 bl_3 br_3 wl_230 vdd gnd cell_6t
Xbit_r231_c3 bl_3 br_3 wl_231 vdd gnd cell_6t
Xbit_r232_c3 bl_3 br_3 wl_232 vdd gnd cell_6t
Xbit_r233_c3 bl_3 br_3 wl_233 vdd gnd cell_6t
Xbit_r234_c3 bl_3 br_3 wl_234 vdd gnd cell_6t
Xbit_r235_c3 bl_3 br_3 wl_235 vdd gnd cell_6t
Xbit_r236_c3 bl_3 br_3 wl_236 vdd gnd cell_6t
Xbit_r237_c3 bl_3 br_3 wl_237 vdd gnd cell_6t
Xbit_r238_c3 bl_3 br_3 wl_238 vdd gnd cell_6t
Xbit_r239_c3 bl_3 br_3 wl_239 vdd gnd cell_6t
Xbit_r240_c3 bl_3 br_3 wl_240 vdd gnd cell_6t
Xbit_r241_c3 bl_3 br_3 wl_241 vdd gnd cell_6t
Xbit_r242_c3 bl_3 br_3 wl_242 vdd gnd cell_6t
Xbit_r243_c3 bl_3 br_3 wl_243 vdd gnd cell_6t
Xbit_r244_c3 bl_3 br_3 wl_244 vdd gnd cell_6t
Xbit_r245_c3 bl_3 br_3 wl_245 vdd gnd cell_6t
Xbit_r246_c3 bl_3 br_3 wl_246 vdd gnd cell_6t
Xbit_r247_c3 bl_3 br_3 wl_247 vdd gnd cell_6t
Xbit_r248_c3 bl_3 br_3 wl_248 vdd gnd cell_6t
Xbit_r249_c3 bl_3 br_3 wl_249 vdd gnd cell_6t
Xbit_r250_c3 bl_3 br_3 wl_250 vdd gnd cell_6t
Xbit_r251_c3 bl_3 br_3 wl_251 vdd gnd cell_6t
Xbit_r252_c3 bl_3 br_3 wl_252 vdd gnd cell_6t
Xbit_r253_c3 bl_3 br_3 wl_253 vdd gnd cell_6t
Xbit_r254_c3 bl_3 br_3 wl_254 vdd gnd cell_6t
Xbit_r255_c3 bl_3 br_3 wl_255 vdd gnd cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd cell_6t
Xbit_r1_c4 bl_4 br_4 wl_1 vdd gnd cell_6t
Xbit_r2_c4 bl_4 br_4 wl_2 vdd gnd cell_6t
Xbit_r3_c4 bl_4 br_4 wl_3 vdd gnd cell_6t
Xbit_r4_c4 bl_4 br_4 wl_4 vdd gnd cell_6t
Xbit_r5_c4 bl_4 br_4 wl_5 vdd gnd cell_6t
Xbit_r6_c4 bl_4 br_4 wl_6 vdd gnd cell_6t
Xbit_r7_c4 bl_4 br_4 wl_7 vdd gnd cell_6t
Xbit_r8_c4 bl_4 br_4 wl_8 vdd gnd cell_6t
Xbit_r9_c4 bl_4 br_4 wl_9 vdd gnd cell_6t
Xbit_r10_c4 bl_4 br_4 wl_10 vdd gnd cell_6t
Xbit_r11_c4 bl_4 br_4 wl_11 vdd gnd cell_6t
Xbit_r12_c4 bl_4 br_4 wl_12 vdd gnd cell_6t
Xbit_r13_c4 bl_4 br_4 wl_13 vdd gnd cell_6t
Xbit_r14_c4 bl_4 br_4 wl_14 vdd gnd cell_6t
Xbit_r15_c4 bl_4 br_4 wl_15 vdd gnd cell_6t
Xbit_r16_c4 bl_4 br_4 wl_16 vdd gnd cell_6t
Xbit_r17_c4 bl_4 br_4 wl_17 vdd gnd cell_6t
Xbit_r18_c4 bl_4 br_4 wl_18 vdd gnd cell_6t
Xbit_r19_c4 bl_4 br_4 wl_19 vdd gnd cell_6t
Xbit_r20_c4 bl_4 br_4 wl_20 vdd gnd cell_6t
Xbit_r21_c4 bl_4 br_4 wl_21 vdd gnd cell_6t
Xbit_r22_c4 bl_4 br_4 wl_22 vdd gnd cell_6t
Xbit_r23_c4 bl_4 br_4 wl_23 vdd gnd cell_6t
Xbit_r24_c4 bl_4 br_4 wl_24 vdd gnd cell_6t
Xbit_r25_c4 bl_4 br_4 wl_25 vdd gnd cell_6t
Xbit_r26_c4 bl_4 br_4 wl_26 vdd gnd cell_6t
Xbit_r27_c4 bl_4 br_4 wl_27 vdd gnd cell_6t
Xbit_r28_c4 bl_4 br_4 wl_28 vdd gnd cell_6t
Xbit_r29_c4 bl_4 br_4 wl_29 vdd gnd cell_6t
Xbit_r30_c4 bl_4 br_4 wl_30 vdd gnd cell_6t
Xbit_r31_c4 bl_4 br_4 wl_31 vdd gnd cell_6t
Xbit_r32_c4 bl_4 br_4 wl_32 vdd gnd cell_6t
Xbit_r33_c4 bl_4 br_4 wl_33 vdd gnd cell_6t
Xbit_r34_c4 bl_4 br_4 wl_34 vdd gnd cell_6t
Xbit_r35_c4 bl_4 br_4 wl_35 vdd gnd cell_6t
Xbit_r36_c4 bl_4 br_4 wl_36 vdd gnd cell_6t
Xbit_r37_c4 bl_4 br_4 wl_37 vdd gnd cell_6t
Xbit_r38_c4 bl_4 br_4 wl_38 vdd gnd cell_6t
Xbit_r39_c4 bl_4 br_4 wl_39 vdd gnd cell_6t
Xbit_r40_c4 bl_4 br_4 wl_40 vdd gnd cell_6t
Xbit_r41_c4 bl_4 br_4 wl_41 vdd gnd cell_6t
Xbit_r42_c4 bl_4 br_4 wl_42 vdd gnd cell_6t
Xbit_r43_c4 bl_4 br_4 wl_43 vdd gnd cell_6t
Xbit_r44_c4 bl_4 br_4 wl_44 vdd gnd cell_6t
Xbit_r45_c4 bl_4 br_4 wl_45 vdd gnd cell_6t
Xbit_r46_c4 bl_4 br_4 wl_46 vdd gnd cell_6t
Xbit_r47_c4 bl_4 br_4 wl_47 vdd gnd cell_6t
Xbit_r48_c4 bl_4 br_4 wl_48 vdd gnd cell_6t
Xbit_r49_c4 bl_4 br_4 wl_49 vdd gnd cell_6t
Xbit_r50_c4 bl_4 br_4 wl_50 vdd gnd cell_6t
Xbit_r51_c4 bl_4 br_4 wl_51 vdd gnd cell_6t
Xbit_r52_c4 bl_4 br_4 wl_52 vdd gnd cell_6t
Xbit_r53_c4 bl_4 br_4 wl_53 vdd gnd cell_6t
Xbit_r54_c4 bl_4 br_4 wl_54 vdd gnd cell_6t
Xbit_r55_c4 bl_4 br_4 wl_55 vdd gnd cell_6t
Xbit_r56_c4 bl_4 br_4 wl_56 vdd gnd cell_6t
Xbit_r57_c4 bl_4 br_4 wl_57 vdd gnd cell_6t
Xbit_r58_c4 bl_4 br_4 wl_58 vdd gnd cell_6t
Xbit_r59_c4 bl_4 br_4 wl_59 vdd gnd cell_6t
Xbit_r60_c4 bl_4 br_4 wl_60 vdd gnd cell_6t
Xbit_r61_c4 bl_4 br_4 wl_61 vdd gnd cell_6t
Xbit_r62_c4 bl_4 br_4 wl_62 vdd gnd cell_6t
Xbit_r63_c4 bl_4 br_4 wl_63 vdd gnd cell_6t
Xbit_r64_c4 bl_4 br_4 wl_64 vdd gnd cell_6t
Xbit_r65_c4 bl_4 br_4 wl_65 vdd gnd cell_6t
Xbit_r66_c4 bl_4 br_4 wl_66 vdd gnd cell_6t
Xbit_r67_c4 bl_4 br_4 wl_67 vdd gnd cell_6t
Xbit_r68_c4 bl_4 br_4 wl_68 vdd gnd cell_6t
Xbit_r69_c4 bl_4 br_4 wl_69 vdd gnd cell_6t
Xbit_r70_c4 bl_4 br_4 wl_70 vdd gnd cell_6t
Xbit_r71_c4 bl_4 br_4 wl_71 vdd gnd cell_6t
Xbit_r72_c4 bl_4 br_4 wl_72 vdd gnd cell_6t
Xbit_r73_c4 bl_4 br_4 wl_73 vdd gnd cell_6t
Xbit_r74_c4 bl_4 br_4 wl_74 vdd gnd cell_6t
Xbit_r75_c4 bl_4 br_4 wl_75 vdd gnd cell_6t
Xbit_r76_c4 bl_4 br_4 wl_76 vdd gnd cell_6t
Xbit_r77_c4 bl_4 br_4 wl_77 vdd gnd cell_6t
Xbit_r78_c4 bl_4 br_4 wl_78 vdd gnd cell_6t
Xbit_r79_c4 bl_4 br_4 wl_79 vdd gnd cell_6t
Xbit_r80_c4 bl_4 br_4 wl_80 vdd gnd cell_6t
Xbit_r81_c4 bl_4 br_4 wl_81 vdd gnd cell_6t
Xbit_r82_c4 bl_4 br_4 wl_82 vdd gnd cell_6t
Xbit_r83_c4 bl_4 br_4 wl_83 vdd gnd cell_6t
Xbit_r84_c4 bl_4 br_4 wl_84 vdd gnd cell_6t
Xbit_r85_c4 bl_4 br_4 wl_85 vdd gnd cell_6t
Xbit_r86_c4 bl_4 br_4 wl_86 vdd gnd cell_6t
Xbit_r87_c4 bl_4 br_4 wl_87 vdd gnd cell_6t
Xbit_r88_c4 bl_4 br_4 wl_88 vdd gnd cell_6t
Xbit_r89_c4 bl_4 br_4 wl_89 vdd gnd cell_6t
Xbit_r90_c4 bl_4 br_4 wl_90 vdd gnd cell_6t
Xbit_r91_c4 bl_4 br_4 wl_91 vdd gnd cell_6t
Xbit_r92_c4 bl_4 br_4 wl_92 vdd gnd cell_6t
Xbit_r93_c4 bl_4 br_4 wl_93 vdd gnd cell_6t
Xbit_r94_c4 bl_4 br_4 wl_94 vdd gnd cell_6t
Xbit_r95_c4 bl_4 br_4 wl_95 vdd gnd cell_6t
Xbit_r96_c4 bl_4 br_4 wl_96 vdd gnd cell_6t
Xbit_r97_c4 bl_4 br_4 wl_97 vdd gnd cell_6t
Xbit_r98_c4 bl_4 br_4 wl_98 vdd gnd cell_6t
Xbit_r99_c4 bl_4 br_4 wl_99 vdd gnd cell_6t
Xbit_r100_c4 bl_4 br_4 wl_100 vdd gnd cell_6t
Xbit_r101_c4 bl_4 br_4 wl_101 vdd gnd cell_6t
Xbit_r102_c4 bl_4 br_4 wl_102 vdd gnd cell_6t
Xbit_r103_c4 bl_4 br_4 wl_103 vdd gnd cell_6t
Xbit_r104_c4 bl_4 br_4 wl_104 vdd gnd cell_6t
Xbit_r105_c4 bl_4 br_4 wl_105 vdd gnd cell_6t
Xbit_r106_c4 bl_4 br_4 wl_106 vdd gnd cell_6t
Xbit_r107_c4 bl_4 br_4 wl_107 vdd gnd cell_6t
Xbit_r108_c4 bl_4 br_4 wl_108 vdd gnd cell_6t
Xbit_r109_c4 bl_4 br_4 wl_109 vdd gnd cell_6t
Xbit_r110_c4 bl_4 br_4 wl_110 vdd gnd cell_6t
Xbit_r111_c4 bl_4 br_4 wl_111 vdd gnd cell_6t
Xbit_r112_c4 bl_4 br_4 wl_112 vdd gnd cell_6t
Xbit_r113_c4 bl_4 br_4 wl_113 vdd gnd cell_6t
Xbit_r114_c4 bl_4 br_4 wl_114 vdd gnd cell_6t
Xbit_r115_c4 bl_4 br_4 wl_115 vdd gnd cell_6t
Xbit_r116_c4 bl_4 br_4 wl_116 vdd gnd cell_6t
Xbit_r117_c4 bl_4 br_4 wl_117 vdd gnd cell_6t
Xbit_r118_c4 bl_4 br_4 wl_118 vdd gnd cell_6t
Xbit_r119_c4 bl_4 br_4 wl_119 vdd gnd cell_6t
Xbit_r120_c4 bl_4 br_4 wl_120 vdd gnd cell_6t
Xbit_r121_c4 bl_4 br_4 wl_121 vdd gnd cell_6t
Xbit_r122_c4 bl_4 br_4 wl_122 vdd gnd cell_6t
Xbit_r123_c4 bl_4 br_4 wl_123 vdd gnd cell_6t
Xbit_r124_c4 bl_4 br_4 wl_124 vdd gnd cell_6t
Xbit_r125_c4 bl_4 br_4 wl_125 vdd gnd cell_6t
Xbit_r126_c4 bl_4 br_4 wl_126 vdd gnd cell_6t
Xbit_r127_c4 bl_4 br_4 wl_127 vdd gnd cell_6t
Xbit_r128_c4 bl_4 br_4 wl_128 vdd gnd cell_6t
Xbit_r129_c4 bl_4 br_4 wl_129 vdd gnd cell_6t
Xbit_r130_c4 bl_4 br_4 wl_130 vdd gnd cell_6t
Xbit_r131_c4 bl_4 br_4 wl_131 vdd gnd cell_6t
Xbit_r132_c4 bl_4 br_4 wl_132 vdd gnd cell_6t
Xbit_r133_c4 bl_4 br_4 wl_133 vdd gnd cell_6t
Xbit_r134_c4 bl_4 br_4 wl_134 vdd gnd cell_6t
Xbit_r135_c4 bl_4 br_4 wl_135 vdd gnd cell_6t
Xbit_r136_c4 bl_4 br_4 wl_136 vdd gnd cell_6t
Xbit_r137_c4 bl_4 br_4 wl_137 vdd gnd cell_6t
Xbit_r138_c4 bl_4 br_4 wl_138 vdd gnd cell_6t
Xbit_r139_c4 bl_4 br_4 wl_139 vdd gnd cell_6t
Xbit_r140_c4 bl_4 br_4 wl_140 vdd gnd cell_6t
Xbit_r141_c4 bl_4 br_4 wl_141 vdd gnd cell_6t
Xbit_r142_c4 bl_4 br_4 wl_142 vdd gnd cell_6t
Xbit_r143_c4 bl_4 br_4 wl_143 vdd gnd cell_6t
Xbit_r144_c4 bl_4 br_4 wl_144 vdd gnd cell_6t
Xbit_r145_c4 bl_4 br_4 wl_145 vdd gnd cell_6t
Xbit_r146_c4 bl_4 br_4 wl_146 vdd gnd cell_6t
Xbit_r147_c4 bl_4 br_4 wl_147 vdd gnd cell_6t
Xbit_r148_c4 bl_4 br_4 wl_148 vdd gnd cell_6t
Xbit_r149_c4 bl_4 br_4 wl_149 vdd gnd cell_6t
Xbit_r150_c4 bl_4 br_4 wl_150 vdd gnd cell_6t
Xbit_r151_c4 bl_4 br_4 wl_151 vdd gnd cell_6t
Xbit_r152_c4 bl_4 br_4 wl_152 vdd gnd cell_6t
Xbit_r153_c4 bl_4 br_4 wl_153 vdd gnd cell_6t
Xbit_r154_c4 bl_4 br_4 wl_154 vdd gnd cell_6t
Xbit_r155_c4 bl_4 br_4 wl_155 vdd gnd cell_6t
Xbit_r156_c4 bl_4 br_4 wl_156 vdd gnd cell_6t
Xbit_r157_c4 bl_4 br_4 wl_157 vdd gnd cell_6t
Xbit_r158_c4 bl_4 br_4 wl_158 vdd gnd cell_6t
Xbit_r159_c4 bl_4 br_4 wl_159 vdd gnd cell_6t
Xbit_r160_c4 bl_4 br_4 wl_160 vdd gnd cell_6t
Xbit_r161_c4 bl_4 br_4 wl_161 vdd gnd cell_6t
Xbit_r162_c4 bl_4 br_4 wl_162 vdd gnd cell_6t
Xbit_r163_c4 bl_4 br_4 wl_163 vdd gnd cell_6t
Xbit_r164_c4 bl_4 br_4 wl_164 vdd gnd cell_6t
Xbit_r165_c4 bl_4 br_4 wl_165 vdd gnd cell_6t
Xbit_r166_c4 bl_4 br_4 wl_166 vdd gnd cell_6t
Xbit_r167_c4 bl_4 br_4 wl_167 vdd gnd cell_6t
Xbit_r168_c4 bl_4 br_4 wl_168 vdd gnd cell_6t
Xbit_r169_c4 bl_4 br_4 wl_169 vdd gnd cell_6t
Xbit_r170_c4 bl_4 br_4 wl_170 vdd gnd cell_6t
Xbit_r171_c4 bl_4 br_4 wl_171 vdd gnd cell_6t
Xbit_r172_c4 bl_4 br_4 wl_172 vdd gnd cell_6t
Xbit_r173_c4 bl_4 br_4 wl_173 vdd gnd cell_6t
Xbit_r174_c4 bl_4 br_4 wl_174 vdd gnd cell_6t
Xbit_r175_c4 bl_4 br_4 wl_175 vdd gnd cell_6t
Xbit_r176_c4 bl_4 br_4 wl_176 vdd gnd cell_6t
Xbit_r177_c4 bl_4 br_4 wl_177 vdd gnd cell_6t
Xbit_r178_c4 bl_4 br_4 wl_178 vdd gnd cell_6t
Xbit_r179_c4 bl_4 br_4 wl_179 vdd gnd cell_6t
Xbit_r180_c4 bl_4 br_4 wl_180 vdd gnd cell_6t
Xbit_r181_c4 bl_4 br_4 wl_181 vdd gnd cell_6t
Xbit_r182_c4 bl_4 br_4 wl_182 vdd gnd cell_6t
Xbit_r183_c4 bl_4 br_4 wl_183 vdd gnd cell_6t
Xbit_r184_c4 bl_4 br_4 wl_184 vdd gnd cell_6t
Xbit_r185_c4 bl_4 br_4 wl_185 vdd gnd cell_6t
Xbit_r186_c4 bl_4 br_4 wl_186 vdd gnd cell_6t
Xbit_r187_c4 bl_4 br_4 wl_187 vdd gnd cell_6t
Xbit_r188_c4 bl_4 br_4 wl_188 vdd gnd cell_6t
Xbit_r189_c4 bl_4 br_4 wl_189 vdd gnd cell_6t
Xbit_r190_c4 bl_4 br_4 wl_190 vdd gnd cell_6t
Xbit_r191_c4 bl_4 br_4 wl_191 vdd gnd cell_6t
Xbit_r192_c4 bl_4 br_4 wl_192 vdd gnd cell_6t
Xbit_r193_c4 bl_4 br_4 wl_193 vdd gnd cell_6t
Xbit_r194_c4 bl_4 br_4 wl_194 vdd gnd cell_6t
Xbit_r195_c4 bl_4 br_4 wl_195 vdd gnd cell_6t
Xbit_r196_c4 bl_4 br_4 wl_196 vdd gnd cell_6t
Xbit_r197_c4 bl_4 br_4 wl_197 vdd gnd cell_6t
Xbit_r198_c4 bl_4 br_4 wl_198 vdd gnd cell_6t
Xbit_r199_c4 bl_4 br_4 wl_199 vdd gnd cell_6t
Xbit_r200_c4 bl_4 br_4 wl_200 vdd gnd cell_6t
Xbit_r201_c4 bl_4 br_4 wl_201 vdd gnd cell_6t
Xbit_r202_c4 bl_4 br_4 wl_202 vdd gnd cell_6t
Xbit_r203_c4 bl_4 br_4 wl_203 vdd gnd cell_6t
Xbit_r204_c4 bl_4 br_4 wl_204 vdd gnd cell_6t
Xbit_r205_c4 bl_4 br_4 wl_205 vdd gnd cell_6t
Xbit_r206_c4 bl_4 br_4 wl_206 vdd gnd cell_6t
Xbit_r207_c4 bl_4 br_4 wl_207 vdd gnd cell_6t
Xbit_r208_c4 bl_4 br_4 wl_208 vdd gnd cell_6t
Xbit_r209_c4 bl_4 br_4 wl_209 vdd gnd cell_6t
Xbit_r210_c4 bl_4 br_4 wl_210 vdd gnd cell_6t
Xbit_r211_c4 bl_4 br_4 wl_211 vdd gnd cell_6t
Xbit_r212_c4 bl_4 br_4 wl_212 vdd gnd cell_6t
Xbit_r213_c4 bl_4 br_4 wl_213 vdd gnd cell_6t
Xbit_r214_c4 bl_4 br_4 wl_214 vdd gnd cell_6t
Xbit_r215_c4 bl_4 br_4 wl_215 vdd gnd cell_6t
Xbit_r216_c4 bl_4 br_4 wl_216 vdd gnd cell_6t
Xbit_r217_c4 bl_4 br_4 wl_217 vdd gnd cell_6t
Xbit_r218_c4 bl_4 br_4 wl_218 vdd gnd cell_6t
Xbit_r219_c4 bl_4 br_4 wl_219 vdd gnd cell_6t
Xbit_r220_c4 bl_4 br_4 wl_220 vdd gnd cell_6t
Xbit_r221_c4 bl_4 br_4 wl_221 vdd gnd cell_6t
Xbit_r222_c4 bl_4 br_4 wl_222 vdd gnd cell_6t
Xbit_r223_c4 bl_4 br_4 wl_223 vdd gnd cell_6t
Xbit_r224_c4 bl_4 br_4 wl_224 vdd gnd cell_6t
Xbit_r225_c4 bl_4 br_4 wl_225 vdd gnd cell_6t
Xbit_r226_c4 bl_4 br_4 wl_226 vdd gnd cell_6t
Xbit_r227_c4 bl_4 br_4 wl_227 vdd gnd cell_6t
Xbit_r228_c4 bl_4 br_4 wl_228 vdd gnd cell_6t
Xbit_r229_c4 bl_4 br_4 wl_229 vdd gnd cell_6t
Xbit_r230_c4 bl_4 br_4 wl_230 vdd gnd cell_6t
Xbit_r231_c4 bl_4 br_4 wl_231 vdd gnd cell_6t
Xbit_r232_c4 bl_4 br_4 wl_232 vdd gnd cell_6t
Xbit_r233_c4 bl_4 br_4 wl_233 vdd gnd cell_6t
Xbit_r234_c4 bl_4 br_4 wl_234 vdd gnd cell_6t
Xbit_r235_c4 bl_4 br_4 wl_235 vdd gnd cell_6t
Xbit_r236_c4 bl_4 br_4 wl_236 vdd gnd cell_6t
Xbit_r237_c4 bl_4 br_4 wl_237 vdd gnd cell_6t
Xbit_r238_c4 bl_4 br_4 wl_238 vdd gnd cell_6t
Xbit_r239_c4 bl_4 br_4 wl_239 vdd gnd cell_6t
Xbit_r240_c4 bl_4 br_4 wl_240 vdd gnd cell_6t
Xbit_r241_c4 bl_4 br_4 wl_241 vdd gnd cell_6t
Xbit_r242_c4 bl_4 br_4 wl_242 vdd gnd cell_6t
Xbit_r243_c4 bl_4 br_4 wl_243 vdd gnd cell_6t
Xbit_r244_c4 bl_4 br_4 wl_244 vdd gnd cell_6t
Xbit_r245_c4 bl_4 br_4 wl_245 vdd gnd cell_6t
Xbit_r246_c4 bl_4 br_4 wl_246 vdd gnd cell_6t
Xbit_r247_c4 bl_4 br_4 wl_247 vdd gnd cell_6t
Xbit_r248_c4 bl_4 br_4 wl_248 vdd gnd cell_6t
Xbit_r249_c4 bl_4 br_4 wl_249 vdd gnd cell_6t
Xbit_r250_c4 bl_4 br_4 wl_250 vdd gnd cell_6t
Xbit_r251_c4 bl_4 br_4 wl_251 vdd gnd cell_6t
Xbit_r252_c4 bl_4 br_4 wl_252 vdd gnd cell_6t
Xbit_r253_c4 bl_4 br_4 wl_253 vdd gnd cell_6t
Xbit_r254_c4 bl_4 br_4 wl_254 vdd gnd cell_6t
Xbit_r255_c4 bl_4 br_4 wl_255 vdd gnd cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd cell_6t
Xbit_r1_c5 bl_5 br_5 wl_1 vdd gnd cell_6t
Xbit_r2_c5 bl_5 br_5 wl_2 vdd gnd cell_6t
Xbit_r3_c5 bl_5 br_5 wl_3 vdd gnd cell_6t
Xbit_r4_c5 bl_5 br_5 wl_4 vdd gnd cell_6t
Xbit_r5_c5 bl_5 br_5 wl_5 vdd gnd cell_6t
Xbit_r6_c5 bl_5 br_5 wl_6 vdd gnd cell_6t
Xbit_r7_c5 bl_5 br_5 wl_7 vdd gnd cell_6t
Xbit_r8_c5 bl_5 br_5 wl_8 vdd gnd cell_6t
Xbit_r9_c5 bl_5 br_5 wl_9 vdd gnd cell_6t
Xbit_r10_c5 bl_5 br_5 wl_10 vdd gnd cell_6t
Xbit_r11_c5 bl_5 br_5 wl_11 vdd gnd cell_6t
Xbit_r12_c5 bl_5 br_5 wl_12 vdd gnd cell_6t
Xbit_r13_c5 bl_5 br_5 wl_13 vdd gnd cell_6t
Xbit_r14_c5 bl_5 br_5 wl_14 vdd gnd cell_6t
Xbit_r15_c5 bl_5 br_5 wl_15 vdd gnd cell_6t
Xbit_r16_c5 bl_5 br_5 wl_16 vdd gnd cell_6t
Xbit_r17_c5 bl_5 br_5 wl_17 vdd gnd cell_6t
Xbit_r18_c5 bl_5 br_5 wl_18 vdd gnd cell_6t
Xbit_r19_c5 bl_5 br_5 wl_19 vdd gnd cell_6t
Xbit_r20_c5 bl_5 br_5 wl_20 vdd gnd cell_6t
Xbit_r21_c5 bl_5 br_5 wl_21 vdd gnd cell_6t
Xbit_r22_c5 bl_5 br_5 wl_22 vdd gnd cell_6t
Xbit_r23_c5 bl_5 br_5 wl_23 vdd gnd cell_6t
Xbit_r24_c5 bl_5 br_5 wl_24 vdd gnd cell_6t
Xbit_r25_c5 bl_5 br_5 wl_25 vdd gnd cell_6t
Xbit_r26_c5 bl_5 br_5 wl_26 vdd gnd cell_6t
Xbit_r27_c5 bl_5 br_5 wl_27 vdd gnd cell_6t
Xbit_r28_c5 bl_5 br_5 wl_28 vdd gnd cell_6t
Xbit_r29_c5 bl_5 br_5 wl_29 vdd gnd cell_6t
Xbit_r30_c5 bl_5 br_5 wl_30 vdd gnd cell_6t
Xbit_r31_c5 bl_5 br_5 wl_31 vdd gnd cell_6t
Xbit_r32_c5 bl_5 br_5 wl_32 vdd gnd cell_6t
Xbit_r33_c5 bl_5 br_5 wl_33 vdd gnd cell_6t
Xbit_r34_c5 bl_5 br_5 wl_34 vdd gnd cell_6t
Xbit_r35_c5 bl_5 br_5 wl_35 vdd gnd cell_6t
Xbit_r36_c5 bl_5 br_5 wl_36 vdd gnd cell_6t
Xbit_r37_c5 bl_5 br_5 wl_37 vdd gnd cell_6t
Xbit_r38_c5 bl_5 br_5 wl_38 vdd gnd cell_6t
Xbit_r39_c5 bl_5 br_5 wl_39 vdd gnd cell_6t
Xbit_r40_c5 bl_5 br_5 wl_40 vdd gnd cell_6t
Xbit_r41_c5 bl_5 br_5 wl_41 vdd gnd cell_6t
Xbit_r42_c5 bl_5 br_5 wl_42 vdd gnd cell_6t
Xbit_r43_c5 bl_5 br_5 wl_43 vdd gnd cell_6t
Xbit_r44_c5 bl_5 br_5 wl_44 vdd gnd cell_6t
Xbit_r45_c5 bl_5 br_5 wl_45 vdd gnd cell_6t
Xbit_r46_c5 bl_5 br_5 wl_46 vdd gnd cell_6t
Xbit_r47_c5 bl_5 br_5 wl_47 vdd gnd cell_6t
Xbit_r48_c5 bl_5 br_5 wl_48 vdd gnd cell_6t
Xbit_r49_c5 bl_5 br_5 wl_49 vdd gnd cell_6t
Xbit_r50_c5 bl_5 br_5 wl_50 vdd gnd cell_6t
Xbit_r51_c5 bl_5 br_5 wl_51 vdd gnd cell_6t
Xbit_r52_c5 bl_5 br_5 wl_52 vdd gnd cell_6t
Xbit_r53_c5 bl_5 br_5 wl_53 vdd gnd cell_6t
Xbit_r54_c5 bl_5 br_5 wl_54 vdd gnd cell_6t
Xbit_r55_c5 bl_5 br_5 wl_55 vdd gnd cell_6t
Xbit_r56_c5 bl_5 br_5 wl_56 vdd gnd cell_6t
Xbit_r57_c5 bl_5 br_5 wl_57 vdd gnd cell_6t
Xbit_r58_c5 bl_5 br_5 wl_58 vdd gnd cell_6t
Xbit_r59_c5 bl_5 br_5 wl_59 vdd gnd cell_6t
Xbit_r60_c5 bl_5 br_5 wl_60 vdd gnd cell_6t
Xbit_r61_c5 bl_5 br_5 wl_61 vdd gnd cell_6t
Xbit_r62_c5 bl_5 br_5 wl_62 vdd gnd cell_6t
Xbit_r63_c5 bl_5 br_5 wl_63 vdd gnd cell_6t
Xbit_r64_c5 bl_5 br_5 wl_64 vdd gnd cell_6t
Xbit_r65_c5 bl_5 br_5 wl_65 vdd gnd cell_6t
Xbit_r66_c5 bl_5 br_5 wl_66 vdd gnd cell_6t
Xbit_r67_c5 bl_5 br_5 wl_67 vdd gnd cell_6t
Xbit_r68_c5 bl_5 br_5 wl_68 vdd gnd cell_6t
Xbit_r69_c5 bl_5 br_5 wl_69 vdd gnd cell_6t
Xbit_r70_c5 bl_5 br_5 wl_70 vdd gnd cell_6t
Xbit_r71_c5 bl_5 br_5 wl_71 vdd gnd cell_6t
Xbit_r72_c5 bl_5 br_5 wl_72 vdd gnd cell_6t
Xbit_r73_c5 bl_5 br_5 wl_73 vdd gnd cell_6t
Xbit_r74_c5 bl_5 br_5 wl_74 vdd gnd cell_6t
Xbit_r75_c5 bl_5 br_5 wl_75 vdd gnd cell_6t
Xbit_r76_c5 bl_5 br_5 wl_76 vdd gnd cell_6t
Xbit_r77_c5 bl_5 br_5 wl_77 vdd gnd cell_6t
Xbit_r78_c5 bl_5 br_5 wl_78 vdd gnd cell_6t
Xbit_r79_c5 bl_5 br_5 wl_79 vdd gnd cell_6t
Xbit_r80_c5 bl_5 br_5 wl_80 vdd gnd cell_6t
Xbit_r81_c5 bl_5 br_5 wl_81 vdd gnd cell_6t
Xbit_r82_c5 bl_5 br_5 wl_82 vdd gnd cell_6t
Xbit_r83_c5 bl_5 br_5 wl_83 vdd gnd cell_6t
Xbit_r84_c5 bl_5 br_5 wl_84 vdd gnd cell_6t
Xbit_r85_c5 bl_5 br_5 wl_85 vdd gnd cell_6t
Xbit_r86_c5 bl_5 br_5 wl_86 vdd gnd cell_6t
Xbit_r87_c5 bl_5 br_5 wl_87 vdd gnd cell_6t
Xbit_r88_c5 bl_5 br_5 wl_88 vdd gnd cell_6t
Xbit_r89_c5 bl_5 br_5 wl_89 vdd gnd cell_6t
Xbit_r90_c5 bl_5 br_5 wl_90 vdd gnd cell_6t
Xbit_r91_c5 bl_5 br_5 wl_91 vdd gnd cell_6t
Xbit_r92_c5 bl_5 br_5 wl_92 vdd gnd cell_6t
Xbit_r93_c5 bl_5 br_5 wl_93 vdd gnd cell_6t
Xbit_r94_c5 bl_5 br_5 wl_94 vdd gnd cell_6t
Xbit_r95_c5 bl_5 br_5 wl_95 vdd gnd cell_6t
Xbit_r96_c5 bl_5 br_5 wl_96 vdd gnd cell_6t
Xbit_r97_c5 bl_5 br_5 wl_97 vdd gnd cell_6t
Xbit_r98_c5 bl_5 br_5 wl_98 vdd gnd cell_6t
Xbit_r99_c5 bl_5 br_5 wl_99 vdd gnd cell_6t
Xbit_r100_c5 bl_5 br_5 wl_100 vdd gnd cell_6t
Xbit_r101_c5 bl_5 br_5 wl_101 vdd gnd cell_6t
Xbit_r102_c5 bl_5 br_5 wl_102 vdd gnd cell_6t
Xbit_r103_c5 bl_5 br_5 wl_103 vdd gnd cell_6t
Xbit_r104_c5 bl_5 br_5 wl_104 vdd gnd cell_6t
Xbit_r105_c5 bl_5 br_5 wl_105 vdd gnd cell_6t
Xbit_r106_c5 bl_5 br_5 wl_106 vdd gnd cell_6t
Xbit_r107_c5 bl_5 br_5 wl_107 vdd gnd cell_6t
Xbit_r108_c5 bl_5 br_5 wl_108 vdd gnd cell_6t
Xbit_r109_c5 bl_5 br_5 wl_109 vdd gnd cell_6t
Xbit_r110_c5 bl_5 br_5 wl_110 vdd gnd cell_6t
Xbit_r111_c5 bl_5 br_5 wl_111 vdd gnd cell_6t
Xbit_r112_c5 bl_5 br_5 wl_112 vdd gnd cell_6t
Xbit_r113_c5 bl_5 br_5 wl_113 vdd gnd cell_6t
Xbit_r114_c5 bl_5 br_5 wl_114 vdd gnd cell_6t
Xbit_r115_c5 bl_5 br_5 wl_115 vdd gnd cell_6t
Xbit_r116_c5 bl_5 br_5 wl_116 vdd gnd cell_6t
Xbit_r117_c5 bl_5 br_5 wl_117 vdd gnd cell_6t
Xbit_r118_c5 bl_5 br_5 wl_118 vdd gnd cell_6t
Xbit_r119_c5 bl_5 br_5 wl_119 vdd gnd cell_6t
Xbit_r120_c5 bl_5 br_5 wl_120 vdd gnd cell_6t
Xbit_r121_c5 bl_5 br_5 wl_121 vdd gnd cell_6t
Xbit_r122_c5 bl_5 br_5 wl_122 vdd gnd cell_6t
Xbit_r123_c5 bl_5 br_5 wl_123 vdd gnd cell_6t
Xbit_r124_c5 bl_5 br_5 wl_124 vdd gnd cell_6t
Xbit_r125_c5 bl_5 br_5 wl_125 vdd gnd cell_6t
Xbit_r126_c5 bl_5 br_5 wl_126 vdd gnd cell_6t
Xbit_r127_c5 bl_5 br_5 wl_127 vdd gnd cell_6t
Xbit_r128_c5 bl_5 br_5 wl_128 vdd gnd cell_6t
Xbit_r129_c5 bl_5 br_5 wl_129 vdd gnd cell_6t
Xbit_r130_c5 bl_5 br_5 wl_130 vdd gnd cell_6t
Xbit_r131_c5 bl_5 br_5 wl_131 vdd gnd cell_6t
Xbit_r132_c5 bl_5 br_5 wl_132 vdd gnd cell_6t
Xbit_r133_c5 bl_5 br_5 wl_133 vdd gnd cell_6t
Xbit_r134_c5 bl_5 br_5 wl_134 vdd gnd cell_6t
Xbit_r135_c5 bl_5 br_5 wl_135 vdd gnd cell_6t
Xbit_r136_c5 bl_5 br_5 wl_136 vdd gnd cell_6t
Xbit_r137_c5 bl_5 br_5 wl_137 vdd gnd cell_6t
Xbit_r138_c5 bl_5 br_5 wl_138 vdd gnd cell_6t
Xbit_r139_c5 bl_5 br_5 wl_139 vdd gnd cell_6t
Xbit_r140_c5 bl_5 br_5 wl_140 vdd gnd cell_6t
Xbit_r141_c5 bl_5 br_5 wl_141 vdd gnd cell_6t
Xbit_r142_c5 bl_5 br_5 wl_142 vdd gnd cell_6t
Xbit_r143_c5 bl_5 br_5 wl_143 vdd gnd cell_6t
Xbit_r144_c5 bl_5 br_5 wl_144 vdd gnd cell_6t
Xbit_r145_c5 bl_5 br_5 wl_145 vdd gnd cell_6t
Xbit_r146_c5 bl_5 br_5 wl_146 vdd gnd cell_6t
Xbit_r147_c5 bl_5 br_5 wl_147 vdd gnd cell_6t
Xbit_r148_c5 bl_5 br_5 wl_148 vdd gnd cell_6t
Xbit_r149_c5 bl_5 br_5 wl_149 vdd gnd cell_6t
Xbit_r150_c5 bl_5 br_5 wl_150 vdd gnd cell_6t
Xbit_r151_c5 bl_5 br_5 wl_151 vdd gnd cell_6t
Xbit_r152_c5 bl_5 br_5 wl_152 vdd gnd cell_6t
Xbit_r153_c5 bl_5 br_5 wl_153 vdd gnd cell_6t
Xbit_r154_c5 bl_5 br_5 wl_154 vdd gnd cell_6t
Xbit_r155_c5 bl_5 br_5 wl_155 vdd gnd cell_6t
Xbit_r156_c5 bl_5 br_5 wl_156 vdd gnd cell_6t
Xbit_r157_c5 bl_5 br_5 wl_157 vdd gnd cell_6t
Xbit_r158_c5 bl_5 br_5 wl_158 vdd gnd cell_6t
Xbit_r159_c5 bl_5 br_5 wl_159 vdd gnd cell_6t
Xbit_r160_c5 bl_5 br_5 wl_160 vdd gnd cell_6t
Xbit_r161_c5 bl_5 br_5 wl_161 vdd gnd cell_6t
Xbit_r162_c5 bl_5 br_5 wl_162 vdd gnd cell_6t
Xbit_r163_c5 bl_5 br_5 wl_163 vdd gnd cell_6t
Xbit_r164_c5 bl_5 br_5 wl_164 vdd gnd cell_6t
Xbit_r165_c5 bl_5 br_5 wl_165 vdd gnd cell_6t
Xbit_r166_c5 bl_5 br_5 wl_166 vdd gnd cell_6t
Xbit_r167_c5 bl_5 br_5 wl_167 vdd gnd cell_6t
Xbit_r168_c5 bl_5 br_5 wl_168 vdd gnd cell_6t
Xbit_r169_c5 bl_5 br_5 wl_169 vdd gnd cell_6t
Xbit_r170_c5 bl_5 br_5 wl_170 vdd gnd cell_6t
Xbit_r171_c5 bl_5 br_5 wl_171 vdd gnd cell_6t
Xbit_r172_c5 bl_5 br_5 wl_172 vdd gnd cell_6t
Xbit_r173_c5 bl_5 br_5 wl_173 vdd gnd cell_6t
Xbit_r174_c5 bl_5 br_5 wl_174 vdd gnd cell_6t
Xbit_r175_c5 bl_5 br_5 wl_175 vdd gnd cell_6t
Xbit_r176_c5 bl_5 br_5 wl_176 vdd gnd cell_6t
Xbit_r177_c5 bl_5 br_5 wl_177 vdd gnd cell_6t
Xbit_r178_c5 bl_5 br_5 wl_178 vdd gnd cell_6t
Xbit_r179_c5 bl_5 br_5 wl_179 vdd gnd cell_6t
Xbit_r180_c5 bl_5 br_5 wl_180 vdd gnd cell_6t
Xbit_r181_c5 bl_5 br_5 wl_181 vdd gnd cell_6t
Xbit_r182_c5 bl_5 br_5 wl_182 vdd gnd cell_6t
Xbit_r183_c5 bl_5 br_5 wl_183 vdd gnd cell_6t
Xbit_r184_c5 bl_5 br_5 wl_184 vdd gnd cell_6t
Xbit_r185_c5 bl_5 br_5 wl_185 vdd gnd cell_6t
Xbit_r186_c5 bl_5 br_5 wl_186 vdd gnd cell_6t
Xbit_r187_c5 bl_5 br_5 wl_187 vdd gnd cell_6t
Xbit_r188_c5 bl_5 br_5 wl_188 vdd gnd cell_6t
Xbit_r189_c5 bl_5 br_5 wl_189 vdd gnd cell_6t
Xbit_r190_c5 bl_5 br_5 wl_190 vdd gnd cell_6t
Xbit_r191_c5 bl_5 br_5 wl_191 vdd gnd cell_6t
Xbit_r192_c5 bl_5 br_5 wl_192 vdd gnd cell_6t
Xbit_r193_c5 bl_5 br_5 wl_193 vdd gnd cell_6t
Xbit_r194_c5 bl_5 br_5 wl_194 vdd gnd cell_6t
Xbit_r195_c5 bl_5 br_5 wl_195 vdd gnd cell_6t
Xbit_r196_c5 bl_5 br_5 wl_196 vdd gnd cell_6t
Xbit_r197_c5 bl_5 br_5 wl_197 vdd gnd cell_6t
Xbit_r198_c5 bl_5 br_5 wl_198 vdd gnd cell_6t
Xbit_r199_c5 bl_5 br_5 wl_199 vdd gnd cell_6t
Xbit_r200_c5 bl_5 br_5 wl_200 vdd gnd cell_6t
Xbit_r201_c5 bl_5 br_5 wl_201 vdd gnd cell_6t
Xbit_r202_c5 bl_5 br_5 wl_202 vdd gnd cell_6t
Xbit_r203_c5 bl_5 br_5 wl_203 vdd gnd cell_6t
Xbit_r204_c5 bl_5 br_5 wl_204 vdd gnd cell_6t
Xbit_r205_c5 bl_5 br_5 wl_205 vdd gnd cell_6t
Xbit_r206_c5 bl_5 br_5 wl_206 vdd gnd cell_6t
Xbit_r207_c5 bl_5 br_5 wl_207 vdd gnd cell_6t
Xbit_r208_c5 bl_5 br_5 wl_208 vdd gnd cell_6t
Xbit_r209_c5 bl_5 br_5 wl_209 vdd gnd cell_6t
Xbit_r210_c5 bl_5 br_5 wl_210 vdd gnd cell_6t
Xbit_r211_c5 bl_5 br_5 wl_211 vdd gnd cell_6t
Xbit_r212_c5 bl_5 br_5 wl_212 vdd gnd cell_6t
Xbit_r213_c5 bl_5 br_5 wl_213 vdd gnd cell_6t
Xbit_r214_c5 bl_5 br_5 wl_214 vdd gnd cell_6t
Xbit_r215_c5 bl_5 br_5 wl_215 vdd gnd cell_6t
Xbit_r216_c5 bl_5 br_5 wl_216 vdd gnd cell_6t
Xbit_r217_c5 bl_5 br_5 wl_217 vdd gnd cell_6t
Xbit_r218_c5 bl_5 br_5 wl_218 vdd gnd cell_6t
Xbit_r219_c5 bl_5 br_5 wl_219 vdd gnd cell_6t
Xbit_r220_c5 bl_5 br_5 wl_220 vdd gnd cell_6t
Xbit_r221_c5 bl_5 br_5 wl_221 vdd gnd cell_6t
Xbit_r222_c5 bl_5 br_5 wl_222 vdd gnd cell_6t
Xbit_r223_c5 bl_5 br_5 wl_223 vdd gnd cell_6t
Xbit_r224_c5 bl_5 br_5 wl_224 vdd gnd cell_6t
Xbit_r225_c5 bl_5 br_5 wl_225 vdd gnd cell_6t
Xbit_r226_c5 bl_5 br_5 wl_226 vdd gnd cell_6t
Xbit_r227_c5 bl_5 br_5 wl_227 vdd gnd cell_6t
Xbit_r228_c5 bl_5 br_5 wl_228 vdd gnd cell_6t
Xbit_r229_c5 bl_5 br_5 wl_229 vdd gnd cell_6t
Xbit_r230_c5 bl_5 br_5 wl_230 vdd gnd cell_6t
Xbit_r231_c5 bl_5 br_5 wl_231 vdd gnd cell_6t
Xbit_r232_c5 bl_5 br_5 wl_232 vdd gnd cell_6t
Xbit_r233_c5 bl_5 br_5 wl_233 vdd gnd cell_6t
Xbit_r234_c5 bl_5 br_5 wl_234 vdd gnd cell_6t
Xbit_r235_c5 bl_5 br_5 wl_235 vdd gnd cell_6t
Xbit_r236_c5 bl_5 br_5 wl_236 vdd gnd cell_6t
Xbit_r237_c5 bl_5 br_5 wl_237 vdd gnd cell_6t
Xbit_r238_c5 bl_5 br_5 wl_238 vdd gnd cell_6t
Xbit_r239_c5 bl_5 br_5 wl_239 vdd gnd cell_6t
Xbit_r240_c5 bl_5 br_5 wl_240 vdd gnd cell_6t
Xbit_r241_c5 bl_5 br_5 wl_241 vdd gnd cell_6t
Xbit_r242_c5 bl_5 br_5 wl_242 vdd gnd cell_6t
Xbit_r243_c5 bl_5 br_5 wl_243 vdd gnd cell_6t
Xbit_r244_c5 bl_5 br_5 wl_244 vdd gnd cell_6t
Xbit_r245_c5 bl_5 br_5 wl_245 vdd gnd cell_6t
Xbit_r246_c5 bl_5 br_5 wl_246 vdd gnd cell_6t
Xbit_r247_c5 bl_5 br_5 wl_247 vdd gnd cell_6t
Xbit_r248_c5 bl_5 br_5 wl_248 vdd gnd cell_6t
Xbit_r249_c5 bl_5 br_5 wl_249 vdd gnd cell_6t
Xbit_r250_c5 bl_5 br_5 wl_250 vdd gnd cell_6t
Xbit_r251_c5 bl_5 br_5 wl_251 vdd gnd cell_6t
Xbit_r252_c5 bl_5 br_5 wl_252 vdd gnd cell_6t
Xbit_r253_c5 bl_5 br_5 wl_253 vdd gnd cell_6t
Xbit_r254_c5 bl_5 br_5 wl_254 vdd gnd cell_6t
Xbit_r255_c5 bl_5 br_5 wl_255 vdd gnd cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd cell_6t
Xbit_r1_c6 bl_6 br_6 wl_1 vdd gnd cell_6t
Xbit_r2_c6 bl_6 br_6 wl_2 vdd gnd cell_6t
Xbit_r3_c6 bl_6 br_6 wl_3 vdd gnd cell_6t
Xbit_r4_c6 bl_6 br_6 wl_4 vdd gnd cell_6t
Xbit_r5_c6 bl_6 br_6 wl_5 vdd gnd cell_6t
Xbit_r6_c6 bl_6 br_6 wl_6 vdd gnd cell_6t
Xbit_r7_c6 bl_6 br_6 wl_7 vdd gnd cell_6t
Xbit_r8_c6 bl_6 br_6 wl_8 vdd gnd cell_6t
Xbit_r9_c6 bl_6 br_6 wl_9 vdd gnd cell_6t
Xbit_r10_c6 bl_6 br_6 wl_10 vdd gnd cell_6t
Xbit_r11_c6 bl_6 br_6 wl_11 vdd gnd cell_6t
Xbit_r12_c6 bl_6 br_6 wl_12 vdd gnd cell_6t
Xbit_r13_c6 bl_6 br_6 wl_13 vdd gnd cell_6t
Xbit_r14_c6 bl_6 br_6 wl_14 vdd gnd cell_6t
Xbit_r15_c6 bl_6 br_6 wl_15 vdd gnd cell_6t
Xbit_r16_c6 bl_6 br_6 wl_16 vdd gnd cell_6t
Xbit_r17_c6 bl_6 br_6 wl_17 vdd gnd cell_6t
Xbit_r18_c6 bl_6 br_6 wl_18 vdd gnd cell_6t
Xbit_r19_c6 bl_6 br_6 wl_19 vdd gnd cell_6t
Xbit_r20_c6 bl_6 br_6 wl_20 vdd gnd cell_6t
Xbit_r21_c6 bl_6 br_6 wl_21 vdd gnd cell_6t
Xbit_r22_c6 bl_6 br_6 wl_22 vdd gnd cell_6t
Xbit_r23_c6 bl_6 br_6 wl_23 vdd gnd cell_6t
Xbit_r24_c6 bl_6 br_6 wl_24 vdd gnd cell_6t
Xbit_r25_c6 bl_6 br_6 wl_25 vdd gnd cell_6t
Xbit_r26_c6 bl_6 br_6 wl_26 vdd gnd cell_6t
Xbit_r27_c6 bl_6 br_6 wl_27 vdd gnd cell_6t
Xbit_r28_c6 bl_6 br_6 wl_28 vdd gnd cell_6t
Xbit_r29_c6 bl_6 br_6 wl_29 vdd gnd cell_6t
Xbit_r30_c6 bl_6 br_6 wl_30 vdd gnd cell_6t
Xbit_r31_c6 bl_6 br_6 wl_31 vdd gnd cell_6t
Xbit_r32_c6 bl_6 br_6 wl_32 vdd gnd cell_6t
Xbit_r33_c6 bl_6 br_6 wl_33 vdd gnd cell_6t
Xbit_r34_c6 bl_6 br_6 wl_34 vdd gnd cell_6t
Xbit_r35_c6 bl_6 br_6 wl_35 vdd gnd cell_6t
Xbit_r36_c6 bl_6 br_6 wl_36 vdd gnd cell_6t
Xbit_r37_c6 bl_6 br_6 wl_37 vdd gnd cell_6t
Xbit_r38_c6 bl_6 br_6 wl_38 vdd gnd cell_6t
Xbit_r39_c6 bl_6 br_6 wl_39 vdd gnd cell_6t
Xbit_r40_c6 bl_6 br_6 wl_40 vdd gnd cell_6t
Xbit_r41_c6 bl_6 br_6 wl_41 vdd gnd cell_6t
Xbit_r42_c6 bl_6 br_6 wl_42 vdd gnd cell_6t
Xbit_r43_c6 bl_6 br_6 wl_43 vdd gnd cell_6t
Xbit_r44_c6 bl_6 br_6 wl_44 vdd gnd cell_6t
Xbit_r45_c6 bl_6 br_6 wl_45 vdd gnd cell_6t
Xbit_r46_c6 bl_6 br_6 wl_46 vdd gnd cell_6t
Xbit_r47_c6 bl_6 br_6 wl_47 vdd gnd cell_6t
Xbit_r48_c6 bl_6 br_6 wl_48 vdd gnd cell_6t
Xbit_r49_c6 bl_6 br_6 wl_49 vdd gnd cell_6t
Xbit_r50_c6 bl_6 br_6 wl_50 vdd gnd cell_6t
Xbit_r51_c6 bl_6 br_6 wl_51 vdd gnd cell_6t
Xbit_r52_c6 bl_6 br_6 wl_52 vdd gnd cell_6t
Xbit_r53_c6 bl_6 br_6 wl_53 vdd gnd cell_6t
Xbit_r54_c6 bl_6 br_6 wl_54 vdd gnd cell_6t
Xbit_r55_c6 bl_6 br_6 wl_55 vdd gnd cell_6t
Xbit_r56_c6 bl_6 br_6 wl_56 vdd gnd cell_6t
Xbit_r57_c6 bl_6 br_6 wl_57 vdd gnd cell_6t
Xbit_r58_c6 bl_6 br_6 wl_58 vdd gnd cell_6t
Xbit_r59_c6 bl_6 br_6 wl_59 vdd gnd cell_6t
Xbit_r60_c6 bl_6 br_6 wl_60 vdd gnd cell_6t
Xbit_r61_c6 bl_6 br_6 wl_61 vdd gnd cell_6t
Xbit_r62_c6 bl_6 br_6 wl_62 vdd gnd cell_6t
Xbit_r63_c6 bl_6 br_6 wl_63 vdd gnd cell_6t
Xbit_r64_c6 bl_6 br_6 wl_64 vdd gnd cell_6t
Xbit_r65_c6 bl_6 br_6 wl_65 vdd gnd cell_6t
Xbit_r66_c6 bl_6 br_6 wl_66 vdd gnd cell_6t
Xbit_r67_c6 bl_6 br_6 wl_67 vdd gnd cell_6t
Xbit_r68_c6 bl_6 br_6 wl_68 vdd gnd cell_6t
Xbit_r69_c6 bl_6 br_6 wl_69 vdd gnd cell_6t
Xbit_r70_c6 bl_6 br_6 wl_70 vdd gnd cell_6t
Xbit_r71_c6 bl_6 br_6 wl_71 vdd gnd cell_6t
Xbit_r72_c6 bl_6 br_6 wl_72 vdd gnd cell_6t
Xbit_r73_c6 bl_6 br_6 wl_73 vdd gnd cell_6t
Xbit_r74_c6 bl_6 br_6 wl_74 vdd gnd cell_6t
Xbit_r75_c6 bl_6 br_6 wl_75 vdd gnd cell_6t
Xbit_r76_c6 bl_6 br_6 wl_76 vdd gnd cell_6t
Xbit_r77_c6 bl_6 br_6 wl_77 vdd gnd cell_6t
Xbit_r78_c6 bl_6 br_6 wl_78 vdd gnd cell_6t
Xbit_r79_c6 bl_6 br_6 wl_79 vdd gnd cell_6t
Xbit_r80_c6 bl_6 br_6 wl_80 vdd gnd cell_6t
Xbit_r81_c6 bl_6 br_6 wl_81 vdd gnd cell_6t
Xbit_r82_c6 bl_6 br_6 wl_82 vdd gnd cell_6t
Xbit_r83_c6 bl_6 br_6 wl_83 vdd gnd cell_6t
Xbit_r84_c6 bl_6 br_6 wl_84 vdd gnd cell_6t
Xbit_r85_c6 bl_6 br_6 wl_85 vdd gnd cell_6t
Xbit_r86_c6 bl_6 br_6 wl_86 vdd gnd cell_6t
Xbit_r87_c6 bl_6 br_6 wl_87 vdd gnd cell_6t
Xbit_r88_c6 bl_6 br_6 wl_88 vdd gnd cell_6t
Xbit_r89_c6 bl_6 br_6 wl_89 vdd gnd cell_6t
Xbit_r90_c6 bl_6 br_6 wl_90 vdd gnd cell_6t
Xbit_r91_c6 bl_6 br_6 wl_91 vdd gnd cell_6t
Xbit_r92_c6 bl_6 br_6 wl_92 vdd gnd cell_6t
Xbit_r93_c6 bl_6 br_6 wl_93 vdd gnd cell_6t
Xbit_r94_c6 bl_6 br_6 wl_94 vdd gnd cell_6t
Xbit_r95_c6 bl_6 br_6 wl_95 vdd gnd cell_6t
Xbit_r96_c6 bl_6 br_6 wl_96 vdd gnd cell_6t
Xbit_r97_c6 bl_6 br_6 wl_97 vdd gnd cell_6t
Xbit_r98_c6 bl_6 br_6 wl_98 vdd gnd cell_6t
Xbit_r99_c6 bl_6 br_6 wl_99 vdd gnd cell_6t
Xbit_r100_c6 bl_6 br_6 wl_100 vdd gnd cell_6t
Xbit_r101_c6 bl_6 br_6 wl_101 vdd gnd cell_6t
Xbit_r102_c6 bl_6 br_6 wl_102 vdd gnd cell_6t
Xbit_r103_c6 bl_6 br_6 wl_103 vdd gnd cell_6t
Xbit_r104_c6 bl_6 br_6 wl_104 vdd gnd cell_6t
Xbit_r105_c6 bl_6 br_6 wl_105 vdd gnd cell_6t
Xbit_r106_c6 bl_6 br_6 wl_106 vdd gnd cell_6t
Xbit_r107_c6 bl_6 br_6 wl_107 vdd gnd cell_6t
Xbit_r108_c6 bl_6 br_6 wl_108 vdd gnd cell_6t
Xbit_r109_c6 bl_6 br_6 wl_109 vdd gnd cell_6t
Xbit_r110_c6 bl_6 br_6 wl_110 vdd gnd cell_6t
Xbit_r111_c6 bl_6 br_6 wl_111 vdd gnd cell_6t
Xbit_r112_c6 bl_6 br_6 wl_112 vdd gnd cell_6t
Xbit_r113_c6 bl_6 br_6 wl_113 vdd gnd cell_6t
Xbit_r114_c6 bl_6 br_6 wl_114 vdd gnd cell_6t
Xbit_r115_c6 bl_6 br_6 wl_115 vdd gnd cell_6t
Xbit_r116_c6 bl_6 br_6 wl_116 vdd gnd cell_6t
Xbit_r117_c6 bl_6 br_6 wl_117 vdd gnd cell_6t
Xbit_r118_c6 bl_6 br_6 wl_118 vdd gnd cell_6t
Xbit_r119_c6 bl_6 br_6 wl_119 vdd gnd cell_6t
Xbit_r120_c6 bl_6 br_6 wl_120 vdd gnd cell_6t
Xbit_r121_c6 bl_6 br_6 wl_121 vdd gnd cell_6t
Xbit_r122_c6 bl_6 br_6 wl_122 vdd gnd cell_6t
Xbit_r123_c6 bl_6 br_6 wl_123 vdd gnd cell_6t
Xbit_r124_c6 bl_6 br_6 wl_124 vdd gnd cell_6t
Xbit_r125_c6 bl_6 br_6 wl_125 vdd gnd cell_6t
Xbit_r126_c6 bl_6 br_6 wl_126 vdd gnd cell_6t
Xbit_r127_c6 bl_6 br_6 wl_127 vdd gnd cell_6t
Xbit_r128_c6 bl_6 br_6 wl_128 vdd gnd cell_6t
Xbit_r129_c6 bl_6 br_6 wl_129 vdd gnd cell_6t
Xbit_r130_c6 bl_6 br_6 wl_130 vdd gnd cell_6t
Xbit_r131_c6 bl_6 br_6 wl_131 vdd gnd cell_6t
Xbit_r132_c6 bl_6 br_6 wl_132 vdd gnd cell_6t
Xbit_r133_c6 bl_6 br_6 wl_133 vdd gnd cell_6t
Xbit_r134_c6 bl_6 br_6 wl_134 vdd gnd cell_6t
Xbit_r135_c6 bl_6 br_6 wl_135 vdd gnd cell_6t
Xbit_r136_c6 bl_6 br_6 wl_136 vdd gnd cell_6t
Xbit_r137_c6 bl_6 br_6 wl_137 vdd gnd cell_6t
Xbit_r138_c6 bl_6 br_6 wl_138 vdd gnd cell_6t
Xbit_r139_c6 bl_6 br_6 wl_139 vdd gnd cell_6t
Xbit_r140_c6 bl_6 br_6 wl_140 vdd gnd cell_6t
Xbit_r141_c6 bl_6 br_6 wl_141 vdd gnd cell_6t
Xbit_r142_c6 bl_6 br_6 wl_142 vdd gnd cell_6t
Xbit_r143_c6 bl_6 br_6 wl_143 vdd gnd cell_6t
Xbit_r144_c6 bl_6 br_6 wl_144 vdd gnd cell_6t
Xbit_r145_c6 bl_6 br_6 wl_145 vdd gnd cell_6t
Xbit_r146_c6 bl_6 br_6 wl_146 vdd gnd cell_6t
Xbit_r147_c6 bl_6 br_6 wl_147 vdd gnd cell_6t
Xbit_r148_c6 bl_6 br_6 wl_148 vdd gnd cell_6t
Xbit_r149_c6 bl_6 br_6 wl_149 vdd gnd cell_6t
Xbit_r150_c6 bl_6 br_6 wl_150 vdd gnd cell_6t
Xbit_r151_c6 bl_6 br_6 wl_151 vdd gnd cell_6t
Xbit_r152_c6 bl_6 br_6 wl_152 vdd gnd cell_6t
Xbit_r153_c6 bl_6 br_6 wl_153 vdd gnd cell_6t
Xbit_r154_c6 bl_6 br_6 wl_154 vdd gnd cell_6t
Xbit_r155_c6 bl_6 br_6 wl_155 vdd gnd cell_6t
Xbit_r156_c6 bl_6 br_6 wl_156 vdd gnd cell_6t
Xbit_r157_c6 bl_6 br_6 wl_157 vdd gnd cell_6t
Xbit_r158_c6 bl_6 br_6 wl_158 vdd gnd cell_6t
Xbit_r159_c6 bl_6 br_6 wl_159 vdd gnd cell_6t
Xbit_r160_c6 bl_6 br_6 wl_160 vdd gnd cell_6t
Xbit_r161_c6 bl_6 br_6 wl_161 vdd gnd cell_6t
Xbit_r162_c6 bl_6 br_6 wl_162 vdd gnd cell_6t
Xbit_r163_c6 bl_6 br_6 wl_163 vdd gnd cell_6t
Xbit_r164_c6 bl_6 br_6 wl_164 vdd gnd cell_6t
Xbit_r165_c6 bl_6 br_6 wl_165 vdd gnd cell_6t
Xbit_r166_c6 bl_6 br_6 wl_166 vdd gnd cell_6t
Xbit_r167_c6 bl_6 br_6 wl_167 vdd gnd cell_6t
Xbit_r168_c6 bl_6 br_6 wl_168 vdd gnd cell_6t
Xbit_r169_c6 bl_6 br_6 wl_169 vdd gnd cell_6t
Xbit_r170_c6 bl_6 br_6 wl_170 vdd gnd cell_6t
Xbit_r171_c6 bl_6 br_6 wl_171 vdd gnd cell_6t
Xbit_r172_c6 bl_6 br_6 wl_172 vdd gnd cell_6t
Xbit_r173_c6 bl_6 br_6 wl_173 vdd gnd cell_6t
Xbit_r174_c6 bl_6 br_6 wl_174 vdd gnd cell_6t
Xbit_r175_c6 bl_6 br_6 wl_175 vdd gnd cell_6t
Xbit_r176_c6 bl_6 br_6 wl_176 vdd gnd cell_6t
Xbit_r177_c6 bl_6 br_6 wl_177 vdd gnd cell_6t
Xbit_r178_c6 bl_6 br_6 wl_178 vdd gnd cell_6t
Xbit_r179_c6 bl_6 br_6 wl_179 vdd gnd cell_6t
Xbit_r180_c6 bl_6 br_6 wl_180 vdd gnd cell_6t
Xbit_r181_c6 bl_6 br_6 wl_181 vdd gnd cell_6t
Xbit_r182_c6 bl_6 br_6 wl_182 vdd gnd cell_6t
Xbit_r183_c6 bl_6 br_6 wl_183 vdd gnd cell_6t
Xbit_r184_c6 bl_6 br_6 wl_184 vdd gnd cell_6t
Xbit_r185_c6 bl_6 br_6 wl_185 vdd gnd cell_6t
Xbit_r186_c6 bl_6 br_6 wl_186 vdd gnd cell_6t
Xbit_r187_c6 bl_6 br_6 wl_187 vdd gnd cell_6t
Xbit_r188_c6 bl_6 br_6 wl_188 vdd gnd cell_6t
Xbit_r189_c6 bl_6 br_6 wl_189 vdd gnd cell_6t
Xbit_r190_c6 bl_6 br_6 wl_190 vdd gnd cell_6t
Xbit_r191_c6 bl_6 br_6 wl_191 vdd gnd cell_6t
Xbit_r192_c6 bl_6 br_6 wl_192 vdd gnd cell_6t
Xbit_r193_c6 bl_6 br_6 wl_193 vdd gnd cell_6t
Xbit_r194_c6 bl_6 br_6 wl_194 vdd gnd cell_6t
Xbit_r195_c6 bl_6 br_6 wl_195 vdd gnd cell_6t
Xbit_r196_c6 bl_6 br_6 wl_196 vdd gnd cell_6t
Xbit_r197_c6 bl_6 br_6 wl_197 vdd gnd cell_6t
Xbit_r198_c6 bl_6 br_6 wl_198 vdd gnd cell_6t
Xbit_r199_c6 bl_6 br_6 wl_199 vdd gnd cell_6t
Xbit_r200_c6 bl_6 br_6 wl_200 vdd gnd cell_6t
Xbit_r201_c6 bl_6 br_6 wl_201 vdd gnd cell_6t
Xbit_r202_c6 bl_6 br_6 wl_202 vdd gnd cell_6t
Xbit_r203_c6 bl_6 br_6 wl_203 vdd gnd cell_6t
Xbit_r204_c6 bl_6 br_6 wl_204 vdd gnd cell_6t
Xbit_r205_c6 bl_6 br_6 wl_205 vdd gnd cell_6t
Xbit_r206_c6 bl_6 br_6 wl_206 vdd gnd cell_6t
Xbit_r207_c6 bl_6 br_6 wl_207 vdd gnd cell_6t
Xbit_r208_c6 bl_6 br_6 wl_208 vdd gnd cell_6t
Xbit_r209_c6 bl_6 br_6 wl_209 vdd gnd cell_6t
Xbit_r210_c6 bl_6 br_6 wl_210 vdd gnd cell_6t
Xbit_r211_c6 bl_6 br_6 wl_211 vdd gnd cell_6t
Xbit_r212_c6 bl_6 br_6 wl_212 vdd gnd cell_6t
Xbit_r213_c6 bl_6 br_6 wl_213 vdd gnd cell_6t
Xbit_r214_c6 bl_6 br_6 wl_214 vdd gnd cell_6t
Xbit_r215_c6 bl_6 br_6 wl_215 vdd gnd cell_6t
Xbit_r216_c6 bl_6 br_6 wl_216 vdd gnd cell_6t
Xbit_r217_c6 bl_6 br_6 wl_217 vdd gnd cell_6t
Xbit_r218_c6 bl_6 br_6 wl_218 vdd gnd cell_6t
Xbit_r219_c6 bl_6 br_6 wl_219 vdd gnd cell_6t
Xbit_r220_c6 bl_6 br_6 wl_220 vdd gnd cell_6t
Xbit_r221_c6 bl_6 br_6 wl_221 vdd gnd cell_6t
Xbit_r222_c6 bl_6 br_6 wl_222 vdd gnd cell_6t
Xbit_r223_c6 bl_6 br_6 wl_223 vdd gnd cell_6t
Xbit_r224_c6 bl_6 br_6 wl_224 vdd gnd cell_6t
Xbit_r225_c6 bl_6 br_6 wl_225 vdd gnd cell_6t
Xbit_r226_c6 bl_6 br_6 wl_226 vdd gnd cell_6t
Xbit_r227_c6 bl_6 br_6 wl_227 vdd gnd cell_6t
Xbit_r228_c6 bl_6 br_6 wl_228 vdd gnd cell_6t
Xbit_r229_c6 bl_6 br_6 wl_229 vdd gnd cell_6t
Xbit_r230_c6 bl_6 br_6 wl_230 vdd gnd cell_6t
Xbit_r231_c6 bl_6 br_6 wl_231 vdd gnd cell_6t
Xbit_r232_c6 bl_6 br_6 wl_232 vdd gnd cell_6t
Xbit_r233_c6 bl_6 br_6 wl_233 vdd gnd cell_6t
Xbit_r234_c6 bl_6 br_6 wl_234 vdd gnd cell_6t
Xbit_r235_c6 bl_6 br_6 wl_235 vdd gnd cell_6t
Xbit_r236_c6 bl_6 br_6 wl_236 vdd gnd cell_6t
Xbit_r237_c6 bl_6 br_6 wl_237 vdd gnd cell_6t
Xbit_r238_c6 bl_6 br_6 wl_238 vdd gnd cell_6t
Xbit_r239_c6 bl_6 br_6 wl_239 vdd gnd cell_6t
Xbit_r240_c6 bl_6 br_6 wl_240 vdd gnd cell_6t
Xbit_r241_c6 bl_6 br_6 wl_241 vdd gnd cell_6t
Xbit_r242_c6 bl_6 br_6 wl_242 vdd gnd cell_6t
Xbit_r243_c6 bl_6 br_6 wl_243 vdd gnd cell_6t
Xbit_r244_c6 bl_6 br_6 wl_244 vdd gnd cell_6t
Xbit_r245_c6 bl_6 br_6 wl_245 vdd gnd cell_6t
Xbit_r246_c6 bl_6 br_6 wl_246 vdd gnd cell_6t
Xbit_r247_c6 bl_6 br_6 wl_247 vdd gnd cell_6t
Xbit_r248_c6 bl_6 br_6 wl_248 vdd gnd cell_6t
Xbit_r249_c6 bl_6 br_6 wl_249 vdd gnd cell_6t
Xbit_r250_c6 bl_6 br_6 wl_250 vdd gnd cell_6t
Xbit_r251_c6 bl_6 br_6 wl_251 vdd gnd cell_6t
Xbit_r252_c6 bl_6 br_6 wl_252 vdd gnd cell_6t
Xbit_r253_c6 bl_6 br_6 wl_253 vdd gnd cell_6t
Xbit_r254_c6 bl_6 br_6 wl_254 vdd gnd cell_6t
Xbit_r255_c6 bl_6 br_6 wl_255 vdd gnd cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd cell_6t
Xbit_r1_c7 bl_7 br_7 wl_1 vdd gnd cell_6t
Xbit_r2_c7 bl_7 br_7 wl_2 vdd gnd cell_6t
Xbit_r3_c7 bl_7 br_7 wl_3 vdd gnd cell_6t
Xbit_r4_c7 bl_7 br_7 wl_4 vdd gnd cell_6t
Xbit_r5_c7 bl_7 br_7 wl_5 vdd gnd cell_6t
Xbit_r6_c7 bl_7 br_7 wl_6 vdd gnd cell_6t
Xbit_r7_c7 bl_7 br_7 wl_7 vdd gnd cell_6t
Xbit_r8_c7 bl_7 br_7 wl_8 vdd gnd cell_6t
Xbit_r9_c7 bl_7 br_7 wl_9 vdd gnd cell_6t
Xbit_r10_c7 bl_7 br_7 wl_10 vdd gnd cell_6t
Xbit_r11_c7 bl_7 br_7 wl_11 vdd gnd cell_6t
Xbit_r12_c7 bl_7 br_7 wl_12 vdd gnd cell_6t
Xbit_r13_c7 bl_7 br_7 wl_13 vdd gnd cell_6t
Xbit_r14_c7 bl_7 br_7 wl_14 vdd gnd cell_6t
Xbit_r15_c7 bl_7 br_7 wl_15 vdd gnd cell_6t
Xbit_r16_c7 bl_7 br_7 wl_16 vdd gnd cell_6t
Xbit_r17_c7 bl_7 br_7 wl_17 vdd gnd cell_6t
Xbit_r18_c7 bl_7 br_7 wl_18 vdd gnd cell_6t
Xbit_r19_c7 bl_7 br_7 wl_19 vdd gnd cell_6t
Xbit_r20_c7 bl_7 br_7 wl_20 vdd gnd cell_6t
Xbit_r21_c7 bl_7 br_7 wl_21 vdd gnd cell_6t
Xbit_r22_c7 bl_7 br_7 wl_22 vdd gnd cell_6t
Xbit_r23_c7 bl_7 br_7 wl_23 vdd gnd cell_6t
Xbit_r24_c7 bl_7 br_7 wl_24 vdd gnd cell_6t
Xbit_r25_c7 bl_7 br_7 wl_25 vdd gnd cell_6t
Xbit_r26_c7 bl_7 br_7 wl_26 vdd gnd cell_6t
Xbit_r27_c7 bl_7 br_7 wl_27 vdd gnd cell_6t
Xbit_r28_c7 bl_7 br_7 wl_28 vdd gnd cell_6t
Xbit_r29_c7 bl_7 br_7 wl_29 vdd gnd cell_6t
Xbit_r30_c7 bl_7 br_7 wl_30 vdd gnd cell_6t
Xbit_r31_c7 bl_7 br_7 wl_31 vdd gnd cell_6t
Xbit_r32_c7 bl_7 br_7 wl_32 vdd gnd cell_6t
Xbit_r33_c7 bl_7 br_7 wl_33 vdd gnd cell_6t
Xbit_r34_c7 bl_7 br_7 wl_34 vdd gnd cell_6t
Xbit_r35_c7 bl_7 br_7 wl_35 vdd gnd cell_6t
Xbit_r36_c7 bl_7 br_7 wl_36 vdd gnd cell_6t
Xbit_r37_c7 bl_7 br_7 wl_37 vdd gnd cell_6t
Xbit_r38_c7 bl_7 br_7 wl_38 vdd gnd cell_6t
Xbit_r39_c7 bl_7 br_7 wl_39 vdd gnd cell_6t
Xbit_r40_c7 bl_7 br_7 wl_40 vdd gnd cell_6t
Xbit_r41_c7 bl_7 br_7 wl_41 vdd gnd cell_6t
Xbit_r42_c7 bl_7 br_7 wl_42 vdd gnd cell_6t
Xbit_r43_c7 bl_7 br_7 wl_43 vdd gnd cell_6t
Xbit_r44_c7 bl_7 br_7 wl_44 vdd gnd cell_6t
Xbit_r45_c7 bl_7 br_7 wl_45 vdd gnd cell_6t
Xbit_r46_c7 bl_7 br_7 wl_46 vdd gnd cell_6t
Xbit_r47_c7 bl_7 br_7 wl_47 vdd gnd cell_6t
Xbit_r48_c7 bl_7 br_7 wl_48 vdd gnd cell_6t
Xbit_r49_c7 bl_7 br_7 wl_49 vdd gnd cell_6t
Xbit_r50_c7 bl_7 br_7 wl_50 vdd gnd cell_6t
Xbit_r51_c7 bl_7 br_7 wl_51 vdd gnd cell_6t
Xbit_r52_c7 bl_7 br_7 wl_52 vdd gnd cell_6t
Xbit_r53_c7 bl_7 br_7 wl_53 vdd gnd cell_6t
Xbit_r54_c7 bl_7 br_7 wl_54 vdd gnd cell_6t
Xbit_r55_c7 bl_7 br_7 wl_55 vdd gnd cell_6t
Xbit_r56_c7 bl_7 br_7 wl_56 vdd gnd cell_6t
Xbit_r57_c7 bl_7 br_7 wl_57 vdd gnd cell_6t
Xbit_r58_c7 bl_7 br_7 wl_58 vdd gnd cell_6t
Xbit_r59_c7 bl_7 br_7 wl_59 vdd gnd cell_6t
Xbit_r60_c7 bl_7 br_7 wl_60 vdd gnd cell_6t
Xbit_r61_c7 bl_7 br_7 wl_61 vdd gnd cell_6t
Xbit_r62_c7 bl_7 br_7 wl_62 vdd gnd cell_6t
Xbit_r63_c7 bl_7 br_7 wl_63 vdd gnd cell_6t
Xbit_r64_c7 bl_7 br_7 wl_64 vdd gnd cell_6t
Xbit_r65_c7 bl_7 br_7 wl_65 vdd gnd cell_6t
Xbit_r66_c7 bl_7 br_7 wl_66 vdd gnd cell_6t
Xbit_r67_c7 bl_7 br_7 wl_67 vdd gnd cell_6t
Xbit_r68_c7 bl_7 br_7 wl_68 vdd gnd cell_6t
Xbit_r69_c7 bl_7 br_7 wl_69 vdd gnd cell_6t
Xbit_r70_c7 bl_7 br_7 wl_70 vdd gnd cell_6t
Xbit_r71_c7 bl_7 br_7 wl_71 vdd gnd cell_6t
Xbit_r72_c7 bl_7 br_7 wl_72 vdd gnd cell_6t
Xbit_r73_c7 bl_7 br_7 wl_73 vdd gnd cell_6t
Xbit_r74_c7 bl_7 br_7 wl_74 vdd gnd cell_6t
Xbit_r75_c7 bl_7 br_7 wl_75 vdd gnd cell_6t
Xbit_r76_c7 bl_7 br_7 wl_76 vdd gnd cell_6t
Xbit_r77_c7 bl_7 br_7 wl_77 vdd gnd cell_6t
Xbit_r78_c7 bl_7 br_7 wl_78 vdd gnd cell_6t
Xbit_r79_c7 bl_7 br_7 wl_79 vdd gnd cell_6t
Xbit_r80_c7 bl_7 br_7 wl_80 vdd gnd cell_6t
Xbit_r81_c7 bl_7 br_7 wl_81 vdd gnd cell_6t
Xbit_r82_c7 bl_7 br_7 wl_82 vdd gnd cell_6t
Xbit_r83_c7 bl_7 br_7 wl_83 vdd gnd cell_6t
Xbit_r84_c7 bl_7 br_7 wl_84 vdd gnd cell_6t
Xbit_r85_c7 bl_7 br_7 wl_85 vdd gnd cell_6t
Xbit_r86_c7 bl_7 br_7 wl_86 vdd gnd cell_6t
Xbit_r87_c7 bl_7 br_7 wl_87 vdd gnd cell_6t
Xbit_r88_c7 bl_7 br_7 wl_88 vdd gnd cell_6t
Xbit_r89_c7 bl_7 br_7 wl_89 vdd gnd cell_6t
Xbit_r90_c7 bl_7 br_7 wl_90 vdd gnd cell_6t
Xbit_r91_c7 bl_7 br_7 wl_91 vdd gnd cell_6t
Xbit_r92_c7 bl_7 br_7 wl_92 vdd gnd cell_6t
Xbit_r93_c7 bl_7 br_7 wl_93 vdd gnd cell_6t
Xbit_r94_c7 bl_7 br_7 wl_94 vdd gnd cell_6t
Xbit_r95_c7 bl_7 br_7 wl_95 vdd gnd cell_6t
Xbit_r96_c7 bl_7 br_7 wl_96 vdd gnd cell_6t
Xbit_r97_c7 bl_7 br_7 wl_97 vdd gnd cell_6t
Xbit_r98_c7 bl_7 br_7 wl_98 vdd gnd cell_6t
Xbit_r99_c7 bl_7 br_7 wl_99 vdd gnd cell_6t
Xbit_r100_c7 bl_7 br_7 wl_100 vdd gnd cell_6t
Xbit_r101_c7 bl_7 br_7 wl_101 vdd gnd cell_6t
Xbit_r102_c7 bl_7 br_7 wl_102 vdd gnd cell_6t
Xbit_r103_c7 bl_7 br_7 wl_103 vdd gnd cell_6t
Xbit_r104_c7 bl_7 br_7 wl_104 vdd gnd cell_6t
Xbit_r105_c7 bl_7 br_7 wl_105 vdd gnd cell_6t
Xbit_r106_c7 bl_7 br_7 wl_106 vdd gnd cell_6t
Xbit_r107_c7 bl_7 br_7 wl_107 vdd gnd cell_6t
Xbit_r108_c7 bl_7 br_7 wl_108 vdd gnd cell_6t
Xbit_r109_c7 bl_7 br_7 wl_109 vdd gnd cell_6t
Xbit_r110_c7 bl_7 br_7 wl_110 vdd gnd cell_6t
Xbit_r111_c7 bl_7 br_7 wl_111 vdd gnd cell_6t
Xbit_r112_c7 bl_7 br_7 wl_112 vdd gnd cell_6t
Xbit_r113_c7 bl_7 br_7 wl_113 vdd gnd cell_6t
Xbit_r114_c7 bl_7 br_7 wl_114 vdd gnd cell_6t
Xbit_r115_c7 bl_7 br_7 wl_115 vdd gnd cell_6t
Xbit_r116_c7 bl_7 br_7 wl_116 vdd gnd cell_6t
Xbit_r117_c7 bl_7 br_7 wl_117 vdd gnd cell_6t
Xbit_r118_c7 bl_7 br_7 wl_118 vdd gnd cell_6t
Xbit_r119_c7 bl_7 br_7 wl_119 vdd gnd cell_6t
Xbit_r120_c7 bl_7 br_7 wl_120 vdd gnd cell_6t
Xbit_r121_c7 bl_7 br_7 wl_121 vdd gnd cell_6t
Xbit_r122_c7 bl_7 br_7 wl_122 vdd gnd cell_6t
Xbit_r123_c7 bl_7 br_7 wl_123 vdd gnd cell_6t
Xbit_r124_c7 bl_7 br_7 wl_124 vdd gnd cell_6t
Xbit_r125_c7 bl_7 br_7 wl_125 vdd gnd cell_6t
Xbit_r126_c7 bl_7 br_7 wl_126 vdd gnd cell_6t
Xbit_r127_c7 bl_7 br_7 wl_127 vdd gnd cell_6t
Xbit_r128_c7 bl_7 br_7 wl_128 vdd gnd cell_6t
Xbit_r129_c7 bl_7 br_7 wl_129 vdd gnd cell_6t
Xbit_r130_c7 bl_7 br_7 wl_130 vdd gnd cell_6t
Xbit_r131_c7 bl_7 br_7 wl_131 vdd gnd cell_6t
Xbit_r132_c7 bl_7 br_7 wl_132 vdd gnd cell_6t
Xbit_r133_c7 bl_7 br_7 wl_133 vdd gnd cell_6t
Xbit_r134_c7 bl_7 br_7 wl_134 vdd gnd cell_6t
Xbit_r135_c7 bl_7 br_7 wl_135 vdd gnd cell_6t
Xbit_r136_c7 bl_7 br_7 wl_136 vdd gnd cell_6t
Xbit_r137_c7 bl_7 br_7 wl_137 vdd gnd cell_6t
Xbit_r138_c7 bl_7 br_7 wl_138 vdd gnd cell_6t
Xbit_r139_c7 bl_7 br_7 wl_139 vdd gnd cell_6t
Xbit_r140_c7 bl_7 br_7 wl_140 vdd gnd cell_6t
Xbit_r141_c7 bl_7 br_7 wl_141 vdd gnd cell_6t
Xbit_r142_c7 bl_7 br_7 wl_142 vdd gnd cell_6t
Xbit_r143_c7 bl_7 br_7 wl_143 vdd gnd cell_6t
Xbit_r144_c7 bl_7 br_7 wl_144 vdd gnd cell_6t
Xbit_r145_c7 bl_7 br_7 wl_145 vdd gnd cell_6t
Xbit_r146_c7 bl_7 br_7 wl_146 vdd gnd cell_6t
Xbit_r147_c7 bl_7 br_7 wl_147 vdd gnd cell_6t
Xbit_r148_c7 bl_7 br_7 wl_148 vdd gnd cell_6t
Xbit_r149_c7 bl_7 br_7 wl_149 vdd gnd cell_6t
Xbit_r150_c7 bl_7 br_7 wl_150 vdd gnd cell_6t
Xbit_r151_c7 bl_7 br_7 wl_151 vdd gnd cell_6t
Xbit_r152_c7 bl_7 br_7 wl_152 vdd gnd cell_6t
Xbit_r153_c7 bl_7 br_7 wl_153 vdd gnd cell_6t
Xbit_r154_c7 bl_7 br_7 wl_154 vdd gnd cell_6t
Xbit_r155_c7 bl_7 br_7 wl_155 vdd gnd cell_6t
Xbit_r156_c7 bl_7 br_7 wl_156 vdd gnd cell_6t
Xbit_r157_c7 bl_7 br_7 wl_157 vdd gnd cell_6t
Xbit_r158_c7 bl_7 br_7 wl_158 vdd gnd cell_6t
Xbit_r159_c7 bl_7 br_7 wl_159 vdd gnd cell_6t
Xbit_r160_c7 bl_7 br_7 wl_160 vdd gnd cell_6t
Xbit_r161_c7 bl_7 br_7 wl_161 vdd gnd cell_6t
Xbit_r162_c7 bl_7 br_7 wl_162 vdd gnd cell_6t
Xbit_r163_c7 bl_7 br_7 wl_163 vdd gnd cell_6t
Xbit_r164_c7 bl_7 br_7 wl_164 vdd gnd cell_6t
Xbit_r165_c7 bl_7 br_7 wl_165 vdd gnd cell_6t
Xbit_r166_c7 bl_7 br_7 wl_166 vdd gnd cell_6t
Xbit_r167_c7 bl_7 br_7 wl_167 vdd gnd cell_6t
Xbit_r168_c7 bl_7 br_7 wl_168 vdd gnd cell_6t
Xbit_r169_c7 bl_7 br_7 wl_169 vdd gnd cell_6t
Xbit_r170_c7 bl_7 br_7 wl_170 vdd gnd cell_6t
Xbit_r171_c7 bl_7 br_7 wl_171 vdd gnd cell_6t
Xbit_r172_c7 bl_7 br_7 wl_172 vdd gnd cell_6t
Xbit_r173_c7 bl_7 br_7 wl_173 vdd gnd cell_6t
Xbit_r174_c7 bl_7 br_7 wl_174 vdd gnd cell_6t
Xbit_r175_c7 bl_7 br_7 wl_175 vdd gnd cell_6t
Xbit_r176_c7 bl_7 br_7 wl_176 vdd gnd cell_6t
Xbit_r177_c7 bl_7 br_7 wl_177 vdd gnd cell_6t
Xbit_r178_c7 bl_7 br_7 wl_178 vdd gnd cell_6t
Xbit_r179_c7 bl_7 br_7 wl_179 vdd gnd cell_6t
Xbit_r180_c7 bl_7 br_7 wl_180 vdd gnd cell_6t
Xbit_r181_c7 bl_7 br_7 wl_181 vdd gnd cell_6t
Xbit_r182_c7 bl_7 br_7 wl_182 vdd gnd cell_6t
Xbit_r183_c7 bl_7 br_7 wl_183 vdd gnd cell_6t
Xbit_r184_c7 bl_7 br_7 wl_184 vdd gnd cell_6t
Xbit_r185_c7 bl_7 br_7 wl_185 vdd gnd cell_6t
Xbit_r186_c7 bl_7 br_7 wl_186 vdd gnd cell_6t
Xbit_r187_c7 bl_7 br_7 wl_187 vdd gnd cell_6t
Xbit_r188_c7 bl_7 br_7 wl_188 vdd gnd cell_6t
Xbit_r189_c7 bl_7 br_7 wl_189 vdd gnd cell_6t
Xbit_r190_c7 bl_7 br_7 wl_190 vdd gnd cell_6t
Xbit_r191_c7 bl_7 br_7 wl_191 vdd gnd cell_6t
Xbit_r192_c7 bl_7 br_7 wl_192 vdd gnd cell_6t
Xbit_r193_c7 bl_7 br_7 wl_193 vdd gnd cell_6t
Xbit_r194_c7 bl_7 br_7 wl_194 vdd gnd cell_6t
Xbit_r195_c7 bl_7 br_7 wl_195 vdd gnd cell_6t
Xbit_r196_c7 bl_7 br_7 wl_196 vdd gnd cell_6t
Xbit_r197_c7 bl_7 br_7 wl_197 vdd gnd cell_6t
Xbit_r198_c7 bl_7 br_7 wl_198 vdd gnd cell_6t
Xbit_r199_c7 bl_7 br_7 wl_199 vdd gnd cell_6t
Xbit_r200_c7 bl_7 br_7 wl_200 vdd gnd cell_6t
Xbit_r201_c7 bl_7 br_7 wl_201 vdd gnd cell_6t
Xbit_r202_c7 bl_7 br_7 wl_202 vdd gnd cell_6t
Xbit_r203_c7 bl_7 br_7 wl_203 vdd gnd cell_6t
Xbit_r204_c7 bl_7 br_7 wl_204 vdd gnd cell_6t
Xbit_r205_c7 bl_7 br_7 wl_205 vdd gnd cell_6t
Xbit_r206_c7 bl_7 br_7 wl_206 vdd gnd cell_6t
Xbit_r207_c7 bl_7 br_7 wl_207 vdd gnd cell_6t
Xbit_r208_c7 bl_7 br_7 wl_208 vdd gnd cell_6t
Xbit_r209_c7 bl_7 br_7 wl_209 vdd gnd cell_6t
Xbit_r210_c7 bl_7 br_7 wl_210 vdd gnd cell_6t
Xbit_r211_c7 bl_7 br_7 wl_211 vdd gnd cell_6t
Xbit_r212_c7 bl_7 br_7 wl_212 vdd gnd cell_6t
Xbit_r213_c7 bl_7 br_7 wl_213 vdd gnd cell_6t
Xbit_r214_c7 bl_7 br_7 wl_214 vdd gnd cell_6t
Xbit_r215_c7 bl_7 br_7 wl_215 vdd gnd cell_6t
Xbit_r216_c7 bl_7 br_7 wl_216 vdd gnd cell_6t
Xbit_r217_c7 bl_7 br_7 wl_217 vdd gnd cell_6t
Xbit_r218_c7 bl_7 br_7 wl_218 vdd gnd cell_6t
Xbit_r219_c7 bl_7 br_7 wl_219 vdd gnd cell_6t
Xbit_r220_c7 bl_7 br_7 wl_220 vdd gnd cell_6t
Xbit_r221_c7 bl_7 br_7 wl_221 vdd gnd cell_6t
Xbit_r222_c7 bl_7 br_7 wl_222 vdd gnd cell_6t
Xbit_r223_c7 bl_7 br_7 wl_223 vdd gnd cell_6t
Xbit_r224_c7 bl_7 br_7 wl_224 vdd gnd cell_6t
Xbit_r225_c7 bl_7 br_7 wl_225 vdd gnd cell_6t
Xbit_r226_c7 bl_7 br_7 wl_226 vdd gnd cell_6t
Xbit_r227_c7 bl_7 br_7 wl_227 vdd gnd cell_6t
Xbit_r228_c7 bl_7 br_7 wl_228 vdd gnd cell_6t
Xbit_r229_c7 bl_7 br_7 wl_229 vdd gnd cell_6t
Xbit_r230_c7 bl_7 br_7 wl_230 vdd gnd cell_6t
Xbit_r231_c7 bl_7 br_7 wl_231 vdd gnd cell_6t
Xbit_r232_c7 bl_7 br_7 wl_232 vdd gnd cell_6t
Xbit_r233_c7 bl_7 br_7 wl_233 vdd gnd cell_6t
Xbit_r234_c7 bl_7 br_7 wl_234 vdd gnd cell_6t
Xbit_r235_c7 bl_7 br_7 wl_235 vdd gnd cell_6t
Xbit_r236_c7 bl_7 br_7 wl_236 vdd gnd cell_6t
Xbit_r237_c7 bl_7 br_7 wl_237 vdd gnd cell_6t
Xbit_r238_c7 bl_7 br_7 wl_238 vdd gnd cell_6t
Xbit_r239_c7 bl_7 br_7 wl_239 vdd gnd cell_6t
Xbit_r240_c7 bl_7 br_7 wl_240 vdd gnd cell_6t
Xbit_r241_c7 bl_7 br_7 wl_241 vdd gnd cell_6t
Xbit_r242_c7 bl_7 br_7 wl_242 vdd gnd cell_6t
Xbit_r243_c7 bl_7 br_7 wl_243 vdd gnd cell_6t
Xbit_r244_c7 bl_7 br_7 wl_244 vdd gnd cell_6t
Xbit_r245_c7 bl_7 br_7 wl_245 vdd gnd cell_6t
Xbit_r246_c7 bl_7 br_7 wl_246 vdd gnd cell_6t
Xbit_r247_c7 bl_7 br_7 wl_247 vdd gnd cell_6t
Xbit_r248_c7 bl_7 br_7 wl_248 vdd gnd cell_6t
Xbit_r249_c7 bl_7 br_7 wl_249 vdd gnd cell_6t
Xbit_r250_c7 bl_7 br_7 wl_250 vdd gnd cell_6t
Xbit_r251_c7 bl_7 br_7 wl_251 vdd gnd cell_6t
Xbit_r252_c7 bl_7 br_7 wl_252 vdd gnd cell_6t
Xbit_r253_c7 bl_7 br_7 wl_253 vdd gnd cell_6t
Xbit_r254_c7 bl_7 br_7 wl_254 vdd gnd cell_6t
Xbit_r255_c7 bl_7 br_7 wl_255 vdd gnd cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd cell_6t
Xbit_r1_c8 bl_8 br_8 wl_1 vdd gnd cell_6t
Xbit_r2_c8 bl_8 br_8 wl_2 vdd gnd cell_6t
Xbit_r3_c8 bl_8 br_8 wl_3 vdd gnd cell_6t
Xbit_r4_c8 bl_8 br_8 wl_4 vdd gnd cell_6t
Xbit_r5_c8 bl_8 br_8 wl_5 vdd gnd cell_6t
Xbit_r6_c8 bl_8 br_8 wl_6 vdd gnd cell_6t
Xbit_r7_c8 bl_8 br_8 wl_7 vdd gnd cell_6t
Xbit_r8_c8 bl_8 br_8 wl_8 vdd gnd cell_6t
Xbit_r9_c8 bl_8 br_8 wl_9 vdd gnd cell_6t
Xbit_r10_c8 bl_8 br_8 wl_10 vdd gnd cell_6t
Xbit_r11_c8 bl_8 br_8 wl_11 vdd gnd cell_6t
Xbit_r12_c8 bl_8 br_8 wl_12 vdd gnd cell_6t
Xbit_r13_c8 bl_8 br_8 wl_13 vdd gnd cell_6t
Xbit_r14_c8 bl_8 br_8 wl_14 vdd gnd cell_6t
Xbit_r15_c8 bl_8 br_8 wl_15 vdd gnd cell_6t
Xbit_r16_c8 bl_8 br_8 wl_16 vdd gnd cell_6t
Xbit_r17_c8 bl_8 br_8 wl_17 vdd gnd cell_6t
Xbit_r18_c8 bl_8 br_8 wl_18 vdd gnd cell_6t
Xbit_r19_c8 bl_8 br_8 wl_19 vdd gnd cell_6t
Xbit_r20_c8 bl_8 br_8 wl_20 vdd gnd cell_6t
Xbit_r21_c8 bl_8 br_8 wl_21 vdd gnd cell_6t
Xbit_r22_c8 bl_8 br_8 wl_22 vdd gnd cell_6t
Xbit_r23_c8 bl_8 br_8 wl_23 vdd gnd cell_6t
Xbit_r24_c8 bl_8 br_8 wl_24 vdd gnd cell_6t
Xbit_r25_c8 bl_8 br_8 wl_25 vdd gnd cell_6t
Xbit_r26_c8 bl_8 br_8 wl_26 vdd gnd cell_6t
Xbit_r27_c8 bl_8 br_8 wl_27 vdd gnd cell_6t
Xbit_r28_c8 bl_8 br_8 wl_28 vdd gnd cell_6t
Xbit_r29_c8 bl_8 br_8 wl_29 vdd gnd cell_6t
Xbit_r30_c8 bl_8 br_8 wl_30 vdd gnd cell_6t
Xbit_r31_c8 bl_8 br_8 wl_31 vdd gnd cell_6t
Xbit_r32_c8 bl_8 br_8 wl_32 vdd gnd cell_6t
Xbit_r33_c8 bl_8 br_8 wl_33 vdd gnd cell_6t
Xbit_r34_c8 bl_8 br_8 wl_34 vdd gnd cell_6t
Xbit_r35_c8 bl_8 br_8 wl_35 vdd gnd cell_6t
Xbit_r36_c8 bl_8 br_8 wl_36 vdd gnd cell_6t
Xbit_r37_c8 bl_8 br_8 wl_37 vdd gnd cell_6t
Xbit_r38_c8 bl_8 br_8 wl_38 vdd gnd cell_6t
Xbit_r39_c8 bl_8 br_8 wl_39 vdd gnd cell_6t
Xbit_r40_c8 bl_8 br_8 wl_40 vdd gnd cell_6t
Xbit_r41_c8 bl_8 br_8 wl_41 vdd gnd cell_6t
Xbit_r42_c8 bl_8 br_8 wl_42 vdd gnd cell_6t
Xbit_r43_c8 bl_8 br_8 wl_43 vdd gnd cell_6t
Xbit_r44_c8 bl_8 br_8 wl_44 vdd gnd cell_6t
Xbit_r45_c8 bl_8 br_8 wl_45 vdd gnd cell_6t
Xbit_r46_c8 bl_8 br_8 wl_46 vdd gnd cell_6t
Xbit_r47_c8 bl_8 br_8 wl_47 vdd gnd cell_6t
Xbit_r48_c8 bl_8 br_8 wl_48 vdd gnd cell_6t
Xbit_r49_c8 bl_8 br_8 wl_49 vdd gnd cell_6t
Xbit_r50_c8 bl_8 br_8 wl_50 vdd gnd cell_6t
Xbit_r51_c8 bl_8 br_8 wl_51 vdd gnd cell_6t
Xbit_r52_c8 bl_8 br_8 wl_52 vdd gnd cell_6t
Xbit_r53_c8 bl_8 br_8 wl_53 vdd gnd cell_6t
Xbit_r54_c8 bl_8 br_8 wl_54 vdd gnd cell_6t
Xbit_r55_c8 bl_8 br_8 wl_55 vdd gnd cell_6t
Xbit_r56_c8 bl_8 br_8 wl_56 vdd gnd cell_6t
Xbit_r57_c8 bl_8 br_8 wl_57 vdd gnd cell_6t
Xbit_r58_c8 bl_8 br_8 wl_58 vdd gnd cell_6t
Xbit_r59_c8 bl_8 br_8 wl_59 vdd gnd cell_6t
Xbit_r60_c8 bl_8 br_8 wl_60 vdd gnd cell_6t
Xbit_r61_c8 bl_8 br_8 wl_61 vdd gnd cell_6t
Xbit_r62_c8 bl_8 br_8 wl_62 vdd gnd cell_6t
Xbit_r63_c8 bl_8 br_8 wl_63 vdd gnd cell_6t
Xbit_r64_c8 bl_8 br_8 wl_64 vdd gnd cell_6t
Xbit_r65_c8 bl_8 br_8 wl_65 vdd gnd cell_6t
Xbit_r66_c8 bl_8 br_8 wl_66 vdd gnd cell_6t
Xbit_r67_c8 bl_8 br_8 wl_67 vdd gnd cell_6t
Xbit_r68_c8 bl_8 br_8 wl_68 vdd gnd cell_6t
Xbit_r69_c8 bl_8 br_8 wl_69 vdd gnd cell_6t
Xbit_r70_c8 bl_8 br_8 wl_70 vdd gnd cell_6t
Xbit_r71_c8 bl_8 br_8 wl_71 vdd gnd cell_6t
Xbit_r72_c8 bl_8 br_8 wl_72 vdd gnd cell_6t
Xbit_r73_c8 bl_8 br_8 wl_73 vdd gnd cell_6t
Xbit_r74_c8 bl_8 br_8 wl_74 vdd gnd cell_6t
Xbit_r75_c8 bl_8 br_8 wl_75 vdd gnd cell_6t
Xbit_r76_c8 bl_8 br_8 wl_76 vdd gnd cell_6t
Xbit_r77_c8 bl_8 br_8 wl_77 vdd gnd cell_6t
Xbit_r78_c8 bl_8 br_8 wl_78 vdd gnd cell_6t
Xbit_r79_c8 bl_8 br_8 wl_79 vdd gnd cell_6t
Xbit_r80_c8 bl_8 br_8 wl_80 vdd gnd cell_6t
Xbit_r81_c8 bl_8 br_8 wl_81 vdd gnd cell_6t
Xbit_r82_c8 bl_8 br_8 wl_82 vdd gnd cell_6t
Xbit_r83_c8 bl_8 br_8 wl_83 vdd gnd cell_6t
Xbit_r84_c8 bl_8 br_8 wl_84 vdd gnd cell_6t
Xbit_r85_c8 bl_8 br_8 wl_85 vdd gnd cell_6t
Xbit_r86_c8 bl_8 br_8 wl_86 vdd gnd cell_6t
Xbit_r87_c8 bl_8 br_8 wl_87 vdd gnd cell_6t
Xbit_r88_c8 bl_8 br_8 wl_88 vdd gnd cell_6t
Xbit_r89_c8 bl_8 br_8 wl_89 vdd gnd cell_6t
Xbit_r90_c8 bl_8 br_8 wl_90 vdd gnd cell_6t
Xbit_r91_c8 bl_8 br_8 wl_91 vdd gnd cell_6t
Xbit_r92_c8 bl_8 br_8 wl_92 vdd gnd cell_6t
Xbit_r93_c8 bl_8 br_8 wl_93 vdd gnd cell_6t
Xbit_r94_c8 bl_8 br_8 wl_94 vdd gnd cell_6t
Xbit_r95_c8 bl_8 br_8 wl_95 vdd gnd cell_6t
Xbit_r96_c8 bl_8 br_8 wl_96 vdd gnd cell_6t
Xbit_r97_c8 bl_8 br_8 wl_97 vdd gnd cell_6t
Xbit_r98_c8 bl_8 br_8 wl_98 vdd gnd cell_6t
Xbit_r99_c8 bl_8 br_8 wl_99 vdd gnd cell_6t
Xbit_r100_c8 bl_8 br_8 wl_100 vdd gnd cell_6t
Xbit_r101_c8 bl_8 br_8 wl_101 vdd gnd cell_6t
Xbit_r102_c8 bl_8 br_8 wl_102 vdd gnd cell_6t
Xbit_r103_c8 bl_8 br_8 wl_103 vdd gnd cell_6t
Xbit_r104_c8 bl_8 br_8 wl_104 vdd gnd cell_6t
Xbit_r105_c8 bl_8 br_8 wl_105 vdd gnd cell_6t
Xbit_r106_c8 bl_8 br_8 wl_106 vdd gnd cell_6t
Xbit_r107_c8 bl_8 br_8 wl_107 vdd gnd cell_6t
Xbit_r108_c8 bl_8 br_8 wl_108 vdd gnd cell_6t
Xbit_r109_c8 bl_8 br_8 wl_109 vdd gnd cell_6t
Xbit_r110_c8 bl_8 br_8 wl_110 vdd gnd cell_6t
Xbit_r111_c8 bl_8 br_8 wl_111 vdd gnd cell_6t
Xbit_r112_c8 bl_8 br_8 wl_112 vdd gnd cell_6t
Xbit_r113_c8 bl_8 br_8 wl_113 vdd gnd cell_6t
Xbit_r114_c8 bl_8 br_8 wl_114 vdd gnd cell_6t
Xbit_r115_c8 bl_8 br_8 wl_115 vdd gnd cell_6t
Xbit_r116_c8 bl_8 br_8 wl_116 vdd gnd cell_6t
Xbit_r117_c8 bl_8 br_8 wl_117 vdd gnd cell_6t
Xbit_r118_c8 bl_8 br_8 wl_118 vdd gnd cell_6t
Xbit_r119_c8 bl_8 br_8 wl_119 vdd gnd cell_6t
Xbit_r120_c8 bl_8 br_8 wl_120 vdd gnd cell_6t
Xbit_r121_c8 bl_8 br_8 wl_121 vdd gnd cell_6t
Xbit_r122_c8 bl_8 br_8 wl_122 vdd gnd cell_6t
Xbit_r123_c8 bl_8 br_8 wl_123 vdd gnd cell_6t
Xbit_r124_c8 bl_8 br_8 wl_124 vdd gnd cell_6t
Xbit_r125_c8 bl_8 br_8 wl_125 vdd gnd cell_6t
Xbit_r126_c8 bl_8 br_8 wl_126 vdd gnd cell_6t
Xbit_r127_c8 bl_8 br_8 wl_127 vdd gnd cell_6t
Xbit_r128_c8 bl_8 br_8 wl_128 vdd gnd cell_6t
Xbit_r129_c8 bl_8 br_8 wl_129 vdd gnd cell_6t
Xbit_r130_c8 bl_8 br_8 wl_130 vdd gnd cell_6t
Xbit_r131_c8 bl_8 br_8 wl_131 vdd gnd cell_6t
Xbit_r132_c8 bl_8 br_8 wl_132 vdd gnd cell_6t
Xbit_r133_c8 bl_8 br_8 wl_133 vdd gnd cell_6t
Xbit_r134_c8 bl_8 br_8 wl_134 vdd gnd cell_6t
Xbit_r135_c8 bl_8 br_8 wl_135 vdd gnd cell_6t
Xbit_r136_c8 bl_8 br_8 wl_136 vdd gnd cell_6t
Xbit_r137_c8 bl_8 br_8 wl_137 vdd gnd cell_6t
Xbit_r138_c8 bl_8 br_8 wl_138 vdd gnd cell_6t
Xbit_r139_c8 bl_8 br_8 wl_139 vdd gnd cell_6t
Xbit_r140_c8 bl_8 br_8 wl_140 vdd gnd cell_6t
Xbit_r141_c8 bl_8 br_8 wl_141 vdd gnd cell_6t
Xbit_r142_c8 bl_8 br_8 wl_142 vdd gnd cell_6t
Xbit_r143_c8 bl_8 br_8 wl_143 vdd gnd cell_6t
Xbit_r144_c8 bl_8 br_8 wl_144 vdd gnd cell_6t
Xbit_r145_c8 bl_8 br_8 wl_145 vdd gnd cell_6t
Xbit_r146_c8 bl_8 br_8 wl_146 vdd gnd cell_6t
Xbit_r147_c8 bl_8 br_8 wl_147 vdd gnd cell_6t
Xbit_r148_c8 bl_8 br_8 wl_148 vdd gnd cell_6t
Xbit_r149_c8 bl_8 br_8 wl_149 vdd gnd cell_6t
Xbit_r150_c8 bl_8 br_8 wl_150 vdd gnd cell_6t
Xbit_r151_c8 bl_8 br_8 wl_151 vdd gnd cell_6t
Xbit_r152_c8 bl_8 br_8 wl_152 vdd gnd cell_6t
Xbit_r153_c8 bl_8 br_8 wl_153 vdd gnd cell_6t
Xbit_r154_c8 bl_8 br_8 wl_154 vdd gnd cell_6t
Xbit_r155_c8 bl_8 br_8 wl_155 vdd gnd cell_6t
Xbit_r156_c8 bl_8 br_8 wl_156 vdd gnd cell_6t
Xbit_r157_c8 bl_8 br_8 wl_157 vdd gnd cell_6t
Xbit_r158_c8 bl_8 br_8 wl_158 vdd gnd cell_6t
Xbit_r159_c8 bl_8 br_8 wl_159 vdd gnd cell_6t
Xbit_r160_c8 bl_8 br_8 wl_160 vdd gnd cell_6t
Xbit_r161_c8 bl_8 br_8 wl_161 vdd gnd cell_6t
Xbit_r162_c8 bl_8 br_8 wl_162 vdd gnd cell_6t
Xbit_r163_c8 bl_8 br_8 wl_163 vdd gnd cell_6t
Xbit_r164_c8 bl_8 br_8 wl_164 vdd gnd cell_6t
Xbit_r165_c8 bl_8 br_8 wl_165 vdd gnd cell_6t
Xbit_r166_c8 bl_8 br_8 wl_166 vdd gnd cell_6t
Xbit_r167_c8 bl_8 br_8 wl_167 vdd gnd cell_6t
Xbit_r168_c8 bl_8 br_8 wl_168 vdd gnd cell_6t
Xbit_r169_c8 bl_8 br_8 wl_169 vdd gnd cell_6t
Xbit_r170_c8 bl_8 br_8 wl_170 vdd gnd cell_6t
Xbit_r171_c8 bl_8 br_8 wl_171 vdd gnd cell_6t
Xbit_r172_c8 bl_8 br_8 wl_172 vdd gnd cell_6t
Xbit_r173_c8 bl_8 br_8 wl_173 vdd gnd cell_6t
Xbit_r174_c8 bl_8 br_8 wl_174 vdd gnd cell_6t
Xbit_r175_c8 bl_8 br_8 wl_175 vdd gnd cell_6t
Xbit_r176_c8 bl_8 br_8 wl_176 vdd gnd cell_6t
Xbit_r177_c8 bl_8 br_8 wl_177 vdd gnd cell_6t
Xbit_r178_c8 bl_8 br_8 wl_178 vdd gnd cell_6t
Xbit_r179_c8 bl_8 br_8 wl_179 vdd gnd cell_6t
Xbit_r180_c8 bl_8 br_8 wl_180 vdd gnd cell_6t
Xbit_r181_c8 bl_8 br_8 wl_181 vdd gnd cell_6t
Xbit_r182_c8 bl_8 br_8 wl_182 vdd gnd cell_6t
Xbit_r183_c8 bl_8 br_8 wl_183 vdd gnd cell_6t
Xbit_r184_c8 bl_8 br_8 wl_184 vdd gnd cell_6t
Xbit_r185_c8 bl_8 br_8 wl_185 vdd gnd cell_6t
Xbit_r186_c8 bl_8 br_8 wl_186 vdd gnd cell_6t
Xbit_r187_c8 bl_8 br_8 wl_187 vdd gnd cell_6t
Xbit_r188_c8 bl_8 br_8 wl_188 vdd gnd cell_6t
Xbit_r189_c8 bl_8 br_8 wl_189 vdd gnd cell_6t
Xbit_r190_c8 bl_8 br_8 wl_190 vdd gnd cell_6t
Xbit_r191_c8 bl_8 br_8 wl_191 vdd gnd cell_6t
Xbit_r192_c8 bl_8 br_8 wl_192 vdd gnd cell_6t
Xbit_r193_c8 bl_8 br_8 wl_193 vdd gnd cell_6t
Xbit_r194_c8 bl_8 br_8 wl_194 vdd gnd cell_6t
Xbit_r195_c8 bl_8 br_8 wl_195 vdd gnd cell_6t
Xbit_r196_c8 bl_8 br_8 wl_196 vdd gnd cell_6t
Xbit_r197_c8 bl_8 br_8 wl_197 vdd gnd cell_6t
Xbit_r198_c8 bl_8 br_8 wl_198 vdd gnd cell_6t
Xbit_r199_c8 bl_8 br_8 wl_199 vdd gnd cell_6t
Xbit_r200_c8 bl_8 br_8 wl_200 vdd gnd cell_6t
Xbit_r201_c8 bl_8 br_8 wl_201 vdd gnd cell_6t
Xbit_r202_c8 bl_8 br_8 wl_202 vdd gnd cell_6t
Xbit_r203_c8 bl_8 br_8 wl_203 vdd gnd cell_6t
Xbit_r204_c8 bl_8 br_8 wl_204 vdd gnd cell_6t
Xbit_r205_c8 bl_8 br_8 wl_205 vdd gnd cell_6t
Xbit_r206_c8 bl_8 br_8 wl_206 vdd gnd cell_6t
Xbit_r207_c8 bl_8 br_8 wl_207 vdd gnd cell_6t
Xbit_r208_c8 bl_8 br_8 wl_208 vdd gnd cell_6t
Xbit_r209_c8 bl_8 br_8 wl_209 vdd gnd cell_6t
Xbit_r210_c8 bl_8 br_8 wl_210 vdd gnd cell_6t
Xbit_r211_c8 bl_8 br_8 wl_211 vdd gnd cell_6t
Xbit_r212_c8 bl_8 br_8 wl_212 vdd gnd cell_6t
Xbit_r213_c8 bl_8 br_8 wl_213 vdd gnd cell_6t
Xbit_r214_c8 bl_8 br_8 wl_214 vdd gnd cell_6t
Xbit_r215_c8 bl_8 br_8 wl_215 vdd gnd cell_6t
Xbit_r216_c8 bl_8 br_8 wl_216 vdd gnd cell_6t
Xbit_r217_c8 bl_8 br_8 wl_217 vdd gnd cell_6t
Xbit_r218_c8 bl_8 br_8 wl_218 vdd gnd cell_6t
Xbit_r219_c8 bl_8 br_8 wl_219 vdd gnd cell_6t
Xbit_r220_c8 bl_8 br_8 wl_220 vdd gnd cell_6t
Xbit_r221_c8 bl_8 br_8 wl_221 vdd gnd cell_6t
Xbit_r222_c8 bl_8 br_8 wl_222 vdd gnd cell_6t
Xbit_r223_c8 bl_8 br_8 wl_223 vdd gnd cell_6t
Xbit_r224_c8 bl_8 br_8 wl_224 vdd gnd cell_6t
Xbit_r225_c8 bl_8 br_8 wl_225 vdd gnd cell_6t
Xbit_r226_c8 bl_8 br_8 wl_226 vdd gnd cell_6t
Xbit_r227_c8 bl_8 br_8 wl_227 vdd gnd cell_6t
Xbit_r228_c8 bl_8 br_8 wl_228 vdd gnd cell_6t
Xbit_r229_c8 bl_8 br_8 wl_229 vdd gnd cell_6t
Xbit_r230_c8 bl_8 br_8 wl_230 vdd gnd cell_6t
Xbit_r231_c8 bl_8 br_8 wl_231 vdd gnd cell_6t
Xbit_r232_c8 bl_8 br_8 wl_232 vdd gnd cell_6t
Xbit_r233_c8 bl_8 br_8 wl_233 vdd gnd cell_6t
Xbit_r234_c8 bl_8 br_8 wl_234 vdd gnd cell_6t
Xbit_r235_c8 bl_8 br_8 wl_235 vdd gnd cell_6t
Xbit_r236_c8 bl_8 br_8 wl_236 vdd gnd cell_6t
Xbit_r237_c8 bl_8 br_8 wl_237 vdd gnd cell_6t
Xbit_r238_c8 bl_8 br_8 wl_238 vdd gnd cell_6t
Xbit_r239_c8 bl_8 br_8 wl_239 vdd gnd cell_6t
Xbit_r240_c8 bl_8 br_8 wl_240 vdd gnd cell_6t
Xbit_r241_c8 bl_8 br_8 wl_241 vdd gnd cell_6t
Xbit_r242_c8 bl_8 br_8 wl_242 vdd gnd cell_6t
Xbit_r243_c8 bl_8 br_8 wl_243 vdd gnd cell_6t
Xbit_r244_c8 bl_8 br_8 wl_244 vdd gnd cell_6t
Xbit_r245_c8 bl_8 br_8 wl_245 vdd gnd cell_6t
Xbit_r246_c8 bl_8 br_8 wl_246 vdd gnd cell_6t
Xbit_r247_c8 bl_8 br_8 wl_247 vdd gnd cell_6t
Xbit_r248_c8 bl_8 br_8 wl_248 vdd gnd cell_6t
Xbit_r249_c8 bl_8 br_8 wl_249 vdd gnd cell_6t
Xbit_r250_c8 bl_8 br_8 wl_250 vdd gnd cell_6t
Xbit_r251_c8 bl_8 br_8 wl_251 vdd gnd cell_6t
Xbit_r252_c8 bl_8 br_8 wl_252 vdd gnd cell_6t
Xbit_r253_c8 bl_8 br_8 wl_253 vdd gnd cell_6t
Xbit_r254_c8 bl_8 br_8 wl_254 vdd gnd cell_6t
Xbit_r255_c8 bl_8 br_8 wl_255 vdd gnd cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd cell_6t
Xbit_r1_c9 bl_9 br_9 wl_1 vdd gnd cell_6t
Xbit_r2_c9 bl_9 br_9 wl_2 vdd gnd cell_6t
Xbit_r3_c9 bl_9 br_9 wl_3 vdd gnd cell_6t
Xbit_r4_c9 bl_9 br_9 wl_4 vdd gnd cell_6t
Xbit_r5_c9 bl_9 br_9 wl_5 vdd gnd cell_6t
Xbit_r6_c9 bl_9 br_9 wl_6 vdd gnd cell_6t
Xbit_r7_c9 bl_9 br_9 wl_7 vdd gnd cell_6t
Xbit_r8_c9 bl_9 br_9 wl_8 vdd gnd cell_6t
Xbit_r9_c9 bl_9 br_9 wl_9 vdd gnd cell_6t
Xbit_r10_c9 bl_9 br_9 wl_10 vdd gnd cell_6t
Xbit_r11_c9 bl_9 br_9 wl_11 vdd gnd cell_6t
Xbit_r12_c9 bl_9 br_9 wl_12 vdd gnd cell_6t
Xbit_r13_c9 bl_9 br_9 wl_13 vdd gnd cell_6t
Xbit_r14_c9 bl_9 br_9 wl_14 vdd gnd cell_6t
Xbit_r15_c9 bl_9 br_9 wl_15 vdd gnd cell_6t
Xbit_r16_c9 bl_9 br_9 wl_16 vdd gnd cell_6t
Xbit_r17_c9 bl_9 br_9 wl_17 vdd gnd cell_6t
Xbit_r18_c9 bl_9 br_9 wl_18 vdd gnd cell_6t
Xbit_r19_c9 bl_9 br_9 wl_19 vdd gnd cell_6t
Xbit_r20_c9 bl_9 br_9 wl_20 vdd gnd cell_6t
Xbit_r21_c9 bl_9 br_9 wl_21 vdd gnd cell_6t
Xbit_r22_c9 bl_9 br_9 wl_22 vdd gnd cell_6t
Xbit_r23_c9 bl_9 br_9 wl_23 vdd gnd cell_6t
Xbit_r24_c9 bl_9 br_9 wl_24 vdd gnd cell_6t
Xbit_r25_c9 bl_9 br_9 wl_25 vdd gnd cell_6t
Xbit_r26_c9 bl_9 br_9 wl_26 vdd gnd cell_6t
Xbit_r27_c9 bl_9 br_9 wl_27 vdd gnd cell_6t
Xbit_r28_c9 bl_9 br_9 wl_28 vdd gnd cell_6t
Xbit_r29_c9 bl_9 br_9 wl_29 vdd gnd cell_6t
Xbit_r30_c9 bl_9 br_9 wl_30 vdd gnd cell_6t
Xbit_r31_c9 bl_9 br_9 wl_31 vdd gnd cell_6t
Xbit_r32_c9 bl_9 br_9 wl_32 vdd gnd cell_6t
Xbit_r33_c9 bl_9 br_9 wl_33 vdd gnd cell_6t
Xbit_r34_c9 bl_9 br_9 wl_34 vdd gnd cell_6t
Xbit_r35_c9 bl_9 br_9 wl_35 vdd gnd cell_6t
Xbit_r36_c9 bl_9 br_9 wl_36 vdd gnd cell_6t
Xbit_r37_c9 bl_9 br_9 wl_37 vdd gnd cell_6t
Xbit_r38_c9 bl_9 br_9 wl_38 vdd gnd cell_6t
Xbit_r39_c9 bl_9 br_9 wl_39 vdd gnd cell_6t
Xbit_r40_c9 bl_9 br_9 wl_40 vdd gnd cell_6t
Xbit_r41_c9 bl_9 br_9 wl_41 vdd gnd cell_6t
Xbit_r42_c9 bl_9 br_9 wl_42 vdd gnd cell_6t
Xbit_r43_c9 bl_9 br_9 wl_43 vdd gnd cell_6t
Xbit_r44_c9 bl_9 br_9 wl_44 vdd gnd cell_6t
Xbit_r45_c9 bl_9 br_9 wl_45 vdd gnd cell_6t
Xbit_r46_c9 bl_9 br_9 wl_46 vdd gnd cell_6t
Xbit_r47_c9 bl_9 br_9 wl_47 vdd gnd cell_6t
Xbit_r48_c9 bl_9 br_9 wl_48 vdd gnd cell_6t
Xbit_r49_c9 bl_9 br_9 wl_49 vdd gnd cell_6t
Xbit_r50_c9 bl_9 br_9 wl_50 vdd gnd cell_6t
Xbit_r51_c9 bl_9 br_9 wl_51 vdd gnd cell_6t
Xbit_r52_c9 bl_9 br_9 wl_52 vdd gnd cell_6t
Xbit_r53_c9 bl_9 br_9 wl_53 vdd gnd cell_6t
Xbit_r54_c9 bl_9 br_9 wl_54 vdd gnd cell_6t
Xbit_r55_c9 bl_9 br_9 wl_55 vdd gnd cell_6t
Xbit_r56_c9 bl_9 br_9 wl_56 vdd gnd cell_6t
Xbit_r57_c9 bl_9 br_9 wl_57 vdd gnd cell_6t
Xbit_r58_c9 bl_9 br_9 wl_58 vdd gnd cell_6t
Xbit_r59_c9 bl_9 br_9 wl_59 vdd gnd cell_6t
Xbit_r60_c9 bl_9 br_9 wl_60 vdd gnd cell_6t
Xbit_r61_c9 bl_9 br_9 wl_61 vdd gnd cell_6t
Xbit_r62_c9 bl_9 br_9 wl_62 vdd gnd cell_6t
Xbit_r63_c9 bl_9 br_9 wl_63 vdd gnd cell_6t
Xbit_r64_c9 bl_9 br_9 wl_64 vdd gnd cell_6t
Xbit_r65_c9 bl_9 br_9 wl_65 vdd gnd cell_6t
Xbit_r66_c9 bl_9 br_9 wl_66 vdd gnd cell_6t
Xbit_r67_c9 bl_9 br_9 wl_67 vdd gnd cell_6t
Xbit_r68_c9 bl_9 br_9 wl_68 vdd gnd cell_6t
Xbit_r69_c9 bl_9 br_9 wl_69 vdd gnd cell_6t
Xbit_r70_c9 bl_9 br_9 wl_70 vdd gnd cell_6t
Xbit_r71_c9 bl_9 br_9 wl_71 vdd gnd cell_6t
Xbit_r72_c9 bl_9 br_9 wl_72 vdd gnd cell_6t
Xbit_r73_c9 bl_9 br_9 wl_73 vdd gnd cell_6t
Xbit_r74_c9 bl_9 br_9 wl_74 vdd gnd cell_6t
Xbit_r75_c9 bl_9 br_9 wl_75 vdd gnd cell_6t
Xbit_r76_c9 bl_9 br_9 wl_76 vdd gnd cell_6t
Xbit_r77_c9 bl_9 br_9 wl_77 vdd gnd cell_6t
Xbit_r78_c9 bl_9 br_9 wl_78 vdd gnd cell_6t
Xbit_r79_c9 bl_9 br_9 wl_79 vdd gnd cell_6t
Xbit_r80_c9 bl_9 br_9 wl_80 vdd gnd cell_6t
Xbit_r81_c9 bl_9 br_9 wl_81 vdd gnd cell_6t
Xbit_r82_c9 bl_9 br_9 wl_82 vdd gnd cell_6t
Xbit_r83_c9 bl_9 br_9 wl_83 vdd gnd cell_6t
Xbit_r84_c9 bl_9 br_9 wl_84 vdd gnd cell_6t
Xbit_r85_c9 bl_9 br_9 wl_85 vdd gnd cell_6t
Xbit_r86_c9 bl_9 br_9 wl_86 vdd gnd cell_6t
Xbit_r87_c9 bl_9 br_9 wl_87 vdd gnd cell_6t
Xbit_r88_c9 bl_9 br_9 wl_88 vdd gnd cell_6t
Xbit_r89_c9 bl_9 br_9 wl_89 vdd gnd cell_6t
Xbit_r90_c9 bl_9 br_9 wl_90 vdd gnd cell_6t
Xbit_r91_c9 bl_9 br_9 wl_91 vdd gnd cell_6t
Xbit_r92_c9 bl_9 br_9 wl_92 vdd gnd cell_6t
Xbit_r93_c9 bl_9 br_9 wl_93 vdd gnd cell_6t
Xbit_r94_c9 bl_9 br_9 wl_94 vdd gnd cell_6t
Xbit_r95_c9 bl_9 br_9 wl_95 vdd gnd cell_6t
Xbit_r96_c9 bl_9 br_9 wl_96 vdd gnd cell_6t
Xbit_r97_c9 bl_9 br_9 wl_97 vdd gnd cell_6t
Xbit_r98_c9 bl_9 br_9 wl_98 vdd gnd cell_6t
Xbit_r99_c9 bl_9 br_9 wl_99 vdd gnd cell_6t
Xbit_r100_c9 bl_9 br_9 wl_100 vdd gnd cell_6t
Xbit_r101_c9 bl_9 br_9 wl_101 vdd gnd cell_6t
Xbit_r102_c9 bl_9 br_9 wl_102 vdd gnd cell_6t
Xbit_r103_c9 bl_9 br_9 wl_103 vdd gnd cell_6t
Xbit_r104_c9 bl_9 br_9 wl_104 vdd gnd cell_6t
Xbit_r105_c9 bl_9 br_9 wl_105 vdd gnd cell_6t
Xbit_r106_c9 bl_9 br_9 wl_106 vdd gnd cell_6t
Xbit_r107_c9 bl_9 br_9 wl_107 vdd gnd cell_6t
Xbit_r108_c9 bl_9 br_9 wl_108 vdd gnd cell_6t
Xbit_r109_c9 bl_9 br_9 wl_109 vdd gnd cell_6t
Xbit_r110_c9 bl_9 br_9 wl_110 vdd gnd cell_6t
Xbit_r111_c9 bl_9 br_9 wl_111 vdd gnd cell_6t
Xbit_r112_c9 bl_9 br_9 wl_112 vdd gnd cell_6t
Xbit_r113_c9 bl_9 br_9 wl_113 vdd gnd cell_6t
Xbit_r114_c9 bl_9 br_9 wl_114 vdd gnd cell_6t
Xbit_r115_c9 bl_9 br_9 wl_115 vdd gnd cell_6t
Xbit_r116_c9 bl_9 br_9 wl_116 vdd gnd cell_6t
Xbit_r117_c9 bl_9 br_9 wl_117 vdd gnd cell_6t
Xbit_r118_c9 bl_9 br_9 wl_118 vdd gnd cell_6t
Xbit_r119_c9 bl_9 br_9 wl_119 vdd gnd cell_6t
Xbit_r120_c9 bl_9 br_9 wl_120 vdd gnd cell_6t
Xbit_r121_c9 bl_9 br_9 wl_121 vdd gnd cell_6t
Xbit_r122_c9 bl_9 br_9 wl_122 vdd gnd cell_6t
Xbit_r123_c9 bl_9 br_9 wl_123 vdd gnd cell_6t
Xbit_r124_c9 bl_9 br_9 wl_124 vdd gnd cell_6t
Xbit_r125_c9 bl_9 br_9 wl_125 vdd gnd cell_6t
Xbit_r126_c9 bl_9 br_9 wl_126 vdd gnd cell_6t
Xbit_r127_c9 bl_9 br_9 wl_127 vdd gnd cell_6t
Xbit_r128_c9 bl_9 br_9 wl_128 vdd gnd cell_6t
Xbit_r129_c9 bl_9 br_9 wl_129 vdd gnd cell_6t
Xbit_r130_c9 bl_9 br_9 wl_130 vdd gnd cell_6t
Xbit_r131_c9 bl_9 br_9 wl_131 vdd gnd cell_6t
Xbit_r132_c9 bl_9 br_9 wl_132 vdd gnd cell_6t
Xbit_r133_c9 bl_9 br_9 wl_133 vdd gnd cell_6t
Xbit_r134_c9 bl_9 br_9 wl_134 vdd gnd cell_6t
Xbit_r135_c9 bl_9 br_9 wl_135 vdd gnd cell_6t
Xbit_r136_c9 bl_9 br_9 wl_136 vdd gnd cell_6t
Xbit_r137_c9 bl_9 br_9 wl_137 vdd gnd cell_6t
Xbit_r138_c9 bl_9 br_9 wl_138 vdd gnd cell_6t
Xbit_r139_c9 bl_9 br_9 wl_139 vdd gnd cell_6t
Xbit_r140_c9 bl_9 br_9 wl_140 vdd gnd cell_6t
Xbit_r141_c9 bl_9 br_9 wl_141 vdd gnd cell_6t
Xbit_r142_c9 bl_9 br_9 wl_142 vdd gnd cell_6t
Xbit_r143_c9 bl_9 br_9 wl_143 vdd gnd cell_6t
Xbit_r144_c9 bl_9 br_9 wl_144 vdd gnd cell_6t
Xbit_r145_c9 bl_9 br_9 wl_145 vdd gnd cell_6t
Xbit_r146_c9 bl_9 br_9 wl_146 vdd gnd cell_6t
Xbit_r147_c9 bl_9 br_9 wl_147 vdd gnd cell_6t
Xbit_r148_c9 bl_9 br_9 wl_148 vdd gnd cell_6t
Xbit_r149_c9 bl_9 br_9 wl_149 vdd gnd cell_6t
Xbit_r150_c9 bl_9 br_9 wl_150 vdd gnd cell_6t
Xbit_r151_c9 bl_9 br_9 wl_151 vdd gnd cell_6t
Xbit_r152_c9 bl_9 br_9 wl_152 vdd gnd cell_6t
Xbit_r153_c9 bl_9 br_9 wl_153 vdd gnd cell_6t
Xbit_r154_c9 bl_9 br_9 wl_154 vdd gnd cell_6t
Xbit_r155_c9 bl_9 br_9 wl_155 vdd gnd cell_6t
Xbit_r156_c9 bl_9 br_9 wl_156 vdd gnd cell_6t
Xbit_r157_c9 bl_9 br_9 wl_157 vdd gnd cell_6t
Xbit_r158_c9 bl_9 br_9 wl_158 vdd gnd cell_6t
Xbit_r159_c9 bl_9 br_9 wl_159 vdd gnd cell_6t
Xbit_r160_c9 bl_9 br_9 wl_160 vdd gnd cell_6t
Xbit_r161_c9 bl_9 br_9 wl_161 vdd gnd cell_6t
Xbit_r162_c9 bl_9 br_9 wl_162 vdd gnd cell_6t
Xbit_r163_c9 bl_9 br_9 wl_163 vdd gnd cell_6t
Xbit_r164_c9 bl_9 br_9 wl_164 vdd gnd cell_6t
Xbit_r165_c9 bl_9 br_9 wl_165 vdd gnd cell_6t
Xbit_r166_c9 bl_9 br_9 wl_166 vdd gnd cell_6t
Xbit_r167_c9 bl_9 br_9 wl_167 vdd gnd cell_6t
Xbit_r168_c9 bl_9 br_9 wl_168 vdd gnd cell_6t
Xbit_r169_c9 bl_9 br_9 wl_169 vdd gnd cell_6t
Xbit_r170_c9 bl_9 br_9 wl_170 vdd gnd cell_6t
Xbit_r171_c9 bl_9 br_9 wl_171 vdd gnd cell_6t
Xbit_r172_c9 bl_9 br_9 wl_172 vdd gnd cell_6t
Xbit_r173_c9 bl_9 br_9 wl_173 vdd gnd cell_6t
Xbit_r174_c9 bl_9 br_9 wl_174 vdd gnd cell_6t
Xbit_r175_c9 bl_9 br_9 wl_175 vdd gnd cell_6t
Xbit_r176_c9 bl_9 br_9 wl_176 vdd gnd cell_6t
Xbit_r177_c9 bl_9 br_9 wl_177 vdd gnd cell_6t
Xbit_r178_c9 bl_9 br_9 wl_178 vdd gnd cell_6t
Xbit_r179_c9 bl_9 br_9 wl_179 vdd gnd cell_6t
Xbit_r180_c9 bl_9 br_9 wl_180 vdd gnd cell_6t
Xbit_r181_c9 bl_9 br_9 wl_181 vdd gnd cell_6t
Xbit_r182_c9 bl_9 br_9 wl_182 vdd gnd cell_6t
Xbit_r183_c9 bl_9 br_9 wl_183 vdd gnd cell_6t
Xbit_r184_c9 bl_9 br_9 wl_184 vdd gnd cell_6t
Xbit_r185_c9 bl_9 br_9 wl_185 vdd gnd cell_6t
Xbit_r186_c9 bl_9 br_9 wl_186 vdd gnd cell_6t
Xbit_r187_c9 bl_9 br_9 wl_187 vdd gnd cell_6t
Xbit_r188_c9 bl_9 br_9 wl_188 vdd gnd cell_6t
Xbit_r189_c9 bl_9 br_9 wl_189 vdd gnd cell_6t
Xbit_r190_c9 bl_9 br_9 wl_190 vdd gnd cell_6t
Xbit_r191_c9 bl_9 br_9 wl_191 vdd gnd cell_6t
Xbit_r192_c9 bl_9 br_9 wl_192 vdd gnd cell_6t
Xbit_r193_c9 bl_9 br_9 wl_193 vdd gnd cell_6t
Xbit_r194_c9 bl_9 br_9 wl_194 vdd gnd cell_6t
Xbit_r195_c9 bl_9 br_9 wl_195 vdd gnd cell_6t
Xbit_r196_c9 bl_9 br_9 wl_196 vdd gnd cell_6t
Xbit_r197_c9 bl_9 br_9 wl_197 vdd gnd cell_6t
Xbit_r198_c9 bl_9 br_9 wl_198 vdd gnd cell_6t
Xbit_r199_c9 bl_9 br_9 wl_199 vdd gnd cell_6t
Xbit_r200_c9 bl_9 br_9 wl_200 vdd gnd cell_6t
Xbit_r201_c9 bl_9 br_9 wl_201 vdd gnd cell_6t
Xbit_r202_c9 bl_9 br_9 wl_202 vdd gnd cell_6t
Xbit_r203_c9 bl_9 br_9 wl_203 vdd gnd cell_6t
Xbit_r204_c9 bl_9 br_9 wl_204 vdd gnd cell_6t
Xbit_r205_c9 bl_9 br_9 wl_205 vdd gnd cell_6t
Xbit_r206_c9 bl_9 br_9 wl_206 vdd gnd cell_6t
Xbit_r207_c9 bl_9 br_9 wl_207 vdd gnd cell_6t
Xbit_r208_c9 bl_9 br_9 wl_208 vdd gnd cell_6t
Xbit_r209_c9 bl_9 br_9 wl_209 vdd gnd cell_6t
Xbit_r210_c9 bl_9 br_9 wl_210 vdd gnd cell_6t
Xbit_r211_c9 bl_9 br_9 wl_211 vdd gnd cell_6t
Xbit_r212_c9 bl_9 br_9 wl_212 vdd gnd cell_6t
Xbit_r213_c9 bl_9 br_9 wl_213 vdd gnd cell_6t
Xbit_r214_c9 bl_9 br_9 wl_214 vdd gnd cell_6t
Xbit_r215_c9 bl_9 br_9 wl_215 vdd gnd cell_6t
Xbit_r216_c9 bl_9 br_9 wl_216 vdd gnd cell_6t
Xbit_r217_c9 bl_9 br_9 wl_217 vdd gnd cell_6t
Xbit_r218_c9 bl_9 br_9 wl_218 vdd gnd cell_6t
Xbit_r219_c9 bl_9 br_9 wl_219 vdd gnd cell_6t
Xbit_r220_c9 bl_9 br_9 wl_220 vdd gnd cell_6t
Xbit_r221_c9 bl_9 br_9 wl_221 vdd gnd cell_6t
Xbit_r222_c9 bl_9 br_9 wl_222 vdd gnd cell_6t
Xbit_r223_c9 bl_9 br_9 wl_223 vdd gnd cell_6t
Xbit_r224_c9 bl_9 br_9 wl_224 vdd gnd cell_6t
Xbit_r225_c9 bl_9 br_9 wl_225 vdd gnd cell_6t
Xbit_r226_c9 bl_9 br_9 wl_226 vdd gnd cell_6t
Xbit_r227_c9 bl_9 br_9 wl_227 vdd gnd cell_6t
Xbit_r228_c9 bl_9 br_9 wl_228 vdd gnd cell_6t
Xbit_r229_c9 bl_9 br_9 wl_229 vdd gnd cell_6t
Xbit_r230_c9 bl_9 br_9 wl_230 vdd gnd cell_6t
Xbit_r231_c9 bl_9 br_9 wl_231 vdd gnd cell_6t
Xbit_r232_c9 bl_9 br_9 wl_232 vdd gnd cell_6t
Xbit_r233_c9 bl_9 br_9 wl_233 vdd gnd cell_6t
Xbit_r234_c9 bl_9 br_9 wl_234 vdd gnd cell_6t
Xbit_r235_c9 bl_9 br_9 wl_235 vdd gnd cell_6t
Xbit_r236_c9 bl_9 br_9 wl_236 vdd gnd cell_6t
Xbit_r237_c9 bl_9 br_9 wl_237 vdd gnd cell_6t
Xbit_r238_c9 bl_9 br_9 wl_238 vdd gnd cell_6t
Xbit_r239_c9 bl_9 br_9 wl_239 vdd gnd cell_6t
Xbit_r240_c9 bl_9 br_9 wl_240 vdd gnd cell_6t
Xbit_r241_c9 bl_9 br_9 wl_241 vdd gnd cell_6t
Xbit_r242_c9 bl_9 br_9 wl_242 vdd gnd cell_6t
Xbit_r243_c9 bl_9 br_9 wl_243 vdd gnd cell_6t
Xbit_r244_c9 bl_9 br_9 wl_244 vdd gnd cell_6t
Xbit_r245_c9 bl_9 br_9 wl_245 vdd gnd cell_6t
Xbit_r246_c9 bl_9 br_9 wl_246 vdd gnd cell_6t
Xbit_r247_c9 bl_9 br_9 wl_247 vdd gnd cell_6t
Xbit_r248_c9 bl_9 br_9 wl_248 vdd gnd cell_6t
Xbit_r249_c9 bl_9 br_9 wl_249 vdd gnd cell_6t
Xbit_r250_c9 bl_9 br_9 wl_250 vdd gnd cell_6t
Xbit_r251_c9 bl_9 br_9 wl_251 vdd gnd cell_6t
Xbit_r252_c9 bl_9 br_9 wl_252 vdd gnd cell_6t
Xbit_r253_c9 bl_9 br_9 wl_253 vdd gnd cell_6t
Xbit_r254_c9 bl_9 br_9 wl_254 vdd gnd cell_6t
Xbit_r255_c9 bl_9 br_9 wl_255 vdd gnd cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd cell_6t
Xbit_r1_c10 bl_10 br_10 wl_1 vdd gnd cell_6t
Xbit_r2_c10 bl_10 br_10 wl_2 vdd gnd cell_6t
Xbit_r3_c10 bl_10 br_10 wl_3 vdd gnd cell_6t
Xbit_r4_c10 bl_10 br_10 wl_4 vdd gnd cell_6t
Xbit_r5_c10 bl_10 br_10 wl_5 vdd gnd cell_6t
Xbit_r6_c10 bl_10 br_10 wl_6 vdd gnd cell_6t
Xbit_r7_c10 bl_10 br_10 wl_7 vdd gnd cell_6t
Xbit_r8_c10 bl_10 br_10 wl_8 vdd gnd cell_6t
Xbit_r9_c10 bl_10 br_10 wl_9 vdd gnd cell_6t
Xbit_r10_c10 bl_10 br_10 wl_10 vdd gnd cell_6t
Xbit_r11_c10 bl_10 br_10 wl_11 vdd gnd cell_6t
Xbit_r12_c10 bl_10 br_10 wl_12 vdd gnd cell_6t
Xbit_r13_c10 bl_10 br_10 wl_13 vdd gnd cell_6t
Xbit_r14_c10 bl_10 br_10 wl_14 vdd gnd cell_6t
Xbit_r15_c10 bl_10 br_10 wl_15 vdd gnd cell_6t
Xbit_r16_c10 bl_10 br_10 wl_16 vdd gnd cell_6t
Xbit_r17_c10 bl_10 br_10 wl_17 vdd gnd cell_6t
Xbit_r18_c10 bl_10 br_10 wl_18 vdd gnd cell_6t
Xbit_r19_c10 bl_10 br_10 wl_19 vdd gnd cell_6t
Xbit_r20_c10 bl_10 br_10 wl_20 vdd gnd cell_6t
Xbit_r21_c10 bl_10 br_10 wl_21 vdd gnd cell_6t
Xbit_r22_c10 bl_10 br_10 wl_22 vdd gnd cell_6t
Xbit_r23_c10 bl_10 br_10 wl_23 vdd gnd cell_6t
Xbit_r24_c10 bl_10 br_10 wl_24 vdd gnd cell_6t
Xbit_r25_c10 bl_10 br_10 wl_25 vdd gnd cell_6t
Xbit_r26_c10 bl_10 br_10 wl_26 vdd gnd cell_6t
Xbit_r27_c10 bl_10 br_10 wl_27 vdd gnd cell_6t
Xbit_r28_c10 bl_10 br_10 wl_28 vdd gnd cell_6t
Xbit_r29_c10 bl_10 br_10 wl_29 vdd gnd cell_6t
Xbit_r30_c10 bl_10 br_10 wl_30 vdd gnd cell_6t
Xbit_r31_c10 bl_10 br_10 wl_31 vdd gnd cell_6t
Xbit_r32_c10 bl_10 br_10 wl_32 vdd gnd cell_6t
Xbit_r33_c10 bl_10 br_10 wl_33 vdd gnd cell_6t
Xbit_r34_c10 bl_10 br_10 wl_34 vdd gnd cell_6t
Xbit_r35_c10 bl_10 br_10 wl_35 vdd gnd cell_6t
Xbit_r36_c10 bl_10 br_10 wl_36 vdd gnd cell_6t
Xbit_r37_c10 bl_10 br_10 wl_37 vdd gnd cell_6t
Xbit_r38_c10 bl_10 br_10 wl_38 vdd gnd cell_6t
Xbit_r39_c10 bl_10 br_10 wl_39 vdd gnd cell_6t
Xbit_r40_c10 bl_10 br_10 wl_40 vdd gnd cell_6t
Xbit_r41_c10 bl_10 br_10 wl_41 vdd gnd cell_6t
Xbit_r42_c10 bl_10 br_10 wl_42 vdd gnd cell_6t
Xbit_r43_c10 bl_10 br_10 wl_43 vdd gnd cell_6t
Xbit_r44_c10 bl_10 br_10 wl_44 vdd gnd cell_6t
Xbit_r45_c10 bl_10 br_10 wl_45 vdd gnd cell_6t
Xbit_r46_c10 bl_10 br_10 wl_46 vdd gnd cell_6t
Xbit_r47_c10 bl_10 br_10 wl_47 vdd gnd cell_6t
Xbit_r48_c10 bl_10 br_10 wl_48 vdd gnd cell_6t
Xbit_r49_c10 bl_10 br_10 wl_49 vdd gnd cell_6t
Xbit_r50_c10 bl_10 br_10 wl_50 vdd gnd cell_6t
Xbit_r51_c10 bl_10 br_10 wl_51 vdd gnd cell_6t
Xbit_r52_c10 bl_10 br_10 wl_52 vdd gnd cell_6t
Xbit_r53_c10 bl_10 br_10 wl_53 vdd gnd cell_6t
Xbit_r54_c10 bl_10 br_10 wl_54 vdd gnd cell_6t
Xbit_r55_c10 bl_10 br_10 wl_55 vdd gnd cell_6t
Xbit_r56_c10 bl_10 br_10 wl_56 vdd gnd cell_6t
Xbit_r57_c10 bl_10 br_10 wl_57 vdd gnd cell_6t
Xbit_r58_c10 bl_10 br_10 wl_58 vdd gnd cell_6t
Xbit_r59_c10 bl_10 br_10 wl_59 vdd gnd cell_6t
Xbit_r60_c10 bl_10 br_10 wl_60 vdd gnd cell_6t
Xbit_r61_c10 bl_10 br_10 wl_61 vdd gnd cell_6t
Xbit_r62_c10 bl_10 br_10 wl_62 vdd gnd cell_6t
Xbit_r63_c10 bl_10 br_10 wl_63 vdd gnd cell_6t
Xbit_r64_c10 bl_10 br_10 wl_64 vdd gnd cell_6t
Xbit_r65_c10 bl_10 br_10 wl_65 vdd gnd cell_6t
Xbit_r66_c10 bl_10 br_10 wl_66 vdd gnd cell_6t
Xbit_r67_c10 bl_10 br_10 wl_67 vdd gnd cell_6t
Xbit_r68_c10 bl_10 br_10 wl_68 vdd gnd cell_6t
Xbit_r69_c10 bl_10 br_10 wl_69 vdd gnd cell_6t
Xbit_r70_c10 bl_10 br_10 wl_70 vdd gnd cell_6t
Xbit_r71_c10 bl_10 br_10 wl_71 vdd gnd cell_6t
Xbit_r72_c10 bl_10 br_10 wl_72 vdd gnd cell_6t
Xbit_r73_c10 bl_10 br_10 wl_73 vdd gnd cell_6t
Xbit_r74_c10 bl_10 br_10 wl_74 vdd gnd cell_6t
Xbit_r75_c10 bl_10 br_10 wl_75 vdd gnd cell_6t
Xbit_r76_c10 bl_10 br_10 wl_76 vdd gnd cell_6t
Xbit_r77_c10 bl_10 br_10 wl_77 vdd gnd cell_6t
Xbit_r78_c10 bl_10 br_10 wl_78 vdd gnd cell_6t
Xbit_r79_c10 bl_10 br_10 wl_79 vdd gnd cell_6t
Xbit_r80_c10 bl_10 br_10 wl_80 vdd gnd cell_6t
Xbit_r81_c10 bl_10 br_10 wl_81 vdd gnd cell_6t
Xbit_r82_c10 bl_10 br_10 wl_82 vdd gnd cell_6t
Xbit_r83_c10 bl_10 br_10 wl_83 vdd gnd cell_6t
Xbit_r84_c10 bl_10 br_10 wl_84 vdd gnd cell_6t
Xbit_r85_c10 bl_10 br_10 wl_85 vdd gnd cell_6t
Xbit_r86_c10 bl_10 br_10 wl_86 vdd gnd cell_6t
Xbit_r87_c10 bl_10 br_10 wl_87 vdd gnd cell_6t
Xbit_r88_c10 bl_10 br_10 wl_88 vdd gnd cell_6t
Xbit_r89_c10 bl_10 br_10 wl_89 vdd gnd cell_6t
Xbit_r90_c10 bl_10 br_10 wl_90 vdd gnd cell_6t
Xbit_r91_c10 bl_10 br_10 wl_91 vdd gnd cell_6t
Xbit_r92_c10 bl_10 br_10 wl_92 vdd gnd cell_6t
Xbit_r93_c10 bl_10 br_10 wl_93 vdd gnd cell_6t
Xbit_r94_c10 bl_10 br_10 wl_94 vdd gnd cell_6t
Xbit_r95_c10 bl_10 br_10 wl_95 vdd gnd cell_6t
Xbit_r96_c10 bl_10 br_10 wl_96 vdd gnd cell_6t
Xbit_r97_c10 bl_10 br_10 wl_97 vdd gnd cell_6t
Xbit_r98_c10 bl_10 br_10 wl_98 vdd gnd cell_6t
Xbit_r99_c10 bl_10 br_10 wl_99 vdd gnd cell_6t
Xbit_r100_c10 bl_10 br_10 wl_100 vdd gnd cell_6t
Xbit_r101_c10 bl_10 br_10 wl_101 vdd gnd cell_6t
Xbit_r102_c10 bl_10 br_10 wl_102 vdd gnd cell_6t
Xbit_r103_c10 bl_10 br_10 wl_103 vdd gnd cell_6t
Xbit_r104_c10 bl_10 br_10 wl_104 vdd gnd cell_6t
Xbit_r105_c10 bl_10 br_10 wl_105 vdd gnd cell_6t
Xbit_r106_c10 bl_10 br_10 wl_106 vdd gnd cell_6t
Xbit_r107_c10 bl_10 br_10 wl_107 vdd gnd cell_6t
Xbit_r108_c10 bl_10 br_10 wl_108 vdd gnd cell_6t
Xbit_r109_c10 bl_10 br_10 wl_109 vdd gnd cell_6t
Xbit_r110_c10 bl_10 br_10 wl_110 vdd gnd cell_6t
Xbit_r111_c10 bl_10 br_10 wl_111 vdd gnd cell_6t
Xbit_r112_c10 bl_10 br_10 wl_112 vdd gnd cell_6t
Xbit_r113_c10 bl_10 br_10 wl_113 vdd gnd cell_6t
Xbit_r114_c10 bl_10 br_10 wl_114 vdd gnd cell_6t
Xbit_r115_c10 bl_10 br_10 wl_115 vdd gnd cell_6t
Xbit_r116_c10 bl_10 br_10 wl_116 vdd gnd cell_6t
Xbit_r117_c10 bl_10 br_10 wl_117 vdd gnd cell_6t
Xbit_r118_c10 bl_10 br_10 wl_118 vdd gnd cell_6t
Xbit_r119_c10 bl_10 br_10 wl_119 vdd gnd cell_6t
Xbit_r120_c10 bl_10 br_10 wl_120 vdd gnd cell_6t
Xbit_r121_c10 bl_10 br_10 wl_121 vdd gnd cell_6t
Xbit_r122_c10 bl_10 br_10 wl_122 vdd gnd cell_6t
Xbit_r123_c10 bl_10 br_10 wl_123 vdd gnd cell_6t
Xbit_r124_c10 bl_10 br_10 wl_124 vdd gnd cell_6t
Xbit_r125_c10 bl_10 br_10 wl_125 vdd gnd cell_6t
Xbit_r126_c10 bl_10 br_10 wl_126 vdd gnd cell_6t
Xbit_r127_c10 bl_10 br_10 wl_127 vdd gnd cell_6t
Xbit_r128_c10 bl_10 br_10 wl_128 vdd gnd cell_6t
Xbit_r129_c10 bl_10 br_10 wl_129 vdd gnd cell_6t
Xbit_r130_c10 bl_10 br_10 wl_130 vdd gnd cell_6t
Xbit_r131_c10 bl_10 br_10 wl_131 vdd gnd cell_6t
Xbit_r132_c10 bl_10 br_10 wl_132 vdd gnd cell_6t
Xbit_r133_c10 bl_10 br_10 wl_133 vdd gnd cell_6t
Xbit_r134_c10 bl_10 br_10 wl_134 vdd gnd cell_6t
Xbit_r135_c10 bl_10 br_10 wl_135 vdd gnd cell_6t
Xbit_r136_c10 bl_10 br_10 wl_136 vdd gnd cell_6t
Xbit_r137_c10 bl_10 br_10 wl_137 vdd gnd cell_6t
Xbit_r138_c10 bl_10 br_10 wl_138 vdd gnd cell_6t
Xbit_r139_c10 bl_10 br_10 wl_139 vdd gnd cell_6t
Xbit_r140_c10 bl_10 br_10 wl_140 vdd gnd cell_6t
Xbit_r141_c10 bl_10 br_10 wl_141 vdd gnd cell_6t
Xbit_r142_c10 bl_10 br_10 wl_142 vdd gnd cell_6t
Xbit_r143_c10 bl_10 br_10 wl_143 vdd gnd cell_6t
Xbit_r144_c10 bl_10 br_10 wl_144 vdd gnd cell_6t
Xbit_r145_c10 bl_10 br_10 wl_145 vdd gnd cell_6t
Xbit_r146_c10 bl_10 br_10 wl_146 vdd gnd cell_6t
Xbit_r147_c10 bl_10 br_10 wl_147 vdd gnd cell_6t
Xbit_r148_c10 bl_10 br_10 wl_148 vdd gnd cell_6t
Xbit_r149_c10 bl_10 br_10 wl_149 vdd gnd cell_6t
Xbit_r150_c10 bl_10 br_10 wl_150 vdd gnd cell_6t
Xbit_r151_c10 bl_10 br_10 wl_151 vdd gnd cell_6t
Xbit_r152_c10 bl_10 br_10 wl_152 vdd gnd cell_6t
Xbit_r153_c10 bl_10 br_10 wl_153 vdd gnd cell_6t
Xbit_r154_c10 bl_10 br_10 wl_154 vdd gnd cell_6t
Xbit_r155_c10 bl_10 br_10 wl_155 vdd gnd cell_6t
Xbit_r156_c10 bl_10 br_10 wl_156 vdd gnd cell_6t
Xbit_r157_c10 bl_10 br_10 wl_157 vdd gnd cell_6t
Xbit_r158_c10 bl_10 br_10 wl_158 vdd gnd cell_6t
Xbit_r159_c10 bl_10 br_10 wl_159 vdd gnd cell_6t
Xbit_r160_c10 bl_10 br_10 wl_160 vdd gnd cell_6t
Xbit_r161_c10 bl_10 br_10 wl_161 vdd gnd cell_6t
Xbit_r162_c10 bl_10 br_10 wl_162 vdd gnd cell_6t
Xbit_r163_c10 bl_10 br_10 wl_163 vdd gnd cell_6t
Xbit_r164_c10 bl_10 br_10 wl_164 vdd gnd cell_6t
Xbit_r165_c10 bl_10 br_10 wl_165 vdd gnd cell_6t
Xbit_r166_c10 bl_10 br_10 wl_166 vdd gnd cell_6t
Xbit_r167_c10 bl_10 br_10 wl_167 vdd gnd cell_6t
Xbit_r168_c10 bl_10 br_10 wl_168 vdd gnd cell_6t
Xbit_r169_c10 bl_10 br_10 wl_169 vdd gnd cell_6t
Xbit_r170_c10 bl_10 br_10 wl_170 vdd gnd cell_6t
Xbit_r171_c10 bl_10 br_10 wl_171 vdd gnd cell_6t
Xbit_r172_c10 bl_10 br_10 wl_172 vdd gnd cell_6t
Xbit_r173_c10 bl_10 br_10 wl_173 vdd gnd cell_6t
Xbit_r174_c10 bl_10 br_10 wl_174 vdd gnd cell_6t
Xbit_r175_c10 bl_10 br_10 wl_175 vdd gnd cell_6t
Xbit_r176_c10 bl_10 br_10 wl_176 vdd gnd cell_6t
Xbit_r177_c10 bl_10 br_10 wl_177 vdd gnd cell_6t
Xbit_r178_c10 bl_10 br_10 wl_178 vdd gnd cell_6t
Xbit_r179_c10 bl_10 br_10 wl_179 vdd gnd cell_6t
Xbit_r180_c10 bl_10 br_10 wl_180 vdd gnd cell_6t
Xbit_r181_c10 bl_10 br_10 wl_181 vdd gnd cell_6t
Xbit_r182_c10 bl_10 br_10 wl_182 vdd gnd cell_6t
Xbit_r183_c10 bl_10 br_10 wl_183 vdd gnd cell_6t
Xbit_r184_c10 bl_10 br_10 wl_184 vdd gnd cell_6t
Xbit_r185_c10 bl_10 br_10 wl_185 vdd gnd cell_6t
Xbit_r186_c10 bl_10 br_10 wl_186 vdd gnd cell_6t
Xbit_r187_c10 bl_10 br_10 wl_187 vdd gnd cell_6t
Xbit_r188_c10 bl_10 br_10 wl_188 vdd gnd cell_6t
Xbit_r189_c10 bl_10 br_10 wl_189 vdd gnd cell_6t
Xbit_r190_c10 bl_10 br_10 wl_190 vdd gnd cell_6t
Xbit_r191_c10 bl_10 br_10 wl_191 vdd gnd cell_6t
Xbit_r192_c10 bl_10 br_10 wl_192 vdd gnd cell_6t
Xbit_r193_c10 bl_10 br_10 wl_193 vdd gnd cell_6t
Xbit_r194_c10 bl_10 br_10 wl_194 vdd gnd cell_6t
Xbit_r195_c10 bl_10 br_10 wl_195 vdd gnd cell_6t
Xbit_r196_c10 bl_10 br_10 wl_196 vdd gnd cell_6t
Xbit_r197_c10 bl_10 br_10 wl_197 vdd gnd cell_6t
Xbit_r198_c10 bl_10 br_10 wl_198 vdd gnd cell_6t
Xbit_r199_c10 bl_10 br_10 wl_199 vdd gnd cell_6t
Xbit_r200_c10 bl_10 br_10 wl_200 vdd gnd cell_6t
Xbit_r201_c10 bl_10 br_10 wl_201 vdd gnd cell_6t
Xbit_r202_c10 bl_10 br_10 wl_202 vdd gnd cell_6t
Xbit_r203_c10 bl_10 br_10 wl_203 vdd gnd cell_6t
Xbit_r204_c10 bl_10 br_10 wl_204 vdd gnd cell_6t
Xbit_r205_c10 bl_10 br_10 wl_205 vdd gnd cell_6t
Xbit_r206_c10 bl_10 br_10 wl_206 vdd gnd cell_6t
Xbit_r207_c10 bl_10 br_10 wl_207 vdd gnd cell_6t
Xbit_r208_c10 bl_10 br_10 wl_208 vdd gnd cell_6t
Xbit_r209_c10 bl_10 br_10 wl_209 vdd gnd cell_6t
Xbit_r210_c10 bl_10 br_10 wl_210 vdd gnd cell_6t
Xbit_r211_c10 bl_10 br_10 wl_211 vdd gnd cell_6t
Xbit_r212_c10 bl_10 br_10 wl_212 vdd gnd cell_6t
Xbit_r213_c10 bl_10 br_10 wl_213 vdd gnd cell_6t
Xbit_r214_c10 bl_10 br_10 wl_214 vdd gnd cell_6t
Xbit_r215_c10 bl_10 br_10 wl_215 vdd gnd cell_6t
Xbit_r216_c10 bl_10 br_10 wl_216 vdd gnd cell_6t
Xbit_r217_c10 bl_10 br_10 wl_217 vdd gnd cell_6t
Xbit_r218_c10 bl_10 br_10 wl_218 vdd gnd cell_6t
Xbit_r219_c10 bl_10 br_10 wl_219 vdd gnd cell_6t
Xbit_r220_c10 bl_10 br_10 wl_220 vdd gnd cell_6t
Xbit_r221_c10 bl_10 br_10 wl_221 vdd gnd cell_6t
Xbit_r222_c10 bl_10 br_10 wl_222 vdd gnd cell_6t
Xbit_r223_c10 bl_10 br_10 wl_223 vdd gnd cell_6t
Xbit_r224_c10 bl_10 br_10 wl_224 vdd gnd cell_6t
Xbit_r225_c10 bl_10 br_10 wl_225 vdd gnd cell_6t
Xbit_r226_c10 bl_10 br_10 wl_226 vdd gnd cell_6t
Xbit_r227_c10 bl_10 br_10 wl_227 vdd gnd cell_6t
Xbit_r228_c10 bl_10 br_10 wl_228 vdd gnd cell_6t
Xbit_r229_c10 bl_10 br_10 wl_229 vdd gnd cell_6t
Xbit_r230_c10 bl_10 br_10 wl_230 vdd gnd cell_6t
Xbit_r231_c10 bl_10 br_10 wl_231 vdd gnd cell_6t
Xbit_r232_c10 bl_10 br_10 wl_232 vdd gnd cell_6t
Xbit_r233_c10 bl_10 br_10 wl_233 vdd gnd cell_6t
Xbit_r234_c10 bl_10 br_10 wl_234 vdd gnd cell_6t
Xbit_r235_c10 bl_10 br_10 wl_235 vdd gnd cell_6t
Xbit_r236_c10 bl_10 br_10 wl_236 vdd gnd cell_6t
Xbit_r237_c10 bl_10 br_10 wl_237 vdd gnd cell_6t
Xbit_r238_c10 bl_10 br_10 wl_238 vdd gnd cell_6t
Xbit_r239_c10 bl_10 br_10 wl_239 vdd gnd cell_6t
Xbit_r240_c10 bl_10 br_10 wl_240 vdd gnd cell_6t
Xbit_r241_c10 bl_10 br_10 wl_241 vdd gnd cell_6t
Xbit_r242_c10 bl_10 br_10 wl_242 vdd gnd cell_6t
Xbit_r243_c10 bl_10 br_10 wl_243 vdd gnd cell_6t
Xbit_r244_c10 bl_10 br_10 wl_244 vdd gnd cell_6t
Xbit_r245_c10 bl_10 br_10 wl_245 vdd gnd cell_6t
Xbit_r246_c10 bl_10 br_10 wl_246 vdd gnd cell_6t
Xbit_r247_c10 bl_10 br_10 wl_247 vdd gnd cell_6t
Xbit_r248_c10 bl_10 br_10 wl_248 vdd gnd cell_6t
Xbit_r249_c10 bl_10 br_10 wl_249 vdd gnd cell_6t
Xbit_r250_c10 bl_10 br_10 wl_250 vdd gnd cell_6t
Xbit_r251_c10 bl_10 br_10 wl_251 vdd gnd cell_6t
Xbit_r252_c10 bl_10 br_10 wl_252 vdd gnd cell_6t
Xbit_r253_c10 bl_10 br_10 wl_253 vdd gnd cell_6t
Xbit_r254_c10 bl_10 br_10 wl_254 vdd gnd cell_6t
Xbit_r255_c10 bl_10 br_10 wl_255 vdd gnd cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd cell_6t
Xbit_r1_c11 bl_11 br_11 wl_1 vdd gnd cell_6t
Xbit_r2_c11 bl_11 br_11 wl_2 vdd gnd cell_6t
Xbit_r3_c11 bl_11 br_11 wl_3 vdd gnd cell_6t
Xbit_r4_c11 bl_11 br_11 wl_4 vdd gnd cell_6t
Xbit_r5_c11 bl_11 br_11 wl_5 vdd gnd cell_6t
Xbit_r6_c11 bl_11 br_11 wl_6 vdd gnd cell_6t
Xbit_r7_c11 bl_11 br_11 wl_7 vdd gnd cell_6t
Xbit_r8_c11 bl_11 br_11 wl_8 vdd gnd cell_6t
Xbit_r9_c11 bl_11 br_11 wl_9 vdd gnd cell_6t
Xbit_r10_c11 bl_11 br_11 wl_10 vdd gnd cell_6t
Xbit_r11_c11 bl_11 br_11 wl_11 vdd gnd cell_6t
Xbit_r12_c11 bl_11 br_11 wl_12 vdd gnd cell_6t
Xbit_r13_c11 bl_11 br_11 wl_13 vdd gnd cell_6t
Xbit_r14_c11 bl_11 br_11 wl_14 vdd gnd cell_6t
Xbit_r15_c11 bl_11 br_11 wl_15 vdd gnd cell_6t
Xbit_r16_c11 bl_11 br_11 wl_16 vdd gnd cell_6t
Xbit_r17_c11 bl_11 br_11 wl_17 vdd gnd cell_6t
Xbit_r18_c11 bl_11 br_11 wl_18 vdd gnd cell_6t
Xbit_r19_c11 bl_11 br_11 wl_19 vdd gnd cell_6t
Xbit_r20_c11 bl_11 br_11 wl_20 vdd gnd cell_6t
Xbit_r21_c11 bl_11 br_11 wl_21 vdd gnd cell_6t
Xbit_r22_c11 bl_11 br_11 wl_22 vdd gnd cell_6t
Xbit_r23_c11 bl_11 br_11 wl_23 vdd gnd cell_6t
Xbit_r24_c11 bl_11 br_11 wl_24 vdd gnd cell_6t
Xbit_r25_c11 bl_11 br_11 wl_25 vdd gnd cell_6t
Xbit_r26_c11 bl_11 br_11 wl_26 vdd gnd cell_6t
Xbit_r27_c11 bl_11 br_11 wl_27 vdd gnd cell_6t
Xbit_r28_c11 bl_11 br_11 wl_28 vdd gnd cell_6t
Xbit_r29_c11 bl_11 br_11 wl_29 vdd gnd cell_6t
Xbit_r30_c11 bl_11 br_11 wl_30 vdd gnd cell_6t
Xbit_r31_c11 bl_11 br_11 wl_31 vdd gnd cell_6t
Xbit_r32_c11 bl_11 br_11 wl_32 vdd gnd cell_6t
Xbit_r33_c11 bl_11 br_11 wl_33 vdd gnd cell_6t
Xbit_r34_c11 bl_11 br_11 wl_34 vdd gnd cell_6t
Xbit_r35_c11 bl_11 br_11 wl_35 vdd gnd cell_6t
Xbit_r36_c11 bl_11 br_11 wl_36 vdd gnd cell_6t
Xbit_r37_c11 bl_11 br_11 wl_37 vdd gnd cell_6t
Xbit_r38_c11 bl_11 br_11 wl_38 vdd gnd cell_6t
Xbit_r39_c11 bl_11 br_11 wl_39 vdd gnd cell_6t
Xbit_r40_c11 bl_11 br_11 wl_40 vdd gnd cell_6t
Xbit_r41_c11 bl_11 br_11 wl_41 vdd gnd cell_6t
Xbit_r42_c11 bl_11 br_11 wl_42 vdd gnd cell_6t
Xbit_r43_c11 bl_11 br_11 wl_43 vdd gnd cell_6t
Xbit_r44_c11 bl_11 br_11 wl_44 vdd gnd cell_6t
Xbit_r45_c11 bl_11 br_11 wl_45 vdd gnd cell_6t
Xbit_r46_c11 bl_11 br_11 wl_46 vdd gnd cell_6t
Xbit_r47_c11 bl_11 br_11 wl_47 vdd gnd cell_6t
Xbit_r48_c11 bl_11 br_11 wl_48 vdd gnd cell_6t
Xbit_r49_c11 bl_11 br_11 wl_49 vdd gnd cell_6t
Xbit_r50_c11 bl_11 br_11 wl_50 vdd gnd cell_6t
Xbit_r51_c11 bl_11 br_11 wl_51 vdd gnd cell_6t
Xbit_r52_c11 bl_11 br_11 wl_52 vdd gnd cell_6t
Xbit_r53_c11 bl_11 br_11 wl_53 vdd gnd cell_6t
Xbit_r54_c11 bl_11 br_11 wl_54 vdd gnd cell_6t
Xbit_r55_c11 bl_11 br_11 wl_55 vdd gnd cell_6t
Xbit_r56_c11 bl_11 br_11 wl_56 vdd gnd cell_6t
Xbit_r57_c11 bl_11 br_11 wl_57 vdd gnd cell_6t
Xbit_r58_c11 bl_11 br_11 wl_58 vdd gnd cell_6t
Xbit_r59_c11 bl_11 br_11 wl_59 vdd gnd cell_6t
Xbit_r60_c11 bl_11 br_11 wl_60 vdd gnd cell_6t
Xbit_r61_c11 bl_11 br_11 wl_61 vdd gnd cell_6t
Xbit_r62_c11 bl_11 br_11 wl_62 vdd gnd cell_6t
Xbit_r63_c11 bl_11 br_11 wl_63 vdd gnd cell_6t
Xbit_r64_c11 bl_11 br_11 wl_64 vdd gnd cell_6t
Xbit_r65_c11 bl_11 br_11 wl_65 vdd gnd cell_6t
Xbit_r66_c11 bl_11 br_11 wl_66 vdd gnd cell_6t
Xbit_r67_c11 bl_11 br_11 wl_67 vdd gnd cell_6t
Xbit_r68_c11 bl_11 br_11 wl_68 vdd gnd cell_6t
Xbit_r69_c11 bl_11 br_11 wl_69 vdd gnd cell_6t
Xbit_r70_c11 bl_11 br_11 wl_70 vdd gnd cell_6t
Xbit_r71_c11 bl_11 br_11 wl_71 vdd gnd cell_6t
Xbit_r72_c11 bl_11 br_11 wl_72 vdd gnd cell_6t
Xbit_r73_c11 bl_11 br_11 wl_73 vdd gnd cell_6t
Xbit_r74_c11 bl_11 br_11 wl_74 vdd gnd cell_6t
Xbit_r75_c11 bl_11 br_11 wl_75 vdd gnd cell_6t
Xbit_r76_c11 bl_11 br_11 wl_76 vdd gnd cell_6t
Xbit_r77_c11 bl_11 br_11 wl_77 vdd gnd cell_6t
Xbit_r78_c11 bl_11 br_11 wl_78 vdd gnd cell_6t
Xbit_r79_c11 bl_11 br_11 wl_79 vdd gnd cell_6t
Xbit_r80_c11 bl_11 br_11 wl_80 vdd gnd cell_6t
Xbit_r81_c11 bl_11 br_11 wl_81 vdd gnd cell_6t
Xbit_r82_c11 bl_11 br_11 wl_82 vdd gnd cell_6t
Xbit_r83_c11 bl_11 br_11 wl_83 vdd gnd cell_6t
Xbit_r84_c11 bl_11 br_11 wl_84 vdd gnd cell_6t
Xbit_r85_c11 bl_11 br_11 wl_85 vdd gnd cell_6t
Xbit_r86_c11 bl_11 br_11 wl_86 vdd gnd cell_6t
Xbit_r87_c11 bl_11 br_11 wl_87 vdd gnd cell_6t
Xbit_r88_c11 bl_11 br_11 wl_88 vdd gnd cell_6t
Xbit_r89_c11 bl_11 br_11 wl_89 vdd gnd cell_6t
Xbit_r90_c11 bl_11 br_11 wl_90 vdd gnd cell_6t
Xbit_r91_c11 bl_11 br_11 wl_91 vdd gnd cell_6t
Xbit_r92_c11 bl_11 br_11 wl_92 vdd gnd cell_6t
Xbit_r93_c11 bl_11 br_11 wl_93 vdd gnd cell_6t
Xbit_r94_c11 bl_11 br_11 wl_94 vdd gnd cell_6t
Xbit_r95_c11 bl_11 br_11 wl_95 vdd gnd cell_6t
Xbit_r96_c11 bl_11 br_11 wl_96 vdd gnd cell_6t
Xbit_r97_c11 bl_11 br_11 wl_97 vdd gnd cell_6t
Xbit_r98_c11 bl_11 br_11 wl_98 vdd gnd cell_6t
Xbit_r99_c11 bl_11 br_11 wl_99 vdd gnd cell_6t
Xbit_r100_c11 bl_11 br_11 wl_100 vdd gnd cell_6t
Xbit_r101_c11 bl_11 br_11 wl_101 vdd gnd cell_6t
Xbit_r102_c11 bl_11 br_11 wl_102 vdd gnd cell_6t
Xbit_r103_c11 bl_11 br_11 wl_103 vdd gnd cell_6t
Xbit_r104_c11 bl_11 br_11 wl_104 vdd gnd cell_6t
Xbit_r105_c11 bl_11 br_11 wl_105 vdd gnd cell_6t
Xbit_r106_c11 bl_11 br_11 wl_106 vdd gnd cell_6t
Xbit_r107_c11 bl_11 br_11 wl_107 vdd gnd cell_6t
Xbit_r108_c11 bl_11 br_11 wl_108 vdd gnd cell_6t
Xbit_r109_c11 bl_11 br_11 wl_109 vdd gnd cell_6t
Xbit_r110_c11 bl_11 br_11 wl_110 vdd gnd cell_6t
Xbit_r111_c11 bl_11 br_11 wl_111 vdd gnd cell_6t
Xbit_r112_c11 bl_11 br_11 wl_112 vdd gnd cell_6t
Xbit_r113_c11 bl_11 br_11 wl_113 vdd gnd cell_6t
Xbit_r114_c11 bl_11 br_11 wl_114 vdd gnd cell_6t
Xbit_r115_c11 bl_11 br_11 wl_115 vdd gnd cell_6t
Xbit_r116_c11 bl_11 br_11 wl_116 vdd gnd cell_6t
Xbit_r117_c11 bl_11 br_11 wl_117 vdd gnd cell_6t
Xbit_r118_c11 bl_11 br_11 wl_118 vdd gnd cell_6t
Xbit_r119_c11 bl_11 br_11 wl_119 vdd gnd cell_6t
Xbit_r120_c11 bl_11 br_11 wl_120 vdd gnd cell_6t
Xbit_r121_c11 bl_11 br_11 wl_121 vdd gnd cell_6t
Xbit_r122_c11 bl_11 br_11 wl_122 vdd gnd cell_6t
Xbit_r123_c11 bl_11 br_11 wl_123 vdd gnd cell_6t
Xbit_r124_c11 bl_11 br_11 wl_124 vdd gnd cell_6t
Xbit_r125_c11 bl_11 br_11 wl_125 vdd gnd cell_6t
Xbit_r126_c11 bl_11 br_11 wl_126 vdd gnd cell_6t
Xbit_r127_c11 bl_11 br_11 wl_127 vdd gnd cell_6t
Xbit_r128_c11 bl_11 br_11 wl_128 vdd gnd cell_6t
Xbit_r129_c11 bl_11 br_11 wl_129 vdd gnd cell_6t
Xbit_r130_c11 bl_11 br_11 wl_130 vdd gnd cell_6t
Xbit_r131_c11 bl_11 br_11 wl_131 vdd gnd cell_6t
Xbit_r132_c11 bl_11 br_11 wl_132 vdd gnd cell_6t
Xbit_r133_c11 bl_11 br_11 wl_133 vdd gnd cell_6t
Xbit_r134_c11 bl_11 br_11 wl_134 vdd gnd cell_6t
Xbit_r135_c11 bl_11 br_11 wl_135 vdd gnd cell_6t
Xbit_r136_c11 bl_11 br_11 wl_136 vdd gnd cell_6t
Xbit_r137_c11 bl_11 br_11 wl_137 vdd gnd cell_6t
Xbit_r138_c11 bl_11 br_11 wl_138 vdd gnd cell_6t
Xbit_r139_c11 bl_11 br_11 wl_139 vdd gnd cell_6t
Xbit_r140_c11 bl_11 br_11 wl_140 vdd gnd cell_6t
Xbit_r141_c11 bl_11 br_11 wl_141 vdd gnd cell_6t
Xbit_r142_c11 bl_11 br_11 wl_142 vdd gnd cell_6t
Xbit_r143_c11 bl_11 br_11 wl_143 vdd gnd cell_6t
Xbit_r144_c11 bl_11 br_11 wl_144 vdd gnd cell_6t
Xbit_r145_c11 bl_11 br_11 wl_145 vdd gnd cell_6t
Xbit_r146_c11 bl_11 br_11 wl_146 vdd gnd cell_6t
Xbit_r147_c11 bl_11 br_11 wl_147 vdd gnd cell_6t
Xbit_r148_c11 bl_11 br_11 wl_148 vdd gnd cell_6t
Xbit_r149_c11 bl_11 br_11 wl_149 vdd gnd cell_6t
Xbit_r150_c11 bl_11 br_11 wl_150 vdd gnd cell_6t
Xbit_r151_c11 bl_11 br_11 wl_151 vdd gnd cell_6t
Xbit_r152_c11 bl_11 br_11 wl_152 vdd gnd cell_6t
Xbit_r153_c11 bl_11 br_11 wl_153 vdd gnd cell_6t
Xbit_r154_c11 bl_11 br_11 wl_154 vdd gnd cell_6t
Xbit_r155_c11 bl_11 br_11 wl_155 vdd gnd cell_6t
Xbit_r156_c11 bl_11 br_11 wl_156 vdd gnd cell_6t
Xbit_r157_c11 bl_11 br_11 wl_157 vdd gnd cell_6t
Xbit_r158_c11 bl_11 br_11 wl_158 vdd gnd cell_6t
Xbit_r159_c11 bl_11 br_11 wl_159 vdd gnd cell_6t
Xbit_r160_c11 bl_11 br_11 wl_160 vdd gnd cell_6t
Xbit_r161_c11 bl_11 br_11 wl_161 vdd gnd cell_6t
Xbit_r162_c11 bl_11 br_11 wl_162 vdd gnd cell_6t
Xbit_r163_c11 bl_11 br_11 wl_163 vdd gnd cell_6t
Xbit_r164_c11 bl_11 br_11 wl_164 vdd gnd cell_6t
Xbit_r165_c11 bl_11 br_11 wl_165 vdd gnd cell_6t
Xbit_r166_c11 bl_11 br_11 wl_166 vdd gnd cell_6t
Xbit_r167_c11 bl_11 br_11 wl_167 vdd gnd cell_6t
Xbit_r168_c11 bl_11 br_11 wl_168 vdd gnd cell_6t
Xbit_r169_c11 bl_11 br_11 wl_169 vdd gnd cell_6t
Xbit_r170_c11 bl_11 br_11 wl_170 vdd gnd cell_6t
Xbit_r171_c11 bl_11 br_11 wl_171 vdd gnd cell_6t
Xbit_r172_c11 bl_11 br_11 wl_172 vdd gnd cell_6t
Xbit_r173_c11 bl_11 br_11 wl_173 vdd gnd cell_6t
Xbit_r174_c11 bl_11 br_11 wl_174 vdd gnd cell_6t
Xbit_r175_c11 bl_11 br_11 wl_175 vdd gnd cell_6t
Xbit_r176_c11 bl_11 br_11 wl_176 vdd gnd cell_6t
Xbit_r177_c11 bl_11 br_11 wl_177 vdd gnd cell_6t
Xbit_r178_c11 bl_11 br_11 wl_178 vdd gnd cell_6t
Xbit_r179_c11 bl_11 br_11 wl_179 vdd gnd cell_6t
Xbit_r180_c11 bl_11 br_11 wl_180 vdd gnd cell_6t
Xbit_r181_c11 bl_11 br_11 wl_181 vdd gnd cell_6t
Xbit_r182_c11 bl_11 br_11 wl_182 vdd gnd cell_6t
Xbit_r183_c11 bl_11 br_11 wl_183 vdd gnd cell_6t
Xbit_r184_c11 bl_11 br_11 wl_184 vdd gnd cell_6t
Xbit_r185_c11 bl_11 br_11 wl_185 vdd gnd cell_6t
Xbit_r186_c11 bl_11 br_11 wl_186 vdd gnd cell_6t
Xbit_r187_c11 bl_11 br_11 wl_187 vdd gnd cell_6t
Xbit_r188_c11 bl_11 br_11 wl_188 vdd gnd cell_6t
Xbit_r189_c11 bl_11 br_11 wl_189 vdd gnd cell_6t
Xbit_r190_c11 bl_11 br_11 wl_190 vdd gnd cell_6t
Xbit_r191_c11 bl_11 br_11 wl_191 vdd gnd cell_6t
Xbit_r192_c11 bl_11 br_11 wl_192 vdd gnd cell_6t
Xbit_r193_c11 bl_11 br_11 wl_193 vdd gnd cell_6t
Xbit_r194_c11 bl_11 br_11 wl_194 vdd gnd cell_6t
Xbit_r195_c11 bl_11 br_11 wl_195 vdd gnd cell_6t
Xbit_r196_c11 bl_11 br_11 wl_196 vdd gnd cell_6t
Xbit_r197_c11 bl_11 br_11 wl_197 vdd gnd cell_6t
Xbit_r198_c11 bl_11 br_11 wl_198 vdd gnd cell_6t
Xbit_r199_c11 bl_11 br_11 wl_199 vdd gnd cell_6t
Xbit_r200_c11 bl_11 br_11 wl_200 vdd gnd cell_6t
Xbit_r201_c11 bl_11 br_11 wl_201 vdd gnd cell_6t
Xbit_r202_c11 bl_11 br_11 wl_202 vdd gnd cell_6t
Xbit_r203_c11 bl_11 br_11 wl_203 vdd gnd cell_6t
Xbit_r204_c11 bl_11 br_11 wl_204 vdd gnd cell_6t
Xbit_r205_c11 bl_11 br_11 wl_205 vdd gnd cell_6t
Xbit_r206_c11 bl_11 br_11 wl_206 vdd gnd cell_6t
Xbit_r207_c11 bl_11 br_11 wl_207 vdd gnd cell_6t
Xbit_r208_c11 bl_11 br_11 wl_208 vdd gnd cell_6t
Xbit_r209_c11 bl_11 br_11 wl_209 vdd gnd cell_6t
Xbit_r210_c11 bl_11 br_11 wl_210 vdd gnd cell_6t
Xbit_r211_c11 bl_11 br_11 wl_211 vdd gnd cell_6t
Xbit_r212_c11 bl_11 br_11 wl_212 vdd gnd cell_6t
Xbit_r213_c11 bl_11 br_11 wl_213 vdd gnd cell_6t
Xbit_r214_c11 bl_11 br_11 wl_214 vdd gnd cell_6t
Xbit_r215_c11 bl_11 br_11 wl_215 vdd gnd cell_6t
Xbit_r216_c11 bl_11 br_11 wl_216 vdd gnd cell_6t
Xbit_r217_c11 bl_11 br_11 wl_217 vdd gnd cell_6t
Xbit_r218_c11 bl_11 br_11 wl_218 vdd gnd cell_6t
Xbit_r219_c11 bl_11 br_11 wl_219 vdd gnd cell_6t
Xbit_r220_c11 bl_11 br_11 wl_220 vdd gnd cell_6t
Xbit_r221_c11 bl_11 br_11 wl_221 vdd gnd cell_6t
Xbit_r222_c11 bl_11 br_11 wl_222 vdd gnd cell_6t
Xbit_r223_c11 bl_11 br_11 wl_223 vdd gnd cell_6t
Xbit_r224_c11 bl_11 br_11 wl_224 vdd gnd cell_6t
Xbit_r225_c11 bl_11 br_11 wl_225 vdd gnd cell_6t
Xbit_r226_c11 bl_11 br_11 wl_226 vdd gnd cell_6t
Xbit_r227_c11 bl_11 br_11 wl_227 vdd gnd cell_6t
Xbit_r228_c11 bl_11 br_11 wl_228 vdd gnd cell_6t
Xbit_r229_c11 bl_11 br_11 wl_229 vdd gnd cell_6t
Xbit_r230_c11 bl_11 br_11 wl_230 vdd gnd cell_6t
Xbit_r231_c11 bl_11 br_11 wl_231 vdd gnd cell_6t
Xbit_r232_c11 bl_11 br_11 wl_232 vdd gnd cell_6t
Xbit_r233_c11 bl_11 br_11 wl_233 vdd gnd cell_6t
Xbit_r234_c11 bl_11 br_11 wl_234 vdd gnd cell_6t
Xbit_r235_c11 bl_11 br_11 wl_235 vdd gnd cell_6t
Xbit_r236_c11 bl_11 br_11 wl_236 vdd gnd cell_6t
Xbit_r237_c11 bl_11 br_11 wl_237 vdd gnd cell_6t
Xbit_r238_c11 bl_11 br_11 wl_238 vdd gnd cell_6t
Xbit_r239_c11 bl_11 br_11 wl_239 vdd gnd cell_6t
Xbit_r240_c11 bl_11 br_11 wl_240 vdd gnd cell_6t
Xbit_r241_c11 bl_11 br_11 wl_241 vdd gnd cell_6t
Xbit_r242_c11 bl_11 br_11 wl_242 vdd gnd cell_6t
Xbit_r243_c11 bl_11 br_11 wl_243 vdd gnd cell_6t
Xbit_r244_c11 bl_11 br_11 wl_244 vdd gnd cell_6t
Xbit_r245_c11 bl_11 br_11 wl_245 vdd gnd cell_6t
Xbit_r246_c11 bl_11 br_11 wl_246 vdd gnd cell_6t
Xbit_r247_c11 bl_11 br_11 wl_247 vdd gnd cell_6t
Xbit_r248_c11 bl_11 br_11 wl_248 vdd gnd cell_6t
Xbit_r249_c11 bl_11 br_11 wl_249 vdd gnd cell_6t
Xbit_r250_c11 bl_11 br_11 wl_250 vdd gnd cell_6t
Xbit_r251_c11 bl_11 br_11 wl_251 vdd gnd cell_6t
Xbit_r252_c11 bl_11 br_11 wl_252 vdd gnd cell_6t
Xbit_r253_c11 bl_11 br_11 wl_253 vdd gnd cell_6t
Xbit_r254_c11 bl_11 br_11 wl_254 vdd gnd cell_6t
Xbit_r255_c11 bl_11 br_11 wl_255 vdd gnd cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd cell_6t
Xbit_r1_c12 bl_12 br_12 wl_1 vdd gnd cell_6t
Xbit_r2_c12 bl_12 br_12 wl_2 vdd gnd cell_6t
Xbit_r3_c12 bl_12 br_12 wl_3 vdd gnd cell_6t
Xbit_r4_c12 bl_12 br_12 wl_4 vdd gnd cell_6t
Xbit_r5_c12 bl_12 br_12 wl_5 vdd gnd cell_6t
Xbit_r6_c12 bl_12 br_12 wl_6 vdd gnd cell_6t
Xbit_r7_c12 bl_12 br_12 wl_7 vdd gnd cell_6t
Xbit_r8_c12 bl_12 br_12 wl_8 vdd gnd cell_6t
Xbit_r9_c12 bl_12 br_12 wl_9 vdd gnd cell_6t
Xbit_r10_c12 bl_12 br_12 wl_10 vdd gnd cell_6t
Xbit_r11_c12 bl_12 br_12 wl_11 vdd gnd cell_6t
Xbit_r12_c12 bl_12 br_12 wl_12 vdd gnd cell_6t
Xbit_r13_c12 bl_12 br_12 wl_13 vdd gnd cell_6t
Xbit_r14_c12 bl_12 br_12 wl_14 vdd gnd cell_6t
Xbit_r15_c12 bl_12 br_12 wl_15 vdd gnd cell_6t
Xbit_r16_c12 bl_12 br_12 wl_16 vdd gnd cell_6t
Xbit_r17_c12 bl_12 br_12 wl_17 vdd gnd cell_6t
Xbit_r18_c12 bl_12 br_12 wl_18 vdd gnd cell_6t
Xbit_r19_c12 bl_12 br_12 wl_19 vdd gnd cell_6t
Xbit_r20_c12 bl_12 br_12 wl_20 vdd gnd cell_6t
Xbit_r21_c12 bl_12 br_12 wl_21 vdd gnd cell_6t
Xbit_r22_c12 bl_12 br_12 wl_22 vdd gnd cell_6t
Xbit_r23_c12 bl_12 br_12 wl_23 vdd gnd cell_6t
Xbit_r24_c12 bl_12 br_12 wl_24 vdd gnd cell_6t
Xbit_r25_c12 bl_12 br_12 wl_25 vdd gnd cell_6t
Xbit_r26_c12 bl_12 br_12 wl_26 vdd gnd cell_6t
Xbit_r27_c12 bl_12 br_12 wl_27 vdd gnd cell_6t
Xbit_r28_c12 bl_12 br_12 wl_28 vdd gnd cell_6t
Xbit_r29_c12 bl_12 br_12 wl_29 vdd gnd cell_6t
Xbit_r30_c12 bl_12 br_12 wl_30 vdd gnd cell_6t
Xbit_r31_c12 bl_12 br_12 wl_31 vdd gnd cell_6t
Xbit_r32_c12 bl_12 br_12 wl_32 vdd gnd cell_6t
Xbit_r33_c12 bl_12 br_12 wl_33 vdd gnd cell_6t
Xbit_r34_c12 bl_12 br_12 wl_34 vdd gnd cell_6t
Xbit_r35_c12 bl_12 br_12 wl_35 vdd gnd cell_6t
Xbit_r36_c12 bl_12 br_12 wl_36 vdd gnd cell_6t
Xbit_r37_c12 bl_12 br_12 wl_37 vdd gnd cell_6t
Xbit_r38_c12 bl_12 br_12 wl_38 vdd gnd cell_6t
Xbit_r39_c12 bl_12 br_12 wl_39 vdd gnd cell_6t
Xbit_r40_c12 bl_12 br_12 wl_40 vdd gnd cell_6t
Xbit_r41_c12 bl_12 br_12 wl_41 vdd gnd cell_6t
Xbit_r42_c12 bl_12 br_12 wl_42 vdd gnd cell_6t
Xbit_r43_c12 bl_12 br_12 wl_43 vdd gnd cell_6t
Xbit_r44_c12 bl_12 br_12 wl_44 vdd gnd cell_6t
Xbit_r45_c12 bl_12 br_12 wl_45 vdd gnd cell_6t
Xbit_r46_c12 bl_12 br_12 wl_46 vdd gnd cell_6t
Xbit_r47_c12 bl_12 br_12 wl_47 vdd gnd cell_6t
Xbit_r48_c12 bl_12 br_12 wl_48 vdd gnd cell_6t
Xbit_r49_c12 bl_12 br_12 wl_49 vdd gnd cell_6t
Xbit_r50_c12 bl_12 br_12 wl_50 vdd gnd cell_6t
Xbit_r51_c12 bl_12 br_12 wl_51 vdd gnd cell_6t
Xbit_r52_c12 bl_12 br_12 wl_52 vdd gnd cell_6t
Xbit_r53_c12 bl_12 br_12 wl_53 vdd gnd cell_6t
Xbit_r54_c12 bl_12 br_12 wl_54 vdd gnd cell_6t
Xbit_r55_c12 bl_12 br_12 wl_55 vdd gnd cell_6t
Xbit_r56_c12 bl_12 br_12 wl_56 vdd gnd cell_6t
Xbit_r57_c12 bl_12 br_12 wl_57 vdd gnd cell_6t
Xbit_r58_c12 bl_12 br_12 wl_58 vdd gnd cell_6t
Xbit_r59_c12 bl_12 br_12 wl_59 vdd gnd cell_6t
Xbit_r60_c12 bl_12 br_12 wl_60 vdd gnd cell_6t
Xbit_r61_c12 bl_12 br_12 wl_61 vdd gnd cell_6t
Xbit_r62_c12 bl_12 br_12 wl_62 vdd gnd cell_6t
Xbit_r63_c12 bl_12 br_12 wl_63 vdd gnd cell_6t
Xbit_r64_c12 bl_12 br_12 wl_64 vdd gnd cell_6t
Xbit_r65_c12 bl_12 br_12 wl_65 vdd gnd cell_6t
Xbit_r66_c12 bl_12 br_12 wl_66 vdd gnd cell_6t
Xbit_r67_c12 bl_12 br_12 wl_67 vdd gnd cell_6t
Xbit_r68_c12 bl_12 br_12 wl_68 vdd gnd cell_6t
Xbit_r69_c12 bl_12 br_12 wl_69 vdd gnd cell_6t
Xbit_r70_c12 bl_12 br_12 wl_70 vdd gnd cell_6t
Xbit_r71_c12 bl_12 br_12 wl_71 vdd gnd cell_6t
Xbit_r72_c12 bl_12 br_12 wl_72 vdd gnd cell_6t
Xbit_r73_c12 bl_12 br_12 wl_73 vdd gnd cell_6t
Xbit_r74_c12 bl_12 br_12 wl_74 vdd gnd cell_6t
Xbit_r75_c12 bl_12 br_12 wl_75 vdd gnd cell_6t
Xbit_r76_c12 bl_12 br_12 wl_76 vdd gnd cell_6t
Xbit_r77_c12 bl_12 br_12 wl_77 vdd gnd cell_6t
Xbit_r78_c12 bl_12 br_12 wl_78 vdd gnd cell_6t
Xbit_r79_c12 bl_12 br_12 wl_79 vdd gnd cell_6t
Xbit_r80_c12 bl_12 br_12 wl_80 vdd gnd cell_6t
Xbit_r81_c12 bl_12 br_12 wl_81 vdd gnd cell_6t
Xbit_r82_c12 bl_12 br_12 wl_82 vdd gnd cell_6t
Xbit_r83_c12 bl_12 br_12 wl_83 vdd gnd cell_6t
Xbit_r84_c12 bl_12 br_12 wl_84 vdd gnd cell_6t
Xbit_r85_c12 bl_12 br_12 wl_85 vdd gnd cell_6t
Xbit_r86_c12 bl_12 br_12 wl_86 vdd gnd cell_6t
Xbit_r87_c12 bl_12 br_12 wl_87 vdd gnd cell_6t
Xbit_r88_c12 bl_12 br_12 wl_88 vdd gnd cell_6t
Xbit_r89_c12 bl_12 br_12 wl_89 vdd gnd cell_6t
Xbit_r90_c12 bl_12 br_12 wl_90 vdd gnd cell_6t
Xbit_r91_c12 bl_12 br_12 wl_91 vdd gnd cell_6t
Xbit_r92_c12 bl_12 br_12 wl_92 vdd gnd cell_6t
Xbit_r93_c12 bl_12 br_12 wl_93 vdd gnd cell_6t
Xbit_r94_c12 bl_12 br_12 wl_94 vdd gnd cell_6t
Xbit_r95_c12 bl_12 br_12 wl_95 vdd gnd cell_6t
Xbit_r96_c12 bl_12 br_12 wl_96 vdd gnd cell_6t
Xbit_r97_c12 bl_12 br_12 wl_97 vdd gnd cell_6t
Xbit_r98_c12 bl_12 br_12 wl_98 vdd gnd cell_6t
Xbit_r99_c12 bl_12 br_12 wl_99 vdd gnd cell_6t
Xbit_r100_c12 bl_12 br_12 wl_100 vdd gnd cell_6t
Xbit_r101_c12 bl_12 br_12 wl_101 vdd gnd cell_6t
Xbit_r102_c12 bl_12 br_12 wl_102 vdd gnd cell_6t
Xbit_r103_c12 bl_12 br_12 wl_103 vdd gnd cell_6t
Xbit_r104_c12 bl_12 br_12 wl_104 vdd gnd cell_6t
Xbit_r105_c12 bl_12 br_12 wl_105 vdd gnd cell_6t
Xbit_r106_c12 bl_12 br_12 wl_106 vdd gnd cell_6t
Xbit_r107_c12 bl_12 br_12 wl_107 vdd gnd cell_6t
Xbit_r108_c12 bl_12 br_12 wl_108 vdd gnd cell_6t
Xbit_r109_c12 bl_12 br_12 wl_109 vdd gnd cell_6t
Xbit_r110_c12 bl_12 br_12 wl_110 vdd gnd cell_6t
Xbit_r111_c12 bl_12 br_12 wl_111 vdd gnd cell_6t
Xbit_r112_c12 bl_12 br_12 wl_112 vdd gnd cell_6t
Xbit_r113_c12 bl_12 br_12 wl_113 vdd gnd cell_6t
Xbit_r114_c12 bl_12 br_12 wl_114 vdd gnd cell_6t
Xbit_r115_c12 bl_12 br_12 wl_115 vdd gnd cell_6t
Xbit_r116_c12 bl_12 br_12 wl_116 vdd gnd cell_6t
Xbit_r117_c12 bl_12 br_12 wl_117 vdd gnd cell_6t
Xbit_r118_c12 bl_12 br_12 wl_118 vdd gnd cell_6t
Xbit_r119_c12 bl_12 br_12 wl_119 vdd gnd cell_6t
Xbit_r120_c12 bl_12 br_12 wl_120 vdd gnd cell_6t
Xbit_r121_c12 bl_12 br_12 wl_121 vdd gnd cell_6t
Xbit_r122_c12 bl_12 br_12 wl_122 vdd gnd cell_6t
Xbit_r123_c12 bl_12 br_12 wl_123 vdd gnd cell_6t
Xbit_r124_c12 bl_12 br_12 wl_124 vdd gnd cell_6t
Xbit_r125_c12 bl_12 br_12 wl_125 vdd gnd cell_6t
Xbit_r126_c12 bl_12 br_12 wl_126 vdd gnd cell_6t
Xbit_r127_c12 bl_12 br_12 wl_127 vdd gnd cell_6t
Xbit_r128_c12 bl_12 br_12 wl_128 vdd gnd cell_6t
Xbit_r129_c12 bl_12 br_12 wl_129 vdd gnd cell_6t
Xbit_r130_c12 bl_12 br_12 wl_130 vdd gnd cell_6t
Xbit_r131_c12 bl_12 br_12 wl_131 vdd gnd cell_6t
Xbit_r132_c12 bl_12 br_12 wl_132 vdd gnd cell_6t
Xbit_r133_c12 bl_12 br_12 wl_133 vdd gnd cell_6t
Xbit_r134_c12 bl_12 br_12 wl_134 vdd gnd cell_6t
Xbit_r135_c12 bl_12 br_12 wl_135 vdd gnd cell_6t
Xbit_r136_c12 bl_12 br_12 wl_136 vdd gnd cell_6t
Xbit_r137_c12 bl_12 br_12 wl_137 vdd gnd cell_6t
Xbit_r138_c12 bl_12 br_12 wl_138 vdd gnd cell_6t
Xbit_r139_c12 bl_12 br_12 wl_139 vdd gnd cell_6t
Xbit_r140_c12 bl_12 br_12 wl_140 vdd gnd cell_6t
Xbit_r141_c12 bl_12 br_12 wl_141 vdd gnd cell_6t
Xbit_r142_c12 bl_12 br_12 wl_142 vdd gnd cell_6t
Xbit_r143_c12 bl_12 br_12 wl_143 vdd gnd cell_6t
Xbit_r144_c12 bl_12 br_12 wl_144 vdd gnd cell_6t
Xbit_r145_c12 bl_12 br_12 wl_145 vdd gnd cell_6t
Xbit_r146_c12 bl_12 br_12 wl_146 vdd gnd cell_6t
Xbit_r147_c12 bl_12 br_12 wl_147 vdd gnd cell_6t
Xbit_r148_c12 bl_12 br_12 wl_148 vdd gnd cell_6t
Xbit_r149_c12 bl_12 br_12 wl_149 vdd gnd cell_6t
Xbit_r150_c12 bl_12 br_12 wl_150 vdd gnd cell_6t
Xbit_r151_c12 bl_12 br_12 wl_151 vdd gnd cell_6t
Xbit_r152_c12 bl_12 br_12 wl_152 vdd gnd cell_6t
Xbit_r153_c12 bl_12 br_12 wl_153 vdd gnd cell_6t
Xbit_r154_c12 bl_12 br_12 wl_154 vdd gnd cell_6t
Xbit_r155_c12 bl_12 br_12 wl_155 vdd gnd cell_6t
Xbit_r156_c12 bl_12 br_12 wl_156 vdd gnd cell_6t
Xbit_r157_c12 bl_12 br_12 wl_157 vdd gnd cell_6t
Xbit_r158_c12 bl_12 br_12 wl_158 vdd gnd cell_6t
Xbit_r159_c12 bl_12 br_12 wl_159 vdd gnd cell_6t
Xbit_r160_c12 bl_12 br_12 wl_160 vdd gnd cell_6t
Xbit_r161_c12 bl_12 br_12 wl_161 vdd gnd cell_6t
Xbit_r162_c12 bl_12 br_12 wl_162 vdd gnd cell_6t
Xbit_r163_c12 bl_12 br_12 wl_163 vdd gnd cell_6t
Xbit_r164_c12 bl_12 br_12 wl_164 vdd gnd cell_6t
Xbit_r165_c12 bl_12 br_12 wl_165 vdd gnd cell_6t
Xbit_r166_c12 bl_12 br_12 wl_166 vdd gnd cell_6t
Xbit_r167_c12 bl_12 br_12 wl_167 vdd gnd cell_6t
Xbit_r168_c12 bl_12 br_12 wl_168 vdd gnd cell_6t
Xbit_r169_c12 bl_12 br_12 wl_169 vdd gnd cell_6t
Xbit_r170_c12 bl_12 br_12 wl_170 vdd gnd cell_6t
Xbit_r171_c12 bl_12 br_12 wl_171 vdd gnd cell_6t
Xbit_r172_c12 bl_12 br_12 wl_172 vdd gnd cell_6t
Xbit_r173_c12 bl_12 br_12 wl_173 vdd gnd cell_6t
Xbit_r174_c12 bl_12 br_12 wl_174 vdd gnd cell_6t
Xbit_r175_c12 bl_12 br_12 wl_175 vdd gnd cell_6t
Xbit_r176_c12 bl_12 br_12 wl_176 vdd gnd cell_6t
Xbit_r177_c12 bl_12 br_12 wl_177 vdd gnd cell_6t
Xbit_r178_c12 bl_12 br_12 wl_178 vdd gnd cell_6t
Xbit_r179_c12 bl_12 br_12 wl_179 vdd gnd cell_6t
Xbit_r180_c12 bl_12 br_12 wl_180 vdd gnd cell_6t
Xbit_r181_c12 bl_12 br_12 wl_181 vdd gnd cell_6t
Xbit_r182_c12 bl_12 br_12 wl_182 vdd gnd cell_6t
Xbit_r183_c12 bl_12 br_12 wl_183 vdd gnd cell_6t
Xbit_r184_c12 bl_12 br_12 wl_184 vdd gnd cell_6t
Xbit_r185_c12 bl_12 br_12 wl_185 vdd gnd cell_6t
Xbit_r186_c12 bl_12 br_12 wl_186 vdd gnd cell_6t
Xbit_r187_c12 bl_12 br_12 wl_187 vdd gnd cell_6t
Xbit_r188_c12 bl_12 br_12 wl_188 vdd gnd cell_6t
Xbit_r189_c12 bl_12 br_12 wl_189 vdd gnd cell_6t
Xbit_r190_c12 bl_12 br_12 wl_190 vdd gnd cell_6t
Xbit_r191_c12 bl_12 br_12 wl_191 vdd gnd cell_6t
Xbit_r192_c12 bl_12 br_12 wl_192 vdd gnd cell_6t
Xbit_r193_c12 bl_12 br_12 wl_193 vdd gnd cell_6t
Xbit_r194_c12 bl_12 br_12 wl_194 vdd gnd cell_6t
Xbit_r195_c12 bl_12 br_12 wl_195 vdd gnd cell_6t
Xbit_r196_c12 bl_12 br_12 wl_196 vdd gnd cell_6t
Xbit_r197_c12 bl_12 br_12 wl_197 vdd gnd cell_6t
Xbit_r198_c12 bl_12 br_12 wl_198 vdd gnd cell_6t
Xbit_r199_c12 bl_12 br_12 wl_199 vdd gnd cell_6t
Xbit_r200_c12 bl_12 br_12 wl_200 vdd gnd cell_6t
Xbit_r201_c12 bl_12 br_12 wl_201 vdd gnd cell_6t
Xbit_r202_c12 bl_12 br_12 wl_202 vdd gnd cell_6t
Xbit_r203_c12 bl_12 br_12 wl_203 vdd gnd cell_6t
Xbit_r204_c12 bl_12 br_12 wl_204 vdd gnd cell_6t
Xbit_r205_c12 bl_12 br_12 wl_205 vdd gnd cell_6t
Xbit_r206_c12 bl_12 br_12 wl_206 vdd gnd cell_6t
Xbit_r207_c12 bl_12 br_12 wl_207 vdd gnd cell_6t
Xbit_r208_c12 bl_12 br_12 wl_208 vdd gnd cell_6t
Xbit_r209_c12 bl_12 br_12 wl_209 vdd gnd cell_6t
Xbit_r210_c12 bl_12 br_12 wl_210 vdd gnd cell_6t
Xbit_r211_c12 bl_12 br_12 wl_211 vdd gnd cell_6t
Xbit_r212_c12 bl_12 br_12 wl_212 vdd gnd cell_6t
Xbit_r213_c12 bl_12 br_12 wl_213 vdd gnd cell_6t
Xbit_r214_c12 bl_12 br_12 wl_214 vdd gnd cell_6t
Xbit_r215_c12 bl_12 br_12 wl_215 vdd gnd cell_6t
Xbit_r216_c12 bl_12 br_12 wl_216 vdd gnd cell_6t
Xbit_r217_c12 bl_12 br_12 wl_217 vdd gnd cell_6t
Xbit_r218_c12 bl_12 br_12 wl_218 vdd gnd cell_6t
Xbit_r219_c12 bl_12 br_12 wl_219 vdd gnd cell_6t
Xbit_r220_c12 bl_12 br_12 wl_220 vdd gnd cell_6t
Xbit_r221_c12 bl_12 br_12 wl_221 vdd gnd cell_6t
Xbit_r222_c12 bl_12 br_12 wl_222 vdd gnd cell_6t
Xbit_r223_c12 bl_12 br_12 wl_223 vdd gnd cell_6t
Xbit_r224_c12 bl_12 br_12 wl_224 vdd gnd cell_6t
Xbit_r225_c12 bl_12 br_12 wl_225 vdd gnd cell_6t
Xbit_r226_c12 bl_12 br_12 wl_226 vdd gnd cell_6t
Xbit_r227_c12 bl_12 br_12 wl_227 vdd gnd cell_6t
Xbit_r228_c12 bl_12 br_12 wl_228 vdd gnd cell_6t
Xbit_r229_c12 bl_12 br_12 wl_229 vdd gnd cell_6t
Xbit_r230_c12 bl_12 br_12 wl_230 vdd gnd cell_6t
Xbit_r231_c12 bl_12 br_12 wl_231 vdd gnd cell_6t
Xbit_r232_c12 bl_12 br_12 wl_232 vdd gnd cell_6t
Xbit_r233_c12 bl_12 br_12 wl_233 vdd gnd cell_6t
Xbit_r234_c12 bl_12 br_12 wl_234 vdd gnd cell_6t
Xbit_r235_c12 bl_12 br_12 wl_235 vdd gnd cell_6t
Xbit_r236_c12 bl_12 br_12 wl_236 vdd gnd cell_6t
Xbit_r237_c12 bl_12 br_12 wl_237 vdd gnd cell_6t
Xbit_r238_c12 bl_12 br_12 wl_238 vdd gnd cell_6t
Xbit_r239_c12 bl_12 br_12 wl_239 vdd gnd cell_6t
Xbit_r240_c12 bl_12 br_12 wl_240 vdd gnd cell_6t
Xbit_r241_c12 bl_12 br_12 wl_241 vdd gnd cell_6t
Xbit_r242_c12 bl_12 br_12 wl_242 vdd gnd cell_6t
Xbit_r243_c12 bl_12 br_12 wl_243 vdd gnd cell_6t
Xbit_r244_c12 bl_12 br_12 wl_244 vdd gnd cell_6t
Xbit_r245_c12 bl_12 br_12 wl_245 vdd gnd cell_6t
Xbit_r246_c12 bl_12 br_12 wl_246 vdd gnd cell_6t
Xbit_r247_c12 bl_12 br_12 wl_247 vdd gnd cell_6t
Xbit_r248_c12 bl_12 br_12 wl_248 vdd gnd cell_6t
Xbit_r249_c12 bl_12 br_12 wl_249 vdd gnd cell_6t
Xbit_r250_c12 bl_12 br_12 wl_250 vdd gnd cell_6t
Xbit_r251_c12 bl_12 br_12 wl_251 vdd gnd cell_6t
Xbit_r252_c12 bl_12 br_12 wl_252 vdd gnd cell_6t
Xbit_r253_c12 bl_12 br_12 wl_253 vdd gnd cell_6t
Xbit_r254_c12 bl_12 br_12 wl_254 vdd gnd cell_6t
Xbit_r255_c12 bl_12 br_12 wl_255 vdd gnd cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd cell_6t
Xbit_r1_c13 bl_13 br_13 wl_1 vdd gnd cell_6t
Xbit_r2_c13 bl_13 br_13 wl_2 vdd gnd cell_6t
Xbit_r3_c13 bl_13 br_13 wl_3 vdd gnd cell_6t
Xbit_r4_c13 bl_13 br_13 wl_4 vdd gnd cell_6t
Xbit_r5_c13 bl_13 br_13 wl_5 vdd gnd cell_6t
Xbit_r6_c13 bl_13 br_13 wl_6 vdd gnd cell_6t
Xbit_r7_c13 bl_13 br_13 wl_7 vdd gnd cell_6t
Xbit_r8_c13 bl_13 br_13 wl_8 vdd gnd cell_6t
Xbit_r9_c13 bl_13 br_13 wl_9 vdd gnd cell_6t
Xbit_r10_c13 bl_13 br_13 wl_10 vdd gnd cell_6t
Xbit_r11_c13 bl_13 br_13 wl_11 vdd gnd cell_6t
Xbit_r12_c13 bl_13 br_13 wl_12 vdd gnd cell_6t
Xbit_r13_c13 bl_13 br_13 wl_13 vdd gnd cell_6t
Xbit_r14_c13 bl_13 br_13 wl_14 vdd gnd cell_6t
Xbit_r15_c13 bl_13 br_13 wl_15 vdd gnd cell_6t
Xbit_r16_c13 bl_13 br_13 wl_16 vdd gnd cell_6t
Xbit_r17_c13 bl_13 br_13 wl_17 vdd gnd cell_6t
Xbit_r18_c13 bl_13 br_13 wl_18 vdd gnd cell_6t
Xbit_r19_c13 bl_13 br_13 wl_19 vdd gnd cell_6t
Xbit_r20_c13 bl_13 br_13 wl_20 vdd gnd cell_6t
Xbit_r21_c13 bl_13 br_13 wl_21 vdd gnd cell_6t
Xbit_r22_c13 bl_13 br_13 wl_22 vdd gnd cell_6t
Xbit_r23_c13 bl_13 br_13 wl_23 vdd gnd cell_6t
Xbit_r24_c13 bl_13 br_13 wl_24 vdd gnd cell_6t
Xbit_r25_c13 bl_13 br_13 wl_25 vdd gnd cell_6t
Xbit_r26_c13 bl_13 br_13 wl_26 vdd gnd cell_6t
Xbit_r27_c13 bl_13 br_13 wl_27 vdd gnd cell_6t
Xbit_r28_c13 bl_13 br_13 wl_28 vdd gnd cell_6t
Xbit_r29_c13 bl_13 br_13 wl_29 vdd gnd cell_6t
Xbit_r30_c13 bl_13 br_13 wl_30 vdd gnd cell_6t
Xbit_r31_c13 bl_13 br_13 wl_31 vdd gnd cell_6t
Xbit_r32_c13 bl_13 br_13 wl_32 vdd gnd cell_6t
Xbit_r33_c13 bl_13 br_13 wl_33 vdd gnd cell_6t
Xbit_r34_c13 bl_13 br_13 wl_34 vdd gnd cell_6t
Xbit_r35_c13 bl_13 br_13 wl_35 vdd gnd cell_6t
Xbit_r36_c13 bl_13 br_13 wl_36 vdd gnd cell_6t
Xbit_r37_c13 bl_13 br_13 wl_37 vdd gnd cell_6t
Xbit_r38_c13 bl_13 br_13 wl_38 vdd gnd cell_6t
Xbit_r39_c13 bl_13 br_13 wl_39 vdd gnd cell_6t
Xbit_r40_c13 bl_13 br_13 wl_40 vdd gnd cell_6t
Xbit_r41_c13 bl_13 br_13 wl_41 vdd gnd cell_6t
Xbit_r42_c13 bl_13 br_13 wl_42 vdd gnd cell_6t
Xbit_r43_c13 bl_13 br_13 wl_43 vdd gnd cell_6t
Xbit_r44_c13 bl_13 br_13 wl_44 vdd gnd cell_6t
Xbit_r45_c13 bl_13 br_13 wl_45 vdd gnd cell_6t
Xbit_r46_c13 bl_13 br_13 wl_46 vdd gnd cell_6t
Xbit_r47_c13 bl_13 br_13 wl_47 vdd gnd cell_6t
Xbit_r48_c13 bl_13 br_13 wl_48 vdd gnd cell_6t
Xbit_r49_c13 bl_13 br_13 wl_49 vdd gnd cell_6t
Xbit_r50_c13 bl_13 br_13 wl_50 vdd gnd cell_6t
Xbit_r51_c13 bl_13 br_13 wl_51 vdd gnd cell_6t
Xbit_r52_c13 bl_13 br_13 wl_52 vdd gnd cell_6t
Xbit_r53_c13 bl_13 br_13 wl_53 vdd gnd cell_6t
Xbit_r54_c13 bl_13 br_13 wl_54 vdd gnd cell_6t
Xbit_r55_c13 bl_13 br_13 wl_55 vdd gnd cell_6t
Xbit_r56_c13 bl_13 br_13 wl_56 vdd gnd cell_6t
Xbit_r57_c13 bl_13 br_13 wl_57 vdd gnd cell_6t
Xbit_r58_c13 bl_13 br_13 wl_58 vdd gnd cell_6t
Xbit_r59_c13 bl_13 br_13 wl_59 vdd gnd cell_6t
Xbit_r60_c13 bl_13 br_13 wl_60 vdd gnd cell_6t
Xbit_r61_c13 bl_13 br_13 wl_61 vdd gnd cell_6t
Xbit_r62_c13 bl_13 br_13 wl_62 vdd gnd cell_6t
Xbit_r63_c13 bl_13 br_13 wl_63 vdd gnd cell_6t
Xbit_r64_c13 bl_13 br_13 wl_64 vdd gnd cell_6t
Xbit_r65_c13 bl_13 br_13 wl_65 vdd gnd cell_6t
Xbit_r66_c13 bl_13 br_13 wl_66 vdd gnd cell_6t
Xbit_r67_c13 bl_13 br_13 wl_67 vdd gnd cell_6t
Xbit_r68_c13 bl_13 br_13 wl_68 vdd gnd cell_6t
Xbit_r69_c13 bl_13 br_13 wl_69 vdd gnd cell_6t
Xbit_r70_c13 bl_13 br_13 wl_70 vdd gnd cell_6t
Xbit_r71_c13 bl_13 br_13 wl_71 vdd gnd cell_6t
Xbit_r72_c13 bl_13 br_13 wl_72 vdd gnd cell_6t
Xbit_r73_c13 bl_13 br_13 wl_73 vdd gnd cell_6t
Xbit_r74_c13 bl_13 br_13 wl_74 vdd gnd cell_6t
Xbit_r75_c13 bl_13 br_13 wl_75 vdd gnd cell_6t
Xbit_r76_c13 bl_13 br_13 wl_76 vdd gnd cell_6t
Xbit_r77_c13 bl_13 br_13 wl_77 vdd gnd cell_6t
Xbit_r78_c13 bl_13 br_13 wl_78 vdd gnd cell_6t
Xbit_r79_c13 bl_13 br_13 wl_79 vdd gnd cell_6t
Xbit_r80_c13 bl_13 br_13 wl_80 vdd gnd cell_6t
Xbit_r81_c13 bl_13 br_13 wl_81 vdd gnd cell_6t
Xbit_r82_c13 bl_13 br_13 wl_82 vdd gnd cell_6t
Xbit_r83_c13 bl_13 br_13 wl_83 vdd gnd cell_6t
Xbit_r84_c13 bl_13 br_13 wl_84 vdd gnd cell_6t
Xbit_r85_c13 bl_13 br_13 wl_85 vdd gnd cell_6t
Xbit_r86_c13 bl_13 br_13 wl_86 vdd gnd cell_6t
Xbit_r87_c13 bl_13 br_13 wl_87 vdd gnd cell_6t
Xbit_r88_c13 bl_13 br_13 wl_88 vdd gnd cell_6t
Xbit_r89_c13 bl_13 br_13 wl_89 vdd gnd cell_6t
Xbit_r90_c13 bl_13 br_13 wl_90 vdd gnd cell_6t
Xbit_r91_c13 bl_13 br_13 wl_91 vdd gnd cell_6t
Xbit_r92_c13 bl_13 br_13 wl_92 vdd gnd cell_6t
Xbit_r93_c13 bl_13 br_13 wl_93 vdd gnd cell_6t
Xbit_r94_c13 bl_13 br_13 wl_94 vdd gnd cell_6t
Xbit_r95_c13 bl_13 br_13 wl_95 vdd gnd cell_6t
Xbit_r96_c13 bl_13 br_13 wl_96 vdd gnd cell_6t
Xbit_r97_c13 bl_13 br_13 wl_97 vdd gnd cell_6t
Xbit_r98_c13 bl_13 br_13 wl_98 vdd gnd cell_6t
Xbit_r99_c13 bl_13 br_13 wl_99 vdd gnd cell_6t
Xbit_r100_c13 bl_13 br_13 wl_100 vdd gnd cell_6t
Xbit_r101_c13 bl_13 br_13 wl_101 vdd gnd cell_6t
Xbit_r102_c13 bl_13 br_13 wl_102 vdd gnd cell_6t
Xbit_r103_c13 bl_13 br_13 wl_103 vdd gnd cell_6t
Xbit_r104_c13 bl_13 br_13 wl_104 vdd gnd cell_6t
Xbit_r105_c13 bl_13 br_13 wl_105 vdd gnd cell_6t
Xbit_r106_c13 bl_13 br_13 wl_106 vdd gnd cell_6t
Xbit_r107_c13 bl_13 br_13 wl_107 vdd gnd cell_6t
Xbit_r108_c13 bl_13 br_13 wl_108 vdd gnd cell_6t
Xbit_r109_c13 bl_13 br_13 wl_109 vdd gnd cell_6t
Xbit_r110_c13 bl_13 br_13 wl_110 vdd gnd cell_6t
Xbit_r111_c13 bl_13 br_13 wl_111 vdd gnd cell_6t
Xbit_r112_c13 bl_13 br_13 wl_112 vdd gnd cell_6t
Xbit_r113_c13 bl_13 br_13 wl_113 vdd gnd cell_6t
Xbit_r114_c13 bl_13 br_13 wl_114 vdd gnd cell_6t
Xbit_r115_c13 bl_13 br_13 wl_115 vdd gnd cell_6t
Xbit_r116_c13 bl_13 br_13 wl_116 vdd gnd cell_6t
Xbit_r117_c13 bl_13 br_13 wl_117 vdd gnd cell_6t
Xbit_r118_c13 bl_13 br_13 wl_118 vdd gnd cell_6t
Xbit_r119_c13 bl_13 br_13 wl_119 vdd gnd cell_6t
Xbit_r120_c13 bl_13 br_13 wl_120 vdd gnd cell_6t
Xbit_r121_c13 bl_13 br_13 wl_121 vdd gnd cell_6t
Xbit_r122_c13 bl_13 br_13 wl_122 vdd gnd cell_6t
Xbit_r123_c13 bl_13 br_13 wl_123 vdd gnd cell_6t
Xbit_r124_c13 bl_13 br_13 wl_124 vdd gnd cell_6t
Xbit_r125_c13 bl_13 br_13 wl_125 vdd gnd cell_6t
Xbit_r126_c13 bl_13 br_13 wl_126 vdd gnd cell_6t
Xbit_r127_c13 bl_13 br_13 wl_127 vdd gnd cell_6t
Xbit_r128_c13 bl_13 br_13 wl_128 vdd gnd cell_6t
Xbit_r129_c13 bl_13 br_13 wl_129 vdd gnd cell_6t
Xbit_r130_c13 bl_13 br_13 wl_130 vdd gnd cell_6t
Xbit_r131_c13 bl_13 br_13 wl_131 vdd gnd cell_6t
Xbit_r132_c13 bl_13 br_13 wl_132 vdd gnd cell_6t
Xbit_r133_c13 bl_13 br_13 wl_133 vdd gnd cell_6t
Xbit_r134_c13 bl_13 br_13 wl_134 vdd gnd cell_6t
Xbit_r135_c13 bl_13 br_13 wl_135 vdd gnd cell_6t
Xbit_r136_c13 bl_13 br_13 wl_136 vdd gnd cell_6t
Xbit_r137_c13 bl_13 br_13 wl_137 vdd gnd cell_6t
Xbit_r138_c13 bl_13 br_13 wl_138 vdd gnd cell_6t
Xbit_r139_c13 bl_13 br_13 wl_139 vdd gnd cell_6t
Xbit_r140_c13 bl_13 br_13 wl_140 vdd gnd cell_6t
Xbit_r141_c13 bl_13 br_13 wl_141 vdd gnd cell_6t
Xbit_r142_c13 bl_13 br_13 wl_142 vdd gnd cell_6t
Xbit_r143_c13 bl_13 br_13 wl_143 vdd gnd cell_6t
Xbit_r144_c13 bl_13 br_13 wl_144 vdd gnd cell_6t
Xbit_r145_c13 bl_13 br_13 wl_145 vdd gnd cell_6t
Xbit_r146_c13 bl_13 br_13 wl_146 vdd gnd cell_6t
Xbit_r147_c13 bl_13 br_13 wl_147 vdd gnd cell_6t
Xbit_r148_c13 bl_13 br_13 wl_148 vdd gnd cell_6t
Xbit_r149_c13 bl_13 br_13 wl_149 vdd gnd cell_6t
Xbit_r150_c13 bl_13 br_13 wl_150 vdd gnd cell_6t
Xbit_r151_c13 bl_13 br_13 wl_151 vdd gnd cell_6t
Xbit_r152_c13 bl_13 br_13 wl_152 vdd gnd cell_6t
Xbit_r153_c13 bl_13 br_13 wl_153 vdd gnd cell_6t
Xbit_r154_c13 bl_13 br_13 wl_154 vdd gnd cell_6t
Xbit_r155_c13 bl_13 br_13 wl_155 vdd gnd cell_6t
Xbit_r156_c13 bl_13 br_13 wl_156 vdd gnd cell_6t
Xbit_r157_c13 bl_13 br_13 wl_157 vdd gnd cell_6t
Xbit_r158_c13 bl_13 br_13 wl_158 vdd gnd cell_6t
Xbit_r159_c13 bl_13 br_13 wl_159 vdd gnd cell_6t
Xbit_r160_c13 bl_13 br_13 wl_160 vdd gnd cell_6t
Xbit_r161_c13 bl_13 br_13 wl_161 vdd gnd cell_6t
Xbit_r162_c13 bl_13 br_13 wl_162 vdd gnd cell_6t
Xbit_r163_c13 bl_13 br_13 wl_163 vdd gnd cell_6t
Xbit_r164_c13 bl_13 br_13 wl_164 vdd gnd cell_6t
Xbit_r165_c13 bl_13 br_13 wl_165 vdd gnd cell_6t
Xbit_r166_c13 bl_13 br_13 wl_166 vdd gnd cell_6t
Xbit_r167_c13 bl_13 br_13 wl_167 vdd gnd cell_6t
Xbit_r168_c13 bl_13 br_13 wl_168 vdd gnd cell_6t
Xbit_r169_c13 bl_13 br_13 wl_169 vdd gnd cell_6t
Xbit_r170_c13 bl_13 br_13 wl_170 vdd gnd cell_6t
Xbit_r171_c13 bl_13 br_13 wl_171 vdd gnd cell_6t
Xbit_r172_c13 bl_13 br_13 wl_172 vdd gnd cell_6t
Xbit_r173_c13 bl_13 br_13 wl_173 vdd gnd cell_6t
Xbit_r174_c13 bl_13 br_13 wl_174 vdd gnd cell_6t
Xbit_r175_c13 bl_13 br_13 wl_175 vdd gnd cell_6t
Xbit_r176_c13 bl_13 br_13 wl_176 vdd gnd cell_6t
Xbit_r177_c13 bl_13 br_13 wl_177 vdd gnd cell_6t
Xbit_r178_c13 bl_13 br_13 wl_178 vdd gnd cell_6t
Xbit_r179_c13 bl_13 br_13 wl_179 vdd gnd cell_6t
Xbit_r180_c13 bl_13 br_13 wl_180 vdd gnd cell_6t
Xbit_r181_c13 bl_13 br_13 wl_181 vdd gnd cell_6t
Xbit_r182_c13 bl_13 br_13 wl_182 vdd gnd cell_6t
Xbit_r183_c13 bl_13 br_13 wl_183 vdd gnd cell_6t
Xbit_r184_c13 bl_13 br_13 wl_184 vdd gnd cell_6t
Xbit_r185_c13 bl_13 br_13 wl_185 vdd gnd cell_6t
Xbit_r186_c13 bl_13 br_13 wl_186 vdd gnd cell_6t
Xbit_r187_c13 bl_13 br_13 wl_187 vdd gnd cell_6t
Xbit_r188_c13 bl_13 br_13 wl_188 vdd gnd cell_6t
Xbit_r189_c13 bl_13 br_13 wl_189 vdd gnd cell_6t
Xbit_r190_c13 bl_13 br_13 wl_190 vdd gnd cell_6t
Xbit_r191_c13 bl_13 br_13 wl_191 vdd gnd cell_6t
Xbit_r192_c13 bl_13 br_13 wl_192 vdd gnd cell_6t
Xbit_r193_c13 bl_13 br_13 wl_193 vdd gnd cell_6t
Xbit_r194_c13 bl_13 br_13 wl_194 vdd gnd cell_6t
Xbit_r195_c13 bl_13 br_13 wl_195 vdd gnd cell_6t
Xbit_r196_c13 bl_13 br_13 wl_196 vdd gnd cell_6t
Xbit_r197_c13 bl_13 br_13 wl_197 vdd gnd cell_6t
Xbit_r198_c13 bl_13 br_13 wl_198 vdd gnd cell_6t
Xbit_r199_c13 bl_13 br_13 wl_199 vdd gnd cell_6t
Xbit_r200_c13 bl_13 br_13 wl_200 vdd gnd cell_6t
Xbit_r201_c13 bl_13 br_13 wl_201 vdd gnd cell_6t
Xbit_r202_c13 bl_13 br_13 wl_202 vdd gnd cell_6t
Xbit_r203_c13 bl_13 br_13 wl_203 vdd gnd cell_6t
Xbit_r204_c13 bl_13 br_13 wl_204 vdd gnd cell_6t
Xbit_r205_c13 bl_13 br_13 wl_205 vdd gnd cell_6t
Xbit_r206_c13 bl_13 br_13 wl_206 vdd gnd cell_6t
Xbit_r207_c13 bl_13 br_13 wl_207 vdd gnd cell_6t
Xbit_r208_c13 bl_13 br_13 wl_208 vdd gnd cell_6t
Xbit_r209_c13 bl_13 br_13 wl_209 vdd gnd cell_6t
Xbit_r210_c13 bl_13 br_13 wl_210 vdd gnd cell_6t
Xbit_r211_c13 bl_13 br_13 wl_211 vdd gnd cell_6t
Xbit_r212_c13 bl_13 br_13 wl_212 vdd gnd cell_6t
Xbit_r213_c13 bl_13 br_13 wl_213 vdd gnd cell_6t
Xbit_r214_c13 bl_13 br_13 wl_214 vdd gnd cell_6t
Xbit_r215_c13 bl_13 br_13 wl_215 vdd gnd cell_6t
Xbit_r216_c13 bl_13 br_13 wl_216 vdd gnd cell_6t
Xbit_r217_c13 bl_13 br_13 wl_217 vdd gnd cell_6t
Xbit_r218_c13 bl_13 br_13 wl_218 vdd gnd cell_6t
Xbit_r219_c13 bl_13 br_13 wl_219 vdd gnd cell_6t
Xbit_r220_c13 bl_13 br_13 wl_220 vdd gnd cell_6t
Xbit_r221_c13 bl_13 br_13 wl_221 vdd gnd cell_6t
Xbit_r222_c13 bl_13 br_13 wl_222 vdd gnd cell_6t
Xbit_r223_c13 bl_13 br_13 wl_223 vdd gnd cell_6t
Xbit_r224_c13 bl_13 br_13 wl_224 vdd gnd cell_6t
Xbit_r225_c13 bl_13 br_13 wl_225 vdd gnd cell_6t
Xbit_r226_c13 bl_13 br_13 wl_226 vdd gnd cell_6t
Xbit_r227_c13 bl_13 br_13 wl_227 vdd gnd cell_6t
Xbit_r228_c13 bl_13 br_13 wl_228 vdd gnd cell_6t
Xbit_r229_c13 bl_13 br_13 wl_229 vdd gnd cell_6t
Xbit_r230_c13 bl_13 br_13 wl_230 vdd gnd cell_6t
Xbit_r231_c13 bl_13 br_13 wl_231 vdd gnd cell_6t
Xbit_r232_c13 bl_13 br_13 wl_232 vdd gnd cell_6t
Xbit_r233_c13 bl_13 br_13 wl_233 vdd gnd cell_6t
Xbit_r234_c13 bl_13 br_13 wl_234 vdd gnd cell_6t
Xbit_r235_c13 bl_13 br_13 wl_235 vdd gnd cell_6t
Xbit_r236_c13 bl_13 br_13 wl_236 vdd gnd cell_6t
Xbit_r237_c13 bl_13 br_13 wl_237 vdd gnd cell_6t
Xbit_r238_c13 bl_13 br_13 wl_238 vdd gnd cell_6t
Xbit_r239_c13 bl_13 br_13 wl_239 vdd gnd cell_6t
Xbit_r240_c13 bl_13 br_13 wl_240 vdd gnd cell_6t
Xbit_r241_c13 bl_13 br_13 wl_241 vdd gnd cell_6t
Xbit_r242_c13 bl_13 br_13 wl_242 vdd gnd cell_6t
Xbit_r243_c13 bl_13 br_13 wl_243 vdd gnd cell_6t
Xbit_r244_c13 bl_13 br_13 wl_244 vdd gnd cell_6t
Xbit_r245_c13 bl_13 br_13 wl_245 vdd gnd cell_6t
Xbit_r246_c13 bl_13 br_13 wl_246 vdd gnd cell_6t
Xbit_r247_c13 bl_13 br_13 wl_247 vdd gnd cell_6t
Xbit_r248_c13 bl_13 br_13 wl_248 vdd gnd cell_6t
Xbit_r249_c13 bl_13 br_13 wl_249 vdd gnd cell_6t
Xbit_r250_c13 bl_13 br_13 wl_250 vdd gnd cell_6t
Xbit_r251_c13 bl_13 br_13 wl_251 vdd gnd cell_6t
Xbit_r252_c13 bl_13 br_13 wl_252 vdd gnd cell_6t
Xbit_r253_c13 bl_13 br_13 wl_253 vdd gnd cell_6t
Xbit_r254_c13 bl_13 br_13 wl_254 vdd gnd cell_6t
Xbit_r255_c13 bl_13 br_13 wl_255 vdd gnd cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd cell_6t
Xbit_r1_c14 bl_14 br_14 wl_1 vdd gnd cell_6t
Xbit_r2_c14 bl_14 br_14 wl_2 vdd gnd cell_6t
Xbit_r3_c14 bl_14 br_14 wl_3 vdd gnd cell_6t
Xbit_r4_c14 bl_14 br_14 wl_4 vdd gnd cell_6t
Xbit_r5_c14 bl_14 br_14 wl_5 vdd gnd cell_6t
Xbit_r6_c14 bl_14 br_14 wl_6 vdd gnd cell_6t
Xbit_r7_c14 bl_14 br_14 wl_7 vdd gnd cell_6t
Xbit_r8_c14 bl_14 br_14 wl_8 vdd gnd cell_6t
Xbit_r9_c14 bl_14 br_14 wl_9 vdd gnd cell_6t
Xbit_r10_c14 bl_14 br_14 wl_10 vdd gnd cell_6t
Xbit_r11_c14 bl_14 br_14 wl_11 vdd gnd cell_6t
Xbit_r12_c14 bl_14 br_14 wl_12 vdd gnd cell_6t
Xbit_r13_c14 bl_14 br_14 wl_13 vdd gnd cell_6t
Xbit_r14_c14 bl_14 br_14 wl_14 vdd gnd cell_6t
Xbit_r15_c14 bl_14 br_14 wl_15 vdd gnd cell_6t
Xbit_r16_c14 bl_14 br_14 wl_16 vdd gnd cell_6t
Xbit_r17_c14 bl_14 br_14 wl_17 vdd gnd cell_6t
Xbit_r18_c14 bl_14 br_14 wl_18 vdd gnd cell_6t
Xbit_r19_c14 bl_14 br_14 wl_19 vdd gnd cell_6t
Xbit_r20_c14 bl_14 br_14 wl_20 vdd gnd cell_6t
Xbit_r21_c14 bl_14 br_14 wl_21 vdd gnd cell_6t
Xbit_r22_c14 bl_14 br_14 wl_22 vdd gnd cell_6t
Xbit_r23_c14 bl_14 br_14 wl_23 vdd gnd cell_6t
Xbit_r24_c14 bl_14 br_14 wl_24 vdd gnd cell_6t
Xbit_r25_c14 bl_14 br_14 wl_25 vdd gnd cell_6t
Xbit_r26_c14 bl_14 br_14 wl_26 vdd gnd cell_6t
Xbit_r27_c14 bl_14 br_14 wl_27 vdd gnd cell_6t
Xbit_r28_c14 bl_14 br_14 wl_28 vdd gnd cell_6t
Xbit_r29_c14 bl_14 br_14 wl_29 vdd gnd cell_6t
Xbit_r30_c14 bl_14 br_14 wl_30 vdd gnd cell_6t
Xbit_r31_c14 bl_14 br_14 wl_31 vdd gnd cell_6t
Xbit_r32_c14 bl_14 br_14 wl_32 vdd gnd cell_6t
Xbit_r33_c14 bl_14 br_14 wl_33 vdd gnd cell_6t
Xbit_r34_c14 bl_14 br_14 wl_34 vdd gnd cell_6t
Xbit_r35_c14 bl_14 br_14 wl_35 vdd gnd cell_6t
Xbit_r36_c14 bl_14 br_14 wl_36 vdd gnd cell_6t
Xbit_r37_c14 bl_14 br_14 wl_37 vdd gnd cell_6t
Xbit_r38_c14 bl_14 br_14 wl_38 vdd gnd cell_6t
Xbit_r39_c14 bl_14 br_14 wl_39 vdd gnd cell_6t
Xbit_r40_c14 bl_14 br_14 wl_40 vdd gnd cell_6t
Xbit_r41_c14 bl_14 br_14 wl_41 vdd gnd cell_6t
Xbit_r42_c14 bl_14 br_14 wl_42 vdd gnd cell_6t
Xbit_r43_c14 bl_14 br_14 wl_43 vdd gnd cell_6t
Xbit_r44_c14 bl_14 br_14 wl_44 vdd gnd cell_6t
Xbit_r45_c14 bl_14 br_14 wl_45 vdd gnd cell_6t
Xbit_r46_c14 bl_14 br_14 wl_46 vdd gnd cell_6t
Xbit_r47_c14 bl_14 br_14 wl_47 vdd gnd cell_6t
Xbit_r48_c14 bl_14 br_14 wl_48 vdd gnd cell_6t
Xbit_r49_c14 bl_14 br_14 wl_49 vdd gnd cell_6t
Xbit_r50_c14 bl_14 br_14 wl_50 vdd gnd cell_6t
Xbit_r51_c14 bl_14 br_14 wl_51 vdd gnd cell_6t
Xbit_r52_c14 bl_14 br_14 wl_52 vdd gnd cell_6t
Xbit_r53_c14 bl_14 br_14 wl_53 vdd gnd cell_6t
Xbit_r54_c14 bl_14 br_14 wl_54 vdd gnd cell_6t
Xbit_r55_c14 bl_14 br_14 wl_55 vdd gnd cell_6t
Xbit_r56_c14 bl_14 br_14 wl_56 vdd gnd cell_6t
Xbit_r57_c14 bl_14 br_14 wl_57 vdd gnd cell_6t
Xbit_r58_c14 bl_14 br_14 wl_58 vdd gnd cell_6t
Xbit_r59_c14 bl_14 br_14 wl_59 vdd gnd cell_6t
Xbit_r60_c14 bl_14 br_14 wl_60 vdd gnd cell_6t
Xbit_r61_c14 bl_14 br_14 wl_61 vdd gnd cell_6t
Xbit_r62_c14 bl_14 br_14 wl_62 vdd gnd cell_6t
Xbit_r63_c14 bl_14 br_14 wl_63 vdd gnd cell_6t
Xbit_r64_c14 bl_14 br_14 wl_64 vdd gnd cell_6t
Xbit_r65_c14 bl_14 br_14 wl_65 vdd gnd cell_6t
Xbit_r66_c14 bl_14 br_14 wl_66 vdd gnd cell_6t
Xbit_r67_c14 bl_14 br_14 wl_67 vdd gnd cell_6t
Xbit_r68_c14 bl_14 br_14 wl_68 vdd gnd cell_6t
Xbit_r69_c14 bl_14 br_14 wl_69 vdd gnd cell_6t
Xbit_r70_c14 bl_14 br_14 wl_70 vdd gnd cell_6t
Xbit_r71_c14 bl_14 br_14 wl_71 vdd gnd cell_6t
Xbit_r72_c14 bl_14 br_14 wl_72 vdd gnd cell_6t
Xbit_r73_c14 bl_14 br_14 wl_73 vdd gnd cell_6t
Xbit_r74_c14 bl_14 br_14 wl_74 vdd gnd cell_6t
Xbit_r75_c14 bl_14 br_14 wl_75 vdd gnd cell_6t
Xbit_r76_c14 bl_14 br_14 wl_76 vdd gnd cell_6t
Xbit_r77_c14 bl_14 br_14 wl_77 vdd gnd cell_6t
Xbit_r78_c14 bl_14 br_14 wl_78 vdd gnd cell_6t
Xbit_r79_c14 bl_14 br_14 wl_79 vdd gnd cell_6t
Xbit_r80_c14 bl_14 br_14 wl_80 vdd gnd cell_6t
Xbit_r81_c14 bl_14 br_14 wl_81 vdd gnd cell_6t
Xbit_r82_c14 bl_14 br_14 wl_82 vdd gnd cell_6t
Xbit_r83_c14 bl_14 br_14 wl_83 vdd gnd cell_6t
Xbit_r84_c14 bl_14 br_14 wl_84 vdd gnd cell_6t
Xbit_r85_c14 bl_14 br_14 wl_85 vdd gnd cell_6t
Xbit_r86_c14 bl_14 br_14 wl_86 vdd gnd cell_6t
Xbit_r87_c14 bl_14 br_14 wl_87 vdd gnd cell_6t
Xbit_r88_c14 bl_14 br_14 wl_88 vdd gnd cell_6t
Xbit_r89_c14 bl_14 br_14 wl_89 vdd gnd cell_6t
Xbit_r90_c14 bl_14 br_14 wl_90 vdd gnd cell_6t
Xbit_r91_c14 bl_14 br_14 wl_91 vdd gnd cell_6t
Xbit_r92_c14 bl_14 br_14 wl_92 vdd gnd cell_6t
Xbit_r93_c14 bl_14 br_14 wl_93 vdd gnd cell_6t
Xbit_r94_c14 bl_14 br_14 wl_94 vdd gnd cell_6t
Xbit_r95_c14 bl_14 br_14 wl_95 vdd gnd cell_6t
Xbit_r96_c14 bl_14 br_14 wl_96 vdd gnd cell_6t
Xbit_r97_c14 bl_14 br_14 wl_97 vdd gnd cell_6t
Xbit_r98_c14 bl_14 br_14 wl_98 vdd gnd cell_6t
Xbit_r99_c14 bl_14 br_14 wl_99 vdd gnd cell_6t
Xbit_r100_c14 bl_14 br_14 wl_100 vdd gnd cell_6t
Xbit_r101_c14 bl_14 br_14 wl_101 vdd gnd cell_6t
Xbit_r102_c14 bl_14 br_14 wl_102 vdd gnd cell_6t
Xbit_r103_c14 bl_14 br_14 wl_103 vdd gnd cell_6t
Xbit_r104_c14 bl_14 br_14 wl_104 vdd gnd cell_6t
Xbit_r105_c14 bl_14 br_14 wl_105 vdd gnd cell_6t
Xbit_r106_c14 bl_14 br_14 wl_106 vdd gnd cell_6t
Xbit_r107_c14 bl_14 br_14 wl_107 vdd gnd cell_6t
Xbit_r108_c14 bl_14 br_14 wl_108 vdd gnd cell_6t
Xbit_r109_c14 bl_14 br_14 wl_109 vdd gnd cell_6t
Xbit_r110_c14 bl_14 br_14 wl_110 vdd gnd cell_6t
Xbit_r111_c14 bl_14 br_14 wl_111 vdd gnd cell_6t
Xbit_r112_c14 bl_14 br_14 wl_112 vdd gnd cell_6t
Xbit_r113_c14 bl_14 br_14 wl_113 vdd gnd cell_6t
Xbit_r114_c14 bl_14 br_14 wl_114 vdd gnd cell_6t
Xbit_r115_c14 bl_14 br_14 wl_115 vdd gnd cell_6t
Xbit_r116_c14 bl_14 br_14 wl_116 vdd gnd cell_6t
Xbit_r117_c14 bl_14 br_14 wl_117 vdd gnd cell_6t
Xbit_r118_c14 bl_14 br_14 wl_118 vdd gnd cell_6t
Xbit_r119_c14 bl_14 br_14 wl_119 vdd gnd cell_6t
Xbit_r120_c14 bl_14 br_14 wl_120 vdd gnd cell_6t
Xbit_r121_c14 bl_14 br_14 wl_121 vdd gnd cell_6t
Xbit_r122_c14 bl_14 br_14 wl_122 vdd gnd cell_6t
Xbit_r123_c14 bl_14 br_14 wl_123 vdd gnd cell_6t
Xbit_r124_c14 bl_14 br_14 wl_124 vdd gnd cell_6t
Xbit_r125_c14 bl_14 br_14 wl_125 vdd gnd cell_6t
Xbit_r126_c14 bl_14 br_14 wl_126 vdd gnd cell_6t
Xbit_r127_c14 bl_14 br_14 wl_127 vdd gnd cell_6t
Xbit_r128_c14 bl_14 br_14 wl_128 vdd gnd cell_6t
Xbit_r129_c14 bl_14 br_14 wl_129 vdd gnd cell_6t
Xbit_r130_c14 bl_14 br_14 wl_130 vdd gnd cell_6t
Xbit_r131_c14 bl_14 br_14 wl_131 vdd gnd cell_6t
Xbit_r132_c14 bl_14 br_14 wl_132 vdd gnd cell_6t
Xbit_r133_c14 bl_14 br_14 wl_133 vdd gnd cell_6t
Xbit_r134_c14 bl_14 br_14 wl_134 vdd gnd cell_6t
Xbit_r135_c14 bl_14 br_14 wl_135 vdd gnd cell_6t
Xbit_r136_c14 bl_14 br_14 wl_136 vdd gnd cell_6t
Xbit_r137_c14 bl_14 br_14 wl_137 vdd gnd cell_6t
Xbit_r138_c14 bl_14 br_14 wl_138 vdd gnd cell_6t
Xbit_r139_c14 bl_14 br_14 wl_139 vdd gnd cell_6t
Xbit_r140_c14 bl_14 br_14 wl_140 vdd gnd cell_6t
Xbit_r141_c14 bl_14 br_14 wl_141 vdd gnd cell_6t
Xbit_r142_c14 bl_14 br_14 wl_142 vdd gnd cell_6t
Xbit_r143_c14 bl_14 br_14 wl_143 vdd gnd cell_6t
Xbit_r144_c14 bl_14 br_14 wl_144 vdd gnd cell_6t
Xbit_r145_c14 bl_14 br_14 wl_145 vdd gnd cell_6t
Xbit_r146_c14 bl_14 br_14 wl_146 vdd gnd cell_6t
Xbit_r147_c14 bl_14 br_14 wl_147 vdd gnd cell_6t
Xbit_r148_c14 bl_14 br_14 wl_148 vdd gnd cell_6t
Xbit_r149_c14 bl_14 br_14 wl_149 vdd gnd cell_6t
Xbit_r150_c14 bl_14 br_14 wl_150 vdd gnd cell_6t
Xbit_r151_c14 bl_14 br_14 wl_151 vdd gnd cell_6t
Xbit_r152_c14 bl_14 br_14 wl_152 vdd gnd cell_6t
Xbit_r153_c14 bl_14 br_14 wl_153 vdd gnd cell_6t
Xbit_r154_c14 bl_14 br_14 wl_154 vdd gnd cell_6t
Xbit_r155_c14 bl_14 br_14 wl_155 vdd gnd cell_6t
Xbit_r156_c14 bl_14 br_14 wl_156 vdd gnd cell_6t
Xbit_r157_c14 bl_14 br_14 wl_157 vdd gnd cell_6t
Xbit_r158_c14 bl_14 br_14 wl_158 vdd gnd cell_6t
Xbit_r159_c14 bl_14 br_14 wl_159 vdd gnd cell_6t
Xbit_r160_c14 bl_14 br_14 wl_160 vdd gnd cell_6t
Xbit_r161_c14 bl_14 br_14 wl_161 vdd gnd cell_6t
Xbit_r162_c14 bl_14 br_14 wl_162 vdd gnd cell_6t
Xbit_r163_c14 bl_14 br_14 wl_163 vdd gnd cell_6t
Xbit_r164_c14 bl_14 br_14 wl_164 vdd gnd cell_6t
Xbit_r165_c14 bl_14 br_14 wl_165 vdd gnd cell_6t
Xbit_r166_c14 bl_14 br_14 wl_166 vdd gnd cell_6t
Xbit_r167_c14 bl_14 br_14 wl_167 vdd gnd cell_6t
Xbit_r168_c14 bl_14 br_14 wl_168 vdd gnd cell_6t
Xbit_r169_c14 bl_14 br_14 wl_169 vdd gnd cell_6t
Xbit_r170_c14 bl_14 br_14 wl_170 vdd gnd cell_6t
Xbit_r171_c14 bl_14 br_14 wl_171 vdd gnd cell_6t
Xbit_r172_c14 bl_14 br_14 wl_172 vdd gnd cell_6t
Xbit_r173_c14 bl_14 br_14 wl_173 vdd gnd cell_6t
Xbit_r174_c14 bl_14 br_14 wl_174 vdd gnd cell_6t
Xbit_r175_c14 bl_14 br_14 wl_175 vdd gnd cell_6t
Xbit_r176_c14 bl_14 br_14 wl_176 vdd gnd cell_6t
Xbit_r177_c14 bl_14 br_14 wl_177 vdd gnd cell_6t
Xbit_r178_c14 bl_14 br_14 wl_178 vdd gnd cell_6t
Xbit_r179_c14 bl_14 br_14 wl_179 vdd gnd cell_6t
Xbit_r180_c14 bl_14 br_14 wl_180 vdd gnd cell_6t
Xbit_r181_c14 bl_14 br_14 wl_181 vdd gnd cell_6t
Xbit_r182_c14 bl_14 br_14 wl_182 vdd gnd cell_6t
Xbit_r183_c14 bl_14 br_14 wl_183 vdd gnd cell_6t
Xbit_r184_c14 bl_14 br_14 wl_184 vdd gnd cell_6t
Xbit_r185_c14 bl_14 br_14 wl_185 vdd gnd cell_6t
Xbit_r186_c14 bl_14 br_14 wl_186 vdd gnd cell_6t
Xbit_r187_c14 bl_14 br_14 wl_187 vdd gnd cell_6t
Xbit_r188_c14 bl_14 br_14 wl_188 vdd gnd cell_6t
Xbit_r189_c14 bl_14 br_14 wl_189 vdd gnd cell_6t
Xbit_r190_c14 bl_14 br_14 wl_190 vdd gnd cell_6t
Xbit_r191_c14 bl_14 br_14 wl_191 vdd gnd cell_6t
Xbit_r192_c14 bl_14 br_14 wl_192 vdd gnd cell_6t
Xbit_r193_c14 bl_14 br_14 wl_193 vdd gnd cell_6t
Xbit_r194_c14 bl_14 br_14 wl_194 vdd gnd cell_6t
Xbit_r195_c14 bl_14 br_14 wl_195 vdd gnd cell_6t
Xbit_r196_c14 bl_14 br_14 wl_196 vdd gnd cell_6t
Xbit_r197_c14 bl_14 br_14 wl_197 vdd gnd cell_6t
Xbit_r198_c14 bl_14 br_14 wl_198 vdd gnd cell_6t
Xbit_r199_c14 bl_14 br_14 wl_199 vdd gnd cell_6t
Xbit_r200_c14 bl_14 br_14 wl_200 vdd gnd cell_6t
Xbit_r201_c14 bl_14 br_14 wl_201 vdd gnd cell_6t
Xbit_r202_c14 bl_14 br_14 wl_202 vdd gnd cell_6t
Xbit_r203_c14 bl_14 br_14 wl_203 vdd gnd cell_6t
Xbit_r204_c14 bl_14 br_14 wl_204 vdd gnd cell_6t
Xbit_r205_c14 bl_14 br_14 wl_205 vdd gnd cell_6t
Xbit_r206_c14 bl_14 br_14 wl_206 vdd gnd cell_6t
Xbit_r207_c14 bl_14 br_14 wl_207 vdd gnd cell_6t
Xbit_r208_c14 bl_14 br_14 wl_208 vdd gnd cell_6t
Xbit_r209_c14 bl_14 br_14 wl_209 vdd gnd cell_6t
Xbit_r210_c14 bl_14 br_14 wl_210 vdd gnd cell_6t
Xbit_r211_c14 bl_14 br_14 wl_211 vdd gnd cell_6t
Xbit_r212_c14 bl_14 br_14 wl_212 vdd gnd cell_6t
Xbit_r213_c14 bl_14 br_14 wl_213 vdd gnd cell_6t
Xbit_r214_c14 bl_14 br_14 wl_214 vdd gnd cell_6t
Xbit_r215_c14 bl_14 br_14 wl_215 vdd gnd cell_6t
Xbit_r216_c14 bl_14 br_14 wl_216 vdd gnd cell_6t
Xbit_r217_c14 bl_14 br_14 wl_217 vdd gnd cell_6t
Xbit_r218_c14 bl_14 br_14 wl_218 vdd gnd cell_6t
Xbit_r219_c14 bl_14 br_14 wl_219 vdd gnd cell_6t
Xbit_r220_c14 bl_14 br_14 wl_220 vdd gnd cell_6t
Xbit_r221_c14 bl_14 br_14 wl_221 vdd gnd cell_6t
Xbit_r222_c14 bl_14 br_14 wl_222 vdd gnd cell_6t
Xbit_r223_c14 bl_14 br_14 wl_223 vdd gnd cell_6t
Xbit_r224_c14 bl_14 br_14 wl_224 vdd gnd cell_6t
Xbit_r225_c14 bl_14 br_14 wl_225 vdd gnd cell_6t
Xbit_r226_c14 bl_14 br_14 wl_226 vdd gnd cell_6t
Xbit_r227_c14 bl_14 br_14 wl_227 vdd gnd cell_6t
Xbit_r228_c14 bl_14 br_14 wl_228 vdd gnd cell_6t
Xbit_r229_c14 bl_14 br_14 wl_229 vdd gnd cell_6t
Xbit_r230_c14 bl_14 br_14 wl_230 vdd gnd cell_6t
Xbit_r231_c14 bl_14 br_14 wl_231 vdd gnd cell_6t
Xbit_r232_c14 bl_14 br_14 wl_232 vdd gnd cell_6t
Xbit_r233_c14 bl_14 br_14 wl_233 vdd gnd cell_6t
Xbit_r234_c14 bl_14 br_14 wl_234 vdd gnd cell_6t
Xbit_r235_c14 bl_14 br_14 wl_235 vdd gnd cell_6t
Xbit_r236_c14 bl_14 br_14 wl_236 vdd gnd cell_6t
Xbit_r237_c14 bl_14 br_14 wl_237 vdd gnd cell_6t
Xbit_r238_c14 bl_14 br_14 wl_238 vdd gnd cell_6t
Xbit_r239_c14 bl_14 br_14 wl_239 vdd gnd cell_6t
Xbit_r240_c14 bl_14 br_14 wl_240 vdd gnd cell_6t
Xbit_r241_c14 bl_14 br_14 wl_241 vdd gnd cell_6t
Xbit_r242_c14 bl_14 br_14 wl_242 vdd gnd cell_6t
Xbit_r243_c14 bl_14 br_14 wl_243 vdd gnd cell_6t
Xbit_r244_c14 bl_14 br_14 wl_244 vdd gnd cell_6t
Xbit_r245_c14 bl_14 br_14 wl_245 vdd gnd cell_6t
Xbit_r246_c14 bl_14 br_14 wl_246 vdd gnd cell_6t
Xbit_r247_c14 bl_14 br_14 wl_247 vdd gnd cell_6t
Xbit_r248_c14 bl_14 br_14 wl_248 vdd gnd cell_6t
Xbit_r249_c14 bl_14 br_14 wl_249 vdd gnd cell_6t
Xbit_r250_c14 bl_14 br_14 wl_250 vdd gnd cell_6t
Xbit_r251_c14 bl_14 br_14 wl_251 vdd gnd cell_6t
Xbit_r252_c14 bl_14 br_14 wl_252 vdd gnd cell_6t
Xbit_r253_c14 bl_14 br_14 wl_253 vdd gnd cell_6t
Xbit_r254_c14 bl_14 br_14 wl_254 vdd gnd cell_6t
Xbit_r255_c14 bl_14 br_14 wl_255 vdd gnd cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd cell_6t
Xbit_r1_c15 bl_15 br_15 wl_1 vdd gnd cell_6t
Xbit_r2_c15 bl_15 br_15 wl_2 vdd gnd cell_6t
Xbit_r3_c15 bl_15 br_15 wl_3 vdd gnd cell_6t
Xbit_r4_c15 bl_15 br_15 wl_4 vdd gnd cell_6t
Xbit_r5_c15 bl_15 br_15 wl_5 vdd gnd cell_6t
Xbit_r6_c15 bl_15 br_15 wl_6 vdd gnd cell_6t
Xbit_r7_c15 bl_15 br_15 wl_7 vdd gnd cell_6t
Xbit_r8_c15 bl_15 br_15 wl_8 vdd gnd cell_6t
Xbit_r9_c15 bl_15 br_15 wl_9 vdd gnd cell_6t
Xbit_r10_c15 bl_15 br_15 wl_10 vdd gnd cell_6t
Xbit_r11_c15 bl_15 br_15 wl_11 vdd gnd cell_6t
Xbit_r12_c15 bl_15 br_15 wl_12 vdd gnd cell_6t
Xbit_r13_c15 bl_15 br_15 wl_13 vdd gnd cell_6t
Xbit_r14_c15 bl_15 br_15 wl_14 vdd gnd cell_6t
Xbit_r15_c15 bl_15 br_15 wl_15 vdd gnd cell_6t
Xbit_r16_c15 bl_15 br_15 wl_16 vdd gnd cell_6t
Xbit_r17_c15 bl_15 br_15 wl_17 vdd gnd cell_6t
Xbit_r18_c15 bl_15 br_15 wl_18 vdd gnd cell_6t
Xbit_r19_c15 bl_15 br_15 wl_19 vdd gnd cell_6t
Xbit_r20_c15 bl_15 br_15 wl_20 vdd gnd cell_6t
Xbit_r21_c15 bl_15 br_15 wl_21 vdd gnd cell_6t
Xbit_r22_c15 bl_15 br_15 wl_22 vdd gnd cell_6t
Xbit_r23_c15 bl_15 br_15 wl_23 vdd gnd cell_6t
Xbit_r24_c15 bl_15 br_15 wl_24 vdd gnd cell_6t
Xbit_r25_c15 bl_15 br_15 wl_25 vdd gnd cell_6t
Xbit_r26_c15 bl_15 br_15 wl_26 vdd gnd cell_6t
Xbit_r27_c15 bl_15 br_15 wl_27 vdd gnd cell_6t
Xbit_r28_c15 bl_15 br_15 wl_28 vdd gnd cell_6t
Xbit_r29_c15 bl_15 br_15 wl_29 vdd gnd cell_6t
Xbit_r30_c15 bl_15 br_15 wl_30 vdd gnd cell_6t
Xbit_r31_c15 bl_15 br_15 wl_31 vdd gnd cell_6t
Xbit_r32_c15 bl_15 br_15 wl_32 vdd gnd cell_6t
Xbit_r33_c15 bl_15 br_15 wl_33 vdd gnd cell_6t
Xbit_r34_c15 bl_15 br_15 wl_34 vdd gnd cell_6t
Xbit_r35_c15 bl_15 br_15 wl_35 vdd gnd cell_6t
Xbit_r36_c15 bl_15 br_15 wl_36 vdd gnd cell_6t
Xbit_r37_c15 bl_15 br_15 wl_37 vdd gnd cell_6t
Xbit_r38_c15 bl_15 br_15 wl_38 vdd gnd cell_6t
Xbit_r39_c15 bl_15 br_15 wl_39 vdd gnd cell_6t
Xbit_r40_c15 bl_15 br_15 wl_40 vdd gnd cell_6t
Xbit_r41_c15 bl_15 br_15 wl_41 vdd gnd cell_6t
Xbit_r42_c15 bl_15 br_15 wl_42 vdd gnd cell_6t
Xbit_r43_c15 bl_15 br_15 wl_43 vdd gnd cell_6t
Xbit_r44_c15 bl_15 br_15 wl_44 vdd gnd cell_6t
Xbit_r45_c15 bl_15 br_15 wl_45 vdd gnd cell_6t
Xbit_r46_c15 bl_15 br_15 wl_46 vdd gnd cell_6t
Xbit_r47_c15 bl_15 br_15 wl_47 vdd gnd cell_6t
Xbit_r48_c15 bl_15 br_15 wl_48 vdd gnd cell_6t
Xbit_r49_c15 bl_15 br_15 wl_49 vdd gnd cell_6t
Xbit_r50_c15 bl_15 br_15 wl_50 vdd gnd cell_6t
Xbit_r51_c15 bl_15 br_15 wl_51 vdd gnd cell_6t
Xbit_r52_c15 bl_15 br_15 wl_52 vdd gnd cell_6t
Xbit_r53_c15 bl_15 br_15 wl_53 vdd gnd cell_6t
Xbit_r54_c15 bl_15 br_15 wl_54 vdd gnd cell_6t
Xbit_r55_c15 bl_15 br_15 wl_55 vdd gnd cell_6t
Xbit_r56_c15 bl_15 br_15 wl_56 vdd gnd cell_6t
Xbit_r57_c15 bl_15 br_15 wl_57 vdd gnd cell_6t
Xbit_r58_c15 bl_15 br_15 wl_58 vdd gnd cell_6t
Xbit_r59_c15 bl_15 br_15 wl_59 vdd gnd cell_6t
Xbit_r60_c15 bl_15 br_15 wl_60 vdd gnd cell_6t
Xbit_r61_c15 bl_15 br_15 wl_61 vdd gnd cell_6t
Xbit_r62_c15 bl_15 br_15 wl_62 vdd gnd cell_6t
Xbit_r63_c15 bl_15 br_15 wl_63 vdd gnd cell_6t
Xbit_r64_c15 bl_15 br_15 wl_64 vdd gnd cell_6t
Xbit_r65_c15 bl_15 br_15 wl_65 vdd gnd cell_6t
Xbit_r66_c15 bl_15 br_15 wl_66 vdd gnd cell_6t
Xbit_r67_c15 bl_15 br_15 wl_67 vdd gnd cell_6t
Xbit_r68_c15 bl_15 br_15 wl_68 vdd gnd cell_6t
Xbit_r69_c15 bl_15 br_15 wl_69 vdd gnd cell_6t
Xbit_r70_c15 bl_15 br_15 wl_70 vdd gnd cell_6t
Xbit_r71_c15 bl_15 br_15 wl_71 vdd gnd cell_6t
Xbit_r72_c15 bl_15 br_15 wl_72 vdd gnd cell_6t
Xbit_r73_c15 bl_15 br_15 wl_73 vdd gnd cell_6t
Xbit_r74_c15 bl_15 br_15 wl_74 vdd gnd cell_6t
Xbit_r75_c15 bl_15 br_15 wl_75 vdd gnd cell_6t
Xbit_r76_c15 bl_15 br_15 wl_76 vdd gnd cell_6t
Xbit_r77_c15 bl_15 br_15 wl_77 vdd gnd cell_6t
Xbit_r78_c15 bl_15 br_15 wl_78 vdd gnd cell_6t
Xbit_r79_c15 bl_15 br_15 wl_79 vdd gnd cell_6t
Xbit_r80_c15 bl_15 br_15 wl_80 vdd gnd cell_6t
Xbit_r81_c15 bl_15 br_15 wl_81 vdd gnd cell_6t
Xbit_r82_c15 bl_15 br_15 wl_82 vdd gnd cell_6t
Xbit_r83_c15 bl_15 br_15 wl_83 vdd gnd cell_6t
Xbit_r84_c15 bl_15 br_15 wl_84 vdd gnd cell_6t
Xbit_r85_c15 bl_15 br_15 wl_85 vdd gnd cell_6t
Xbit_r86_c15 bl_15 br_15 wl_86 vdd gnd cell_6t
Xbit_r87_c15 bl_15 br_15 wl_87 vdd gnd cell_6t
Xbit_r88_c15 bl_15 br_15 wl_88 vdd gnd cell_6t
Xbit_r89_c15 bl_15 br_15 wl_89 vdd gnd cell_6t
Xbit_r90_c15 bl_15 br_15 wl_90 vdd gnd cell_6t
Xbit_r91_c15 bl_15 br_15 wl_91 vdd gnd cell_6t
Xbit_r92_c15 bl_15 br_15 wl_92 vdd gnd cell_6t
Xbit_r93_c15 bl_15 br_15 wl_93 vdd gnd cell_6t
Xbit_r94_c15 bl_15 br_15 wl_94 vdd gnd cell_6t
Xbit_r95_c15 bl_15 br_15 wl_95 vdd gnd cell_6t
Xbit_r96_c15 bl_15 br_15 wl_96 vdd gnd cell_6t
Xbit_r97_c15 bl_15 br_15 wl_97 vdd gnd cell_6t
Xbit_r98_c15 bl_15 br_15 wl_98 vdd gnd cell_6t
Xbit_r99_c15 bl_15 br_15 wl_99 vdd gnd cell_6t
Xbit_r100_c15 bl_15 br_15 wl_100 vdd gnd cell_6t
Xbit_r101_c15 bl_15 br_15 wl_101 vdd gnd cell_6t
Xbit_r102_c15 bl_15 br_15 wl_102 vdd gnd cell_6t
Xbit_r103_c15 bl_15 br_15 wl_103 vdd gnd cell_6t
Xbit_r104_c15 bl_15 br_15 wl_104 vdd gnd cell_6t
Xbit_r105_c15 bl_15 br_15 wl_105 vdd gnd cell_6t
Xbit_r106_c15 bl_15 br_15 wl_106 vdd gnd cell_6t
Xbit_r107_c15 bl_15 br_15 wl_107 vdd gnd cell_6t
Xbit_r108_c15 bl_15 br_15 wl_108 vdd gnd cell_6t
Xbit_r109_c15 bl_15 br_15 wl_109 vdd gnd cell_6t
Xbit_r110_c15 bl_15 br_15 wl_110 vdd gnd cell_6t
Xbit_r111_c15 bl_15 br_15 wl_111 vdd gnd cell_6t
Xbit_r112_c15 bl_15 br_15 wl_112 vdd gnd cell_6t
Xbit_r113_c15 bl_15 br_15 wl_113 vdd gnd cell_6t
Xbit_r114_c15 bl_15 br_15 wl_114 vdd gnd cell_6t
Xbit_r115_c15 bl_15 br_15 wl_115 vdd gnd cell_6t
Xbit_r116_c15 bl_15 br_15 wl_116 vdd gnd cell_6t
Xbit_r117_c15 bl_15 br_15 wl_117 vdd gnd cell_6t
Xbit_r118_c15 bl_15 br_15 wl_118 vdd gnd cell_6t
Xbit_r119_c15 bl_15 br_15 wl_119 vdd gnd cell_6t
Xbit_r120_c15 bl_15 br_15 wl_120 vdd gnd cell_6t
Xbit_r121_c15 bl_15 br_15 wl_121 vdd gnd cell_6t
Xbit_r122_c15 bl_15 br_15 wl_122 vdd gnd cell_6t
Xbit_r123_c15 bl_15 br_15 wl_123 vdd gnd cell_6t
Xbit_r124_c15 bl_15 br_15 wl_124 vdd gnd cell_6t
Xbit_r125_c15 bl_15 br_15 wl_125 vdd gnd cell_6t
Xbit_r126_c15 bl_15 br_15 wl_126 vdd gnd cell_6t
Xbit_r127_c15 bl_15 br_15 wl_127 vdd gnd cell_6t
Xbit_r128_c15 bl_15 br_15 wl_128 vdd gnd cell_6t
Xbit_r129_c15 bl_15 br_15 wl_129 vdd gnd cell_6t
Xbit_r130_c15 bl_15 br_15 wl_130 vdd gnd cell_6t
Xbit_r131_c15 bl_15 br_15 wl_131 vdd gnd cell_6t
Xbit_r132_c15 bl_15 br_15 wl_132 vdd gnd cell_6t
Xbit_r133_c15 bl_15 br_15 wl_133 vdd gnd cell_6t
Xbit_r134_c15 bl_15 br_15 wl_134 vdd gnd cell_6t
Xbit_r135_c15 bl_15 br_15 wl_135 vdd gnd cell_6t
Xbit_r136_c15 bl_15 br_15 wl_136 vdd gnd cell_6t
Xbit_r137_c15 bl_15 br_15 wl_137 vdd gnd cell_6t
Xbit_r138_c15 bl_15 br_15 wl_138 vdd gnd cell_6t
Xbit_r139_c15 bl_15 br_15 wl_139 vdd gnd cell_6t
Xbit_r140_c15 bl_15 br_15 wl_140 vdd gnd cell_6t
Xbit_r141_c15 bl_15 br_15 wl_141 vdd gnd cell_6t
Xbit_r142_c15 bl_15 br_15 wl_142 vdd gnd cell_6t
Xbit_r143_c15 bl_15 br_15 wl_143 vdd gnd cell_6t
Xbit_r144_c15 bl_15 br_15 wl_144 vdd gnd cell_6t
Xbit_r145_c15 bl_15 br_15 wl_145 vdd gnd cell_6t
Xbit_r146_c15 bl_15 br_15 wl_146 vdd gnd cell_6t
Xbit_r147_c15 bl_15 br_15 wl_147 vdd gnd cell_6t
Xbit_r148_c15 bl_15 br_15 wl_148 vdd gnd cell_6t
Xbit_r149_c15 bl_15 br_15 wl_149 vdd gnd cell_6t
Xbit_r150_c15 bl_15 br_15 wl_150 vdd gnd cell_6t
Xbit_r151_c15 bl_15 br_15 wl_151 vdd gnd cell_6t
Xbit_r152_c15 bl_15 br_15 wl_152 vdd gnd cell_6t
Xbit_r153_c15 bl_15 br_15 wl_153 vdd gnd cell_6t
Xbit_r154_c15 bl_15 br_15 wl_154 vdd gnd cell_6t
Xbit_r155_c15 bl_15 br_15 wl_155 vdd gnd cell_6t
Xbit_r156_c15 bl_15 br_15 wl_156 vdd gnd cell_6t
Xbit_r157_c15 bl_15 br_15 wl_157 vdd gnd cell_6t
Xbit_r158_c15 bl_15 br_15 wl_158 vdd gnd cell_6t
Xbit_r159_c15 bl_15 br_15 wl_159 vdd gnd cell_6t
Xbit_r160_c15 bl_15 br_15 wl_160 vdd gnd cell_6t
Xbit_r161_c15 bl_15 br_15 wl_161 vdd gnd cell_6t
Xbit_r162_c15 bl_15 br_15 wl_162 vdd gnd cell_6t
Xbit_r163_c15 bl_15 br_15 wl_163 vdd gnd cell_6t
Xbit_r164_c15 bl_15 br_15 wl_164 vdd gnd cell_6t
Xbit_r165_c15 bl_15 br_15 wl_165 vdd gnd cell_6t
Xbit_r166_c15 bl_15 br_15 wl_166 vdd gnd cell_6t
Xbit_r167_c15 bl_15 br_15 wl_167 vdd gnd cell_6t
Xbit_r168_c15 bl_15 br_15 wl_168 vdd gnd cell_6t
Xbit_r169_c15 bl_15 br_15 wl_169 vdd gnd cell_6t
Xbit_r170_c15 bl_15 br_15 wl_170 vdd gnd cell_6t
Xbit_r171_c15 bl_15 br_15 wl_171 vdd gnd cell_6t
Xbit_r172_c15 bl_15 br_15 wl_172 vdd gnd cell_6t
Xbit_r173_c15 bl_15 br_15 wl_173 vdd gnd cell_6t
Xbit_r174_c15 bl_15 br_15 wl_174 vdd gnd cell_6t
Xbit_r175_c15 bl_15 br_15 wl_175 vdd gnd cell_6t
Xbit_r176_c15 bl_15 br_15 wl_176 vdd gnd cell_6t
Xbit_r177_c15 bl_15 br_15 wl_177 vdd gnd cell_6t
Xbit_r178_c15 bl_15 br_15 wl_178 vdd gnd cell_6t
Xbit_r179_c15 bl_15 br_15 wl_179 vdd gnd cell_6t
Xbit_r180_c15 bl_15 br_15 wl_180 vdd gnd cell_6t
Xbit_r181_c15 bl_15 br_15 wl_181 vdd gnd cell_6t
Xbit_r182_c15 bl_15 br_15 wl_182 vdd gnd cell_6t
Xbit_r183_c15 bl_15 br_15 wl_183 vdd gnd cell_6t
Xbit_r184_c15 bl_15 br_15 wl_184 vdd gnd cell_6t
Xbit_r185_c15 bl_15 br_15 wl_185 vdd gnd cell_6t
Xbit_r186_c15 bl_15 br_15 wl_186 vdd gnd cell_6t
Xbit_r187_c15 bl_15 br_15 wl_187 vdd gnd cell_6t
Xbit_r188_c15 bl_15 br_15 wl_188 vdd gnd cell_6t
Xbit_r189_c15 bl_15 br_15 wl_189 vdd gnd cell_6t
Xbit_r190_c15 bl_15 br_15 wl_190 vdd gnd cell_6t
Xbit_r191_c15 bl_15 br_15 wl_191 vdd gnd cell_6t
Xbit_r192_c15 bl_15 br_15 wl_192 vdd gnd cell_6t
Xbit_r193_c15 bl_15 br_15 wl_193 vdd gnd cell_6t
Xbit_r194_c15 bl_15 br_15 wl_194 vdd gnd cell_6t
Xbit_r195_c15 bl_15 br_15 wl_195 vdd gnd cell_6t
Xbit_r196_c15 bl_15 br_15 wl_196 vdd gnd cell_6t
Xbit_r197_c15 bl_15 br_15 wl_197 vdd gnd cell_6t
Xbit_r198_c15 bl_15 br_15 wl_198 vdd gnd cell_6t
Xbit_r199_c15 bl_15 br_15 wl_199 vdd gnd cell_6t
Xbit_r200_c15 bl_15 br_15 wl_200 vdd gnd cell_6t
Xbit_r201_c15 bl_15 br_15 wl_201 vdd gnd cell_6t
Xbit_r202_c15 bl_15 br_15 wl_202 vdd gnd cell_6t
Xbit_r203_c15 bl_15 br_15 wl_203 vdd gnd cell_6t
Xbit_r204_c15 bl_15 br_15 wl_204 vdd gnd cell_6t
Xbit_r205_c15 bl_15 br_15 wl_205 vdd gnd cell_6t
Xbit_r206_c15 bl_15 br_15 wl_206 vdd gnd cell_6t
Xbit_r207_c15 bl_15 br_15 wl_207 vdd gnd cell_6t
Xbit_r208_c15 bl_15 br_15 wl_208 vdd gnd cell_6t
Xbit_r209_c15 bl_15 br_15 wl_209 vdd gnd cell_6t
Xbit_r210_c15 bl_15 br_15 wl_210 vdd gnd cell_6t
Xbit_r211_c15 bl_15 br_15 wl_211 vdd gnd cell_6t
Xbit_r212_c15 bl_15 br_15 wl_212 vdd gnd cell_6t
Xbit_r213_c15 bl_15 br_15 wl_213 vdd gnd cell_6t
Xbit_r214_c15 bl_15 br_15 wl_214 vdd gnd cell_6t
Xbit_r215_c15 bl_15 br_15 wl_215 vdd gnd cell_6t
Xbit_r216_c15 bl_15 br_15 wl_216 vdd gnd cell_6t
Xbit_r217_c15 bl_15 br_15 wl_217 vdd gnd cell_6t
Xbit_r218_c15 bl_15 br_15 wl_218 vdd gnd cell_6t
Xbit_r219_c15 bl_15 br_15 wl_219 vdd gnd cell_6t
Xbit_r220_c15 bl_15 br_15 wl_220 vdd gnd cell_6t
Xbit_r221_c15 bl_15 br_15 wl_221 vdd gnd cell_6t
Xbit_r222_c15 bl_15 br_15 wl_222 vdd gnd cell_6t
Xbit_r223_c15 bl_15 br_15 wl_223 vdd gnd cell_6t
Xbit_r224_c15 bl_15 br_15 wl_224 vdd gnd cell_6t
Xbit_r225_c15 bl_15 br_15 wl_225 vdd gnd cell_6t
Xbit_r226_c15 bl_15 br_15 wl_226 vdd gnd cell_6t
Xbit_r227_c15 bl_15 br_15 wl_227 vdd gnd cell_6t
Xbit_r228_c15 bl_15 br_15 wl_228 vdd gnd cell_6t
Xbit_r229_c15 bl_15 br_15 wl_229 vdd gnd cell_6t
Xbit_r230_c15 bl_15 br_15 wl_230 vdd gnd cell_6t
Xbit_r231_c15 bl_15 br_15 wl_231 vdd gnd cell_6t
Xbit_r232_c15 bl_15 br_15 wl_232 vdd gnd cell_6t
Xbit_r233_c15 bl_15 br_15 wl_233 vdd gnd cell_6t
Xbit_r234_c15 bl_15 br_15 wl_234 vdd gnd cell_6t
Xbit_r235_c15 bl_15 br_15 wl_235 vdd gnd cell_6t
Xbit_r236_c15 bl_15 br_15 wl_236 vdd gnd cell_6t
Xbit_r237_c15 bl_15 br_15 wl_237 vdd gnd cell_6t
Xbit_r238_c15 bl_15 br_15 wl_238 vdd gnd cell_6t
Xbit_r239_c15 bl_15 br_15 wl_239 vdd gnd cell_6t
Xbit_r240_c15 bl_15 br_15 wl_240 vdd gnd cell_6t
Xbit_r241_c15 bl_15 br_15 wl_241 vdd gnd cell_6t
Xbit_r242_c15 bl_15 br_15 wl_242 vdd gnd cell_6t
Xbit_r243_c15 bl_15 br_15 wl_243 vdd gnd cell_6t
Xbit_r244_c15 bl_15 br_15 wl_244 vdd gnd cell_6t
Xbit_r245_c15 bl_15 br_15 wl_245 vdd gnd cell_6t
Xbit_r246_c15 bl_15 br_15 wl_246 vdd gnd cell_6t
Xbit_r247_c15 bl_15 br_15 wl_247 vdd gnd cell_6t
Xbit_r248_c15 bl_15 br_15 wl_248 vdd gnd cell_6t
Xbit_r249_c15 bl_15 br_15 wl_249 vdd gnd cell_6t
Xbit_r250_c15 bl_15 br_15 wl_250 vdd gnd cell_6t
Xbit_r251_c15 bl_15 br_15 wl_251 vdd gnd cell_6t
Xbit_r252_c15 bl_15 br_15 wl_252 vdd gnd cell_6t
Xbit_r253_c15 bl_15 br_15 wl_253 vdd gnd cell_6t
Xbit_r254_c15 bl_15 br_15 wl_254 vdd gnd cell_6t
Xbit_r255_c15 bl_15 br_15 wl_255 vdd gnd cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd cell_6t
Xbit_r1_c16 bl_16 br_16 wl_1 vdd gnd cell_6t
Xbit_r2_c16 bl_16 br_16 wl_2 vdd gnd cell_6t
Xbit_r3_c16 bl_16 br_16 wl_3 vdd gnd cell_6t
Xbit_r4_c16 bl_16 br_16 wl_4 vdd gnd cell_6t
Xbit_r5_c16 bl_16 br_16 wl_5 vdd gnd cell_6t
Xbit_r6_c16 bl_16 br_16 wl_6 vdd gnd cell_6t
Xbit_r7_c16 bl_16 br_16 wl_7 vdd gnd cell_6t
Xbit_r8_c16 bl_16 br_16 wl_8 vdd gnd cell_6t
Xbit_r9_c16 bl_16 br_16 wl_9 vdd gnd cell_6t
Xbit_r10_c16 bl_16 br_16 wl_10 vdd gnd cell_6t
Xbit_r11_c16 bl_16 br_16 wl_11 vdd gnd cell_6t
Xbit_r12_c16 bl_16 br_16 wl_12 vdd gnd cell_6t
Xbit_r13_c16 bl_16 br_16 wl_13 vdd gnd cell_6t
Xbit_r14_c16 bl_16 br_16 wl_14 vdd gnd cell_6t
Xbit_r15_c16 bl_16 br_16 wl_15 vdd gnd cell_6t
Xbit_r16_c16 bl_16 br_16 wl_16 vdd gnd cell_6t
Xbit_r17_c16 bl_16 br_16 wl_17 vdd gnd cell_6t
Xbit_r18_c16 bl_16 br_16 wl_18 vdd gnd cell_6t
Xbit_r19_c16 bl_16 br_16 wl_19 vdd gnd cell_6t
Xbit_r20_c16 bl_16 br_16 wl_20 vdd gnd cell_6t
Xbit_r21_c16 bl_16 br_16 wl_21 vdd gnd cell_6t
Xbit_r22_c16 bl_16 br_16 wl_22 vdd gnd cell_6t
Xbit_r23_c16 bl_16 br_16 wl_23 vdd gnd cell_6t
Xbit_r24_c16 bl_16 br_16 wl_24 vdd gnd cell_6t
Xbit_r25_c16 bl_16 br_16 wl_25 vdd gnd cell_6t
Xbit_r26_c16 bl_16 br_16 wl_26 vdd gnd cell_6t
Xbit_r27_c16 bl_16 br_16 wl_27 vdd gnd cell_6t
Xbit_r28_c16 bl_16 br_16 wl_28 vdd gnd cell_6t
Xbit_r29_c16 bl_16 br_16 wl_29 vdd gnd cell_6t
Xbit_r30_c16 bl_16 br_16 wl_30 vdd gnd cell_6t
Xbit_r31_c16 bl_16 br_16 wl_31 vdd gnd cell_6t
Xbit_r32_c16 bl_16 br_16 wl_32 vdd gnd cell_6t
Xbit_r33_c16 bl_16 br_16 wl_33 vdd gnd cell_6t
Xbit_r34_c16 bl_16 br_16 wl_34 vdd gnd cell_6t
Xbit_r35_c16 bl_16 br_16 wl_35 vdd gnd cell_6t
Xbit_r36_c16 bl_16 br_16 wl_36 vdd gnd cell_6t
Xbit_r37_c16 bl_16 br_16 wl_37 vdd gnd cell_6t
Xbit_r38_c16 bl_16 br_16 wl_38 vdd gnd cell_6t
Xbit_r39_c16 bl_16 br_16 wl_39 vdd gnd cell_6t
Xbit_r40_c16 bl_16 br_16 wl_40 vdd gnd cell_6t
Xbit_r41_c16 bl_16 br_16 wl_41 vdd gnd cell_6t
Xbit_r42_c16 bl_16 br_16 wl_42 vdd gnd cell_6t
Xbit_r43_c16 bl_16 br_16 wl_43 vdd gnd cell_6t
Xbit_r44_c16 bl_16 br_16 wl_44 vdd gnd cell_6t
Xbit_r45_c16 bl_16 br_16 wl_45 vdd gnd cell_6t
Xbit_r46_c16 bl_16 br_16 wl_46 vdd gnd cell_6t
Xbit_r47_c16 bl_16 br_16 wl_47 vdd gnd cell_6t
Xbit_r48_c16 bl_16 br_16 wl_48 vdd gnd cell_6t
Xbit_r49_c16 bl_16 br_16 wl_49 vdd gnd cell_6t
Xbit_r50_c16 bl_16 br_16 wl_50 vdd gnd cell_6t
Xbit_r51_c16 bl_16 br_16 wl_51 vdd gnd cell_6t
Xbit_r52_c16 bl_16 br_16 wl_52 vdd gnd cell_6t
Xbit_r53_c16 bl_16 br_16 wl_53 vdd gnd cell_6t
Xbit_r54_c16 bl_16 br_16 wl_54 vdd gnd cell_6t
Xbit_r55_c16 bl_16 br_16 wl_55 vdd gnd cell_6t
Xbit_r56_c16 bl_16 br_16 wl_56 vdd gnd cell_6t
Xbit_r57_c16 bl_16 br_16 wl_57 vdd gnd cell_6t
Xbit_r58_c16 bl_16 br_16 wl_58 vdd gnd cell_6t
Xbit_r59_c16 bl_16 br_16 wl_59 vdd gnd cell_6t
Xbit_r60_c16 bl_16 br_16 wl_60 vdd gnd cell_6t
Xbit_r61_c16 bl_16 br_16 wl_61 vdd gnd cell_6t
Xbit_r62_c16 bl_16 br_16 wl_62 vdd gnd cell_6t
Xbit_r63_c16 bl_16 br_16 wl_63 vdd gnd cell_6t
Xbit_r64_c16 bl_16 br_16 wl_64 vdd gnd cell_6t
Xbit_r65_c16 bl_16 br_16 wl_65 vdd gnd cell_6t
Xbit_r66_c16 bl_16 br_16 wl_66 vdd gnd cell_6t
Xbit_r67_c16 bl_16 br_16 wl_67 vdd gnd cell_6t
Xbit_r68_c16 bl_16 br_16 wl_68 vdd gnd cell_6t
Xbit_r69_c16 bl_16 br_16 wl_69 vdd gnd cell_6t
Xbit_r70_c16 bl_16 br_16 wl_70 vdd gnd cell_6t
Xbit_r71_c16 bl_16 br_16 wl_71 vdd gnd cell_6t
Xbit_r72_c16 bl_16 br_16 wl_72 vdd gnd cell_6t
Xbit_r73_c16 bl_16 br_16 wl_73 vdd gnd cell_6t
Xbit_r74_c16 bl_16 br_16 wl_74 vdd gnd cell_6t
Xbit_r75_c16 bl_16 br_16 wl_75 vdd gnd cell_6t
Xbit_r76_c16 bl_16 br_16 wl_76 vdd gnd cell_6t
Xbit_r77_c16 bl_16 br_16 wl_77 vdd gnd cell_6t
Xbit_r78_c16 bl_16 br_16 wl_78 vdd gnd cell_6t
Xbit_r79_c16 bl_16 br_16 wl_79 vdd gnd cell_6t
Xbit_r80_c16 bl_16 br_16 wl_80 vdd gnd cell_6t
Xbit_r81_c16 bl_16 br_16 wl_81 vdd gnd cell_6t
Xbit_r82_c16 bl_16 br_16 wl_82 vdd gnd cell_6t
Xbit_r83_c16 bl_16 br_16 wl_83 vdd gnd cell_6t
Xbit_r84_c16 bl_16 br_16 wl_84 vdd gnd cell_6t
Xbit_r85_c16 bl_16 br_16 wl_85 vdd gnd cell_6t
Xbit_r86_c16 bl_16 br_16 wl_86 vdd gnd cell_6t
Xbit_r87_c16 bl_16 br_16 wl_87 vdd gnd cell_6t
Xbit_r88_c16 bl_16 br_16 wl_88 vdd gnd cell_6t
Xbit_r89_c16 bl_16 br_16 wl_89 vdd gnd cell_6t
Xbit_r90_c16 bl_16 br_16 wl_90 vdd gnd cell_6t
Xbit_r91_c16 bl_16 br_16 wl_91 vdd gnd cell_6t
Xbit_r92_c16 bl_16 br_16 wl_92 vdd gnd cell_6t
Xbit_r93_c16 bl_16 br_16 wl_93 vdd gnd cell_6t
Xbit_r94_c16 bl_16 br_16 wl_94 vdd gnd cell_6t
Xbit_r95_c16 bl_16 br_16 wl_95 vdd gnd cell_6t
Xbit_r96_c16 bl_16 br_16 wl_96 vdd gnd cell_6t
Xbit_r97_c16 bl_16 br_16 wl_97 vdd gnd cell_6t
Xbit_r98_c16 bl_16 br_16 wl_98 vdd gnd cell_6t
Xbit_r99_c16 bl_16 br_16 wl_99 vdd gnd cell_6t
Xbit_r100_c16 bl_16 br_16 wl_100 vdd gnd cell_6t
Xbit_r101_c16 bl_16 br_16 wl_101 vdd gnd cell_6t
Xbit_r102_c16 bl_16 br_16 wl_102 vdd gnd cell_6t
Xbit_r103_c16 bl_16 br_16 wl_103 vdd gnd cell_6t
Xbit_r104_c16 bl_16 br_16 wl_104 vdd gnd cell_6t
Xbit_r105_c16 bl_16 br_16 wl_105 vdd gnd cell_6t
Xbit_r106_c16 bl_16 br_16 wl_106 vdd gnd cell_6t
Xbit_r107_c16 bl_16 br_16 wl_107 vdd gnd cell_6t
Xbit_r108_c16 bl_16 br_16 wl_108 vdd gnd cell_6t
Xbit_r109_c16 bl_16 br_16 wl_109 vdd gnd cell_6t
Xbit_r110_c16 bl_16 br_16 wl_110 vdd gnd cell_6t
Xbit_r111_c16 bl_16 br_16 wl_111 vdd gnd cell_6t
Xbit_r112_c16 bl_16 br_16 wl_112 vdd gnd cell_6t
Xbit_r113_c16 bl_16 br_16 wl_113 vdd gnd cell_6t
Xbit_r114_c16 bl_16 br_16 wl_114 vdd gnd cell_6t
Xbit_r115_c16 bl_16 br_16 wl_115 vdd gnd cell_6t
Xbit_r116_c16 bl_16 br_16 wl_116 vdd gnd cell_6t
Xbit_r117_c16 bl_16 br_16 wl_117 vdd gnd cell_6t
Xbit_r118_c16 bl_16 br_16 wl_118 vdd gnd cell_6t
Xbit_r119_c16 bl_16 br_16 wl_119 vdd gnd cell_6t
Xbit_r120_c16 bl_16 br_16 wl_120 vdd gnd cell_6t
Xbit_r121_c16 bl_16 br_16 wl_121 vdd gnd cell_6t
Xbit_r122_c16 bl_16 br_16 wl_122 vdd gnd cell_6t
Xbit_r123_c16 bl_16 br_16 wl_123 vdd gnd cell_6t
Xbit_r124_c16 bl_16 br_16 wl_124 vdd gnd cell_6t
Xbit_r125_c16 bl_16 br_16 wl_125 vdd gnd cell_6t
Xbit_r126_c16 bl_16 br_16 wl_126 vdd gnd cell_6t
Xbit_r127_c16 bl_16 br_16 wl_127 vdd gnd cell_6t
Xbit_r128_c16 bl_16 br_16 wl_128 vdd gnd cell_6t
Xbit_r129_c16 bl_16 br_16 wl_129 vdd gnd cell_6t
Xbit_r130_c16 bl_16 br_16 wl_130 vdd gnd cell_6t
Xbit_r131_c16 bl_16 br_16 wl_131 vdd gnd cell_6t
Xbit_r132_c16 bl_16 br_16 wl_132 vdd gnd cell_6t
Xbit_r133_c16 bl_16 br_16 wl_133 vdd gnd cell_6t
Xbit_r134_c16 bl_16 br_16 wl_134 vdd gnd cell_6t
Xbit_r135_c16 bl_16 br_16 wl_135 vdd gnd cell_6t
Xbit_r136_c16 bl_16 br_16 wl_136 vdd gnd cell_6t
Xbit_r137_c16 bl_16 br_16 wl_137 vdd gnd cell_6t
Xbit_r138_c16 bl_16 br_16 wl_138 vdd gnd cell_6t
Xbit_r139_c16 bl_16 br_16 wl_139 vdd gnd cell_6t
Xbit_r140_c16 bl_16 br_16 wl_140 vdd gnd cell_6t
Xbit_r141_c16 bl_16 br_16 wl_141 vdd gnd cell_6t
Xbit_r142_c16 bl_16 br_16 wl_142 vdd gnd cell_6t
Xbit_r143_c16 bl_16 br_16 wl_143 vdd gnd cell_6t
Xbit_r144_c16 bl_16 br_16 wl_144 vdd gnd cell_6t
Xbit_r145_c16 bl_16 br_16 wl_145 vdd gnd cell_6t
Xbit_r146_c16 bl_16 br_16 wl_146 vdd gnd cell_6t
Xbit_r147_c16 bl_16 br_16 wl_147 vdd gnd cell_6t
Xbit_r148_c16 bl_16 br_16 wl_148 vdd gnd cell_6t
Xbit_r149_c16 bl_16 br_16 wl_149 vdd gnd cell_6t
Xbit_r150_c16 bl_16 br_16 wl_150 vdd gnd cell_6t
Xbit_r151_c16 bl_16 br_16 wl_151 vdd gnd cell_6t
Xbit_r152_c16 bl_16 br_16 wl_152 vdd gnd cell_6t
Xbit_r153_c16 bl_16 br_16 wl_153 vdd gnd cell_6t
Xbit_r154_c16 bl_16 br_16 wl_154 vdd gnd cell_6t
Xbit_r155_c16 bl_16 br_16 wl_155 vdd gnd cell_6t
Xbit_r156_c16 bl_16 br_16 wl_156 vdd gnd cell_6t
Xbit_r157_c16 bl_16 br_16 wl_157 vdd gnd cell_6t
Xbit_r158_c16 bl_16 br_16 wl_158 vdd gnd cell_6t
Xbit_r159_c16 bl_16 br_16 wl_159 vdd gnd cell_6t
Xbit_r160_c16 bl_16 br_16 wl_160 vdd gnd cell_6t
Xbit_r161_c16 bl_16 br_16 wl_161 vdd gnd cell_6t
Xbit_r162_c16 bl_16 br_16 wl_162 vdd gnd cell_6t
Xbit_r163_c16 bl_16 br_16 wl_163 vdd gnd cell_6t
Xbit_r164_c16 bl_16 br_16 wl_164 vdd gnd cell_6t
Xbit_r165_c16 bl_16 br_16 wl_165 vdd gnd cell_6t
Xbit_r166_c16 bl_16 br_16 wl_166 vdd gnd cell_6t
Xbit_r167_c16 bl_16 br_16 wl_167 vdd gnd cell_6t
Xbit_r168_c16 bl_16 br_16 wl_168 vdd gnd cell_6t
Xbit_r169_c16 bl_16 br_16 wl_169 vdd gnd cell_6t
Xbit_r170_c16 bl_16 br_16 wl_170 vdd gnd cell_6t
Xbit_r171_c16 bl_16 br_16 wl_171 vdd gnd cell_6t
Xbit_r172_c16 bl_16 br_16 wl_172 vdd gnd cell_6t
Xbit_r173_c16 bl_16 br_16 wl_173 vdd gnd cell_6t
Xbit_r174_c16 bl_16 br_16 wl_174 vdd gnd cell_6t
Xbit_r175_c16 bl_16 br_16 wl_175 vdd gnd cell_6t
Xbit_r176_c16 bl_16 br_16 wl_176 vdd gnd cell_6t
Xbit_r177_c16 bl_16 br_16 wl_177 vdd gnd cell_6t
Xbit_r178_c16 bl_16 br_16 wl_178 vdd gnd cell_6t
Xbit_r179_c16 bl_16 br_16 wl_179 vdd gnd cell_6t
Xbit_r180_c16 bl_16 br_16 wl_180 vdd gnd cell_6t
Xbit_r181_c16 bl_16 br_16 wl_181 vdd gnd cell_6t
Xbit_r182_c16 bl_16 br_16 wl_182 vdd gnd cell_6t
Xbit_r183_c16 bl_16 br_16 wl_183 vdd gnd cell_6t
Xbit_r184_c16 bl_16 br_16 wl_184 vdd gnd cell_6t
Xbit_r185_c16 bl_16 br_16 wl_185 vdd gnd cell_6t
Xbit_r186_c16 bl_16 br_16 wl_186 vdd gnd cell_6t
Xbit_r187_c16 bl_16 br_16 wl_187 vdd gnd cell_6t
Xbit_r188_c16 bl_16 br_16 wl_188 vdd gnd cell_6t
Xbit_r189_c16 bl_16 br_16 wl_189 vdd gnd cell_6t
Xbit_r190_c16 bl_16 br_16 wl_190 vdd gnd cell_6t
Xbit_r191_c16 bl_16 br_16 wl_191 vdd gnd cell_6t
Xbit_r192_c16 bl_16 br_16 wl_192 vdd gnd cell_6t
Xbit_r193_c16 bl_16 br_16 wl_193 vdd gnd cell_6t
Xbit_r194_c16 bl_16 br_16 wl_194 vdd gnd cell_6t
Xbit_r195_c16 bl_16 br_16 wl_195 vdd gnd cell_6t
Xbit_r196_c16 bl_16 br_16 wl_196 vdd gnd cell_6t
Xbit_r197_c16 bl_16 br_16 wl_197 vdd gnd cell_6t
Xbit_r198_c16 bl_16 br_16 wl_198 vdd gnd cell_6t
Xbit_r199_c16 bl_16 br_16 wl_199 vdd gnd cell_6t
Xbit_r200_c16 bl_16 br_16 wl_200 vdd gnd cell_6t
Xbit_r201_c16 bl_16 br_16 wl_201 vdd gnd cell_6t
Xbit_r202_c16 bl_16 br_16 wl_202 vdd gnd cell_6t
Xbit_r203_c16 bl_16 br_16 wl_203 vdd gnd cell_6t
Xbit_r204_c16 bl_16 br_16 wl_204 vdd gnd cell_6t
Xbit_r205_c16 bl_16 br_16 wl_205 vdd gnd cell_6t
Xbit_r206_c16 bl_16 br_16 wl_206 vdd gnd cell_6t
Xbit_r207_c16 bl_16 br_16 wl_207 vdd gnd cell_6t
Xbit_r208_c16 bl_16 br_16 wl_208 vdd gnd cell_6t
Xbit_r209_c16 bl_16 br_16 wl_209 vdd gnd cell_6t
Xbit_r210_c16 bl_16 br_16 wl_210 vdd gnd cell_6t
Xbit_r211_c16 bl_16 br_16 wl_211 vdd gnd cell_6t
Xbit_r212_c16 bl_16 br_16 wl_212 vdd gnd cell_6t
Xbit_r213_c16 bl_16 br_16 wl_213 vdd gnd cell_6t
Xbit_r214_c16 bl_16 br_16 wl_214 vdd gnd cell_6t
Xbit_r215_c16 bl_16 br_16 wl_215 vdd gnd cell_6t
Xbit_r216_c16 bl_16 br_16 wl_216 vdd gnd cell_6t
Xbit_r217_c16 bl_16 br_16 wl_217 vdd gnd cell_6t
Xbit_r218_c16 bl_16 br_16 wl_218 vdd gnd cell_6t
Xbit_r219_c16 bl_16 br_16 wl_219 vdd gnd cell_6t
Xbit_r220_c16 bl_16 br_16 wl_220 vdd gnd cell_6t
Xbit_r221_c16 bl_16 br_16 wl_221 vdd gnd cell_6t
Xbit_r222_c16 bl_16 br_16 wl_222 vdd gnd cell_6t
Xbit_r223_c16 bl_16 br_16 wl_223 vdd gnd cell_6t
Xbit_r224_c16 bl_16 br_16 wl_224 vdd gnd cell_6t
Xbit_r225_c16 bl_16 br_16 wl_225 vdd gnd cell_6t
Xbit_r226_c16 bl_16 br_16 wl_226 vdd gnd cell_6t
Xbit_r227_c16 bl_16 br_16 wl_227 vdd gnd cell_6t
Xbit_r228_c16 bl_16 br_16 wl_228 vdd gnd cell_6t
Xbit_r229_c16 bl_16 br_16 wl_229 vdd gnd cell_6t
Xbit_r230_c16 bl_16 br_16 wl_230 vdd gnd cell_6t
Xbit_r231_c16 bl_16 br_16 wl_231 vdd gnd cell_6t
Xbit_r232_c16 bl_16 br_16 wl_232 vdd gnd cell_6t
Xbit_r233_c16 bl_16 br_16 wl_233 vdd gnd cell_6t
Xbit_r234_c16 bl_16 br_16 wl_234 vdd gnd cell_6t
Xbit_r235_c16 bl_16 br_16 wl_235 vdd gnd cell_6t
Xbit_r236_c16 bl_16 br_16 wl_236 vdd gnd cell_6t
Xbit_r237_c16 bl_16 br_16 wl_237 vdd gnd cell_6t
Xbit_r238_c16 bl_16 br_16 wl_238 vdd gnd cell_6t
Xbit_r239_c16 bl_16 br_16 wl_239 vdd gnd cell_6t
Xbit_r240_c16 bl_16 br_16 wl_240 vdd gnd cell_6t
Xbit_r241_c16 bl_16 br_16 wl_241 vdd gnd cell_6t
Xbit_r242_c16 bl_16 br_16 wl_242 vdd gnd cell_6t
Xbit_r243_c16 bl_16 br_16 wl_243 vdd gnd cell_6t
Xbit_r244_c16 bl_16 br_16 wl_244 vdd gnd cell_6t
Xbit_r245_c16 bl_16 br_16 wl_245 vdd gnd cell_6t
Xbit_r246_c16 bl_16 br_16 wl_246 vdd gnd cell_6t
Xbit_r247_c16 bl_16 br_16 wl_247 vdd gnd cell_6t
Xbit_r248_c16 bl_16 br_16 wl_248 vdd gnd cell_6t
Xbit_r249_c16 bl_16 br_16 wl_249 vdd gnd cell_6t
Xbit_r250_c16 bl_16 br_16 wl_250 vdd gnd cell_6t
Xbit_r251_c16 bl_16 br_16 wl_251 vdd gnd cell_6t
Xbit_r252_c16 bl_16 br_16 wl_252 vdd gnd cell_6t
Xbit_r253_c16 bl_16 br_16 wl_253 vdd gnd cell_6t
Xbit_r254_c16 bl_16 br_16 wl_254 vdd gnd cell_6t
Xbit_r255_c16 bl_16 br_16 wl_255 vdd gnd cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd cell_6t
Xbit_r1_c17 bl_17 br_17 wl_1 vdd gnd cell_6t
Xbit_r2_c17 bl_17 br_17 wl_2 vdd gnd cell_6t
Xbit_r3_c17 bl_17 br_17 wl_3 vdd gnd cell_6t
Xbit_r4_c17 bl_17 br_17 wl_4 vdd gnd cell_6t
Xbit_r5_c17 bl_17 br_17 wl_5 vdd gnd cell_6t
Xbit_r6_c17 bl_17 br_17 wl_6 vdd gnd cell_6t
Xbit_r7_c17 bl_17 br_17 wl_7 vdd gnd cell_6t
Xbit_r8_c17 bl_17 br_17 wl_8 vdd gnd cell_6t
Xbit_r9_c17 bl_17 br_17 wl_9 vdd gnd cell_6t
Xbit_r10_c17 bl_17 br_17 wl_10 vdd gnd cell_6t
Xbit_r11_c17 bl_17 br_17 wl_11 vdd gnd cell_6t
Xbit_r12_c17 bl_17 br_17 wl_12 vdd gnd cell_6t
Xbit_r13_c17 bl_17 br_17 wl_13 vdd gnd cell_6t
Xbit_r14_c17 bl_17 br_17 wl_14 vdd gnd cell_6t
Xbit_r15_c17 bl_17 br_17 wl_15 vdd gnd cell_6t
Xbit_r16_c17 bl_17 br_17 wl_16 vdd gnd cell_6t
Xbit_r17_c17 bl_17 br_17 wl_17 vdd gnd cell_6t
Xbit_r18_c17 bl_17 br_17 wl_18 vdd gnd cell_6t
Xbit_r19_c17 bl_17 br_17 wl_19 vdd gnd cell_6t
Xbit_r20_c17 bl_17 br_17 wl_20 vdd gnd cell_6t
Xbit_r21_c17 bl_17 br_17 wl_21 vdd gnd cell_6t
Xbit_r22_c17 bl_17 br_17 wl_22 vdd gnd cell_6t
Xbit_r23_c17 bl_17 br_17 wl_23 vdd gnd cell_6t
Xbit_r24_c17 bl_17 br_17 wl_24 vdd gnd cell_6t
Xbit_r25_c17 bl_17 br_17 wl_25 vdd gnd cell_6t
Xbit_r26_c17 bl_17 br_17 wl_26 vdd gnd cell_6t
Xbit_r27_c17 bl_17 br_17 wl_27 vdd gnd cell_6t
Xbit_r28_c17 bl_17 br_17 wl_28 vdd gnd cell_6t
Xbit_r29_c17 bl_17 br_17 wl_29 vdd gnd cell_6t
Xbit_r30_c17 bl_17 br_17 wl_30 vdd gnd cell_6t
Xbit_r31_c17 bl_17 br_17 wl_31 vdd gnd cell_6t
Xbit_r32_c17 bl_17 br_17 wl_32 vdd gnd cell_6t
Xbit_r33_c17 bl_17 br_17 wl_33 vdd gnd cell_6t
Xbit_r34_c17 bl_17 br_17 wl_34 vdd gnd cell_6t
Xbit_r35_c17 bl_17 br_17 wl_35 vdd gnd cell_6t
Xbit_r36_c17 bl_17 br_17 wl_36 vdd gnd cell_6t
Xbit_r37_c17 bl_17 br_17 wl_37 vdd gnd cell_6t
Xbit_r38_c17 bl_17 br_17 wl_38 vdd gnd cell_6t
Xbit_r39_c17 bl_17 br_17 wl_39 vdd gnd cell_6t
Xbit_r40_c17 bl_17 br_17 wl_40 vdd gnd cell_6t
Xbit_r41_c17 bl_17 br_17 wl_41 vdd gnd cell_6t
Xbit_r42_c17 bl_17 br_17 wl_42 vdd gnd cell_6t
Xbit_r43_c17 bl_17 br_17 wl_43 vdd gnd cell_6t
Xbit_r44_c17 bl_17 br_17 wl_44 vdd gnd cell_6t
Xbit_r45_c17 bl_17 br_17 wl_45 vdd gnd cell_6t
Xbit_r46_c17 bl_17 br_17 wl_46 vdd gnd cell_6t
Xbit_r47_c17 bl_17 br_17 wl_47 vdd gnd cell_6t
Xbit_r48_c17 bl_17 br_17 wl_48 vdd gnd cell_6t
Xbit_r49_c17 bl_17 br_17 wl_49 vdd gnd cell_6t
Xbit_r50_c17 bl_17 br_17 wl_50 vdd gnd cell_6t
Xbit_r51_c17 bl_17 br_17 wl_51 vdd gnd cell_6t
Xbit_r52_c17 bl_17 br_17 wl_52 vdd gnd cell_6t
Xbit_r53_c17 bl_17 br_17 wl_53 vdd gnd cell_6t
Xbit_r54_c17 bl_17 br_17 wl_54 vdd gnd cell_6t
Xbit_r55_c17 bl_17 br_17 wl_55 vdd gnd cell_6t
Xbit_r56_c17 bl_17 br_17 wl_56 vdd gnd cell_6t
Xbit_r57_c17 bl_17 br_17 wl_57 vdd gnd cell_6t
Xbit_r58_c17 bl_17 br_17 wl_58 vdd gnd cell_6t
Xbit_r59_c17 bl_17 br_17 wl_59 vdd gnd cell_6t
Xbit_r60_c17 bl_17 br_17 wl_60 vdd gnd cell_6t
Xbit_r61_c17 bl_17 br_17 wl_61 vdd gnd cell_6t
Xbit_r62_c17 bl_17 br_17 wl_62 vdd gnd cell_6t
Xbit_r63_c17 bl_17 br_17 wl_63 vdd gnd cell_6t
Xbit_r64_c17 bl_17 br_17 wl_64 vdd gnd cell_6t
Xbit_r65_c17 bl_17 br_17 wl_65 vdd gnd cell_6t
Xbit_r66_c17 bl_17 br_17 wl_66 vdd gnd cell_6t
Xbit_r67_c17 bl_17 br_17 wl_67 vdd gnd cell_6t
Xbit_r68_c17 bl_17 br_17 wl_68 vdd gnd cell_6t
Xbit_r69_c17 bl_17 br_17 wl_69 vdd gnd cell_6t
Xbit_r70_c17 bl_17 br_17 wl_70 vdd gnd cell_6t
Xbit_r71_c17 bl_17 br_17 wl_71 vdd gnd cell_6t
Xbit_r72_c17 bl_17 br_17 wl_72 vdd gnd cell_6t
Xbit_r73_c17 bl_17 br_17 wl_73 vdd gnd cell_6t
Xbit_r74_c17 bl_17 br_17 wl_74 vdd gnd cell_6t
Xbit_r75_c17 bl_17 br_17 wl_75 vdd gnd cell_6t
Xbit_r76_c17 bl_17 br_17 wl_76 vdd gnd cell_6t
Xbit_r77_c17 bl_17 br_17 wl_77 vdd gnd cell_6t
Xbit_r78_c17 bl_17 br_17 wl_78 vdd gnd cell_6t
Xbit_r79_c17 bl_17 br_17 wl_79 vdd gnd cell_6t
Xbit_r80_c17 bl_17 br_17 wl_80 vdd gnd cell_6t
Xbit_r81_c17 bl_17 br_17 wl_81 vdd gnd cell_6t
Xbit_r82_c17 bl_17 br_17 wl_82 vdd gnd cell_6t
Xbit_r83_c17 bl_17 br_17 wl_83 vdd gnd cell_6t
Xbit_r84_c17 bl_17 br_17 wl_84 vdd gnd cell_6t
Xbit_r85_c17 bl_17 br_17 wl_85 vdd gnd cell_6t
Xbit_r86_c17 bl_17 br_17 wl_86 vdd gnd cell_6t
Xbit_r87_c17 bl_17 br_17 wl_87 vdd gnd cell_6t
Xbit_r88_c17 bl_17 br_17 wl_88 vdd gnd cell_6t
Xbit_r89_c17 bl_17 br_17 wl_89 vdd gnd cell_6t
Xbit_r90_c17 bl_17 br_17 wl_90 vdd gnd cell_6t
Xbit_r91_c17 bl_17 br_17 wl_91 vdd gnd cell_6t
Xbit_r92_c17 bl_17 br_17 wl_92 vdd gnd cell_6t
Xbit_r93_c17 bl_17 br_17 wl_93 vdd gnd cell_6t
Xbit_r94_c17 bl_17 br_17 wl_94 vdd gnd cell_6t
Xbit_r95_c17 bl_17 br_17 wl_95 vdd gnd cell_6t
Xbit_r96_c17 bl_17 br_17 wl_96 vdd gnd cell_6t
Xbit_r97_c17 bl_17 br_17 wl_97 vdd gnd cell_6t
Xbit_r98_c17 bl_17 br_17 wl_98 vdd gnd cell_6t
Xbit_r99_c17 bl_17 br_17 wl_99 vdd gnd cell_6t
Xbit_r100_c17 bl_17 br_17 wl_100 vdd gnd cell_6t
Xbit_r101_c17 bl_17 br_17 wl_101 vdd gnd cell_6t
Xbit_r102_c17 bl_17 br_17 wl_102 vdd gnd cell_6t
Xbit_r103_c17 bl_17 br_17 wl_103 vdd gnd cell_6t
Xbit_r104_c17 bl_17 br_17 wl_104 vdd gnd cell_6t
Xbit_r105_c17 bl_17 br_17 wl_105 vdd gnd cell_6t
Xbit_r106_c17 bl_17 br_17 wl_106 vdd gnd cell_6t
Xbit_r107_c17 bl_17 br_17 wl_107 vdd gnd cell_6t
Xbit_r108_c17 bl_17 br_17 wl_108 vdd gnd cell_6t
Xbit_r109_c17 bl_17 br_17 wl_109 vdd gnd cell_6t
Xbit_r110_c17 bl_17 br_17 wl_110 vdd gnd cell_6t
Xbit_r111_c17 bl_17 br_17 wl_111 vdd gnd cell_6t
Xbit_r112_c17 bl_17 br_17 wl_112 vdd gnd cell_6t
Xbit_r113_c17 bl_17 br_17 wl_113 vdd gnd cell_6t
Xbit_r114_c17 bl_17 br_17 wl_114 vdd gnd cell_6t
Xbit_r115_c17 bl_17 br_17 wl_115 vdd gnd cell_6t
Xbit_r116_c17 bl_17 br_17 wl_116 vdd gnd cell_6t
Xbit_r117_c17 bl_17 br_17 wl_117 vdd gnd cell_6t
Xbit_r118_c17 bl_17 br_17 wl_118 vdd gnd cell_6t
Xbit_r119_c17 bl_17 br_17 wl_119 vdd gnd cell_6t
Xbit_r120_c17 bl_17 br_17 wl_120 vdd gnd cell_6t
Xbit_r121_c17 bl_17 br_17 wl_121 vdd gnd cell_6t
Xbit_r122_c17 bl_17 br_17 wl_122 vdd gnd cell_6t
Xbit_r123_c17 bl_17 br_17 wl_123 vdd gnd cell_6t
Xbit_r124_c17 bl_17 br_17 wl_124 vdd gnd cell_6t
Xbit_r125_c17 bl_17 br_17 wl_125 vdd gnd cell_6t
Xbit_r126_c17 bl_17 br_17 wl_126 vdd gnd cell_6t
Xbit_r127_c17 bl_17 br_17 wl_127 vdd gnd cell_6t
Xbit_r128_c17 bl_17 br_17 wl_128 vdd gnd cell_6t
Xbit_r129_c17 bl_17 br_17 wl_129 vdd gnd cell_6t
Xbit_r130_c17 bl_17 br_17 wl_130 vdd gnd cell_6t
Xbit_r131_c17 bl_17 br_17 wl_131 vdd gnd cell_6t
Xbit_r132_c17 bl_17 br_17 wl_132 vdd gnd cell_6t
Xbit_r133_c17 bl_17 br_17 wl_133 vdd gnd cell_6t
Xbit_r134_c17 bl_17 br_17 wl_134 vdd gnd cell_6t
Xbit_r135_c17 bl_17 br_17 wl_135 vdd gnd cell_6t
Xbit_r136_c17 bl_17 br_17 wl_136 vdd gnd cell_6t
Xbit_r137_c17 bl_17 br_17 wl_137 vdd gnd cell_6t
Xbit_r138_c17 bl_17 br_17 wl_138 vdd gnd cell_6t
Xbit_r139_c17 bl_17 br_17 wl_139 vdd gnd cell_6t
Xbit_r140_c17 bl_17 br_17 wl_140 vdd gnd cell_6t
Xbit_r141_c17 bl_17 br_17 wl_141 vdd gnd cell_6t
Xbit_r142_c17 bl_17 br_17 wl_142 vdd gnd cell_6t
Xbit_r143_c17 bl_17 br_17 wl_143 vdd gnd cell_6t
Xbit_r144_c17 bl_17 br_17 wl_144 vdd gnd cell_6t
Xbit_r145_c17 bl_17 br_17 wl_145 vdd gnd cell_6t
Xbit_r146_c17 bl_17 br_17 wl_146 vdd gnd cell_6t
Xbit_r147_c17 bl_17 br_17 wl_147 vdd gnd cell_6t
Xbit_r148_c17 bl_17 br_17 wl_148 vdd gnd cell_6t
Xbit_r149_c17 bl_17 br_17 wl_149 vdd gnd cell_6t
Xbit_r150_c17 bl_17 br_17 wl_150 vdd gnd cell_6t
Xbit_r151_c17 bl_17 br_17 wl_151 vdd gnd cell_6t
Xbit_r152_c17 bl_17 br_17 wl_152 vdd gnd cell_6t
Xbit_r153_c17 bl_17 br_17 wl_153 vdd gnd cell_6t
Xbit_r154_c17 bl_17 br_17 wl_154 vdd gnd cell_6t
Xbit_r155_c17 bl_17 br_17 wl_155 vdd gnd cell_6t
Xbit_r156_c17 bl_17 br_17 wl_156 vdd gnd cell_6t
Xbit_r157_c17 bl_17 br_17 wl_157 vdd gnd cell_6t
Xbit_r158_c17 bl_17 br_17 wl_158 vdd gnd cell_6t
Xbit_r159_c17 bl_17 br_17 wl_159 vdd gnd cell_6t
Xbit_r160_c17 bl_17 br_17 wl_160 vdd gnd cell_6t
Xbit_r161_c17 bl_17 br_17 wl_161 vdd gnd cell_6t
Xbit_r162_c17 bl_17 br_17 wl_162 vdd gnd cell_6t
Xbit_r163_c17 bl_17 br_17 wl_163 vdd gnd cell_6t
Xbit_r164_c17 bl_17 br_17 wl_164 vdd gnd cell_6t
Xbit_r165_c17 bl_17 br_17 wl_165 vdd gnd cell_6t
Xbit_r166_c17 bl_17 br_17 wl_166 vdd gnd cell_6t
Xbit_r167_c17 bl_17 br_17 wl_167 vdd gnd cell_6t
Xbit_r168_c17 bl_17 br_17 wl_168 vdd gnd cell_6t
Xbit_r169_c17 bl_17 br_17 wl_169 vdd gnd cell_6t
Xbit_r170_c17 bl_17 br_17 wl_170 vdd gnd cell_6t
Xbit_r171_c17 bl_17 br_17 wl_171 vdd gnd cell_6t
Xbit_r172_c17 bl_17 br_17 wl_172 vdd gnd cell_6t
Xbit_r173_c17 bl_17 br_17 wl_173 vdd gnd cell_6t
Xbit_r174_c17 bl_17 br_17 wl_174 vdd gnd cell_6t
Xbit_r175_c17 bl_17 br_17 wl_175 vdd gnd cell_6t
Xbit_r176_c17 bl_17 br_17 wl_176 vdd gnd cell_6t
Xbit_r177_c17 bl_17 br_17 wl_177 vdd gnd cell_6t
Xbit_r178_c17 bl_17 br_17 wl_178 vdd gnd cell_6t
Xbit_r179_c17 bl_17 br_17 wl_179 vdd gnd cell_6t
Xbit_r180_c17 bl_17 br_17 wl_180 vdd gnd cell_6t
Xbit_r181_c17 bl_17 br_17 wl_181 vdd gnd cell_6t
Xbit_r182_c17 bl_17 br_17 wl_182 vdd gnd cell_6t
Xbit_r183_c17 bl_17 br_17 wl_183 vdd gnd cell_6t
Xbit_r184_c17 bl_17 br_17 wl_184 vdd gnd cell_6t
Xbit_r185_c17 bl_17 br_17 wl_185 vdd gnd cell_6t
Xbit_r186_c17 bl_17 br_17 wl_186 vdd gnd cell_6t
Xbit_r187_c17 bl_17 br_17 wl_187 vdd gnd cell_6t
Xbit_r188_c17 bl_17 br_17 wl_188 vdd gnd cell_6t
Xbit_r189_c17 bl_17 br_17 wl_189 vdd gnd cell_6t
Xbit_r190_c17 bl_17 br_17 wl_190 vdd gnd cell_6t
Xbit_r191_c17 bl_17 br_17 wl_191 vdd gnd cell_6t
Xbit_r192_c17 bl_17 br_17 wl_192 vdd gnd cell_6t
Xbit_r193_c17 bl_17 br_17 wl_193 vdd gnd cell_6t
Xbit_r194_c17 bl_17 br_17 wl_194 vdd gnd cell_6t
Xbit_r195_c17 bl_17 br_17 wl_195 vdd gnd cell_6t
Xbit_r196_c17 bl_17 br_17 wl_196 vdd gnd cell_6t
Xbit_r197_c17 bl_17 br_17 wl_197 vdd gnd cell_6t
Xbit_r198_c17 bl_17 br_17 wl_198 vdd gnd cell_6t
Xbit_r199_c17 bl_17 br_17 wl_199 vdd gnd cell_6t
Xbit_r200_c17 bl_17 br_17 wl_200 vdd gnd cell_6t
Xbit_r201_c17 bl_17 br_17 wl_201 vdd gnd cell_6t
Xbit_r202_c17 bl_17 br_17 wl_202 vdd gnd cell_6t
Xbit_r203_c17 bl_17 br_17 wl_203 vdd gnd cell_6t
Xbit_r204_c17 bl_17 br_17 wl_204 vdd gnd cell_6t
Xbit_r205_c17 bl_17 br_17 wl_205 vdd gnd cell_6t
Xbit_r206_c17 bl_17 br_17 wl_206 vdd gnd cell_6t
Xbit_r207_c17 bl_17 br_17 wl_207 vdd gnd cell_6t
Xbit_r208_c17 bl_17 br_17 wl_208 vdd gnd cell_6t
Xbit_r209_c17 bl_17 br_17 wl_209 vdd gnd cell_6t
Xbit_r210_c17 bl_17 br_17 wl_210 vdd gnd cell_6t
Xbit_r211_c17 bl_17 br_17 wl_211 vdd gnd cell_6t
Xbit_r212_c17 bl_17 br_17 wl_212 vdd gnd cell_6t
Xbit_r213_c17 bl_17 br_17 wl_213 vdd gnd cell_6t
Xbit_r214_c17 bl_17 br_17 wl_214 vdd gnd cell_6t
Xbit_r215_c17 bl_17 br_17 wl_215 vdd gnd cell_6t
Xbit_r216_c17 bl_17 br_17 wl_216 vdd gnd cell_6t
Xbit_r217_c17 bl_17 br_17 wl_217 vdd gnd cell_6t
Xbit_r218_c17 bl_17 br_17 wl_218 vdd gnd cell_6t
Xbit_r219_c17 bl_17 br_17 wl_219 vdd gnd cell_6t
Xbit_r220_c17 bl_17 br_17 wl_220 vdd gnd cell_6t
Xbit_r221_c17 bl_17 br_17 wl_221 vdd gnd cell_6t
Xbit_r222_c17 bl_17 br_17 wl_222 vdd gnd cell_6t
Xbit_r223_c17 bl_17 br_17 wl_223 vdd gnd cell_6t
Xbit_r224_c17 bl_17 br_17 wl_224 vdd gnd cell_6t
Xbit_r225_c17 bl_17 br_17 wl_225 vdd gnd cell_6t
Xbit_r226_c17 bl_17 br_17 wl_226 vdd gnd cell_6t
Xbit_r227_c17 bl_17 br_17 wl_227 vdd gnd cell_6t
Xbit_r228_c17 bl_17 br_17 wl_228 vdd gnd cell_6t
Xbit_r229_c17 bl_17 br_17 wl_229 vdd gnd cell_6t
Xbit_r230_c17 bl_17 br_17 wl_230 vdd gnd cell_6t
Xbit_r231_c17 bl_17 br_17 wl_231 vdd gnd cell_6t
Xbit_r232_c17 bl_17 br_17 wl_232 vdd gnd cell_6t
Xbit_r233_c17 bl_17 br_17 wl_233 vdd gnd cell_6t
Xbit_r234_c17 bl_17 br_17 wl_234 vdd gnd cell_6t
Xbit_r235_c17 bl_17 br_17 wl_235 vdd gnd cell_6t
Xbit_r236_c17 bl_17 br_17 wl_236 vdd gnd cell_6t
Xbit_r237_c17 bl_17 br_17 wl_237 vdd gnd cell_6t
Xbit_r238_c17 bl_17 br_17 wl_238 vdd gnd cell_6t
Xbit_r239_c17 bl_17 br_17 wl_239 vdd gnd cell_6t
Xbit_r240_c17 bl_17 br_17 wl_240 vdd gnd cell_6t
Xbit_r241_c17 bl_17 br_17 wl_241 vdd gnd cell_6t
Xbit_r242_c17 bl_17 br_17 wl_242 vdd gnd cell_6t
Xbit_r243_c17 bl_17 br_17 wl_243 vdd gnd cell_6t
Xbit_r244_c17 bl_17 br_17 wl_244 vdd gnd cell_6t
Xbit_r245_c17 bl_17 br_17 wl_245 vdd gnd cell_6t
Xbit_r246_c17 bl_17 br_17 wl_246 vdd gnd cell_6t
Xbit_r247_c17 bl_17 br_17 wl_247 vdd gnd cell_6t
Xbit_r248_c17 bl_17 br_17 wl_248 vdd gnd cell_6t
Xbit_r249_c17 bl_17 br_17 wl_249 vdd gnd cell_6t
Xbit_r250_c17 bl_17 br_17 wl_250 vdd gnd cell_6t
Xbit_r251_c17 bl_17 br_17 wl_251 vdd gnd cell_6t
Xbit_r252_c17 bl_17 br_17 wl_252 vdd gnd cell_6t
Xbit_r253_c17 bl_17 br_17 wl_253 vdd gnd cell_6t
Xbit_r254_c17 bl_17 br_17 wl_254 vdd gnd cell_6t
Xbit_r255_c17 bl_17 br_17 wl_255 vdd gnd cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd cell_6t
Xbit_r1_c18 bl_18 br_18 wl_1 vdd gnd cell_6t
Xbit_r2_c18 bl_18 br_18 wl_2 vdd gnd cell_6t
Xbit_r3_c18 bl_18 br_18 wl_3 vdd gnd cell_6t
Xbit_r4_c18 bl_18 br_18 wl_4 vdd gnd cell_6t
Xbit_r5_c18 bl_18 br_18 wl_5 vdd gnd cell_6t
Xbit_r6_c18 bl_18 br_18 wl_6 vdd gnd cell_6t
Xbit_r7_c18 bl_18 br_18 wl_7 vdd gnd cell_6t
Xbit_r8_c18 bl_18 br_18 wl_8 vdd gnd cell_6t
Xbit_r9_c18 bl_18 br_18 wl_9 vdd gnd cell_6t
Xbit_r10_c18 bl_18 br_18 wl_10 vdd gnd cell_6t
Xbit_r11_c18 bl_18 br_18 wl_11 vdd gnd cell_6t
Xbit_r12_c18 bl_18 br_18 wl_12 vdd gnd cell_6t
Xbit_r13_c18 bl_18 br_18 wl_13 vdd gnd cell_6t
Xbit_r14_c18 bl_18 br_18 wl_14 vdd gnd cell_6t
Xbit_r15_c18 bl_18 br_18 wl_15 vdd gnd cell_6t
Xbit_r16_c18 bl_18 br_18 wl_16 vdd gnd cell_6t
Xbit_r17_c18 bl_18 br_18 wl_17 vdd gnd cell_6t
Xbit_r18_c18 bl_18 br_18 wl_18 vdd gnd cell_6t
Xbit_r19_c18 bl_18 br_18 wl_19 vdd gnd cell_6t
Xbit_r20_c18 bl_18 br_18 wl_20 vdd gnd cell_6t
Xbit_r21_c18 bl_18 br_18 wl_21 vdd gnd cell_6t
Xbit_r22_c18 bl_18 br_18 wl_22 vdd gnd cell_6t
Xbit_r23_c18 bl_18 br_18 wl_23 vdd gnd cell_6t
Xbit_r24_c18 bl_18 br_18 wl_24 vdd gnd cell_6t
Xbit_r25_c18 bl_18 br_18 wl_25 vdd gnd cell_6t
Xbit_r26_c18 bl_18 br_18 wl_26 vdd gnd cell_6t
Xbit_r27_c18 bl_18 br_18 wl_27 vdd gnd cell_6t
Xbit_r28_c18 bl_18 br_18 wl_28 vdd gnd cell_6t
Xbit_r29_c18 bl_18 br_18 wl_29 vdd gnd cell_6t
Xbit_r30_c18 bl_18 br_18 wl_30 vdd gnd cell_6t
Xbit_r31_c18 bl_18 br_18 wl_31 vdd gnd cell_6t
Xbit_r32_c18 bl_18 br_18 wl_32 vdd gnd cell_6t
Xbit_r33_c18 bl_18 br_18 wl_33 vdd gnd cell_6t
Xbit_r34_c18 bl_18 br_18 wl_34 vdd gnd cell_6t
Xbit_r35_c18 bl_18 br_18 wl_35 vdd gnd cell_6t
Xbit_r36_c18 bl_18 br_18 wl_36 vdd gnd cell_6t
Xbit_r37_c18 bl_18 br_18 wl_37 vdd gnd cell_6t
Xbit_r38_c18 bl_18 br_18 wl_38 vdd gnd cell_6t
Xbit_r39_c18 bl_18 br_18 wl_39 vdd gnd cell_6t
Xbit_r40_c18 bl_18 br_18 wl_40 vdd gnd cell_6t
Xbit_r41_c18 bl_18 br_18 wl_41 vdd gnd cell_6t
Xbit_r42_c18 bl_18 br_18 wl_42 vdd gnd cell_6t
Xbit_r43_c18 bl_18 br_18 wl_43 vdd gnd cell_6t
Xbit_r44_c18 bl_18 br_18 wl_44 vdd gnd cell_6t
Xbit_r45_c18 bl_18 br_18 wl_45 vdd gnd cell_6t
Xbit_r46_c18 bl_18 br_18 wl_46 vdd gnd cell_6t
Xbit_r47_c18 bl_18 br_18 wl_47 vdd gnd cell_6t
Xbit_r48_c18 bl_18 br_18 wl_48 vdd gnd cell_6t
Xbit_r49_c18 bl_18 br_18 wl_49 vdd gnd cell_6t
Xbit_r50_c18 bl_18 br_18 wl_50 vdd gnd cell_6t
Xbit_r51_c18 bl_18 br_18 wl_51 vdd gnd cell_6t
Xbit_r52_c18 bl_18 br_18 wl_52 vdd gnd cell_6t
Xbit_r53_c18 bl_18 br_18 wl_53 vdd gnd cell_6t
Xbit_r54_c18 bl_18 br_18 wl_54 vdd gnd cell_6t
Xbit_r55_c18 bl_18 br_18 wl_55 vdd gnd cell_6t
Xbit_r56_c18 bl_18 br_18 wl_56 vdd gnd cell_6t
Xbit_r57_c18 bl_18 br_18 wl_57 vdd gnd cell_6t
Xbit_r58_c18 bl_18 br_18 wl_58 vdd gnd cell_6t
Xbit_r59_c18 bl_18 br_18 wl_59 vdd gnd cell_6t
Xbit_r60_c18 bl_18 br_18 wl_60 vdd gnd cell_6t
Xbit_r61_c18 bl_18 br_18 wl_61 vdd gnd cell_6t
Xbit_r62_c18 bl_18 br_18 wl_62 vdd gnd cell_6t
Xbit_r63_c18 bl_18 br_18 wl_63 vdd gnd cell_6t
Xbit_r64_c18 bl_18 br_18 wl_64 vdd gnd cell_6t
Xbit_r65_c18 bl_18 br_18 wl_65 vdd gnd cell_6t
Xbit_r66_c18 bl_18 br_18 wl_66 vdd gnd cell_6t
Xbit_r67_c18 bl_18 br_18 wl_67 vdd gnd cell_6t
Xbit_r68_c18 bl_18 br_18 wl_68 vdd gnd cell_6t
Xbit_r69_c18 bl_18 br_18 wl_69 vdd gnd cell_6t
Xbit_r70_c18 bl_18 br_18 wl_70 vdd gnd cell_6t
Xbit_r71_c18 bl_18 br_18 wl_71 vdd gnd cell_6t
Xbit_r72_c18 bl_18 br_18 wl_72 vdd gnd cell_6t
Xbit_r73_c18 bl_18 br_18 wl_73 vdd gnd cell_6t
Xbit_r74_c18 bl_18 br_18 wl_74 vdd gnd cell_6t
Xbit_r75_c18 bl_18 br_18 wl_75 vdd gnd cell_6t
Xbit_r76_c18 bl_18 br_18 wl_76 vdd gnd cell_6t
Xbit_r77_c18 bl_18 br_18 wl_77 vdd gnd cell_6t
Xbit_r78_c18 bl_18 br_18 wl_78 vdd gnd cell_6t
Xbit_r79_c18 bl_18 br_18 wl_79 vdd gnd cell_6t
Xbit_r80_c18 bl_18 br_18 wl_80 vdd gnd cell_6t
Xbit_r81_c18 bl_18 br_18 wl_81 vdd gnd cell_6t
Xbit_r82_c18 bl_18 br_18 wl_82 vdd gnd cell_6t
Xbit_r83_c18 bl_18 br_18 wl_83 vdd gnd cell_6t
Xbit_r84_c18 bl_18 br_18 wl_84 vdd gnd cell_6t
Xbit_r85_c18 bl_18 br_18 wl_85 vdd gnd cell_6t
Xbit_r86_c18 bl_18 br_18 wl_86 vdd gnd cell_6t
Xbit_r87_c18 bl_18 br_18 wl_87 vdd gnd cell_6t
Xbit_r88_c18 bl_18 br_18 wl_88 vdd gnd cell_6t
Xbit_r89_c18 bl_18 br_18 wl_89 vdd gnd cell_6t
Xbit_r90_c18 bl_18 br_18 wl_90 vdd gnd cell_6t
Xbit_r91_c18 bl_18 br_18 wl_91 vdd gnd cell_6t
Xbit_r92_c18 bl_18 br_18 wl_92 vdd gnd cell_6t
Xbit_r93_c18 bl_18 br_18 wl_93 vdd gnd cell_6t
Xbit_r94_c18 bl_18 br_18 wl_94 vdd gnd cell_6t
Xbit_r95_c18 bl_18 br_18 wl_95 vdd gnd cell_6t
Xbit_r96_c18 bl_18 br_18 wl_96 vdd gnd cell_6t
Xbit_r97_c18 bl_18 br_18 wl_97 vdd gnd cell_6t
Xbit_r98_c18 bl_18 br_18 wl_98 vdd gnd cell_6t
Xbit_r99_c18 bl_18 br_18 wl_99 vdd gnd cell_6t
Xbit_r100_c18 bl_18 br_18 wl_100 vdd gnd cell_6t
Xbit_r101_c18 bl_18 br_18 wl_101 vdd gnd cell_6t
Xbit_r102_c18 bl_18 br_18 wl_102 vdd gnd cell_6t
Xbit_r103_c18 bl_18 br_18 wl_103 vdd gnd cell_6t
Xbit_r104_c18 bl_18 br_18 wl_104 vdd gnd cell_6t
Xbit_r105_c18 bl_18 br_18 wl_105 vdd gnd cell_6t
Xbit_r106_c18 bl_18 br_18 wl_106 vdd gnd cell_6t
Xbit_r107_c18 bl_18 br_18 wl_107 vdd gnd cell_6t
Xbit_r108_c18 bl_18 br_18 wl_108 vdd gnd cell_6t
Xbit_r109_c18 bl_18 br_18 wl_109 vdd gnd cell_6t
Xbit_r110_c18 bl_18 br_18 wl_110 vdd gnd cell_6t
Xbit_r111_c18 bl_18 br_18 wl_111 vdd gnd cell_6t
Xbit_r112_c18 bl_18 br_18 wl_112 vdd gnd cell_6t
Xbit_r113_c18 bl_18 br_18 wl_113 vdd gnd cell_6t
Xbit_r114_c18 bl_18 br_18 wl_114 vdd gnd cell_6t
Xbit_r115_c18 bl_18 br_18 wl_115 vdd gnd cell_6t
Xbit_r116_c18 bl_18 br_18 wl_116 vdd gnd cell_6t
Xbit_r117_c18 bl_18 br_18 wl_117 vdd gnd cell_6t
Xbit_r118_c18 bl_18 br_18 wl_118 vdd gnd cell_6t
Xbit_r119_c18 bl_18 br_18 wl_119 vdd gnd cell_6t
Xbit_r120_c18 bl_18 br_18 wl_120 vdd gnd cell_6t
Xbit_r121_c18 bl_18 br_18 wl_121 vdd gnd cell_6t
Xbit_r122_c18 bl_18 br_18 wl_122 vdd gnd cell_6t
Xbit_r123_c18 bl_18 br_18 wl_123 vdd gnd cell_6t
Xbit_r124_c18 bl_18 br_18 wl_124 vdd gnd cell_6t
Xbit_r125_c18 bl_18 br_18 wl_125 vdd gnd cell_6t
Xbit_r126_c18 bl_18 br_18 wl_126 vdd gnd cell_6t
Xbit_r127_c18 bl_18 br_18 wl_127 vdd gnd cell_6t
Xbit_r128_c18 bl_18 br_18 wl_128 vdd gnd cell_6t
Xbit_r129_c18 bl_18 br_18 wl_129 vdd gnd cell_6t
Xbit_r130_c18 bl_18 br_18 wl_130 vdd gnd cell_6t
Xbit_r131_c18 bl_18 br_18 wl_131 vdd gnd cell_6t
Xbit_r132_c18 bl_18 br_18 wl_132 vdd gnd cell_6t
Xbit_r133_c18 bl_18 br_18 wl_133 vdd gnd cell_6t
Xbit_r134_c18 bl_18 br_18 wl_134 vdd gnd cell_6t
Xbit_r135_c18 bl_18 br_18 wl_135 vdd gnd cell_6t
Xbit_r136_c18 bl_18 br_18 wl_136 vdd gnd cell_6t
Xbit_r137_c18 bl_18 br_18 wl_137 vdd gnd cell_6t
Xbit_r138_c18 bl_18 br_18 wl_138 vdd gnd cell_6t
Xbit_r139_c18 bl_18 br_18 wl_139 vdd gnd cell_6t
Xbit_r140_c18 bl_18 br_18 wl_140 vdd gnd cell_6t
Xbit_r141_c18 bl_18 br_18 wl_141 vdd gnd cell_6t
Xbit_r142_c18 bl_18 br_18 wl_142 vdd gnd cell_6t
Xbit_r143_c18 bl_18 br_18 wl_143 vdd gnd cell_6t
Xbit_r144_c18 bl_18 br_18 wl_144 vdd gnd cell_6t
Xbit_r145_c18 bl_18 br_18 wl_145 vdd gnd cell_6t
Xbit_r146_c18 bl_18 br_18 wl_146 vdd gnd cell_6t
Xbit_r147_c18 bl_18 br_18 wl_147 vdd gnd cell_6t
Xbit_r148_c18 bl_18 br_18 wl_148 vdd gnd cell_6t
Xbit_r149_c18 bl_18 br_18 wl_149 vdd gnd cell_6t
Xbit_r150_c18 bl_18 br_18 wl_150 vdd gnd cell_6t
Xbit_r151_c18 bl_18 br_18 wl_151 vdd gnd cell_6t
Xbit_r152_c18 bl_18 br_18 wl_152 vdd gnd cell_6t
Xbit_r153_c18 bl_18 br_18 wl_153 vdd gnd cell_6t
Xbit_r154_c18 bl_18 br_18 wl_154 vdd gnd cell_6t
Xbit_r155_c18 bl_18 br_18 wl_155 vdd gnd cell_6t
Xbit_r156_c18 bl_18 br_18 wl_156 vdd gnd cell_6t
Xbit_r157_c18 bl_18 br_18 wl_157 vdd gnd cell_6t
Xbit_r158_c18 bl_18 br_18 wl_158 vdd gnd cell_6t
Xbit_r159_c18 bl_18 br_18 wl_159 vdd gnd cell_6t
Xbit_r160_c18 bl_18 br_18 wl_160 vdd gnd cell_6t
Xbit_r161_c18 bl_18 br_18 wl_161 vdd gnd cell_6t
Xbit_r162_c18 bl_18 br_18 wl_162 vdd gnd cell_6t
Xbit_r163_c18 bl_18 br_18 wl_163 vdd gnd cell_6t
Xbit_r164_c18 bl_18 br_18 wl_164 vdd gnd cell_6t
Xbit_r165_c18 bl_18 br_18 wl_165 vdd gnd cell_6t
Xbit_r166_c18 bl_18 br_18 wl_166 vdd gnd cell_6t
Xbit_r167_c18 bl_18 br_18 wl_167 vdd gnd cell_6t
Xbit_r168_c18 bl_18 br_18 wl_168 vdd gnd cell_6t
Xbit_r169_c18 bl_18 br_18 wl_169 vdd gnd cell_6t
Xbit_r170_c18 bl_18 br_18 wl_170 vdd gnd cell_6t
Xbit_r171_c18 bl_18 br_18 wl_171 vdd gnd cell_6t
Xbit_r172_c18 bl_18 br_18 wl_172 vdd gnd cell_6t
Xbit_r173_c18 bl_18 br_18 wl_173 vdd gnd cell_6t
Xbit_r174_c18 bl_18 br_18 wl_174 vdd gnd cell_6t
Xbit_r175_c18 bl_18 br_18 wl_175 vdd gnd cell_6t
Xbit_r176_c18 bl_18 br_18 wl_176 vdd gnd cell_6t
Xbit_r177_c18 bl_18 br_18 wl_177 vdd gnd cell_6t
Xbit_r178_c18 bl_18 br_18 wl_178 vdd gnd cell_6t
Xbit_r179_c18 bl_18 br_18 wl_179 vdd gnd cell_6t
Xbit_r180_c18 bl_18 br_18 wl_180 vdd gnd cell_6t
Xbit_r181_c18 bl_18 br_18 wl_181 vdd gnd cell_6t
Xbit_r182_c18 bl_18 br_18 wl_182 vdd gnd cell_6t
Xbit_r183_c18 bl_18 br_18 wl_183 vdd gnd cell_6t
Xbit_r184_c18 bl_18 br_18 wl_184 vdd gnd cell_6t
Xbit_r185_c18 bl_18 br_18 wl_185 vdd gnd cell_6t
Xbit_r186_c18 bl_18 br_18 wl_186 vdd gnd cell_6t
Xbit_r187_c18 bl_18 br_18 wl_187 vdd gnd cell_6t
Xbit_r188_c18 bl_18 br_18 wl_188 vdd gnd cell_6t
Xbit_r189_c18 bl_18 br_18 wl_189 vdd gnd cell_6t
Xbit_r190_c18 bl_18 br_18 wl_190 vdd gnd cell_6t
Xbit_r191_c18 bl_18 br_18 wl_191 vdd gnd cell_6t
Xbit_r192_c18 bl_18 br_18 wl_192 vdd gnd cell_6t
Xbit_r193_c18 bl_18 br_18 wl_193 vdd gnd cell_6t
Xbit_r194_c18 bl_18 br_18 wl_194 vdd gnd cell_6t
Xbit_r195_c18 bl_18 br_18 wl_195 vdd gnd cell_6t
Xbit_r196_c18 bl_18 br_18 wl_196 vdd gnd cell_6t
Xbit_r197_c18 bl_18 br_18 wl_197 vdd gnd cell_6t
Xbit_r198_c18 bl_18 br_18 wl_198 vdd gnd cell_6t
Xbit_r199_c18 bl_18 br_18 wl_199 vdd gnd cell_6t
Xbit_r200_c18 bl_18 br_18 wl_200 vdd gnd cell_6t
Xbit_r201_c18 bl_18 br_18 wl_201 vdd gnd cell_6t
Xbit_r202_c18 bl_18 br_18 wl_202 vdd gnd cell_6t
Xbit_r203_c18 bl_18 br_18 wl_203 vdd gnd cell_6t
Xbit_r204_c18 bl_18 br_18 wl_204 vdd gnd cell_6t
Xbit_r205_c18 bl_18 br_18 wl_205 vdd gnd cell_6t
Xbit_r206_c18 bl_18 br_18 wl_206 vdd gnd cell_6t
Xbit_r207_c18 bl_18 br_18 wl_207 vdd gnd cell_6t
Xbit_r208_c18 bl_18 br_18 wl_208 vdd gnd cell_6t
Xbit_r209_c18 bl_18 br_18 wl_209 vdd gnd cell_6t
Xbit_r210_c18 bl_18 br_18 wl_210 vdd gnd cell_6t
Xbit_r211_c18 bl_18 br_18 wl_211 vdd gnd cell_6t
Xbit_r212_c18 bl_18 br_18 wl_212 vdd gnd cell_6t
Xbit_r213_c18 bl_18 br_18 wl_213 vdd gnd cell_6t
Xbit_r214_c18 bl_18 br_18 wl_214 vdd gnd cell_6t
Xbit_r215_c18 bl_18 br_18 wl_215 vdd gnd cell_6t
Xbit_r216_c18 bl_18 br_18 wl_216 vdd gnd cell_6t
Xbit_r217_c18 bl_18 br_18 wl_217 vdd gnd cell_6t
Xbit_r218_c18 bl_18 br_18 wl_218 vdd gnd cell_6t
Xbit_r219_c18 bl_18 br_18 wl_219 vdd gnd cell_6t
Xbit_r220_c18 bl_18 br_18 wl_220 vdd gnd cell_6t
Xbit_r221_c18 bl_18 br_18 wl_221 vdd gnd cell_6t
Xbit_r222_c18 bl_18 br_18 wl_222 vdd gnd cell_6t
Xbit_r223_c18 bl_18 br_18 wl_223 vdd gnd cell_6t
Xbit_r224_c18 bl_18 br_18 wl_224 vdd gnd cell_6t
Xbit_r225_c18 bl_18 br_18 wl_225 vdd gnd cell_6t
Xbit_r226_c18 bl_18 br_18 wl_226 vdd gnd cell_6t
Xbit_r227_c18 bl_18 br_18 wl_227 vdd gnd cell_6t
Xbit_r228_c18 bl_18 br_18 wl_228 vdd gnd cell_6t
Xbit_r229_c18 bl_18 br_18 wl_229 vdd gnd cell_6t
Xbit_r230_c18 bl_18 br_18 wl_230 vdd gnd cell_6t
Xbit_r231_c18 bl_18 br_18 wl_231 vdd gnd cell_6t
Xbit_r232_c18 bl_18 br_18 wl_232 vdd gnd cell_6t
Xbit_r233_c18 bl_18 br_18 wl_233 vdd gnd cell_6t
Xbit_r234_c18 bl_18 br_18 wl_234 vdd gnd cell_6t
Xbit_r235_c18 bl_18 br_18 wl_235 vdd gnd cell_6t
Xbit_r236_c18 bl_18 br_18 wl_236 vdd gnd cell_6t
Xbit_r237_c18 bl_18 br_18 wl_237 vdd gnd cell_6t
Xbit_r238_c18 bl_18 br_18 wl_238 vdd gnd cell_6t
Xbit_r239_c18 bl_18 br_18 wl_239 vdd gnd cell_6t
Xbit_r240_c18 bl_18 br_18 wl_240 vdd gnd cell_6t
Xbit_r241_c18 bl_18 br_18 wl_241 vdd gnd cell_6t
Xbit_r242_c18 bl_18 br_18 wl_242 vdd gnd cell_6t
Xbit_r243_c18 bl_18 br_18 wl_243 vdd gnd cell_6t
Xbit_r244_c18 bl_18 br_18 wl_244 vdd gnd cell_6t
Xbit_r245_c18 bl_18 br_18 wl_245 vdd gnd cell_6t
Xbit_r246_c18 bl_18 br_18 wl_246 vdd gnd cell_6t
Xbit_r247_c18 bl_18 br_18 wl_247 vdd gnd cell_6t
Xbit_r248_c18 bl_18 br_18 wl_248 vdd gnd cell_6t
Xbit_r249_c18 bl_18 br_18 wl_249 vdd gnd cell_6t
Xbit_r250_c18 bl_18 br_18 wl_250 vdd gnd cell_6t
Xbit_r251_c18 bl_18 br_18 wl_251 vdd gnd cell_6t
Xbit_r252_c18 bl_18 br_18 wl_252 vdd gnd cell_6t
Xbit_r253_c18 bl_18 br_18 wl_253 vdd gnd cell_6t
Xbit_r254_c18 bl_18 br_18 wl_254 vdd gnd cell_6t
Xbit_r255_c18 bl_18 br_18 wl_255 vdd gnd cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd cell_6t
Xbit_r1_c19 bl_19 br_19 wl_1 vdd gnd cell_6t
Xbit_r2_c19 bl_19 br_19 wl_2 vdd gnd cell_6t
Xbit_r3_c19 bl_19 br_19 wl_3 vdd gnd cell_6t
Xbit_r4_c19 bl_19 br_19 wl_4 vdd gnd cell_6t
Xbit_r5_c19 bl_19 br_19 wl_5 vdd gnd cell_6t
Xbit_r6_c19 bl_19 br_19 wl_6 vdd gnd cell_6t
Xbit_r7_c19 bl_19 br_19 wl_7 vdd gnd cell_6t
Xbit_r8_c19 bl_19 br_19 wl_8 vdd gnd cell_6t
Xbit_r9_c19 bl_19 br_19 wl_9 vdd gnd cell_6t
Xbit_r10_c19 bl_19 br_19 wl_10 vdd gnd cell_6t
Xbit_r11_c19 bl_19 br_19 wl_11 vdd gnd cell_6t
Xbit_r12_c19 bl_19 br_19 wl_12 vdd gnd cell_6t
Xbit_r13_c19 bl_19 br_19 wl_13 vdd gnd cell_6t
Xbit_r14_c19 bl_19 br_19 wl_14 vdd gnd cell_6t
Xbit_r15_c19 bl_19 br_19 wl_15 vdd gnd cell_6t
Xbit_r16_c19 bl_19 br_19 wl_16 vdd gnd cell_6t
Xbit_r17_c19 bl_19 br_19 wl_17 vdd gnd cell_6t
Xbit_r18_c19 bl_19 br_19 wl_18 vdd gnd cell_6t
Xbit_r19_c19 bl_19 br_19 wl_19 vdd gnd cell_6t
Xbit_r20_c19 bl_19 br_19 wl_20 vdd gnd cell_6t
Xbit_r21_c19 bl_19 br_19 wl_21 vdd gnd cell_6t
Xbit_r22_c19 bl_19 br_19 wl_22 vdd gnd cell_6t
Xbit_r23_c19 bl_19 br_19 wl_23 vdd gnd cell_6t
Xbit_r24_c19 bl_19 br_19 wl_24 vdd gnd cell_6t
Xbit_r25_c19 bl_19 br_19 wl_25 vdd gnd cell_6t
Xbit_r26_c19 bl_19 br_19 wl_26 vdd gnd cell_6t
Xbit_r27_c19 bl_19 br_19 wl_27 vdd gnd cell_6t
Xbit_r28_c19 bl_19 br_19 wl_28 vdd gnd cell_6t
Xbit_r29_c19 bl_19 br_19 wl_29 vdd gnd cell_6t
Xbit_r30_c19 bl_19 br_19 wl_30 vdd gnd cell_6t
Xbit_r31_c19 bl_19 br_19 wl_31 vdd gnd cell_6t
Xbit_r32_c19 bl_19 br_19 wl_32 vdd gnd cell_6t
Xbit_r33_c19 bl_19 br_19 wl_33 vdd gnd cell_6t
Xbit_r34_c19 bl_19 br_19 wl_34 vdd gnd cell_6t
Xbit_r35_c19 bl_19 br_19 wl_35 vdd gnd cell_6t
Xbit_r36_c19 bl_19 br_19 wl_36 vdd gnd cell_6t
Xbit_r37_c19 bl_19 br_19 wl_37 vdd gnd cell_6t
Xbit_r38_c19 bl_19 br_19 wl_38 vdd gnd cell_6t
Xbit_r39_c19 bl_19 br_19 wl_39 vdd gnd cell_6t
Xbit_r40_c19 bl_19 br_19 wl_40 vdd gnd cell_6t
Xbit_r41_c19 bl_19 br_19 wl_41 vdd gnd cell_6t
Xbit_r42_c19 bl_19 br_19 wl_42 vdd gnd cell_6t
Xbit_r43_c19 bl_19 br_19 wl_43 vdd gnd cell_6t
Xbit_r44_c19 bl_19 br_19 wl_44 vdd gnd cell_6t
Xbit_r45_c19 bl_19 br_19 wl_45 vdd gnd cell_6t
Xbit_r46_c19 bl_19 br_19 wl_46 vdd gnd cell_6t
Xbit_r47_c19 bl_19 br_19 wl_47 vdd gnd cell_6t
Xbit_r48_c19 bl_19 br_19 wl_48 vdd gnd cell_6t
Xbit_r49_c19 bl_19 br_19 wl_49 vdd gnd cell_6t
Xbit_r50_c19 bl_19 br_19 wl_50 vdd gnd cell_6t
Xbit_r51_c19 bl_19 br_19 wl_51 vdd gnd cell_6t
Xbit_r52_c19 bl_19 br_19 wl_52 vdd gnd cell_6t
Xbit_r53_c19 bl_19 br_19 wl_53 vdd gnd cell_6t
Xbit_r54_c19 bl_19 br_19 wl_54 vdd gnd cell_6t
Xbit_r55_c19 bl_19 br_19 wl_55 vdd gnd cell_6t
Xbit_r56_c19 bl_19 br_19 wl_56 vdd gnd cell_6t
Xbit_r57_c19 bl_19 br_19 wl_57 vdd gnd cell_6t
Xbit_r58_c19 bl_19 br_19 wl_58 vdd gnd cell_6t
Xbit_r59_c19 bl_19 br_19 wl_59 vdd gnd cell_6t
Xbit_r60_c19 bl_19 br_19 wl_60 vdd gnd cell_6t
Xbit_r61_c19 bl_19 br_19 wl_61 vdd gnd cell_6t
Xbit_r62_c19 bl_19 br_19 wl_62 vdd gnd cell_6t
Xbit_r63_c19 bl_19 br_19 wl_63 vdd gnd cell_6t
Xbit_r64_c19 bl_19 br_19 wl_64 vdd gnd cell_6t
Xbit_r65_c19 bl_19 br_19 wl_65 vdd gnd cell_6t
Xbit_r66_c19 bl_19 br_19 wl_66 vdd gnd cell_6t
Xbit_r67_c19 bl_19 br_19 wl_67 vdd gnd cell_6t
Xbit_r68_c19 bl_19 br_19 wl_68 vdd gnd cell_6t
Xbit_r69_c19 bl_19 br_19 wl_69 vdd gnd cell_6t
Xbit_r70_c19 bl_19 br_19 wl_70 vdd gnd cell_6t
Xbit_r71_c19 bl_19 br_19 wl_71 vdd gnd cell_6t
Xbit_r72_c19 bl_19 br_19 wl_72 vdd gnd cell_6t
Xbit_r73_c19 bl_19 br_19 wl_73 vdd gnd cell_6t
Xbit_r74_c19 bl_19 br_19 wl_74 vdd gnd cell_6t
Xbit_r75_c19 bl_19 br_19 wl_75 vdd gnd cell_6t
Xbit_r76_c19 bl_19 br_19 wl_76 vdd gnd cell_6t
Xbit_r77_c19 bl_19 br_19 wl_77 vdd gnd cell_6t
Xbit_r78_c19 bl_19 br_19 wl_78 vdd gnd cell_6t
Xbit_r79_c19 bl_19 br_19 wl_79 vdd gnd cell_6t
Xbit_r80_c19 bl_19 br_19 wl_80 vdd gnd cell_6t
Xbit_r81_c19 bl_19 br_19 wl_81 vdd gnd cell_6t
Xbit_r82_c19 bl_19 br_19 wl_82 vdd gnd cell_6t
Xbit_r83_c19 bl_19 br_19 wl_83 vdd gnd cell_6t
Xbit_r84_c19 bl_19 br_19 wl_84 vdd gnd cell_6t
Xbit_r85_c19 bl_19 br_19 wl_85 vdd gnd cell_6t
Xbit_r86_c19 bl_19 br_19 wl_86 vdd gnd cell_6t
Xbit_r87_c19 bl_19 br_19 wl_87 vdd gnd cell_6t
Xbit_r88_c19 bl_19 br_19 wl_88 vdd gnd cell_6t
Xbit_r89_c19 bl_19 br_19 wl_89 vdd gnd cell_6t
Xbit_r90_c19 bl_19 br_19 wl_90 vdd gnd cell_6t
Xbit_r91_c19 bl_19 br_19 wl_91 vdd gnd cell_6t
Xbit_r92_c19 bl_19 br_19 wl_92 vdd gnd cell_6t
Xbit_r93_c19 bl_19 br_19 wl_93 vdd gnd cell_6t
Xbit_r94_c19 bl_19 br_19 wl_94 vdd gnd cell_6t
Xbit_r95_c19 bl_19 br_19 wl_95 vdd gnd cell_6t
Xbit_r96_c19 bl_19 br_19 wl_96 vdd gnd cell_6t
Xbit_r97_c19 bl_19 br_19 wl_97 vdd gnd cell_6t
Xbit_r98_c19 bl_19 br_19 wl_98 vdd gnd cell_6t
Xbit_r99_c19 bl_19 br_19 wl_99 vdd gnd cell_6t
Xbit_r100_c19 bl_19 br_19 wl_100 vdd gnd cell_6t
Xbit_r101_c19 bl_19 br_19 wl_101 vdd gnd cell_6t
Xbit_r102_c19 bl_19 br_19 wl_102 vdd gnd cell_6t
Xbit_r103_c19 bl_19 br_19 wl_103 vdd gnd cell_6t
Xbit_r104_c19 bl_19 br_19 wl_104 vdd gnd cell_6t
Xbit_r105_c19 bl_19 br_19 wl_105 vdd gnd cell_6t
Xbit_r106_c19 bl_19 br_19 wl_106 vdd gnd cell_6t
Xbit_r107_c19 bl_19 br_19 wl_107 vdd gnd cell_6t
Xbit_r108_c19 bl_19 br_19 wl_108 vdd gnd cell_6t
Xbit_r109_c19 bl_19 br_19 wl_109 vdd gnd cell_6t
Xbit_r110_c19 bl_19 br_19 wl_110 vdd gnd cell_6t
Xbit_r111_c19 bl_19 br_19 wl_111 vdd gnd cell_6t
Xbit_r112_c19 bl_19 br_19 wl_112 vdd gnd cell_6t
Xbit_r113_c19 bl_19 br_19 wl_113 vdd gnd cell_6t
Xbit_r114_c19 bl_19 br_19 wl_114 vdd gnd cell_6t
Xbit_r115_c19 bl_19 br_19 wl_115 vdd gnd cell_6t
Xbit_r116_c19 bl_19 br_19 wl_116 vdd gnd cell_6t
Xbit_r117_c19 bl_19 br_19 wl_117 vdd gnd cell_6t
Xbit_r118_c19 bl_19 br_19 wl_118 vdd gnd cell_6t
Xbit_r119_c19 bl_19 br_19 wl_119 vdd gnd cell_6t
Xbit_r120_c19 bl_19 br_19 wl_120 vdd gnd cell_6t
Xbit_r121_c19 bl_19 br_19 wl_121 vdd gnd cell_6t
Xbit_r122_c19 bl_19 br_19 wl_122 vdd gnd cell_6t
Xbit_r123_c19 bl_19 br_19 wl_123 vdd gnd cell_6t
Xbit_r124_c19 bl_19 br_19 wl_124 vdd gnd cell_6t
Xbit_r125_c19 bl_19 br_19 wl_125 vdd gnd cell_6t
Xbit_r126_c19 bl_19 br_19 wl_126 vdd gnd cell_6t
Xbit_r127_c19 bl_19 br_19 wl_127 vdd gnd cell_6t
Xbit_r128_c19 bl_19 br_19 wl_128 vdd gnd cell_6t
Xbit_r129_c19 bl_19 br_19 wl_129 vdd gnd cell_6t
Xbit_r130_c19 bl_19 br_19 wl_130 vdd gnd cell_6t
Xbit_r131_c19 bl_19 br_19 wl_131 vdd gnd cell_6t
Xbit_r132_c19 bl_19 br_19 wl_132 vdd gnd cell_6t
Xbit_r133_c19 bl_19 br_19 wl_133 vdd gnd cell_6t
Xbit_r134_c19 bl_19 br_19 wl_134 vdd gnd cell_6t
Xbit_r135_c19 bl_19 br_19 wl_135 vdd gnd cell_6t
Xbit_r136_c19 bl_19 br_19 wl_136 vdd gnd cell_6t
Xbit_r137_c19 bl_19 br_19 wl_137 vdd gnd cell_6t
Xbit_r138_c19 bl_19 br_19 wl_138 vdd gnd cell_6t
Xbit_r139_c19 bl_19 br_19 wl_139 vdd gnd cell_6t
Xbit_r140_c19 bl_19 br_19 wl_140 vdd gnd cell_6t
Xbit_r141_c19 bl_19 br_19 wl_141 vdd gnd cell_6t
Xbit_r142_c19 bl_19 br_19 wl_142 vdd gnd cell_6t
Xbit_r143_c19 bl_19 br_19 wl_143 vdd gnd cell_6t
Xbit_r144_c19 bl_19 br_19 wl_144 vdd gnd cell_6t
Xbit_r145_c19 bl_19 br_19 wl_145 vdd gnd cell_6t
Xbit_r146_c19 bl_19 br_19 wl_146 vdd gnd cell_6t
Xbit_r147_c19 bl_19 br_19 wl_147 vdd gnd cell_6t
Xbit_r148_c19 bl_19 br_19 wl_148 vdd gnd cell_6t
Xbit_r149_c19 bl_19 br_19 wl_149 vdd gnd cell_6t
Xbit_r150_c19 bl_19 br_19 wl_150 vdd gnd cell_6t
Xbit_r151_c19 bl_19 br_19 wl_151 vdd gnd cell_6t
Xbit_r152_c19 bl_19 br_19 wl_152 vdd gnd cell_6t
Xbit_r153_c19 bl_19 br_19 wl_153 vdd gnd cell_6t
Xbit_r154_c19 bl_19 br_19 wl_154 vdd gnd cell_6t
Xbit_r155_c19 bl_19 br_19 wl_155 vdd gnd cell_6t
Xbit_r156_c19 bl_19 br_19 wl_156 vdd gnd cell_6t
Xbit_r157_c19 bl_19 br_19 wl_157 vdd gnd cell_6t
Xbit_r158_c19 bl_19 br_19 wl_158 vdd gnd cell_6t
Xbit_r159_c19 bl_19 br_19 wl_159 vdd gnd cell_6t
Xbit_r160_c19 bl_19 br_19 wl_160 vdd gnd cell_6t
Xbit_r161_c19 bl_19 br_19 wl_161 vdd gnd cell_6t
Xbit_r162_c19 bl_19 br_19 wl_162 vdd gnd cell_6t
Xbit_r163_c19 bl_19 br_19 wl_163 vdd gnd cell_6t
Xbit_r164_c19 bl_19 br_19 wl_164 vdd gnd cell_6t
Xbit_r165_c19 bl_19 br_19 wl_165 vdd gnd cell_6t
Xbit_r166_c19 bl_19 br_19 wl_166 vdd gnd cell_6t
Xbit_r167_c19 bl_19 br_19 wl_167 vdd gnd cell_6t
Xbit_r168_c19 bl_19 br_19 wl_168 vdd gnd cell_6t
Xbit_r169_c19 bl_19 br_19 wl_169 vdd gnd cell_6t
Xbit_r170_c19 bl_19 br_19 wl_170 vdd gnd cell_6t
Xbit_r171_c19 bl_19 br_19 wl_171 vdd gnd cell_6t
Xbit_r172_c19 bl_19 br_19 wl_172 vdd gnd cell_6t
Xbit_r173_c19 bl_19 br_19 wl_173 vdd gnd cell_6t
Xbit_r174_c19 bl_19 br_19 wl_174 vdd gnd cell_6t
Xbit_r175_c19 bl_19 br_19 wl_175 vdd gnd cell_6t
Xbit_r176_c19 bl_19 br_19 wl_176 vdd gnd cell_6t
Xbit_r177_c19 bl_19 br_19 wl_177 vdd gnd cell_6t
Xbit_r178_c19 bl_19 br_19 wl_178 vdd gnd cell_6t
Xbit_r179_c19 bl_19 br_19 wl_179 vdd gnd cell_6t
Xbit_r180_c19 bl_19 br_19 wl_180 vdd gnd cell_6t
Xbit_r181_c19 bl_19 br_19 wl_181 vdd gnd cell_6t
Xbit_r182_c19 bl_19 br_19 wl_182 vdd gnd cell_6t
Xbit_r183_c19 bl_19 br_19 wl_183 vdd gnd cell_6t
Xbit_r184_c19 bl_19 br_19 wl_184 vdd gnd cell_6t
Xbit_r185_c19 bl_19 br_19 wl_185 vdd gnd cell_6t
Xbit_r186_c19 bl_19 br_19 wl_186 vdd gnd cell_6t
Xbit_r187_c19 bl_19 br_19 wl_187 vdd gnd cell_6t
Xbit_r188_c19 bl_19 br_19 wl_188 vdd gnd cell_6t
Xbit_r189_c19 bl_19 br_19 wl_189 vdd gnd cell_6t
Xbit_r190_c19 bl_19 br_19 wl_190 vdd gnd cell_6t
Xbit_r191_c19 bl_19 br_19 wl_191 vdd gnd cell_6t
Xbit_r192_c19 bl_19 br_19 wl_192 vdd gnd cell_6t
Xbit_r193_c19 bl_19 br_19 wl_193 vdd gnd cell_6t
Xbit_r194_c19 bl_19 br_19 wl_194 vdd gnd cell_6t
Xbit_r195_c19 bl_19 br_19 wl_195 vdd gnd cell_6t
Xbit_r196_c19 bl_19 br_19 wl_196 vdd gnd cell_6t
Xbit_r197_c19 bl_19 br_19 wl_197 vdd gnd cell_6t
Xbit_r198_c19 bl_19 br_19 wl_198 vdd gnd cell_6t
Xbit_r199_c19 bl_19 br_19 wl_199 vdd gnd cell_6t
Xbit_r200_c19 bl_19 br_19 wl_200 vdd gnd cell_6t
Xbit_r201_c19 bl_19 br_19 wl_201 vdd gnd cell_6t
Xbit_r202_c19 bl_19 br_19 wl_202 vdd gnd cell_6t
Xbit_r203_c19 bl_19 br_19 wl_203 vdd gnd cell_6t
Xbit_r204_c19 bl_19 br_19 wl_204 vdd gnd cell_6t
Xbit_r205_c19 bl_19 br_19 wl_205 vdd gnd cell_6t
Xbit_r206_c19 bl_19 br_19 wl_206 vdd gnd cell_6t
Xbit_r207_c19 bl_19 br_19 wl_207 vdd gnd cell_6t
Xbit_r208_c19 bl_19 br_19 wl_208 vdd gnd cell_6t
Xbit_r209_c19 bl_19 br_19 wl_209 vdd gnd cell_6t
Xbit_r210_c19 bl_19 br_19 wl_210 vdd gnd cell_6t
Xbit_r211_c19 bl_19 br_19 wl_211 vdd gnd cell_6t
Xbit_r212_c19 bl_19 br_19 wl_212 vdd gnd cell_6t
Xbit_r213_c19 bl_19 br_19 wl_213 vdd gnd cell_6t
Xbit_r214_c19 bl_19 br_19 wl_214 vdd gnd cell_6t
Xbit_r215_c19 bl_19 br_19 wl_215 vdd gnd cell_6t
Xbit_r216_c19 bl_19 br_19 wl_216 vdd gnd cell_6t
Xbit_r217_c19 bl_19 br_19 wl_217 vdd gnd cell_6t
Xbit_r218_c19 bl_19 br_19 wl_218 vdd gnd cell_6t
Xbit_r219_c19 bl_19 br_19 wl_219 vdd gnd cell_6t
Xbit_r220_c19 bl_19 br_19 wl_220 vdd gnd cell_6t
Xbit_r221_c19 bl_19 br_19 wl_221 vdd gnd cell_6t
Xbit_r222_c19 bl_19 br_19 wl_222 vdd gnd cell_6t
Xbit_r223_c19 bl_19 br_19 wl_223 vdd gnd cell_6t
Xbit_r224_c19 bl_19 br_19 wl_224 vdd gnd cell_6t
Xbit_r225_c19 bl_19 br_19 wl_225 vdd gnd cell_6t
Xbit_r226_c19 bl_19 br_19 wl_226 vdd gnd cell_6t
Xbit_r227_c19 bl_19 br_19 wl_227 vdd gnd cell_6t
Xbit_r228_c19 bl_19 br_19 wl_228 vdd gnd cell_6t
Xbit_r229_c19 bl_19 br_19 wl_229 vdd gnd cell_6t
Xbit_r230_c19 bl_19 br_19 wl_230 vdd gnd cell_6t
Xbit_r231_c19 bl_19 br_19 wl_231 vdd gnd cell_6t
Xbit_r232_c19 bl_19 br_19 wl_232 vdd gnd cell_6t
Xbit_r233_c19 bl_19 br_19 wl_233 vdd gnd cell_6t
Xbit_r234_c19 bl_19 br_19 wl_234 vdd gnd cell_6t
Xbit_r235_c19 bl_19 br_19 wl_235 vdd gnd cell_6t
Xbit_r236_c19 bl_19 br_19 wl_236 vdd gnd cell_6t
Xbit_r237_c19 bl_19 br_19 wl_237 vdd gnd cell_6t
Xbit_r238_c19 bl_19 br_19 wl_238 vdd gnd cell_6t
Xbit_r239_c19 bl_19 br_19 wl_239 vdd gnd cell_6t
Xbit_r240_c19 bl_19 br_19 wl_240 vdd gnd cell_6t
Xbit_r241_c19 bl_19 br_19 wl_241 vdd gnd cell_6t
Xbit_r242_c19 bl_19 br_19 wl_242 vdd gnd cell_6t
Xbit_r243_c19 bl_19 br_19 wl_243 vdd gnd cell_6t
Xbit_r244_c19 bl_19 br_19 wl_244 vdd gnd cell_6t
Xbit_r245_c19 bl_19 br_19 wl_245 vdd gnd cell_6t
Xbit_r246_c19 bl_19 br_19 wl_246 vdd gnd cell_6t
Xbit_r247_c19 bl_19 br_19 wl_247 vdd gnd cell_6t
Xbit_r248_c19 bl_19 br_19 wl_248 vdd gnd cell_6t
Xbit_r249_c19 bl_19 br_19 wl_249 vdd gnd cell_6t
Xbit_r250_c19 bl_19 br_19 wl_250 vdd gnd cell_6t
Xbit_r251_c19 bl_19 br_19 wl_251 vdd gnd cell_6t
Xbit_r252_c19 bl_19 br_19 wl_252 vdd gnd cell_6t
Xbit_r253_c19 bl_19 br_19 wl_253 vdd gnd cell_6t
Xbit_r254_c19 bl_19 br_19 wl_254 vdd gnd cell_6t
Xbit_r255_c19 bl_19 br_19 wl_255 vdd gnd cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd cell_6t
Xbit_r1_c20 bl_20 br_20 wl_1 vdd gnd cell_6t
Xbit_r2_c20 bl_20 br_20 wl_2 vdd gnd cell_6t
Xbit_r3_c20 bl_20 br_20 wl_3 vdd gnd cell_6t
Xbit_r4_c20 bl_20 br_20 wl_4 vdd gnd cell_6t
Xbit_r5_c20 bl_20 br_20 wl_5 vdd gnd cell_6t
Xbit_r6_c20 bl_20 br_20 wl_6 vdd gnd cell_6t
Xbit_r7_c20 bl_20 br_20 wl_7 vdd gnd cell_6t
Xbit_r8_c20 bl_20 br_20 wl_8 vdd gnd cell_6t
Xbit_r9_c20 bl_20 br_20 wl_9 vdd gnd cell_6t
Xbit_r10_c20 bl_20 br_20 wl_10 vdd gnd cell_6t
Xbit_r11_c20 bl_20 br_20 wl_11 vdd gnd cell_6t
Xbit_r12_c20 bl_20 br_20 wl_12 vdd gnd cell_6t
Xbit_r13_c20 bl_20 br_20 wl_13 vdd gnd cell_6t
Xbit_r14_c20 bl_20 br_20 wl_14 vdd gnd cell_6t
Xbit_r15_c20 bl_20 br_20 wl_15 vdd gnd cell_6t
Xbit_r16_c20 bl_20 br_20 wl_16 vdd gnd cell_6t
Xbit_r17_c20 bl_20 br_20 wl_17 vdd gnd cell_6t
Xbit_r18_c20 bl_20 br_20 wl_18 vdd gnd cell_6t
Xbit_r19_c20 bl_20 br_20 wl_19 vdd gnd cell_6t
Xbit_r20_c20 bl_20 br_20 wl_20 vdd gnd cell_6t
Xbit_r21_c20 bl_20 br_20 wl_21 vdd gnd cell_6t
Xbit_r22_c20 bl_20 br_20 wl_22 vdd gnd cell_6t
Xbit_r23_c20 bl_20 br_20 wl_23 vdd gnd cell_6t
Xbit_r24_c20 bl_20 br_20 wl_24 vdd gnd cell_6t
Xbit_r25_c20 bl_20 br_20 wl_25 vdd gnd cell_6t
Xbit_r26_c20 bl_20 br_20 wl_26 vdd gnd cell_6t
Xbit_r27_c20 bl_20 br_20 wl_27 vdd gnd cell_6t
Xbit_r28_c20 bl_20 br_20 wl_28 vdd gnd cell_6t
Xbit_r29_c20 bl_20 br_20 wl_29 vdd gnd cell_6t
Xbit_r30_c20 bl_20 br_20 wl_30 vdd gnd cell_6t
Xbit_r31_c20 bl_20 br_20 wl_31 vdd gnd cell_6t
Xbit_r32_c20 bl_20 br_20 wl_32 vdd gnd cell_6t
Xbit_r33_c20 bl_20 br_20 wl_33 vdd gnd cell_6t
Xbit_r34_c20 bl_20 br_20 wl_34 vdd gnd cell_6t
Xbit_r35_c20 bl_20 br_20 wl_35 vdd gnd cell_6t
Xbit_r36_c20 bl_20 br_20 wl_36 vdd gnd cell_6t
Xbit_r37_c20 bl_20 br_20 wl_37 vdd gnd cell_6t
Xbit_r38_c20 bl_20 br_20 wl_38 vdd gnd cell_6t
Xbit_r39_c20 bl_20 br_20 wl_39 vdd gnd cell_6t
Xbit_r40_c20 bl_20 br_20 wl_40 vdd gnd cell_6t
Xbit_r41_c20 bl_20 br_20 wl_41 vdd gnd cell_6t
Xbit_r42_c20 bl_20 br_20 wl_42 vdd gnd cell_6t
Xbit_r43_c20 bl_20 br_20 wl_43 vdd gnd cell_6t
Xbit_r44_c20 bl_20 br_20 wl_44 vdd gnd cell_6t
Xbit_r45_c20 bl_20 br_20 wl_45 vdd gnd cell_6t
Xbit_r46_c20 bl_20 br_20 wl_46 vdd gnd cell_6t
Xbit_r47_c20 bl_20 br_20 wl_47 vdd gnd cell_6t
Xbit_r48_c20 bl_20 br_20 wl_48 vdd gnd cell_6t
Xbit_r49_c20 bl_20 br_20 wl_49 vdd gnd cell_6t
Xbit_r50_c20 bl_20 br_20 wl_50 vdd gnd cell_6t
Xbit_r51_c20 bl_20 br_20 wl_51 vdd gnd cell_6t
Xbit_r52_c20 bl_20 br_20 wl_52 vdd gnd cell_6t
Xbit_r53_c20 bl_20 br_20 wl_53 vdd gnd cell_6t
Xbit_r54_c20 bl_20 br_20 wl_54 vdd gnd cell_6t
Xbit_r55_c20 bl_20 br_20 wl_55 vdd gnd cell_6t
Xbit_r56_c20 bl_20 br_20 wl_56 vdd gnd cell_6t
Xbit_r57_c20 bl_20 br_20 wl_57 vdd gnd cell_6t
Xbit_r58_c20 bl_20 br_20 wl_58 vdd gnd cell_6t
Xbit_r59_c20 bl_20 br_20 wl_59 vdd gnd cell_6t
Xbit_r60_c20 bl_20 br_20 wl_60 vdd gnd cell_6t
Xbit_r61_c20 bl_20 br_20 wl_61 vdd gnd cell_6t
Xbit_r62_c20 bl_20 br_20 wl_62 vdd gnd cell_6t
Xbit_r63_c20 bl_20 br_20 wl_63 vdd gnd cell_6t
Xbit_r64_c20 bl_20 br_20 wl_64 vdd gnd cell_6t
Xbit_r65_c20 bl_20 br_20 wl_65 vdd gnd cell_6t
Xbit_r66_c20 bl_20 br_20 wl_66 vdd gnd cell_6t
Xbit_r67_c20 bl_20 br_20 wl_67 vdd gnd cell_6t
Xbit_r68_c20 bl_20 br_20 wl_68 vdd gnd cell_6t
Xbit_r69_c20 bl_20 br_20 wl_69 vdd gnd cell_6t
Xbit_r70_c20 bl_20 br_20 wl_70 vdd gnd cell_6t
Xbit_r71_c20 bl_20 br_20 wl_71 vdd gnd cell_6t
Xbit_r72_c20 bl_20 br_20 wl_72 vdd gnd cell_6t
Xbit_r73_c20 bl_20 br_20 wl_73 vdd gnd cell_6t
Xbit_r74_c20 bl_20 br_20 wl_74 vdd gnd cell_6t
Xbit_r75_c20 bl_20 br_20 wl_75 vdd gnd cell_6t
Xbit_r76_c20 bl_20 br_20 wl_76 vdd gnd cell_6t
Xbit_r77_c20 bl_20 br_20 wl_77 vdd gnd cell_6t
Xbit_r78_c20 bl_20 br_20 wl_78 vdd gnd cell_6t
Xbit_r79_c20 bl_20 br_20 wl_79 vdd gnd cell_6t
Xbit_r80_c20 bl_20 br_20 wl_80 vdd gnd cell_6t
Xbit_r81_c20 bl_20 br_20 wl_81 vdd gnd cell_6t
Xbit_r82_c20 bl_20 br_20 wl_82 vdd gnd cell_6t
Xbit_r83_c20 bl_20 br_20 wl_83 vdd gnd cell_6t
Xbit_r84_c20 bl_20 br_20 wl_84 vdd gnd cell_6t
Xbit_r85_c20 bl_20 br_20 wl_85 vdd gnd cell_6t
Xbit_r86_c20 bl_20 br_20 wl_86 vdd gnd cell_6t
Xbit_r87_c20 bl_20 br_20 wl_87 vdd gnd cell_6t
Xbit_r88_c20 bl_20 br_20 wl_88 vdd gnd cell_6t
Xbit_r89_c20 bl_20 br_20 wl_89 vdd gnd cell_6t
Xbit_r90_c20 bl_20 br_20 wl_90 vdd gnd cell_6t
Xbit_r91_c20 bl_20 br_20 wl_91 vdd gnd cell_6t
Xbit_r92_c20 bl_20 br_20 wl_92 vdd gnd cell_6t
Xbit_r93_c20 bl_20 br_20 wl_93 vdd gnd cell_6t
Xbit_r94_c20 bl_20 br_20 wl_94 vdd gnd cell_6t
Xbit_r95_c20 bl_20 br_20 wl_95 vdd gnd cell_6t
Xbit_r96_c20 bl_20 br_20 wl_96 vdd gnd cell_6t
Xbit_r97_c20 bl_20 br_20 wl_97 vdd gnd cell_6t
Xbit_r98_c20 bl_20 br_20 wl_98 vdd gnd cell_6t
Xbit_r99_c20 bl_20 br_20 wl_99 vdd gnd cell_6t
Xbit_r100_c20 bl_20 br_20 wl_100 vdd gnd cell_6t
Xbit_r101_c20 bl_20 br_20 wl_101 vdd gnd cell_6t
Xbit_r102_c20 bl_20 br_20 wl_102 vdd gnd cell_6t
Xbit_r103_c20 bl_20 br_20 wl_103 vdd gnd cell_6t
Xbit_r104_c20 bl_20 br_20 wl_104 vdd gnd cell_6t
Xbit_r105_c20 bl_20 br_20 wl_105 vdd gnd cell_6t
Xbit_r106_c20 bl_20 br_20 wl_106 vdd gnd cell_6t
Xbit_r107_c20 bl_20 br_20 wl_107 vdd gnd cell_6t
Xbit_r108_c20 bl_20 br_20 wl_108 vdd gnd cell_6t
Xbit_r109_c20 bl_20 br_20 wl_109 vdd gnd cell_6t
Xbit_r110_c20 bl_20 br_20 wl_110 vdd gnd cell_6t
Xbit_r111_c20 bl_20 br_20 wl_111 vdd gnd cell_6t
Xbit_r112_c20 bl_20 br_20 wl_112 vdd gnd cell_6t
Xbit_r113_c20 bl_20 br_20 wl_113 vdd gnd cell_6t
Xbit_r114_c20 bl_20 br_20 wl_114 vdd gnd cell_6t
Xbit_r115_c20 bl_20 br_20 wl_115 vdd gnd cell_6t
Xbit_r116_c20 bl_20 br_20 wl_116 vdd gnd cell_6t
Xbit_r117_c20 bl_20 br_20 wl_117 vdd gnd cell_6t
Xbit_r118_c20 bl_20 br_20 wl_118 vdd gnd cell_6t
Xbit_r119_c20 bl_20 br_20 wl_119 vdd gnd cell_6t
Xbit_r120_c20 bl_20 br_20 wl_120 vdd gnd cell_6t
Xbit_r121_c20 bl_20 br_20 wl_121 vdd gnd cell_6t
Xbit_r122_c20 bl_20 br_20 wl_122 vdd gnd cell_6t
Xbit_r123_c20 bl_20 br_20 wl_123 vdd gnd cell_6t
Xbit_r124_c20 bl_20 br_20 wl_124 vdd gnd cell_6t
Xbit_r125_c20 bl_20 br_20 wl_125 vdd gnd cell_6t
Xbit_r126_c20 bl_20 br_20 wl_126 vdd gnd cell_6t
Xbit_r127_c20 bl_20 br_20 wl_127 vdd gnd cell_6t
Xbit_r128_c20 bl_20 br_20 wl_128 vdd gnd cell_6t
Xbit_r129_c20 bl_20 br_20 wl_129 vdd gnd cell_6t
Xbit_r130_c20 bl_20 br_20 wl_130 vdd gnd cell_6t
Xbit_r131_c20 bl_20 br_20 wl_131 vdd gnd cell_6t
Xbit_r132_c20 bl_20 br_20 wl_132 vdd gnd cell_6t
Xbit_r133_c20 bl_20 br_20 wl_133 vdd gnd cell_6t
Xbit_r134_c20 bl_20 br_20 wl_134 vdd gnd cell_6t
Xbit_r135_c20 bl_20 br_20 wl_135 vdd gnd cell_6t
Xbit_r136_c20 bl_20 br_20 wl_136 vdd gnd cell_6t
Xbit_r137_c20 bl_20 br_20 wl_137 vdd gnd cell_6t
Xbit_r138_c20 bl_20 br_20 wl_138 vdd gnd cell_6t
Xbit_r139_c20 bl_20 br_20 wl_139 vdd gnd cell_6t
Xbit_r140_c20 bl_20 br_20 wl_140 vdd gnd cell_6t
Xbit_r141_c20 bl_20 br_20 wl_141 vdd gnd cell_6t
Xbit_r142_c20 bl_20 br_20 wl_142 vdd gnd cell_6t
Xbit_r143_c20 bl_20 br_20 wl_143 vdd gnd cell_6t
Xbit_r144_c20 bl_20 br_20 wl_144 vdd gnd cell_6t
Xbit_r145_c20 bl_20 br_20 wl_145 vdd gnd cell_6t
Xbit_r146_c20 bl_20 br_20 wl_146 vdd gnd cell_6t
Xbit_r147_c20 bl_20 br_20 wl_147 vdd gnd cell_6t
Xbit_r148_c20 bl_20 br_20 wl_148 vdd gnd cell_6t
Xbit_r149_c20 bl_20 br_20 wl_149 vdd gnd cell_6t
Xbit_r150_c20 bl_20 br_20 wl_150 vdd gnd cell_6t
Xbit_r151_c20 bl_20 br_20 wl_151 vdd gnd cell_6t
Xbit_r152_c20 bl_20 br_20 wl_152 vdd gnd cell_6t
Xbit_r153_c20 bl_20 br_20 wl_153 vdd gnd cell_6t
Xbit_r154_c20 bl_20 br_20 wl_154 vdd gnd cell_6t
Xbit_r155_c20 bl_20 br_20 wl_155 vdd gnd cell_6t
Xbit_r156_c20 bl_20 br_20 wl_156 vdd gnd cell_6t
Xbit_r157_c20 bl_20 br_20 wl_157 vdd gnd cell_6t
Xbit_r158_c20 bl_20 br_20 wl_158 vdd gnd cell_6t
Xbit_r159_c20 bl_20 br_20 wl_159 vdd gnd cell_6t
Xbit_r160_c20 bl_20 br_20 wl_160 vdd gnd cell_6t
Xbit_r161_c20 bl_20 br_20 wl_161 vdd gnd cell_6t
Xbit_r162_c20 bl_20 br_20 wl_162 vdd gnd cell_6t
Xbit_r163_c20 bl_20 br_20 wl_163 vdd gnd cell_6t
Xbit_r164_c20 bl_20 br_20 wl_164 vdd gnd cell_6t
Xbit_r165_c20 bl_20 br_20 wl_165 vdd gnd cell_6t
Xbit_r166_c20 bl_20 br_20 wl_166 vdd gnd cell_6t
Xbit_r167_c20 bl_20 br_20 wl_167 vdd gnd cell_6t
Xbit_r168_c20 bl_20 br_20 wl_168 vdd gnd cell_6t
Xbit_r169_c20 bl_20 br_20 wl_169 vdd gnd cell_6t
Xbit_r170_c20 bl_20 br_20 wl_170 vdd gnd cell_6t
Xbit_r171_c20 bl_20 br_20 wl_171 vdd gnd cell_6t
Xbit_r172_c20 bl_20 br_20 wl_172 vdd gnd cell_6t
Xbit_r173_c20 bl_20 br_20 wl_173 vdd gnd cell_6t
Xbit_r174_c20 bl_20 br_20 wl_174 vdd gnd cell_6t
Xbit_r175_c20 bl_20 br_20 wl_175 vdd gnd cell_6t
Xbit_r176_c20 bl_20 br_20 wl_176 vdd gnd cell_6t
Xbit_r177_c20 bl_20 br_20 wl_177 vdd gnd cell_6t
Xbit_r178_c20 bl_20 br_20 wl_178 vdd gnd cell_6t
Xbit_r179_c20 bl_20 br_20 wl_179 vdd gnd cell_6t
Xbit_r180_c20 bl_20 br_20 wl_180 vdd gnd cell_6t
Xbit_r181_c20 bl_20 br_20 wl_181 vdd gnd cell_6t
Xbit_r182_c20 bl_20 br_20 wl_182 vdd gnd cell_6t
Xbit_r183_c20 bl_20 br_20 wl_183 vdd gnd cell_6t
Xbit_r184_c20 bl_20 br_20 wl_184 vdd gnd cell_6t
Xbit_r185_c20 bl_20 br_20 wl_185 vdd gnd cell_6t
Xbit_r186_c20 bl_20 br_20 wl_186 vdd gnd cell_6t
Xbit_r187_c20 bl_20 br_20 wl_187 vdd gnd cell_6t
Xbit_r188_c20 bl_20 br_20 wl_188 vdd gnd cell_6t
Xbit_r189_c20 bl_20 br_20 wl_189 vdd gnd cell_6t
Xbit_r190_c20 bl_20 br_20 wl_190 vdd gnd cell_6t
Xbit_r191_c20 bl_20 br_20 wl_191 vdd gnd cell_6t
Xbit_r192_c20 bl_20 br_20 wl_192 vdd gnd cell_6t
Xbit_r193_c20 bl_20 br_20 wl_193 vdd gnd cell_6t
Xbit_r194_c20 bl_20 br_20 wl_194 vdd gnd cell_6t
Xbit_r195_c20 bl_20 br_20 wl_195 vdd gnd cell_6t
Xbit_r196_c20 bl_20 br_20 wl_196 vdd gnd cell_6t
Xbit_r197_c20 bl_20 br_20 wl_197 vdd gnd cell_6t
Xbit_r198_c20 bl_20 br_20 wl_198 vdd gnd cell_6t
Xbit_r199_c20 bl_20 br_20 wl_199 vdd gnd cell_6t
Xbit_r200_c20 bl_20 br_20 wl_200 vdd gnd cell_6t
Xbit_r201_c20 bl_20 br_20 wl_201 vdd gnd cell_6t
Xbit_r202_c20 bl_20 br_20 wl_202 vdd gnd cell_6t
Xbit_r203_c20 bl_20 br_20 wl_203 vdd gnd cell_6t
Xbit_r204_c20 bl_20 br_20 wl_204 vdd gnd cell_6t
Xbit_r205_c20 bl_20 br_20 wl_205 vdd gnd cell_6t
Xbit_r206_c20 bl_20 br_20 wl_206 vdd gnd cell_6t
Xbit_r207_c20 bl_20 br_20 wl_207 vdd gnd cell_6t
Xbit_r208_c20 bl_20 br_20 wl_208 vdd gnd cell_6t
Xbit_r209_c20 bl_20 br_20 wl_209 vdd gnd cell_6t
Xbit_r210_c20 bl_20 br_20 wl_210 vdd gnd cell_6t
Xbit_r211_c20 bl_20 br_20 wl_211 vdd gnd cell_6t
Xbit_r212_c20 bl_20 br_20 wl_212 vdd gnd cell_6t
Xbit_r213_c20 bl_20 br_20 wl_213 vdd gnd cell_6t
Xbit_r214_c20 bl_20 br_20 wl_214 vdd gnd cell_6t
Xbit_r215_c20 bl_20 br_20 wl_215 vdd gnd cell_6t
Xbit_r216_c20 bl_20 br_20 wl_216 vdd gnd cell_6t
Xbit_r217_c20 bl_20 br_20 wl_217 vdd gnd cell_6t
Xbit_r218_c20 bl_20 br_20 wl_218 vdd gnd cell_6t
Xbit_r219_c20 bl_20 br_20 wl_219 vdd gnd cell_6t
Xbit_r220_c20 bl_20 br_20 wl_220 vdd gnd cell_6t
Xbit_r221_c20 bl_20 br_20 wl_221 vdd gnd cell_6t
Xbit_r222_c20 bl_20 br_20 wl_222 vdd gnd cell_6t
Xbit_r223_c20 bl_20 br_20 wl_223 vdd gnd cell_6t
Xbit_r224_c20 bl_20 br_20 wl_224 vdd gnd cell_6t
Xbit_r225_c20 bl_20 br_20 wl_225 vdd gnd cell_6t
Xbit_r226_c20 bl_20 br_20 wl_226 vdd gnd cell_6t
Xbit_r227_c20 bl_20 br_20 wl_227 vdd gnd cell_6t
Xbit_r228_c20 bl_20 br_20 wl_228 vdd gnd cell_6t
Xbit_r229_c20 bl_20 br_20 wl_229 vdd gnd cell_6t
Xbit_r230_c20 bl_20 br_20 wl_230 vdd gnd cell_6t
Xbit_r231_c20 bl_20 br_20 wl_231 vdd gnd cell_6t
Xbit_r232_c20 bl_20 br_20 wl_232 vdd gnd cell_6t
Xbit_r233_c20 bl_20 br_20 wl_233 vdd gnd cell_6t
Xbit_r234_c20 bl_20 br_20 wl_234 vdd gnd cell_6t
Xbit_r235_c20 bl_20 br_20 wl_235 vdd gnd cell_6t
Xbit_r236_c20 bl_20 br_20 wl_236 vdd gnd cell_6t
Xbit_r237_c20 bl_20 br_20 wl_237 vdd gnd cell_6t
Xbit_r238_c20 bl_20 br_20 wl_238 vdd gnd cell_6t
Xbit_r239_c20 bl_20 br_20 wl_239 vdd gnd cell_6t
Xbit_r240_c20 bl_20 br_20 wl_240 vdd gnd cell_6t
Xbit_r241_c20 bl_20 br_20 wl_241 vdd gnd cell_6t
Xbit_r242_c20 bl_20 br_20 wl_242 vdd gnd cell_6t
Xbit_r243_c20 bl_20 br_20 wl_243 vdd gnd cell_6t
Xbit_r244_c20 bl_20 br_20 wl_244 vdd gnd cell_6t
Xbit_r245_c20 bl_20 br_20 wl_245 vdd gnd cell_6t
Xbit_r246_c20 bl_20 br_20 wl_246 vdd gnd cell_6t
Xbit_r247_c20 bl_20 br_20 wl_247 vdd gnd cell_6t
Xbit_r248_c20 bl_20 br_20 wl_248 vdd gnd cell_6t
Xbit_r249_c20 bl_20 br_20 wl_249 vdd gnd cell_6t
Xbit_r250_c20 bl_20 br_20 wl_250 vdd gnd cell_6t
Xbit_r251_c20 bl_20 br_20 wl_251 vdd gnd cell_6t
Xbit_r252_c20 bl_20 br_20 wl_252 vdd gnd cell_6t
Xbit_r253_c20 bl_20 br_20 wl_253 vdd gnd cell_6t
Xbit_r254_c20 bl_20 br_20 wl_254 vdd gnd cell_6t
Xbit_r255_c20 bl_20 br_20 wl_255 vdd gnd cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd cell_6t
Xbit_r1_c21 bl_21 br_21 wl_1 vdd gnd cell_6t
Xbit_r2_c21 bl_21 br_21 wl_2 vdd gnd cell_6t
Xbit_r3_c21 bl_21 br_21 wl_3 vdd gnd cell_6t
Xbit_r4_c21 bl_21 br_21 wl_4 vdd gnd cell_6t
Xbit_r5_c21 bl_21 br_21 wl_5 vdd gnd cell_6t
Xbit_r6_c21 bl_21 br_21 wl_6 vdd gnd cell_6t
Xbit_r7_c21 bl_21 br_21 wl_7 vdd gnd cell_6t
Xbit_r8_c21 bl_21 br_21 wl_8 vdd gnd cell_6t
Xbit_r9_c21 bl_21 br_21 wl_9 vdd gnd cell_6t
Xbit_r10_c21 bl_21 br_21 wl_10 vdd gnd cell_6t
Xbit_r11_c21 bl_21 br_21 wl_11 vdd gnd cell_6t
Xbit_r12_c21 bl_21 br_21 wl_12 vdd gnd cell_6t
Xbit_r13_c21 bl_21 br_21 wl_13 vdd gnd cell_6t
Xbit_r14_c21 bl_21 br_21 wl_14 vdd gnd cell_6t
Xbit_r15_c21 bl_21 br_21 wl_15 vdd gnd cell_6t
Xbit_r16_c21 bl_21 br_21 wl_16 vdd gnd cell_6t
Xbit_r17_c21 bl_21 br_21 wl_17 vdd gnd cell_6t
Xbit_r18_c21 bl_21 br_21 wl_18 vdd gnd cell_6t
Xbit_r19_c21 bl_21 br_21 wl_19 vdd gnd cell_6t
Xbit_r20_c21 bl_21 br_21 wl_20 vdd gnd cell_6t
Xbit_r21_c21 bl_21 br_21 wl_21 vdd gnd cell_6t
Xbit_r22_c21 bl_21 br_21 wl_22 vdd gnd cell_6t
Xbit_r23_c21 bl_21 br_21 wl_23 vdd gnd cell_6t
Xbit_r24_c21 bl_21 br_21 wl_24 vdd gnd cell_6t
Xbit_r25_c21 bl_21 br_21 wl_25 vdd gnd cell_6t
Xbit_r26_c21 bl_21 br_21 wl_26 vdd gnd cell_6t
Xbit_r27_c21 bl_21 br_21 wl_27 vdd gnd cell_6t
Xbit_r28_c21 bl_21 br_21 wl_28 vdd gnd cell_6t
Xbit_r29_c21 bl_21 br_21 wl_29 vdd gnd cell_6t
Xbit_r30_c21 bl_21 br_21 wl_30 vdd gnd cell_6t
Xbit_r31_c21 bl_21 br_21 wl_31 vdd gnd cell_6t
Xbit_r32_c21 bl_21 br_21 wl_32 vdd gnd cell_6t
Xbit_r33_c21 bl_21 br_21 wl_33 vdd gnd cell_6t
Xbit_r34_c21 bl_21 br_21 wl_34 vdd gnd cell_6t
Xbit_r35_c21 bl_21 br_21 wl_35 vdd gnd cell_6t
Xbit_r36_c21 bl_21 br_21 wl_36 vdd gnd cell_6t
Xbit_r37_c21 bl_21 br_21 wl_37 vdd gnd cell_6t
Xbit_r38_c21 bl_21 br_21 wl_38 vdd gnd cell_6t
Xbit_r39_c21 bl_21 br_21 wl_39 vdd gnd cell_6t
Xbit_r40_c21 bl_21 br_21 wl_40 vdd gnd cell_6t
Xbit_r41_c21 bl_21 br_21 wl_41 vdd gnd cell_6t
Xbit_r42_c21 bl_21 br_21 wl_42 vdd gnd cell_6t
Xbit_r43_c21 bl_21 br_21 wl_43 vdd gnd cell_6t
Xbit_r44_c21 bl_21 br_21 wl_44 vdd gnd cell_6t
Xbit_r45_c21 bl_21 br_21 wl_45 vdd gnd cell_6t
Xbit_r46_c21 bl_21 br_21 wl_46 vdd gnd cell_6t
Xbit_r47_c21 bl_21 br_21 wl_47 vdd gnd cell_6t
Xbit_r48_c21 bl_21 br_21 wl_48 vdd gnd cell_6t
Xbit_r49_c21 bl_21 br_21 wl_49 vdd gnd cell_6t
Xbit_r50_c21 bl_21 br_21 wl_50 vdd gnd cell_6t
Xbit_r51_c21 bl_21 br_21 wl_51 vdd gnd cell_6t
Xbit_r52_c21 bl_21 br_21 wl_52 vdd gnd cell_6t
Xbit_r53_c21 bl_21 br_21 wl_53 vdd gnd cell_6t
Xbit_r54_c21 bl_21 br_21 wl_54 vdd gnd cell_6t
Xbit_r55_c21 bl_21 br_21 wl_55 vdd gnd cell_6t
Xbit_r56_c21 bl_21 br_21 wl_56 vdd gnd cell_6t
Xbit_r57_c21 bl_21 br_21 wl_57 vdd gnd cell_6t
Xbit_r58_c21 bl_21 br_21 wl_58 vdd gnd cell_6t
Xbit_r59_c21 bl_21 br_21 wl_59 vdd gnd cell_6t
Xbit_r60_c21 bl_21 br_21 wl_60 vdd gnd cell_6t
Xbit_r61_c21 bl_21 br_21 wl_61 vdd gnd cell_6t
Xbit_r62_c21 bl_21 br_21 wl_62 vdd gnd cell_6t
Xbit_r63_c21 bl_21 br_21 wl_63 vdd gnd cell_6t
Xbit_r64_c21 bl_21 br_21 wl_64 vdd gnd cell_6t
Xbit_r65_c21 bl_21 br_21 wl_65 vdd gnd cell_6t
Xbit_r66_c21 bl_21 br_21 wl_66 vdd gnd cell_6t
Xbit_r67_c21 bl_21 br_21 wl_67 vdd gnd cell_6t
Xbit_r68_c21 bl_21 br_21 wl_68 vdd gnd cell_6t
Xbit_r69_c21 bl_21 br_21 wl_69 vdd gnd cell_6t
Xbit_r70_c21 bl_21 br_21 wl_70 vdd gnd cell_6t
Xbit_r71_c21 bl_21 br_21 wl_71 vdd gnd cell_6t
Xbit_r72_c21 bl_21 br_21 wl_72 vdd gnd cell_6t
Xbit_r73_c21 bl_21 br_21 wl_73 vdd gnd cell_6t
Xbit_r74_c21 bl_21 br_21 wl_74 vdd gnd cell_6t
Xbit_r75_c21 bl_21 br_21 wl_75 vdd gnd cell_6t
Xbit_r76_c21 bl_21 br_21 wl_76 vdd gnd cell_6t
Xbit_r77_c21 bl_21 br_21 wl_77 vdd gnd cell_6t
Xbit_r78_c21 bl_21 br_21 wl_78 vdd gnd cell_6t
Xbit_r79_c21 bl_21 br_21 wl_79 vdd gnd cell_6t
Xbit_r80_c21 bl_21 br_21 wl_80 vdd gnd cell_6t
Xbit_r81_c21 bl_21 br_21 wl_81 vdd gnd cell_6t
Xbit_r82_c21 bl_21 br_21 wl_82 vdd gnd cell_6t
Xbit_r83_c21 bl_21 br_21 wl_83 vdd gnd cell_6t
Xbit_r84_c21 bl_21 br_21 wl_84 vdd gnd cell_6t
Xbit_r85_c21 bl_21 br_21 wl_85 vdd gnd cell_6t
Xbit_r86_c21 bl_21 br_21 wl_86 vdd gnd cell_6t
Xbit_r87_c21 bl_21 br_21 wl_87 vdd gnd cell_6t
Xbit_r88_c21 bl_21 br_21 wl_88 vdd gnd cell_6t
Xbit_r89_c21 bl_21 br_21 wl_89 vdd gnd cell_6t
Xbit_r90_c21 bl_21 br_21 wl_90 vdd gnd cell_6t
Xbit_r91_c21 bl_21 br_21 wl_91 vdd gnd cell_6t
Xbit_r92_c21 bl_21 br_21 wl_92 vdd gnd cell_6t
Xbit_r93_c21 bl_21 br_21 wl_93 vdd gnd cell_6t
Xbit_r94_c21 bl_21 br_21 wl_94 vdd gnd cell_6t
Xbit_r95_c21 bl_21 br_21 wl_95 vdd gnd cell_6t
Xbit_r96_c21 bl_21 br_21 wl_96 vdd gnd cell_6t
Xbit_r97_c21 bl_21 br_21 wl_97 vdd gnd cell_6t
Xbit_r98_c21 bl_21 br_21 wl_98 vdd gnd cell_6t
Xbit_r99_c21 bl_21 br_21 wl_99 vdd gnd cell_6t
Xbit_r100_c21 bl_21 br_21 wl_100 vdd gnd cell_6t
Xbit_r101_c21 bl_21 br_21 wl_101 vdd gnd cell_6t
Xbit_r102_c21 bl_21 br_21 wl_102 vdd gnd cell_6t
Xbit_r103_c21 bl_21 br_21 wl_103 vdd gnd cell_6t
Xbit_r104_c21 bl_21 br_21 wl_104 vdd gnd cell_6t
Xbit_r105_c21 bl_21 br_21 wl_105 vdd gnd cell_6t
Xbit_r106_c21 bl_21 br_21 wl_106 vdd gnd cell_6t
Xbit_r107_c21 bl_21 br_21 wl_107 vdd gnd cell_6t
Xbit_r108_c21 bl_21 br_21 wl_108 vdd gnd cell_6t
Xbit_r109_c21 bl_21 br_21 wl_109 vdd gnd cell_6t
Xbit_r110_c21 bl_21 br_21 wl_110 vdd gnd cell_6t
Xbit_r111_c21 bl_21 br_21 wl_111 vdd gnd cell_6t
Xbit_r112_c21 bl_21 br_21 wl_112 vdd gnd cell_6t
Xbit_r113_c21 bl_21 br_21 wl_113 vdd gnd cell_6t
Xbit_r114_c21 bl_21 br_21 wl_114 vdd gnd cell_6t
Xbit_r115_c21 bl_21 br_21 wl_115 vdd gnd cell_6t
Xbit_r116_c21 bl_21 br_21 wl_116 vdd gnd cell_6t
Xbit_r117_c21 bl_21 br_21 wl_117 vdd gnd cell_6t
Xbit_r118_c21 bl_21 br_21 wl_118 vdd gnd cell_6t
Xbit_r119_c21 bl_21 br_21 wl_119 vdd gnd cell_6t
Xbit_r120_c21 bl_21 br_21 wl_120 vdd gnd cell_6t
Xbit_r121_c21 bl_21 br_21 wl_121 vdd gnd cell_6t
Xbit_r122_c21 bl_21 br_21 wl_122 vdd gnd cell_6t
Xbit_r123_c21 bl_21 br_21 wl_123 vdd gnd cell_6t
Xbit_r124_c21 bl_21 br_21 wl_124 vdd gnd cell_6t
Xbit_r125_c21 bl_21 br_21 wl_125 vdd gnd cell_6t
Xbit_r126_c21 bl_21 br_21 wl_126 vdd gnd cell_6t
Xbit_r127_c21 bl_21 br_21 wl_127 vdd gnd cell_6t
Xbit_r128_c21 bl_21 br_21 wl_128 vdd gnd cell_6t
Xbit_r129_c21 bl_21 br_21 wl_129 vdd gnd cell_6t
Xbit_r130_c21 bl_21 br_21 wl_130 vdd gnd cell_6t
Xbit_r131_c21 bl_21 br_21 wl_131 vdd gnd cell_6t
Xbit_r132_c21 bl_21 br_21 wl_132 vdd gnd cell_6t
Xbit_r133_c21 bl_21 br_21 wl_133 vdd gnd cell_6t
Xbit_r134_c21 bl_21 br_21 wl_134 vdd gnd cell_6t
Xbit_r135_c21 bl_21 br_21 wl_135 vdd gnd cell_6t
Xbit_r136_c21 bl_21 br_21 wl_136 vdd gnd cell_6t
Xbit_r137_c21 bl_21 br_21 wl_137 vdd gnd cell_6t
Xbit_r138_c21 bl_21 br_21 wl_138 vdd gnd cell_6t
Xbit_r139_c21 bl_21 br_21 wl_139 vdd gnd cell_6t
Xbit_r140_c21 bl_21 br_21 wl_140 vdd gnd cell_6t
Xbit_r141_c21 bl_21 br_21 wl_141 vdd gnd cell_6t
Xbit_r142_c21 bl_21 br_21 wl_142 vdd gnd cell_6t
Xbit_r143_c21 bl_21 br_21 wl_143 vdd gnd cell_6t
Xbit_r144_c21 bl_21 br_21 wl_144 vdd gnd cell_6t
Xbit_r145_c21 bl_21 br_21 wl_145 vdd gnd cell_6t
Xbit_r146_c21 bl_21 br_21 wl_146 vdd gnd cell_6t
Xbit_r147_c21 bl_21 br_21 wl_147 vdd gnd cell_6t
Xbit_r148_c21 bl_21 br_21 wl_148 vdd gnd cell_6t
Xbit_r149_c21 bl_21 br_21 wl_149 vdd gnd cell_6t
Xbit_r150_c21 bl_21 br_21 wl_150 vdd gnd cell_6t
Xbit_r151_c21 bl_21 br_21 wl_151 vdd gnd cell_6t
Xbit_r152_c21 bl_21 br_21 wl_152 vdd gnd cell_6t
Xbit_r153_c21 bl_21 br_21 wl_153 vdd gnd cell_6t
Xbit_r154_c21 bl_21 br_21 wl_154 vdd gnd cell_6t
Xbit_r155_c21 bl_21 br_21 wl_155 vdd gnd cell_6t
Xbit_r156_c21 bl_21 br_21 wl_156 vdd gnd cell_6t
Xbit_r157_c21 bl_21 br_21 wl_157 vdd gnd cell_6t
Xbit_r158_c21 bl_21 br_21 wl_158 vdd gnd cell_6t
Xbit_r159_c21 bl_21 br_21 wl_159 vdd gnd cell_6t
Xbit_r160_c21 bl_21 br_21 wl_160 vdd gnd cell_6t
Xbit_r161_c21 bl_21 br_21 wl_161 vdd gnd cell_6t
Xbit_r162_c21 bl_21 br_21 wl_162 vdd gnd cell_6t
Xbit_r163_c21 bl_21 br_21 wl_163 vdd gnd cell_6t
Xbit_r164_c21 bl_21 br_21 wl_164 vdd gnd cell_6t
Xbit_r165_c21 bl_21 br_21 wl_165 vdd gnd cell_6t
Xbit_r166_c21 bl_21 br_21 wl_166 vdd gnd cell_6t
Xbit_r167_c21 bl_21 br_21 wl_167 vdd gnd cell_6t
Xbit_r168_c21 bl_21 br_21 wl_168 vdd gnd cell_6t
Xbit_r169_c21 bl_21 br_21 wl_169 vdd gnd cell_6t
Xbit_r170_c21 bl_21 br_21 wl_170 vdd gnd cell_6t
Xbit_r171_c21 bl_21 br_21 wl_171 vdd gnd cell_6t
Xbit_r172_c21 bl_21 br_21 wl_172 vdd gnd cell_6t
Xbit_r173_c21 bl_21 br_21 wl_173 vdd gnd cell_6t
Xbit_r174_c21 bl_21 br_21 wl_174 vdd gnd cell_6t
Xbit_r175_c21 bl_21 br_21 wl_175 vdd gnd cell_6t
Xbit_r176_c21 bl_21 br_21 wl_176 vdd gnd cell_6t
Xbit_r177_c21 bl_21 br_21 wl_177 vdd gnd cell_6t
Xbit_r178_c21 bl_21 br_21 wl_178 vdd gnd cell_6t
Xbit_r179_c21 bl_21 br_21 wl_179 vdd gnd cell_6t
Xbit_r180_c21 bl_21 br_21 wl_180 vdd gnd cell_6t
Xbit_r181_c21 bl_21 br_21 wl_181 vdd gnd cell_6t
Xbit_r182_c21 bl_21 br_21 wl_182 vdd gnd cell_6t
Xbit_r183_c21 bl_21 br_21 wl_183 vdd gnd cell_6t
Xbit_r184_c21 bl_21 br_21 wl_184 vdd gnd cell_6t
Xbit_r185_c21 bl_21 br_21 wl_185 vdd gnd cell_6t
Xbit_r186_c21 bl_21 br_21 wl_186 vdd gnd cell_6t
Xbit_r187_c21 bl_21 br_21 wl_187 vdd gnd cell_6t
Xbit_r188_c21 bl_21 br_21 wl_188 vdd gnd cell_6t
Xbit_r189_c21 bl_21 br_21 wl_189 vdd gnd cell_6t
Xbit_r190_c21 bl_21 br_21 wl_190 vdd gnd cell_6t
Xbit_r191_c21 bl_21 br_21 wl_191 vdd gnd cell_6t
Xbit_r192_c21 bl_21 br_21 wl_192 vdd gnd cell_6t
Xbit_r193_c21 bl_21 br_21 wl_193 vdd gnd cell_6t
Xbit_r194_c21 bl_21 br_21 wl_194 vdd gnd cell_6t
Xbit_r195_c21 bl_21 br_21 wl_195 vdd gnd cell_6t
Xbit_r196_c21 bl_21 br_21 wl_196 vdd gnd cell_6t
Xbit_r197_c21 bl_21 br_21 wl_197 vdd gnd cell_6t
Xbit_r198_c21 bl_21 br_21 wl_198 vdd gnd cell_6t
Xbit_r199_c21 bl_21 br_21 wl_199 vdd gnd cell_6t
Xbit_r200_c21 bl_21 br_21 wl_200 vdd gnd cell_6t
Xbit_r201_c21 bl_21 br_21 wl_201 vdd gnd cell_6t
Xbit_r202_c21 bl_21 br_21 wl_202 vdd gnd cell_6t
Xbit_r203_c21 bl_21 br_21 wl_203 vdd gnd cell_6t
Xbit_r204_c21 bl_21 br_21 wl_204 vdd gnd cell_6t
Xbit_r205_c21 bl_21 br_21 wl_205 vdd gnd cell_6t
Xbit_r206_c21 bl_21 br_21 wl_206 vdd gnd cell_6t
Xbit_r207_c21 bl_21 br_21 wl_207 vdd gnd cell_6t
Xbit_r208_c21 bl_21 br_21 wl_208 vdd gnd cell_6t
Xbit_r209_c21 bl_21 br_21 wl_209 vdd gnd cell_6t
Xbit_r210_c21 bl_21 br_21 wl_210 vdd gnd cell_6t
Xbit_r211_c21 bl_21 br_21 wl_211 vdd gnd cell_6t
Xbit_r212_c21 bl_21 br_21 wl_212 vdd gnd cell_6t
Xbit_r213_c21 bl_21 br_21 wl_213 vdd gnd cell_6t
Xbit_r214_c21 bl_21 br_21 wl_214 vdd gnd cell_6t
Xbit_r215_c21 bl_21 br_21 wl_215 vdd gnd cell_6t
Xbit_r216_c21 bl_21 br_21 wl_216 vdd gnd cell_6t
Xbit_r217_c21 bl_21 br_21 wl_217 vdd gnd cell_6t
Xbit_r218_c21 bl_21 br_21 wl_218 vdd gnd cell_6t
Xbit_r219_c21 bl_21 br_21 wl_219 vdd gnd cell_6t
Xbit_r220_c21 bl_21 br_21 wl_220 vdd gnd cell_6t
Xbit_r221_c21 bl_21 br_21 wl_221 vdd gnd cell_6t
Xbit_r222_c21 bl_21 br_21 wl_222 vdd gnd cell_6t
Xbit_r223_c21 bl_21 br_21 wl_223 vdd gnd cell_6t
Xbit_r224_c21 bl_21 br_21 wl_224 vdd gnd cell_6t
Xbit_r225_c21 bl_21 br_21 wl_225 vdd gnd cell_6t
Xbit_r226_c21 bl_21 br_21 wl_226 vdd gnd cell_6t
Xbit_r227_c21 bl_21 br_21 wl_227 vdd gnd cell_6t
Xbit_r228_c21 bl_21 br_21 wl_228 vdd gnd cell_6t
Xbit_r229_c21 bl_21 br_21 wl_229 vdd gnd cell_6t
Xbit_r230_c21 bl_21 br_21 wl_230 vdd gnd cell_6t
Xbit_r231_c21 bl_21 br_21 wl_231 vdd gnd cell_6t
Xbit_r232_c21 bl_21 br_21 wl_232 vdd gnd cell_6t
Xbit_r233_c21 bl_21 br_21 wl_233 vdd gnd cell_6t
Xbit_r234_c21 bl_21 br_21 wl_234 vdd gnd cell_6t
Xbit_r235_c21 bl_21 br_21 wl_235 vdd gnd cell_6t
Xbit_r236_c21 bl_21 br_21 wl_236 vdd gnd cell_6t
Xbit_r237_c21 bl_21 br_21 wl_237 vdd gnd cell_6t
Xbit_r238_c21 bl_21 br_21 wl_238 vdd gnd cell_6t
Xbit_r239_c21 bl_21 br_21 wl_239 vdd gnd cell_6t
Xbit_r240_c21 bl_21 br_21 wl_240 vdd gnd cell_6t
Xbit_r241_c21 bl_21 br_21 wl_241 vdd gnd cell_6t
Xbit_r242_c21 bl_21 br_21 wl_242 vdd gnd cell_6t
Xbit_r243_c21 bl_21 br_21 wl_243 vdd gnd cell_6t
Xbit_r244_c21 bl_21 br_21 wl_244 vdd gnd cell_6t
Xbit_r245_c21 bl_21 br_21 wl_245 vdd gnd cell_6t
Xbit_r246_c21 bl_21 br_21 wl_246 vdd gnd cell_6t
Xbit_r247_c21 bl_21 br_21 wl_247 vdd gnd cell_6t
Xbit_r248_c21 bl_21 br_21 wl_248 vdd gnd cell_6t
Xbit_r249_c21 bl_21 br_21 wl_249 vdd gnd cell_6t
Xbit_r250_c21 bl_21 br_21 wl_250 vdd gnd cell_6t
Xbit_r251_c21 bl_21 br_21 wl_251 vdd gnd cell_6t
Xbit_r252_c21 bl_21 br_21 wl_252 vdd gnd cell_6t
Xbit_r253_c21 bl_21 br_21 wl_253 vdd gnd cell_6t
Xbit_r254_c21 bl_21 br_21 wl_254 vdd gnd cell_6t
Xbit_r255_c21 bl_21 br_21 wl_255 vdd gnd cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd cell_6t
Xbit_r1_c22 bl_22 br_22 wl_1 vdd gnd cell_6t
Xbit_r2_c22 bl_22 br_22 wl_2 vdd gnd cell_6t
Xbit_r3_c22 bl_22 br_22 wl_3 vdd gnd cell_6t
Xbit_r4_c22 bl_22 br_22 wl_4 vdd gnd cell_6t
Xbit_r5_c22 bl_22 br_22 wl_5 vdd gnd cell_6t
Xbit_r6_c22 bl_22 br_22 wl_6 vdd gnd cell_6t
Xbit_r7_c22 bl_22 br_22 wl_7 vdd gnd cell_6t
Xbit_r8_c22 bl_22 br_22 wl_8 vdd gnd cell_6t
Xbit_r9_c22 bl_22 br_22 wl_9 vdd gnd cell_6t
Xbit_r10_c22 bl_22 br_22 wl_10 vdd gnd cell_6t
Xbit_r11_c22 bl_22 br_22 wl_11 vdd gnd cell_6t
Xbit_r12_c22 bl_22 br_22 wl_12 vdd gnd cell_6t
Xbit_r13_c22 bl_22 br_22 wl_13 vdd gnd cell_6t
Xbit_r14_c22 bl_22 br_22 wl_14 vdd gnd cell_6t
Xbit_r15_c22 bl_22 br_22 wl_15 vdd gnd cell_6t
Xbit_r16_c22 bl_22 br_22 wl_16 vdd gnd cell_6t
Xbit_r17_c22 bl_22 br_22 wl_17 vdd gnd cell_6t
Xbit_r18_c22 bl_22 br_22 wl_18 vdd gnd cell_6t
Xbit_r19_c22 bl_22 br_22 wl_19 vdd gnd cell_6t
Xbit_r20_c22 bl_22 br_22 wl_20 vdd gnd cell_6t
Xbit_r21_c22 bl_22 br_22 wl_21 vdd gnd cell_6t
Xbit_r22_c22 bl_22 br_22 wl_22 vdd gnd cell_6t
Xbit_r23_c22 bl_22 br_22 wl_23 vdd gnd cell_6t
Xbit_r24_c22 bl_22 br_22 wl_24 vdd gnd cell_6t
Xbit_r25_c22 bl_22 br_22 wl_25 vdd gnd cell_6t
Xbit_r26_c22 bl_22 br_22 wl_26 vdd gnd cell_6t
Xbit_r27_c22 bl_22 br_22 wl_27 vdd gnd cell_6t
Xbit_r28_c22 bl_22 br_22 wl_28 vdd gnd cell_6t
Xbit_r29_c22 bl_22 br_22 wl_29 vdd gnd cell_6t
Xbit_r30_c22 bl_22 br_22 wl_30 vdd gnd cell_6t
Xbit_r31_c22 bl_22 br_22 wl_31 vdd gnd cell_6t
Xbit_r32_c22 bl_22 br_22 wl_32 vdd gnd cell_6t
Xbit_r33_c22 bl_22 br_22 wl_33 vdd gnd cell_6t
Xbit_r34_c22 bl_22 br_22 wl_34 vdd gnd cell_6t
Xbit_r35_c22 bl_22 br_22 wl_35 vdd gnd cell_6t
Xbit_r36_c22 bl_22 br_22 wl_36 vdd gnd cell_6t
Xbit_r37_c22 bl_22 br_22 wl_37 vdd gnd cell_6t
Xbit_r38_c22 bl_22 br_22 wl_38 vdd gnd cell_6t
Xbit_r39_c22 bl_22 br_22 wl_39 vdd gnd cell_6t
Xbit_r40_c22 bl_22 br_22 wl_40 vdd gnd cell_6t
Xbit_r41_c22 bl_22 br_22 wl_41 vdd gnd cell_6t
Xbit_r42_c22 bl_22 br_22 wl_42 vdd gnd cell_6t
Xbit_r43_c22 bl_22 br_22 wl_43 vdd gnd cell_6t
Xbit_r44_c22 bl_22 br_22 wl_44 vdd gnd cell_6t
Xbit_r45_c22 bl_22 br_22 wl_45 vdd gnd cell_6t
Xbit_r46_c22 bl_22 br_22 wl_46 vdd gnd cell_6t
Xbit_r47_c22 bl_22 br_22 wl_47 vdd gnd cell_6t
Xbit_r48_c22 bl_22 br_22 wl_48 vdd gnd cell_6t
Xbit_r49_c22 bl_22 br_22 wl_49 vdd gnd cell_6t
Xbit_r50_c22 bl_22 br_22 wl_50 vdd gnd cell_6t
Xbit_r51_c22 bl_22 br_22 wl_51 vdd gnd cell_6t
Xbit_r52_c22 bl_22 br_22 wl_52 vdd gnd cell_6t
Xbit_r53_c22 bl_22 br_22 wl_53 vdd gnd cell_6t
Xbit_r54_c22 bl_22 br_22 wl_54 vdd gnd cell_6t
Xbit_r55_c22 bl_22 br_22 wl_55 vdd gnd cell_6t
Xbit_r56_c22 bl_22 br_22 wl_56 vdd gnd cell_6t
Xbit_r57_c22 bl_22 br_22 wl_57 vdd gnd cell_6t
Xbit_r58_c22 bl_22 br_22 wl_58 vdd gnd cell_6t
Xbit_r59_c22 bl_22 br_22 wl_59 vdd gnd cell_6t
Xbit_r60_c22 bl_22 br_22 wl_60 vdd gnd cell_6t
Xbit_r61_c22 bl_22 br_22 wl_61 vdd gnd cell_6t
Xbit_r62_c22 bl_22 br_22 wl_62 vdd gnd cell_6t
Xbit_r63_c22 bl_22 br_22 wl_63 vdd gnd cell_6t
Xbit_r64_c22 bl_22 br_22 wl_64 vdd gnd cell_6t
Xbit_r65_c22 bl_22 br_22 wl_65 vdd gnd cell_6t
Xbit_r66_c22 bl_22 br_22 wl_66 vdd gnd cell_6t
Xbit_r67_c22 bl_22 br_22 wl_67 vdd gnd cell_6t
Xbit_r68_c22 bl_22 br_22 wl_68 vdd gnd cell_6t
Xbit_r69_c22 bl_22 br_22 wl_69 vdd gnd cell_6t
Xbit_r70_c22 bl_22 br_22 wl_70 vdd gnd cell_6t
Xbit_r71_c22 bl_22 br_22 wl_71 vdd gnd cell_6t
Xbit_r72_c22 bl_22 br_22 wl_72 vdd gnd cell_6t
Xbit_r73_c22 bl_22 br_22 wl_73 vdd gnd cell_6t
Xbit_r74_c22 bl_22 br_22 wl_74 vdd gnd cell_6t
Xbit_r75_c22 bl_22 br_22 wl_75 vdd gnd cell_6t
Xbit_r76_c22 bl_22 br_22 wl_76 vdd gnd cell_6t
Xbit_r77_c22 bl_22 br_22 wl_77 vdd gnd cell_6t
Xbit_r78_c22 bl_22 br_22 wl_78 vdd gnd cell_6t
Xbit_r79_c22 bl_22 br_22 wl_79 vdd gnd cell_6t
Xbit_r80_c22 bl_22 br_22 wl_80 vdd gnd cell_6t
Xbit_r81_c22 bl_22 br_22 wl_81 vdd gnd cell_6t
Xbit_r82_c22 bl_22 br_22 wl_82 vdd gnd cell_6t
Xbit_r83_c22 bl_22 br_22 wl_83 vdd gnd cell_6t
Xbit_r84_c22 bl_22 br_22 wl_84 vdd gnd cell_6t
Xbit_r85_c22 bl_22 br_22 wl_85 vdd gnd cell_6t
Xbit_r86_c22 bl_22 br_22 wl_86 vdd gnd cell_6t
Xbit_r87_c22 bl_22 br_22 wl_87 vdd gnd cell_6t
Xbit_r88_c22 bl_22 br_22 wl_88 vdd gnd cell_6t
Xbit_r89_c22 bl_22 br_22 wl_89 vdd gnd cell_6t
Xbit_r90_c22 bl_22 br_22 wl_90 vdd gnd cell_6t
Xbit_r91_c22 bl_22 br_22 wl_91 vdd gnd cell_6t
Xbit_r92_c22 bl_22 br_22 wl_92 vdd gnd cell_6t
Xbit_r93_c22 bl_22 br_22 wl_93 vdd gnd cell_6t
Xbit_r94_c22 bl_22 br_22 wl_94 vdd gnd cell_6t
Xbit_r95_c22 bl_22 br_22 wl_95 vdd gnd cell_6t
Xbit_r96_c22 bl_22 br_22 wl_96 vdd gnd cell_6t
Xbit_r97_c22 bl_22 br_22 wl_97 vdd gnd cell_6t
Xbit_r98_c22 bl_22 br_22 wl_98 vdd gnd cell_6t
Xbit_r99_c22 bl_22 br_22 wl_99 vdd gnd cell_6t
Xbit_r100_c22 bl_22 br_22 wl_100 vdd gnd cell_6t
Xbit_r101_c22 bl_22 br_22 wl_101 vdd gnd cell_6t
Xbit_r102_c22 bl_22 br_22 wl_102 vdd gnd cell_6t
Xbit_r103_c22 bl_22 br_22 wl_103 vdd gnd cell_6t
Xbit_r104_c22 bl_22 br_22 wl_104 vdd gnd cell_6t
Xbit_r105_c22 bl_22 br_22 wl_105 vdd gnd cell_6t
Xbit_r106_c22 bl_22 br_22 wl_106 vdd gnd cell_6t
Xbit_r107_c22 bl_22 br_22 wl_107 vdd gnd cell_6t
Xbit_r108_c22 bl_22 br_22 wl_108 vdd gnd cell_6t
Xbit_r109_c22 bl_22 br_22 wl_109 vdd gnd cell_6t
Xbit_r110_c22 bl_22 br_22 wl_110 vdd gnd cell_6t
Xbit_r111_c22 bl_22 br_22 wl_111 vdd gnd cell_6t
Xbit_r112_c22 bl_22 br_22 wl_112 vdd gnd cell_6t
Xbit_r113_c22 bl_22 br_22 wl_113 vdd gnd cell_6t
Xbit_r114_c22 bl_22 br_22 wl_114 vdd gnd cell_6t
Xbit_r115_c22 bl_22 br_22 wl_115 vdd gnd cell_6t
Xbit_r116_c22 bl_22 br_22 wl_116 vdd gnd cell_6t
Xbit_r117_c22 bl_22 br_22 wl_117 vdd gnd cell_6t
Xbit_r118_c22 bl_22 br_22 wl_118 vdd gnd cell_6t
Xbit_r119_c22 bl_22 br_22 wl_119 vdd gnd cell_6t
Xbit_r120_c22 bl_22 br_22 wl_120 vdd gnd cell_6t
Xbit_r121_c22 bl_22 br_22 wl_121 vdd gnd cell_6t
Xbit_r122_c22 bl_22 br_22 wl_122 vdd gnd cell_6t
Xbit_r123_c22 bl_22 br_22 wl_123 vdd gnd cell_6t
Xbit_r124_c22 bl_22 br_22 wl_124 vdd gnd cell_6t
Xbit_r125_c22 bl_22 br_22 wl_125 vdd gnd cell_6t
Xbit_r126_c22 bl_22 br_22 wl_126 vdd gnd cell_6t
Xbit_r127_c22 bl_22 br_22 wl_127 vdd gnd cell_6t
Xbit_r128_c22 bl_22 br_22 wl_128 vdd gnd cell_6t
Xbit_r129_c22 bl_22 br_22 wl_129 vdd gnd cell_6t
Xbit_r130_c22 bl_22 br_22 wl_130 vdd gnd cell_6t
Xbit_r131_c22 bl_22 br_22 wl_131 vdd gnd cell_6t
Xbit_r132_c22 bl_22 br_22 wl_132 vdd gnd cell_6t
Xbit_r133_c22 bl_22 br_22 wl_133 vdd gnd cell_6t
Xbit_r134_c22 bl_22 br_22 wl_134 vdd gnd cell_6t
Xbit_r135_c22 bl_22 br_22 wl_135 vdd gnd cell_6t
Xbit_r136_c22 bl_22 br_22 wl_136 vdd gnd cell_6t
Xbit_r137_c22 bl_22 br_22 wl_137 vdd gnd cell_6t
Xbit_r138_c22 bl_22 br_22 wl_138 vdd gnd cell_6t
Xbit_r139_c22 bl_22 br_22 wl_139 vdd gnd cell_6t
Xbit_r140_c22 bl_22 br_22 wl_140 vdd gnd cell_6t
Xbit_r141_c22 bl_22 br_22 wl_141 vdd gnd cell_6t
Xbit_r142_c22 bl_22 br_22 wl_142 vdd gnd cell_6t
Xbit_r143_c22 bl_22 br_22 wl_143 vdd gnd cell_6t
Xbit_r144_c22 bl_22 br_22 wl_144 vdd gnd cell_6t
Xbit_r145_c22 bl_22 br_22 wl_145 vdd gnd cell_6t
Xbit_r146_c22 bl_22 br_22 wl_146 vdd gnd cell_6t
Xbit_r147_c22 bl_22 br_22 wl_147 vdd gnd cell_6t
Xbit_r148_c22 bl_22 br_22 wl_148 vdd gnd cell_6t
Xbit_r149_c22 bl_22 br_22 wl_149 vdd gnd cell_6t
Xbit_r150_c22 bl_22 br_22 wl_150 vdd gnd cell_6t
Xbit_r151_c22 bl_22 br_22 wl_151 vdd gnd cell_6t
Xbit_r152_c22 bl_22 br_22 wl_152 vdd gnd cell_6t
Xbit_r153_c22 bl_22 br_22 wl_153 vdd gnd cell_6t
Xbit_r154_c22 bl_22 br_22 wl_154 vdd gnd cell_6t
Xbit_r155_c22 bl_22 br_22 wl_155 vdd gnd cell_6t
Xbit_r156_c22 bl_22 br_22 wl_156 vdd gnd cell_6t
Xbit_r157_c22 bl_22 br_22 wl_157 vdd gnd cell_6t
Xbit_r158_c22 bl_22 br_22 wl_158 vdd gnd cell_6t
Xbit_r159_c22 bl_22 br_22 wl_159 vdd gnd cell_6t
Xbit_r160_c22 bl_22 br_22 wl_160 vdd gnd cell_6t
Xbit_r161_c22 bl_22 br_22 wl_161 vdd gnd cell_6t
Xbit_r162_c22 bl_22 br_22 wl_162 vdd gnd cell_6t
Xbit_r163_c22 bl_22 br_22 wl_163 vdd gnd cell_6t
Xbit_r164_c22 bl_22 br_22 wl_164 vdd gnd cell_6t
Xbit_r165_c22 bl_22 br_22 wl_165 vdd gnd cell_6t
Xbit_r166_c22 bl_22 br_22 wl_166 vdd gnd cell_6t
Xbit_r167_c22 bl_22 br_22 wl_167 vdd gnd cell_6t
Xbit_r168_c22 bl_22 br_22 wl_168 vdd gnd cell_6t
Xbit_r169_c22 bl_22 br_22 wl_169 vdd gnd cell_6t
Xbit_r170_c22 bl_22 br_22 wl_170 vdd gnd cell_6t
Xbit_r171_c22 bl_22 br_22 wl_171 vdd gnd cell_6t
Xbit_r172_c22 bl_22 br_22 wl_172 vdd gnd cell_6t
Xbit_r173_c22 bl_22 br_22 wl_173 vdd gnd cell_6t
Xbit_r174_c22 bl_22 br_22 wl_174 vdd gnd cell_6t
Xbit_r175_c22 bl_22 br_22 wl_175 vdd gnd cell_6t
Xbit_r176_c22 bl_22 br_22 wl_176 vdd gnd cell_6t
Xbit_r177_c22 bl_22 br_22 wl_177 vdd gnd cell_6t
Xbit_r178_c22 bl_22 br_22 wl_178 vdd gnd cell_6t
Xbit_r179_c22 bl_22 br_22 wl_179 vdd gnd cell_6t
Xbit_r180_c22 bl_22 br_22 wl_180 vdd gnd cell_6t
Xbit_r181_c22 bl_22 br_22 wl_181 vdd gnd cell_6t
Xbit_r182_c22 bl_22 br_22 wl_182 vdd gnd cell_6t
Xbit_r183_c22 bl_22 br_22 wl_183 vdd gnd cell_6t
Xbit_r184_c22 bl_22 br_22 wl_184 vdd gnd cell_6t
Xbit_r185_c22 bl_22 br_22 wl_185 vdd gnd cell_6t
Xbit_r186_c22 bl_22 br_22 wl_186 vdd gnd cell_6t
Xbit_r187_c22 bl_22 br_22 wl_187 vdd gnd cell_6t
Xbit_r188_c22 bl_22 br_22 wl_188 vdd gnd cell_6t
Xbit_r189_c22 bl_22 br_22 wl_189 vdd gnd cell_6t
Xbit_r190_c22 bl_22 br_22 wl_190 vdd gnd cell_6t
Xbit_r191_c22 bl_22 br_22 wl_191 vdd gnd cell_6t
Xbit_r192_c22 bl_22 br_22 wl_192 vdd gnd cell_6t
Xbit_r193_c22 bl_22 br_22 wl_193 vdd gnd cell_6t
Xbit_r194_c22 bl_22 br_22 wl_194 vdd gnd cell_6t
Xbit_r195_c22 bl_22 br_22 wl_195 vdd gnd cell_6t
Xbit_r196_c22 bl_22 br_22 wl_196 vdd gnd cell_6t
Xbit_r197_c22 bl_22 br_22 wl_197 vdd gnd cell_6t
Xbit_r198_c22 bl_22 br_22 wl_198 vdd gnd cell_6t
Xbit_r199_c22 bl_22 br_22 wl_199 vdd gnd cell_6t
Xbit_r200_c22 bl_22 br_22 wl_200 vdd gnd cell_6t
Xbit_r201_c22 bl_22 br_22 wl_201 vdd gnd cell_6t
Xbit_r202_c22 bl_22 br_22 wl_202 vdd gnd cell_6t
Xbit_r203_c22 bl_22 br_22 wl_203 vdd gnd cell_6t
Xbit_r204_c22 bl_22 br_22 wl_204 vdd gnd cell_6t
Xbit_r205_c22 bl_22 br_22 wl_205 vdd gnd cell_6t
Xbit_r206_c22 bl_22 br_22 wl_206 vdd gnd cell_6t
Xbit_r207_c22 bl_22 br_22 wl_207 vdd gnd cell_6t
Xbit_r208_c22 bl_22 br_22 wl_208 vdd gnd cell_6t
Xbit_r209_c22 bl_22 br_22 wl_209 vdd gnd cell_6t
Xbit_r210_c22 bl_22 br_22 wl_210 vdd gnd cell_6t
Xbit_r211_c22 bl_22 br_22 wl_211 vdd gnd cell_6t
Xbit_r212_c22 bl_22 br_22 wl_212 vdd gnd cell_6t
Xbit_r213_c22 bl_22 br_22 wl_213 vdd gnd cell_6t
Xbit_r214_c22 bl_22 br_22 wl_214 vdd gnd cell_6t
Xbit_r215_c22 bl_22 br_22 wl_215 vdd gnd cell_6t
Xbit_r216_c22 bl_22 br_22 wl_216 vdd gnd cell_6t
Xbit_r217_c22 bl_22 br_22 wl_217 vdd gnd cell_6t
Xbit_r218_c22 bl_22 br_22 wl_218 vdd gnd cell_6t
Xbit_r219_c22 bl_22 br_22 wl_219 vdd gnd cell_6t
Xbit_r220_c22 bl_22 br_22 wl_220 vdd gnd cell_6t
Xbit_r221_c22 bl_22 br_22 wl_221 vdd gnd cell_6t
Xbit_r222_c22 bl_22 br_22 wl_222 vdd gnd cell_6t
Xbit_r223_c22 bl_22 br_22 wl_223 vdd gnd cell_6t
Xbit_r224_c22 bl_22 br_22 wl_224 vdd gnd cell_6t
Xbit_r225_c22 bl_22 br_22 wl_225 vdd gnd cell_6t
Xbit_r226_c22 bl_22 br_22 wl_226 vdd gnd cell_6t
Xbit_r227_c22 bl_22 br_22 wl_227 vdd gnd cell_6t
Xbit_r228_c22 bl_22 br_22 wl_228 vdd gnd cell_6t
Xbit_r229_c22 bl_22 br_22 wl_229 vdd gnd cell_6t
Xbit_r230_c22 bl_22 br_22 wl_230 vdd gnd cell_6t
Xbit_r231_c22 bl_22 br_22 wl_231 vdd gnd cell_6t
Xbit_r232_c22 bl_22 br_22 wl_232 vdd gnd cell_6t
Xbit_r233_c22 bl_22 br_22 wl_233 vdd gnd cell_6t
Xbit_r234_c22 bl_22 br_22 wl_234 vdd gnd cell_6t
Xbit_r235_c22 bl_22 br_22 wl_235 vdd gnd cell_6t
Xbit_r236_c22 bl_22 br_22 wl_236 vdd gnd cell_6t
Xbit_r237_c22 bl_22 br_22 wl_237 vdd gnd cell_6t
Xbit_r238_c22 bl_22 br_22 wl_238 vdd gnd cell_6t
Xbit_r239_c22 bl_22 br_22 wl_239 vdd gnd cell_6t
Xbit_r240_c22 bl_22 br_22 wl_240 vdd gnd cell_6t
Xbit_r241_c22 bl_22 br_22 wl_241 vdd gnd cell_6t
Xbit_r242_c22 bl_22 br_22 wl_242 vdd gnd cell_6t
Xbit_r243_c22 bl_22 br_22 wl_243 vdd gnd cell_6t
Xbit_r244_c22 bl_22 br_22 wl_244 vdd gnd cell_6t
Xbit_r245_c22 bl_22 br_22 wl_245 vdd gnd cell_6t
Xbit_r246_c22 bl_22 br_22 wl_246 vdd gnd cell_6t
Xbit_r247_c22 bl_22 br_22 wl_247 vdd gnd cell_6t
Xbit_r248_c22 bl_22 br_22 wl_248 vdd gnd cell_6t
Xbit_r249_c22 bl_22 br_22 wl_249 vdd gnd cell_6t
Xbit_r250_c22 bl_22 br_22 wl_250 vdd gnd cell_6t
Xbit_r251_c22 bl_22 br_22 wl_251 vdd gnd cell_6t
Xbit_r252_c22 bl_22 br_22 wl_252 vdd gnd cell_6t
Xbit_r253_c22 bl_22 br_22 wl_253 vdd gnd cell_6t
Xbit_r254_c22 bl_22 br_22 wl_254 vdd gnd cell_6t
Xbit_r255_c22 bl_22 br_22 wl_255 vdd gnd cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd cell_6t
Xbit_r1_c23 bl_23 br_23 wl_1 vdd gnd cell_6t
Xbit_r2_c23 bl_23 br_23 wl_2 vdd gnd cell_6t
Xbit_r3_c23 bl_23 br_23 wl_3 vdd gnd cell_6t
Xbit_r4_c23 bl_23 br_23 wl_4 vdd gnd cell_6t
Xbit_r5_c23 bl_23 br_23 wl_5 vdd gnd cell_6t
Xbit_r6_c23 bl_23 br_23 wl_6 vdd gnd cell_6t
Xbit_r7_c23 bl_23 br_23 wl_7 vdd gnd cell_6t
Xbit_r8_c23 bl_23 br_23 wl_8 vdd gnd cell_6t
Xbit_r9_c23 bl_23 br_23 wl_9 vdd gnd cell_6t
Xbit_r10_c23 bl_23 br_23 wl_10 vdd gnd cell_6t
Xbit_r11_c23 bl_23 br_23 wl_11 vdd gnd cell_6t
Xbit_r12_c23 bl_23 br_23 wl_12 vdd gnd cell_6t
Xbit_r13_c23 bl_23 br_23 wl_13 vdd gnd cell_6t
Xbit_r14_c23 bl_23 br_23 wl_14 vdd gnd cell_6t
Xbit_r15_c23 bl_23 br_23 wl_15 vdd gnd cell_6t
Xbit_r16_c23 bl_23 br_23 wl_16 vdd gnd cell_6t
Xbit_r17_c23 bl_23 br_23 wl_17 vdd gnd cell_6t
Xbit_r18_c23 bl_23 br_23 wl_18 vdd gnd cell_6t
Xbit_r19_c23 bl_23 br_23 wl_19 vdd gnd cell_6t
Xbit_r20_c23 bl_23 br_23 wl_20 vdd gnd cell_6t
Xbit_r21_c23 bl_23 br_23 wl_21 vdd gnd cell_6t
Xbit_r22_c23 bl_23 br_23 wl_22 vdd gnd cell_6t
Xbit_r23_c23 bl_23 br_23 wl_23 vdd gnd cell_6t
Xbit_r24_c23 bl_23 br_23 wl_24 vdd gnd cell_6t
Xbit_r25_c23 bl_23 br_23 wl_25 vdd gnd cell_6t
Xbit_r26_c23 bl_23 br_23 wl_26 vdd gnd cell_6t
Xbit_r27_c23 bl_23 br_23 wl_27 vdd gnd cell_6t
Xbit_r28_c23 bl_23 br_23 wl_28 vdd gnd cell_6t
Xbit_r29_c23 bl_23 br_23 wl_29 vdd gnd cell_6t
Xbit_r30_c23 bl_23 br_23 wl_30 vdd gnd cell_6t
Xbit_r31_c23 bl_23 br_23 wl_31 vdd gnd cell_6t
Xbit_r32_c23 bl_23 br_23 wl_32 vdd gnd cell_6t
Xbit_r33_c23 bl_23 br_23 wl_33 vdd gnd cell_6t
Xbit_r34_c23 bl_23 br_23 wl_34 vdd gnd cell_6t
Xbit_r35_c23 bl_23 br_23 wl_35 vdd gnd cell_6t
Xbit_r36_c23 bl_23 br_23 wl_36 vdd gnd cell_6t
Xbit_r37_c23 bl_23 br_23 wl_37 vdd gnd cell_6t
Xbit_r38_c23 bl_23 br_23 wl_38 vdd gnd cell_6t
Xbit_r39_c23 bl_23 br_23 wl_39 vdd gnd cell_6t
Xbit_r40_c23 bl_23 br_23 wl_40 vdd gnd cell_6t
Xbit_r41_c23 bl_23 br_23 wl_41 vdd gnd cell_6t
Xbit_r42_c23 bl_23 br_23 wl_42 vdd gnd cell_6t
Xbit_r43_c23 bl_23 br_23 wl_43 vdd gnd cell_6t
Xbit_r44_c23 bl_23 br_23 wl_44 vdd gnd cell_6t
Xbit_r45_c23 bl_23 br_23 wl_45 vdd gnd cell_6t
Xbit_r46_c23 bl_23 br_23 wl_46 vdd gnd cell_6t
Xbit_r47_c23 bl_23 br_23 wl_47 vdd gnd cell_6t
Xbit_r48_c23 bl_23 br_23 wl_48 vdd gnd cell_6t
Xbit_r49_c23 bl_23 br_23 wl_49 vdd gnd cell_6t
Xbit_r50_c23 bl_23 br_23 wl_50 vdd gnd cell_6t
Xbit_r51_c23 bl_23 br_23 wl_51 vdd gnd cell_6t
Xbit_r52_c23 bl_23 br_23 wl_52 vdd gnd cell_6t
Xbit_r53_c23 bl_23 br_23 wl_53 vdd gnd cell_6t
Xbit_r54_c23 bl_23 br_23 wl_54 vdd gnd cell_6t
Xbit_r55_c23 bl_23 br_23 wl_55 vdd gnd cell_6t
Xbit_r56_c23 bl_23 br_23 wl_56 vdd gnd cell_6t
Xbit_r57_c23 bl_23 br_23 wl_57 vdd gnd cell_6t
Xbit_r58_c23 bl_23 br_23 wl_58 vdd gnd cell_6t
Xbit_r59_c23 bl_23 br_23 wl_59 vdd gnd cell_6t
Xbit_r60_c23 bl_23 br_23 wl_60 vdd gnd cell_6t
Xbit_r61_c23 bl_23 br_23 wl_61 vdd gnd cell_6t
Xbit_r62_c23 bl_23 br_23 wl_62 vdd gnd cell_6t
Xbit_r63_c23 bl_23 br_23 wl_63 vdd gnd cell_6t
Xbit_r64_c23 bl_23 br_23 wl_64 vdd gnd cell_6t
Xbit_r65_c23 bl_23 br_23 wl_65 vdd gnd cell_6t
Xbit_r66_c23 bl_23 br_23 wl_66 vdd gnd cell_6t
Xbit_r67_c23 bl_23 br_23 wl_67 vdd gnd cell_6t
Xbit_r68_c23 bl_23 br_23 wl_68 vdd gnd cell_6t
Xbit_r69_c23 bl_23 br_23 wl_69 vdd gnd cell_6t
Xbit_r70_c23 bl_23 br_23 wl_70 vdd gnd cell_6t
Xbit_r71_c23 bl_23 br_23 wl_71 vdd gnd cell_6t
Xbit_r72_c23 bl_23 br_23 wl_72 vdd gnd cell_6t
Xbit_r73_c23 bl_23 br_23 wl_73 vdd gnd cell_6t
Xbit_r74_c23 bl_23 br_23 wl_74 vdd gnd cell_6t
Xbit_r75_c23 bl_23 br_23 wl_75 vdd gnd cell_6t
Xbit_r76_c23 bl_23 br_23 wl_76 vdd gnd cell_6t
Xbit_r77_c23 bl_23 br_23 wl_77 vdd gnd cell_6t
Xbit_r78_c23 bl_23 br_23 wl_78 vdd gnd cell_6t
Xbit_r79_c23 bl_23 br_23 wl_79 vdd gnd cell_6t
Xbit_r80_c23 bl_23 br_23 wl_80 vdd gnd cell_6t
Xbit_r81_c23 bl_23 br_23 wl_81 vdd gnd cell_6t
Xbit_r82_c23 bl_23 br_23 wl_82 vdd gnd cell_6t
Xbit_r83_c23 bl_23 br_23 wl_83 vdd gnd cell_6t
Xbit_r84_c23 bl_23 br_23 wl_84 vdd gnd cell_6t
Xbit_r85_c23 bl_23 br_23 wl_85 vdd gnd cell_6t
Xbit_r86_c23 bl_23 br_23 wl_86 vdd gnd cell_6t
Xbit_r87_c23 bl_23 br_23 wl_87 vdd gnd cell_6t
Xbit_r88_c23 bl_23 br_23 wl_88 vdd gnd cell_6t
Xbit_r89_c23 bl_23 br_23 wl_89 vdd gnd cell_6t
Xbit_r90_c23 bl_23 br_23 wl_90 vdd gnd cell_6t
Xbit_r91_c23 bl_23 br_23 wl_91 vdd gnd cell_6t
Xbit_r92_c23 bl_23 br_23 wl_92 vdd gnd cell_6t
Xbit_r93_c23 bl_23 br_23 wl_93 vdd gnd cell_6t
Xbit_r94_c23 bl_23 br_23 wl_94 vdd gnd cell_6t
Xbit_r95_c23 bl_23 br_23 wl_95 vdd gnd cell_6t
Xbit_r96_c23 bl_23 br_23 wl_96 vdd gnd cell_6t
Xbit_r97_c23 bl_23 br_23 wl_97 vdd gnd cell_6t
Xbit_r98_c23 bl_23 br_23 wl_98 vdd gnd cell_6t
Xbit_r99_c23 bl_23 br_23 wl_99 vdd gnd cell_6t
Xbit_r100_c23 bl_23 br_23 wl_100 vdd gnd cell_6t
Xbit_r101_c23 bl_23 br_23 wl_101 vdd gnd cell_6t
Xbit_r102_c23 bl_23 br_23 wl_102 vdd gnd cell_6t
Xbit_r103_c23 bl_23 br_23 wl_103 vdd gnd cell_6t
Xbit_r104_c23 bl_23 br_23 wl_104 vdd gnd cell_6t
Xbit_r105_c23 bl_23 br_23 wl_105 vdd gnd cell_6t
Xbit_r106_c23 bl_23 br_23 wl_106 vdd gnd cell_6t
Xbit_r107_c23 bl_23 br_23 wl_107 vdd gnd cell_6t
Xbit_r108_c23 bl_23 br_23 wl_108 vdd gnd cell_6t
Xbit_r109_c23 bl_23 br_23 wl_109 vdd gnd cell_6t
Xbit_r110_c23 bl_23 br_23 wl_110 vdd gnd cell_6t
Xbit_r111_c23 bl_23 br_23 wl_111 vdd gnd cell_6t
Xbit_r112_c23 bl_23 br_23 wl_112 vdd gnd cell_6t
Xbit_r113_c23 bl_23 br_23 wl_113 vdd gnd cell_6t
Xbit_r114_c23 bl_23 br_23 wl_114 vdd gnd cell_6t
Xbit_r115_c23 bl_23 br_23 wl_115 vdd gnd cell_6t
Xbit_r116_c23 bl_23 br_23 wl_116 vdd gnd cell_6t
Xbit_r117_c23 bl_23 br_23 wl_117 vdd gnd cell_6t
Xbit_r118_c23 bl_23 br_23 wl_118 vdd gnd cell_6t
Xbit_r119_c23 bl_23 br_23 wl_119 vdd gnd cell_6t
Xbit_r120_c23 bl_23 br_23 wl_120 vdd gnd cell_6t
Xbit_r121_c23 bl_23 br_23 wl_121 vdd gnd cell_6t
Xbit_r122_c23 bl_23 br_23 wl_122 vdd gnd cell_6t
Xbit_r123_c23 bl_23 br_23 wl_123 vdd gnd cell_6t
Xbit_r124_c23 bl_23 br_23 wl_124 vdd gnd cell_6t
Xbit_r125_c23 bl_23 br_23 wl_125 vdd gnd cell_6t
Xbit_r126_c23 bl_23 br_23 wl_126 vdd gnd cell_6t
Xbit_r127_c23 bl_23 br_23 wl_127 vdd gnd cell_6t
Xbit_r128_c23 bl_23 br_23 wl_128 vdd gnd cell_6t
Xbit_r129_c23 bl_23 br_23 wl_129 vdd gnd cell_6t
Xbit_r130_c23 bl_23 br_23 wl_130 vdd gnd cell_6t
Xbit_r131_c23 bl_23 br_23 wl_131 vdd gnd cell_6t
Xbit_r132_c23 bl_23 br_23 wl_132 vdd gnd cell_6t
Xbit_r133_c23 bl_23 br_23 wl_133 vdd gnd cell_6t
Xbit_r134_c23 bl_23 br_23 wl_134 vdd gnd cell_6t
Xbit_r135_c23 bl_23 br_23 wl_135 vdd gnd cell_6t
Xbit_r136_c23 bl_23 br_23 wl_136 vdd gnd cell_6t
Xbit_r137_c23 bl_23 br_23 wl_137 vdd gnd cell_6t
Xbit_r138_c23 bl_23 br_23 wl_138 vdd gnd cell_6t
Xbit_r139_c23 bl_23 br_23 wl_139 vdd gnd cell_6t
Xbit_r140_c23 bl_23 br_23 wl_140 vdd gnd cell_6t
Xbit_r141_c23 bl_23 br_23 wl_141 vdd gnd cell_6t
Xbit_r142_c23 bl_23 br_23 wl_142 vdd gnd cell_6t
Xbit_r143_c23 bl_23 br_23 wl_143 vdd gnd cell_6t
Xbit_r144_c23 bl_23 br_23 wl_144 vdd gnd cell_6t
Xbit_r145_c23 bl_23 br_23 wl_145 vdd gnd cell_6t
Xbit_r146_c23 bl_23 br_23 wl_146 vdd gnd cell_6t
Xbit_r147_c23 bl_23 br_23 wl_147 vdd gnd cell_6t
Xbit_r148_c23 bl_23 br_23 wl_148 vdd gnd cell_6t
Xbit_r149_c23 bl_23 br_23 wl_149 vdd gnd cell_6t
Xbit_r150_c23 bl_23 br_23 wl_150 vdd gnd cell_6t
Xbit_r151_c23 bl_23 br_23 wl_151 vdd gnd cell_6t
Xbit_r152_c23 bl_23 br_23 wl_152 vdd gnd cell_6t
Xbit_r153_c23 bl_23 br_23 wl_153 vdd gnd cell_6t
Xbit_r154_c23 bl_23 br_23 wl_154 vdd gnd cell_6t
Xbit_r155_c23 bl_23 br_23 wl_155 vdd gnd cell_6t
Xbit_r156_c23 bl_23 br_23 wl_156 vdd gnd cell_6t
Xbit_r157_c23 bl_23 br_23 wl_157 vdd gnd cell_6t
Xbit_r158_c23 bl_23 br_23 wl_158 vdd gnd cell_6t
Xbit_r159_c23 bl_23 br_23 wl_159 vdd gnd cell_6t
Xbit_r160_c23 bl_23 br_23 wl_160 vdd gnd cell_6t
Xbit_r161_c23 bl_23 br_23 wl_161 vdd gnd cell_6t
Xbit_r162_c23 bl_23 br_23 wl_162 vdd gnd cell_6t
Xbit_r163_c23 bl_23 br_23 wl_163 vdd gnd cell_6t
Xbit_r164_c23 bl_23 br_23 wl_164 vdd gnd cell_6t
Xbit_r165_c23 bl_23 br_23 wl_165 vdd gnd cell_6t
Xbit_r166_c23 bl_23 br_23 wl_166 vdd gnd cell_6t
Xbit_r167_c23 bl_23 br_23 wl_167 vdd gnd cell_6t
Xbit_r168_c23 bl_23 br_23 wl_168 vdd gnd cell_6t
Xbit_r169_c23 bl_23 br_23 wl_169 vdd gnd cell_6t
Xbit_r170_c23 bl_23 br_23 wl_170 vdd gnd cell_6t
Xbit_r171_c23 bl_23 br_23 wl_171 vdd gnd cell_6t
Xbit_r172_c23 bl_23 br_23 wl_172 vdd gnd cell_6t
Xbit_r173_c23 bl_23 br_23 wl_173 vdd gnd cell_6t
Xbit_r174_c23 bl_23 br_23 wl_174 vdd gnd cell_6t
Xbit_r175_c23 bl_23 br_23 wl_175 vdd gnd cell_6t
Xbit_r176_c23 bl_23 br_23 wl_176 vdd gnd cell_6t
Xbit_r177_c23 bl_23 br_23 wl_177 vdd gnd cell_6t
Xbit_r178_c23 bl_23 br_23 wl_178 vdd gnd cell_6t
Xbit_r179_c23 bl_23 br_23 wl_179 vdd gnd cell_6t
Xbit_r180_c23 bl_23 br_23 wl_180 vdd gnd cell_6t
Xbit_r181_c23 bl_23 br_23 wl_181 vdd gnd cell_6t
Xbit_r182_c23 bl_23 br_23 wl_182 vdd gnd cell_6t
Xbit_r183_c23 bl_23 br_23 wl_183 vdd gnd cell_6t
Xbit_r184_c23 bl_23 br_23 wl_184 vdd gnd cell_6t
Xbit_r185_c23 bl_23 br_23 wl_185 vdd gnd cell_6t
Xbit_r186_c23 bl_23 br_23 wl_186 vdd gnd cell_6t
Xbit_r187_c23 bl_23 br_23 wl_187 vdd gnd cell_6t
Xbit_r188_c23 bl_23 br_23 wl_188 vdd gnd cell_6t
Xbit_r189_c23 bl_23 br_23 wl_189 vdd gnd cell_6t
Xbit_r190_c23 bl_23 br_23 wl_190 vdd gnd cell_6t
Xbit_r191_c23 bl_23 br_23 wl_191 vdd gnd cell_6t
Xbit_r192_c23 bl_23 br_23 wl_192 vdd gnd cell_6t
Xbit_r193_c23 bl_23 br_23 wl_193 vdd gnd cell_6t
Xbit_r194_c23 bl_23 br_23 wl_194 vdd gnd cell_6t
Xbit_r195_c23 bl_23 br_23 wl_195 vdd gnd cell_6t
Xbit_r196_c23 bl_23 br_23 wl_196 vdd gnd cell_6t
Xbit_r197_c23 bl_23 br_23 wl_197 vdd gnd cell_6t
Xbit_r198_c23 bl_23 br_23 wl_198 vdd gnd cell_6t
Xbit_r199_c23 bl_23 br_23 wl_199 vdd gnd cell_6t
Xbit_r200_c23 bl_23 br_23 wl_200 vdd gnd cell_6t
Xbit_r201_c23 bl_23 br_23 wl_201 vdd gnd cell_6t
Xbit_r202_c23 bl_23 br_23 wl_202 vdd gnd cell_6t
Xbit_r203_c23 bl_23 br_23 wl_203 vdd gnd cell_6t
Xbit_r204_c23 bl_23 br_23 wl_204 vdd gnd cell_6t
Xbit_r205_c23 bl_23 br_23 wl_205 vdd gnd cell_6t
Xbit_r206_c23 bl_23 br_23 wl_206 vdd gnd cell_6t
Xbit_r207_c23 bl_23 br_23 wl_207 vdd gnd cell_6t
Xbit_r208_c23 bl_23 br_23 wl_208 vdd gnd cell_6t
Xbit_r209_c23 bl_23 br_23 wl_209 vdd gnd cell_6t
Xbit_r210_c23 bl_23 br_23 wl_210 vdd gnd cell_6t
Xbit_r211_c23 bl_23 br_23 wl_211 vdd gnd cell_6t
Xbit_r212_c23 bl_23 br_23 wl_212 vdd gnd cell_6t
Xbit_r213_c23 bl_23 br_23 wl_213 vdd gnd cell_6t
Xbit_r214_c23 bl_23 br_23 wl_214 vdd gnd cell_6t
Xbit_r215_c23 bl_23 br_23 wl_215 vdd gnd cell_6t
Xbit_r216_c23 bl_23 br_23 wl_216 vdd gnd cell_6t
Xbit_r217_c23 bl_23 br_23 wl_217 vdd gnd cell_6t
Xbit_r218_c23 bl_23 br_23 wl_218 vdd gnd cell_6t
Xbit_r219_c23 bl_23 br_23 wl_219 vdd gnd cell_6t
Xbit_r220_c23 bl_23 br_23 wl_220 vdd gnd cell_6t
Xbit_r221_c23 bl_23 br_23 wl_221 vdd gnd cell_6t
Xbit_r222_c23 bl_23 br_23 wl_222 vdd gnd cell_6t
Xbit_r223_c23 bl_23 br_23 wl_223 vdd gnd cell_6t
Xbit_r224_c23 bl_23 br_23 wl_224 vdd gnd cell_6t
Xbit_r225_c23 bl_23 br_23 wl_225 vdd gnd cell_6t
Xbit_r226_c23 bl_23 br_23 wl_226 vdd gnd cell_6t
Xbit_r227_c23 bl_23 br_23 wl_227 vdd gnd cell_6t
Xbit_r228_c23 bl_23 br_23 wl_228 vdd gnd cell_6t
Xbit_r229_c23 bl_23 br_23 wl_229 vdd gnd cell_6t
Xbit_r230_c23 bl_23 br_23 wl_230 vdd gnd cell_6t
Xbit_r231_c23 bl_23 br_23 wl_231 vdd gnd cell_6t
Xbit_r232_c23 bl_23 br_23 wl_232 vdd gnd cell_6t
Xbit_r233_c23 bl_23 br_23 wl_233 vdd gnd cell_6t
Xbit_r234_c23 bl_23 br_23 wl_234 vdd gnd cell_6t
Xbit_r235_c23 bl_23 br_23 wl_235 vdd gnd cell_6t
Xbit_r236_c23 bl_23 br_23 wl_236 vdd gnd cell_6t
Xbit_r237_c23 bl_23 br_23 wl_237 vdd gnd cell_6t
Xbit_r238_c23 bl_23 br_23 wl_238 vdd gnd cell_6t
Xbit_r239_c23 bl_23 br_23 wl_239 vdd gnd cell_6t
Xbit_r240_c23 bl_23 br_23 wl_240 vdd gnd cell_6t
Xbit_r241_c23 bl_23 br_23 wl_241 vdd gnd cell_6t
Xbit_r242_c23 bl_23 br_23 wl_242 vdd gnd cell_6t
Xbit_r243_c23 bl_23 br_23 wl_243 vdd gnd cell_6t
Xbit_r244_c23 bl_23 br_23 wl_244 vdd gnd cell_6t
Xbit_r245_c23 bl_23 br_23 wl_245 vdd gnd cell_6t
Xbit_r246_c23 bl_23 br_23 wl_246 vdd gnd cell_6t
Xbit_r247_c23 bl_23 br_23 wl_247 vdd gnd cell_6t
Xbit_r248_c23 bl_23 br_23 wl_248 vdd gnd cell_6t
Xbit_r249_c23 bl_23 br_23 wl_249 vdd gnd cell_6t
Xbit_r250_c23 bl_23 br_23 wl_250 vdd gnd cell_6t
Xbit_r251_c23 bl_23 br_23 wl_251 vdd gnd cell_6t
Xbit_r252_c23 bl_23 br_23 wl_252 vdd gnd cell_6t
Xbit_r253_c23 bl_23 br_23 wl_253 vdd gnd cell_6t
Xbit_r254_c23 bl_23 br_23 wl_254 vdd gnd cell_6t
Xbit_r255_c23 bl_23 br_23 wl_255 vdd gnd cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd cell_6t
Xbit_r1_c24 bl_24 br_24 wl_1 vdd gnd cell_6t
Xbit_r2_c24 bl_24 br_24 wl_2 vdd gnd cell_6t
Xbit_r3_c24 bl_24 br_24 wl_3 vdd gnd cell_6t
Xbit_r4_c24 bl_24 br_24 wl_4 vdd gnd cell_6t
Xbit_r5_c24 bl_24 br_24 wl_5 vdd gnd cell_6t
Xbit_r6_c24 bl_24 br_24 wl_6 vdd gnd cell_6t
Xbit_r7_c24 bl_24 br_24 wl_7 vdd gnd cell_6t
Xbit_r8_c24 bl_24 br_24 wl_8 vdd gnd cell_6t
Xbit_r9_c24 bl_24 br_24 wl_9 vdd gnd cell_6t
Xbit_r10_c24 bl_24 br_24 wl_10 vdd gnd cell_6t
Xbit_r11_c24 bl_24 br_24 wl_11 vdd gnd cell_6t
Xbit_r12_c24 bl_24 br_24 wl_12 vdd gnd cell_6t
Xbit_r13_c24 bl_24 br_24 wl_13 vdd gnd cell_6t
Xbit_r14_c24 bl_24 br_24 wl_14 vdd gnd cell_6t
Xbit_r15_c24 bl_24 br_24 wl_15 vdd gnd cell_6t
Xbit_r16_c24 bl_24 br_24 wl_16 vdd gnd cell_6t
Xbit_r17_c24 bl_24 br_24 wl_17 vdd gnd cell_6t
Xbit_r18_c24 bl_24 br_24 wl_18 vdd gnd cell_6t
Xbit_r19_c24 bl_24 br_24 wl_19 vdd gnd cell_6t
Xbit_r20_c24 bl_24 br_24 wl_20 vdd gnd cell_6t
Xbit_r21_c24 bl_24 br_24 wl_21 vdd gnd cell_6t
Xbit_r22_c24 bl_24 br_24 wl_22 vdd gnd cell_6t
Xbit_r23_c24 bl_24 br_24 wl_23 vdd gnd cell_6t
Xbit_r24_c24 bl_24 br_24 wl_24 vdd gnd cell_6t
Xbit_r25_c24 bl_24 br_24 wl_25 vdd gnd cell_6t
Xbit_r26_c24 bl_24 br_24 wl_26 vdd gnd cell_6t
Xbit_r27_c24 bl_24 br_24 wl_27 vdd gnd cell_6t
Xbit_r28_c24 bl_24 br_24 wl_28 vdd gnd cell_6t
Xbit_r29_c24 bl_24 br_24 wl_29 vdd gnd cell_6t
Xbit_r30_c24 bl_24 br_24 wl_30 vdd gnd cell_6t
Xbit_r31_c24 bl_24 br_24 wl_31 vdd gnd cell_6t
Xbit_r32_c24 bl_24 br_24 wl_32 vdd gnd cell_6t
Xbit_r33_c24 bl_24 br_24 wl_33 vdd gnd cell_6t
Xbit_r34_c24 bl_24 br_24 wl_34 vdd gnd cell_6t
Xbit_r35_c24 bl_24 br_24 wl_35 vdd gnd cell_6t
Xbit_r36_c24 bl_24 br_24 wl_36 vdd gnd cell_6t
Xbit_r37_c24 bl_24 br_24 wl_37 vdd gnd cell_6t
Xbit_r38_c24 bl_24 br_24 wl_38 vdd gnd cell_6t
Xbit_r39_c24 bl_24 br_24 wl_39 vdd gnd cell_6t
Xbit_r40_c24 bl_24 br_24 wl_40 vdd gnd cell_6t
Xbit_r41_c24 bl_24 br_24 wl_41 vdd gnd cell_6t
Xbit_r42_c24 bl_24 br_24 wl_42 vdd gnd cell_6t
Xbit_r43_c24 bl_24 br_24 wl_43 vdd gnd cell_6t
Xbit_r44_c24 bl_24 br_24 wl_44 vdd gnd cell_6t
Xbit_r45_c24 bl_24 br_24 wl_45 vdd gnd cell_6t
Xbit_r46_c24 bl_24 br_24 wl_46 vdd gnd cell_6t
Xbit_r47_c24 bl_24 br_24 wl_47 vdd gnd cell_6t
Xbit_r48_c24 bl_24 br_24 wl_48 vdd gnd cell_6t
Xbit_r49_c24 bl_24 br_24 wl_49 vdd gnd cell_6t
Xbit_r50_c24 bl_24 br_24 wl_50 vdd gnd cell_6t
Xbit_r51_c24 bl_24 br_24 wl_51 vdd gnd cell_6t
Xbit_r52_c24 bl_24 br_24 wl_52 vdd gnd cell_6t
Xbit_r53_c24 bl_24 br_24 wl_53 vdd gnd cell_6t
Xbit_r54_c24 bl_24 br_24 wl_54 vdd gnd cell_6t
Xbit_r55_c24 bl_24 br_24 wl_55 vdd gnd cell_6t
Xbit_r56_c24 bl_24 br_24 wl_56 vdd gnd cell_6t
Xbit_r57_c24 bl_24 br_24 wl_57 vdd gnd cell_6t
Xbit_r58_c24 bl_24 br_24 wl_58 vdd gnd cell_6t
Xbit_r59_c24 bl_24 br_24 wl_59 vdd gnd cell_6t
Xbit_r60_c24 bl_24 br_24 wl_60 vdd gnd cell_6t
Xbit_r61_c24 bl_24 br_24 wl_61 vdd gnd cell_6t
Xbit_r62_c24 bl_24 br_24 wl_62 vdd gnd cell_6t
Xbit_r63_c24 bl_24 br_24 wl_63 vdd gnd cell_6t
Xbit_r64_c24 bl_24 br_24 wl_64 vdd gnd cell_6t
Xbit_r65_c24 bl_24 br_24 wl_65 vdd gnd cell_6t
Xbit_r66_c24 bl_24 br_24 wl_66 vdd gnd cell_6t
Xbit_r67_c24 bl_24 br_24 wl_67 vdd gnd cell_6t
Xbit_r68_c24 bl_24 br_24 wl_68 vdd gnd cell_6t
Xbit_r69_c24 bl_24 br_24 wl_69 vdd gnd cell_6t
Xbit_r70_c24 bl_24 br_24 wl_70 vdd gnd cell_6t
Xbit_r71_c24 bl_24 br_24 wl_71 vdd gnd cell_6t
Xbit_r72_c24 bl_24 br_24 wl_72 vdd gnd cell_6t
Xbit_r73_c24 bl_24 br_24 wl_73 vdd gnd cell_6t
Xbit_r74_c24 bl_24 br_24 wl_74 vdd gnd cell_6t
Xbit_r75_c24 bl_24 br_24 wl_75 vdd gnd cell_6t
Xbit_r76_c24 bl_24 br_24 wl_76 vdd gnd cell_6t
Xbit_r77_c24 bl_24 br_24 wl_77 vdd gnd cell_6t
Xbit_r78_c24 bl_24 br_24 wl_78 vdd gnd cell_6t
Xbit_r79_c24 bl_24 br_24 wl_79 vdd gnd cell_6t
Xbit_r80_c24 bl_24 br_24 wl_80 vdd gnd cell_6t
Xbit_r81_c24 bl_24 br_24 wl_81 vdd gnd cell_6t
Xbit_r82_c24 bl_24 br_24 wl_82 vdd gnd cell_6t
Xbit_r83_c24 bl_24 br_24 wl_83 vdd gnd cell_6t
Xbit_r84_c24 bl_24 br_24 wl_84 vdd gnd cell_6t
Xbit_r85_c24 bl_24 br_24 wl_85 vdd gnd cell_6t
Xbit_r86_c24 bl_24 br_24 wl_86 vdd gnd cell_6t
Xbit_r87_c24 bl_24 br_24 wl_87 vdd gnd cell_6t
Xbit_r88_c24 bl_24 br_24 wl_88 vdd gnd cell_6t
Xbit_r89_c24 bl_24 br_24 wl_89 vdd gnd cell_6t
Xbit_r90_c24 bl_24 br_24 wl_90 vdd gnd cell_6t
Xbit_r91_c24 bl_24 br_24 wl_91 vdd gnd cell_6t
Xbit_r92_c24 bl_24 br_24 wl_92 vdd gnd cell_6t
Xbit_r93_c24 bl_24 br_24 wl_93 vdd gnd cell_6t
Xbit_r94_c24 bl_24 br_24 wl_94 vdd gnd cell_6t
Xbit_r95_c24 bl_24 br_24 wl_95 vdd gnd cell_6t
Xbit_r96_c24 bl_24 br_24 wl_96 vdd gnd cell_6t
Xbit_r97_c24 bl_24 br_24 wl_97 vdd gnd cell_6t
Xbit_r98_c24 bl_24 br_24 wl_98 vdd gnd cell_6t
Xbit_r99_c24 bl_24 br_24 wl_99 vdd gnd cell_6t
Xbit_r100_c24 bl_24 br_24 wl_100 vdd gnd cell_6t
Xbit_r101_c24 bl_24 br_24 wl_101 vdd gnd cell_6t
Xbit_r102_c24 bl_24 br_24 wl_102 vdd gnd cell_6t
Xbit_r103_c24 bl_24 br_24 wl_103 vdd gnd cell_6t
Xbit_r104_c24 bl_24 br_24 wl_104 vdd gnd cell_6t
Xbit_r105_c24 bl_24 br_24 wl_105 vdd gnd cell_6t
Xbit_r106_c24 bl_24 br_24 wl_106 vdd gnd cell_6t
Xbit_r107_c24 bl_24 br_24 wl_107 vdd gnd cell_6t
Xbit_r108_c24 bl_24 br_24 wl_108 vdd gnd cell_6t
Xbit_r109_c24 bl_24 br_24 wl_109 vdd gnd cell_6t
Xbit_r110_c24 bl_24 br_24 wl_110 vdd gnd cell_6t
Xbit_r111_c24 bl_24 br_24 wl_111 vdd gnd cell_6t
Xbit_r112_c24 bl_24 br_24 wl_112 vdd gnd cell_6t
Xbit_r113_c24 bl_24 br_24 wl_113 vdd gnd cell_6t
Xbit_r114_c24 bl_24 br_24 wl_114 vdd gnd cell_6t
Xbit_r115_c24 bl_24 br_24 wl_115 vdd gnd cell_6t
Xbit_r116_c24 bl_24 br_24 wl_116 vdd gnd cell_6t
Xbit_r117_c24 bl_24 br_24 wl_117 vdd gnd cell_6t
Xbit_r118_c24 bl_24 br_24 wl_118 vdd gnd cell_6t
Xbit_r119_c24 bl_24 br_24 wl_119 vdd gnd cell_6t
Xbit_r120_c24 bl_24 br_24 wl_120 vdd gnd cell_6t
Xbit_r121_c24 bl_24 br_24 wl_121 vdd gnd cell_6t
Xbit_r122_c24 bl_24 br_24 wl_122 vdd gnd cell_6t
Xbit_r123_c24 bl_24 br_24 wl_123 vdd gnd cell_6t
Xbit_r124_c24 bl_24 br_24 wl_124 vdd gnd cell_6t
Xbit_r125_c24 bl_24 br_24 wl_125 vdd gnd cell_6t
Xbit_r126_c24 bl_24 br_24 wl_126 vdd gnd cell_6t
Xbit_r127_c24 bl_24 br_24 wl_127 vdd gnd cell_6t
Xbit_r128_c24 bl_24 br_24 wl_128 vdd gnd cell_6t
Xbit_r129_c24 bl_24 br_24 wl_129 vdd gnd cell_6t
Xbit_r130_c24 bl_24 br_24 wl_130 vdd gnd cell_6t
Xbit_r131_c24 bl_24 br_24 wl_131 vdd gnd cell_6t
Xbit_r132_c24 bl_24 br_24 wl_132 vdd gnd cell_6t
Xbit_r133_c24 bl_24 br_24 wl_133 vdd gnd cell_6t
Xbit_r134_c24 bl_24 br_24 wl_134 vdd gnd cell_6t
Xbit_r135_c24 bl_24 br_24 wl_135 vdd gnd cell_6t
Xbit_r136_c24 bl_24 br_24 wl_136 vdd gnd cell_6t
Xbit_r137_c24 bl_24 br_24 wl_137 vdd gnd cell_6t
Xbit_r138_c24 bl_24 br_24 wl_138 vdd gnd cell_6t
Xbit_r139_c24 bl_24 br_24 wl_139 vdd gnd cell_6t
Xbit_r140_c24 bl_24 br_24 wl_140 vdd gnd cell_6t
Xbit_r141_c24 bl_24 br_24 wl_141 vdd gnd cell_6t
Xbit_r142_c24 bl_24 br_24 wl_142 vdd gnd cell_6t
Xbit_r143_c24 bl_24 br_24 wl_143 vdd gnd cell_6t
Xbit_r144_c24 bl_24 br_24 wl_144 vdd gnd cell_6t
Xbit_r145_c24 bl_24 br_24 wl_145 vdd gnd cell_6t
Xbit_r146_c24 bl_24 br_24 wl_146 vdd gnd cell_6t
Xbit_r147_c24 bl_24 br_24 wl_147 vdd gnd cell_6t
Xbit_r148_c24 bl_24 br_24 wl_148 vdd gnd cell_6t
Xbit_r149_c24 bl_24 br_24 wl_149 vdd gnd cell_6t
Xbit_r150_c24 bl_24 br_24 wl_150 vdd gnd cell_6t
Xbit_r151_c24 bl_24 br_24 wl_151 vdd gnd cell_6t
Xbit_r152_c24 bl_24 br_24 wl_152 vdd gnd cell_6t
Xbit_r153_c24 bl_24 br_24 wl_153 vdd gnd cell_6t
Xbit_r154_c24 bl_24 br_24 wl_154 vdd gnd cell_6t
Xbit_r155_c24 bl_24 br_24 wl_155 vdd gnd cell_6t
Xbit_r156_c24 bl_24 br_24 wl_156 vdd gnd cell_6t
Xbit_r157_c24 bl_24 br_24 wl_157 vdd gnd cell_6t
Xbit_r158_c24 bl_24 br_24 wl_158 vdd gnd cell_6t
Xbit_r159_c24 bl_24 br_24 wl_159 vdd gnd cell_6t
Xbit_r160_c24 bl_24 br_24 wl_160 vdd gnd cell_6t
Xbit_r161_c24 bl_24 br_24 wl_161 vdd gnd cell_6t
Xbit_r162_c24 bl_24 br_24 wl_162 vdd gnd cell_6t
Xbit_r163_c24 bl_24 br_24 wl_163 vdd gnd cell_6t
Xbit_r164_c24 bl_24 br_24 wl_164 vdd gnd cell_6t
Xbit_r165_c24 bl_24 br_24 wl_165 vdd gnd cell_6t
Xbit_r166_c24 bl_24 br_24 wl_166 vdd gnd cell_6t
Xbit_r167_c24 bl_24 br_24 wl_167 vdd gnd cell_6t
Xbit_r168_c24 bl_24 br_24 wl_168 vdd gnd cell_6t
Xbit_r169_c24 bl_24 br_24 wl_169 vdd gnd cell_6t
Xbit_r170_c24 bl_24 br_24 wl_170 vdd gnd cell_6t
Xbit_r171_c24 bl_24 br_24 wl_171 vdd gnd cell_6t
Xbit_r172_c24 bl_24 br_24 wl_172 vdd gnd cell_6t
Xbit_r173_c24 bl_24 br_24 wl_173 vdd gnd cell_6t
Xbit_r174_c24 bl_24 br_24 wl_174 vdd gnd cell_6t
Xbit_r175_c24 bl_24 br_24 wl_175 vdd gnd cell_6t
Xbit_r176_c24 bl_24 br_24 wl_176 vdd gnd cell_6t
Xbit_r177_c24 bl_24 br_24 wl_177 vdd gnd cell_6t
Xbit_r178_c24 bl_24 br_24 wl_178 vdd gnd cell_6t
Xbit_r179_c24 bl_24 br_24 wl_179 vdd gnd cell_6t
Xbit_r180_c24 bl_24 br_24 wl_180 vdd gnd cell_6t
Xbit_r181_c24 bl_24 br_24 wl_181 vdd gnd cell_6t
Xbit_r182_c24 bl_24 br_24 wl_182 vdd gnd cell_6t
Xbit_r183_c24 bl_24 br_24 wl_183 vdd gnd cell_6t
Xbit_r184_c24 bl_24 br_24 wl_184 vdd gnd cell_6t
Xbit_r185_c24 bl_24 br_24 wl_185 vdd gnd cell_6t
Xbit_r186_c24 bl_24 br_24 wl_186 vdd gnd cell_6t
Xbit_r187_c24 bl_24 br_24 wl_187 vdd gnd cell_6t
Xbit_r188_c24 bl_24 br_24 wl_188 vdd gnd cell_6t
Xbit_r189_c24 bl_24 br_24 wl_189 vdd gnd cell_6t
Xbit_r190_c24 bl_24 br_24 wl_190 vdd gnd cell_6t
Xbit_r191_c24 bl_24 br_24 wl_191 vdd gnd cell_6t
Xbit_r192_c24 bl_24 br_24 wl_192 vdd gnd cell_6t
Xbit_r193_c24 bl_24 br_24 wl_193 vdd gnd cell_6t
Xbit_r194_c24 bl_24 br_24 wl_194 vdd gnd cell_6t
Xbit_r195_c24 bl_24 br_24 wl_195 vdd gnd cell_6t
Xbit_r196_c24 bl_24 br_24 wl_196 vdd gnd cell_6t
Xbit_r197_c24 bl_24 br_24 wl_197 vdd gnd cell_6t
Xbit_r198_c24 bl_24 br_24 wl_198 vdd gnd cell_6t
Xbit_r199_c24 bl_24 br_24 wl_199 vdd gnd cell_6t
Xbit_r200_c24 bl_24 br_24 wl_200 vdd gnd cell_6t
Xbit_r201_c24 bl_24 br_24 wl_201 vdd gnd cell_6t
Xbit_r202_c24 bl_24 br_24 wl_202 vdd gnd cell_6t
Xbit_r203_c24 bl_24 br_24 wl_203 vdd gnd cell_6t
Xbit_r204_c24 bl_24 br_24 wl_204 vdd gnd cell_6t
Xbit_r205_c24 bl_24 br_24 wl_205 vdd gnd cell_6t
Xbit_r206_c24 bl_24 br_24 wl_206 vdd gnd cell_6t
Xbit_r207_c24 bl_24 br_24 wl_207 vdd gnd cell_6t
Xbit_r208_c24 bl_24 br_24 wl_208 vdd gnd cell_6t
Xbit_r209_c24 bl_24 br_24 wl_209 vdd gnd cell_6t
Xbit_r210_c24 bl_24 br_24 wl_210 vdd gnd cell_6t
Xbit_r211_c24 bl_24 br_24 wl_211 vdd gnd cell_6t
Xbit_r212_c24 bl_24 br_24 wl_212 vdd gnd cell_6t
Xbit_r213_c24 bl_24 br_24 wl_213 vdd gnd cell_6t
Xbit_r214_c24 bl_24 br_24 wl_214 vdd gnd cell_6t
Xbit_r215_c24 bl_24 br_24 wl_215 vdd gnd cell_6t
Xbit_r216_c24 bl_24 br_24 wl_216 vdd gnd cell_6t
Xbit_r217_c24 bl_24 br_24 wl_217 vdd gnd cell_6t
Xbit_r218_c24 bl_24 br_24 wl_218 vdd gnd cell_6t
Xbit_r219_c24 bl_24 br_24 wl_219 vdd gnd cell_6t
Xbit_r220_c24 bl_24 br_24 wl_220 vdd gnd cell_6t
Xbit_r221_c24 bl_24 br_24 wl_221 vdd gnd cell_6t
Xbit_r222_c24 bl_24 br_24 wl_222 vdd gnd cell_6t
Xbit_r223_c24 bl_24 br_24 wl_223 vdd gnd cell_6t
Xbit_r224_c24 bl_24 br_24 wl_224 vdd gnd cell_6t
Xbit_r225_c24 bl_24 br_24 wl_225 vdd gnd cell_6t
Xbit_r226_c24 bl_24 br_24 wl_226 vdd gnd cell_6t
Xbit_r227_c24 bl_24 br_24 wl_227 vdd gnd cell_6t
Xbit_r228_c24 bl_24 br_24 wl_228 vdd gnd cell_6t
Xbit_r229_c24 bl_24 br_24 wl_229 vdd gnd cell_6t
Xbit_r230_c24 bl_24 br_24 wl_230 vdd gnd cell_6t
Xbit_r231_c24 bl_24 br_24 wl_231 vdd gnd cell_6t
Xbit_r232_c24 bl_24 br_24 wl_232 vdd gnd cell_6t
Xbit_r233_c24 bl_24 br_24 wl_233 vdd gnd cell_6t
Xbit_r234_c24 bl_24 br_24 wl_234 vdd gnd cell_6t
Xbit_r235_c24 bl_24 br_24 wl_235 vdd gnd cell_6t
Xbit_r236_c24 bl_24 br_24 wl_236 vdd gnd cell_6t
Xbit_r237_c24 bl_24 br_24 wl_237 vdd gnd cell_6t
Xbit_r238_c24 bl_24 br_24 wl_238 vdd gnd cell_6t
Xbit_r239_c24 bl_24 br_24 wl_239 vdd gnd cell_6t
Xbit_r240_c24 bl_24 br_24 wl_240 vdd gnd cell_6t
Xbit_r241_c24 bl_24 br_24 wl_241 vdd gnd cell_6t
Xbit_r242_c24 bl_24 br_24 wl_242 vdd gnd cell_6t
Xbit_r243_c24 bl_24 br_24 wl_243 vdd gnd cell_6t
Xbit_r244_c24 bl_24 br_24 wl_244 vdd gnd cell_6t
Xbit_r245_c24 bl_24 br_24 wl_245 vdd gnd cell_6t
Xbit_r246_c24 bl_24 br_24 wl_246 vdd gnd cell_6t
Xbit_r247_c24 bl_24 br_24 wl_247 vdd gnd cell_6t
Xbit_r248_c24 bl_24 br_24 wl_248 vdd gnd cell_6t
Xbit_r249_c24 bl_24 br_24 wl_249 vdd gnd cell_6t
Xbit_r250_c24 bl_24 br_24 wl_250 vdd gnd cell_6t
Xbit_r251_c24 bl_24 br_24 wl_251 vdd gnd cell_6t
Xbit_r252_c24 bl_24 br_24 wl_252 vdd gnd cell_6t
Xbit_r253_c24 bl_24 br_24 wl_253 vdd gnd cell_6t
Xbit_r254_c24 bl_24 br_24 wl_254 vdd gnd cell_6t
Xbit_r255_c24 bl_24 br_24 wl_255 vdd gnd cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd cell_6t
Xbit_r1_c25 bl_25 br_25 wl_1 vdd gnd cell_6t
Xbit_r2_c25 bl_25 br_25 wl_2 vdd gnd cell_6t
Xbit_r3_c25 bl_25 br_25 wl_3 vdd gnd cell_6t
Xbit_r4_c25 bl_25 br_25 wl_4 vdd gnd cell_6t
Xbit_r5_c25 bl_25 br_25 wl_5 vdd gnd cell_6t
Xbit_r6_c25 bl_25 br_25 wl_6 vdd gnd cell_6t
Xbit_r7_c25 bl_25 br_25 wl_7 vdd gnd cell_6t
Xbit_r8_c25 bl_25 br_25 wl_8 vdd gnd cell_6t
Xbit_r9_c25 bl_25 br_25 wl_9 vdd gnd cell_6t
Xbit_r10_c25 bl_25 br_25 wl_10 vdd gnd cell_6t
Xbit_r11_c25 bl_25 br_25 wl_11 vdd gnd cell_6t
Xbit_r12_c25 bl_25 br_25 wl_12 vdd gnd cell_6t
Xbit_r13_c25 bl_25 br_25 wl_13 vdd gnd cell_6t
Xbit_r14_c25 bl_25 br_25 wl_14 vdd gnd cell_6t
Xbit_r15_c25 bl_25 br_25 wl_15 vdd gnd cell_6t
Xbit_r16_c25 bl_25 br_25 wl_16 vdd gnd cell_6t
Xbit_r17_c25 bl_25 br_25 wl_17 vdd gnd cell_6t
Xbit_r18_c25 bl_25 br_25 wl_18 vdd gnd cell_6t
Xbit_r19_c25 bl_25 br_25 wl_19 vdd gnd cell_6t
Xbit_r20_c25 bl_25 br_25 wl_20 vdd gnd cell_6t
Xbit_r21_c25 bl_25 br_25 wl_21 vdd gnd cell_6t
Xbit_r22_c25 bl_25 br_25 wl_22 vdd gnd cell_6t
Xbit_r23_c25 bl_25 br_25 wl_23 vdd gnd cell_6t
Xbit_r24_c25 bl_25 br_25 wl_24 vdd gnd cell_6t
Xbit_r25_c25 bl_25 br_25 wl_25 vdd gnd cell_6t
Xbit_r26_c25 bl_25 br_25 wl_26 vdd gnd cell_6t
Xbit_r27_c25 bl_25 br_25 wl_27 vdd gnd cell_6t
Xbit_r28_c25 bl_25 br_25 wl_28 vdd gnd cell_6t
Xbit_r29_c25 bl_25 br_25 wl_29 vdd gnd cell_6t
Xbit_r30_c25 bl_25 br_25 wl_30 vdd gnd cell_6t
Xbit_r31_c25 bl_25 br_25 wl_31 vdd gnd cell_6t
Xbit_r32_c25 bl_25 br_25 wl_32 vdd gnd cell_6t
Xbit_r33_c25 bl_25 br_25 wl_33 vdd gnd cell_6t
Xbit_r34_c25 bl_25 br_25 wl_34 vdd gnd cell_6t
Xbit_r35_c25 bl_25 br_25 wl_35 vdd gnd cell_6t
Xbit_r36_c25 bl_25 br_25 wl_36 vdd gnd cell_6t
Xbit_r37_c25 bl_25 br_25 wl_37 vdd gnd cell_6t
Xbit_r38_c25 bl_25 br_25 wl_38 vdd gnd cell_6t
Xbit_r39_c25 bl_25 br_25 wl_39 vdd gnd cell_6t
Xbit_r40_c25 bl_25 br_25 wl_40 vdd gnd cell_6t
Xbit_r41_c25 bl_25 br_25 wl_41 vdd gnd cell_6t
Xbit_r42_c25 bl_25 br_25 wl_42 vdd gnd cell_6t
Xbit_r43_c25 bl_25 br_25 wl_43 vdd gnd cell_6t
Xbit_r44_c25 bl_25 br_25 wl_44 vdd gnd cell_6t
Xbit_r45_c25 bl_25 br_25 wl_45 vdd gnd cell_6t
Xbit_r46_c25 bl_25 br_25 wl_46 vdd gnd cell_6t
Xbit_r47_c25 bl_25 br_25 wl_47 vdd gnd cell_6t
Xbit_r48_c25 bl_25 br_25 wl_48 vdd gnd cell_6t
Xbit_r49_c25 bl_25 br_25 wl_49 vdd gnd cell_6t
Xbit_r50_c25 bl_25 br_25 wl_50 vdd gnd cell_6t
Xbit_r51_c25 bl_25 br_25 wl_51 vdd gnd cell_6t
Xbit_r52_c25 bl_25 br_25 wl_52 vdd gnd cell_6t
Xbit_r53_c25 bl_25 br_25 wl_53 vdd gnd cell_6t
Xbit_r54_c25 bl_25 br_25 wl_54 vdd gnd cell_6t
Xbit_r55_c25 bl_25 br_25 wl_55 vdd gnd cell_6t
Xbit_r56_c25 bl_25 br_25 wl_56 vdd gnd cell_6t
Xbit_r57_c25 bl_25 br_25 wl_57 vdd gnd cell_6t
Xbit_r58_c25 bl_25 br_25 wl_58 vdd gnd cell_6t
Xbit_r59_c25 bl_25 br_25 wl_59 vdd gnd cell_6t
Xbit_r60_c25 bl_25 br_25 wl_60 vdd gnd cell_6t
Xbit_r61_c25 bl_25 br_25 wl_61 vdd gnd cell_6t
Xbit_r62_c25 bl_25 br_25 wl_62 vdd gnd cell_6t
Xbit_r63_c25 bl_25 br_25 wl_63 vdd gnd cell_6t
Xbit_r64_c25 bl_25 br_25 wl_64 vdd gnd cell_6t
Xbit_r65_c25 bl_25 br_25 wl_65 vdd gnd cell_6t
Xbit_r66_c25 bl_25 br_25 wl_66 vdd gnd cell_6t
Xbit_r67_c25 bl_25 br_25 wl_67 vdd gnd cell_6t
Xbit_r68_c25 bl_25 br_25 wl_68 vdd gnd cell_6t
Xbit_r69_c25 bl_25 br_25 wl_69 vdd gnd cell_6t
Xbit_r70_c25 bl_25 br_25 wl_70 vdd gnd cell_6t
Xbit_r71_c25 bl_25 br_25 wl_71 vdd gnd cell_6t
Xbit_r72_c25 bl_25 br_25 wl_72 vdd gnd cell_6t
Xbit_r73_c25 bl_25 br_25 wl_73 vdd gnd cell_6t
Xbit_r74_c25 bl_25 br_25 wl_74 vdd gnd cell_6t
Xbit_r75_c25 bl_25 br_25 wl_75 vdd gnd cell_6t
Xbit_r76_c25 bl_25 br_25 wl_76 vdd gnd cell_6t
Xbit_r77_c25 bl_25 br_25 wl_77 vdd gnd cell_6t
Xbit_r78_c25 bl_25 br_25 wl_78 vdd gnd cell_6t
Xbit_r79_c25 bl_25 br_25 wl_79 vdd gnd cell_6t
Xbit_r80_c25 bl_25 br_25 wl_80 vdd gnd cell_6t
Xbit_r81_c25 bl_25 br_25 wl_81 vdd gnd cell_6t
Xbit_r82_c25 bl_25 br_25 wl_82 vdd gnd cell_6t
Xbit_r83_c25 bl_25 br_25 wl_83 vdd gnd cell_6t
Xbit_r84_c25 bl_25 br_25 wl_84 vdd gnd cell_6t
Xbit_r85_c25 bl_25 br_25 wl_85 vdd gnd cell_6t
Xbit_r86_c25 bl_25 br_25 wl_86 vdd gnd cell_6t
Xbit_r87_c25 bl_25 br_25 wl_87 vdd gnd cell_6t
Xbit_r88_c25 bl_25 br_25 wl_88 vdd gnd cell_6t
Xbit_r89_c25 bl_25 br_25 wl_89 vdd gnd cell_6t
Xbit_r90_c25 bl_25 br_25 wl_90 vdd gnd cell_6t
Xbit_r91_c25 bl_25 br_25 wl_91 vdd gnd cell_6t
Xbit_r92_c25 bl_25 br_25 wl_92 vdd gnd cell_6t
Xbit_r93_c25 bl_25 br_25 wl_93 vdd gnd cell_6t
Xbit_r94_c25 bl_25 br_25 wl_94 vdd gnd cell_6t
Xbit_r95_c25 bl_25 br_25 wl_95 vdd gnd cell_6t
Xbit_r96_c25 bl_25 br_25 wl_96 vdd gnd cell_6t
Xbit_r97_c25 bl_25 br_25 wl_97 vdd gnd cell_6t
Xbit_r98_c25 bl_25 br_25 wl_98 vdd gnd cell_6t
Xbit_r99_c25 bl_25 br_25 wl_99 vdd gnd cell_6t
Xbit_r100_c25 bl_25 br_25 wl_100 vdd gnd cell_6t
Xbit_r101_c25 bl_25 br_25 wl_101 vdd gnd cell_6t
Xbit_r102_c25 bl_25 br_25 wl_102 vdd gnd cell_6t
Xbit_r103_c25 bl_25 br_25 wl_103 vdd gnd cell_6t
Xbit_r104_c25 bl_25 br_25 wl_104 vdd gnd cell_6t
Xbit_r105_c25 bl_25 br_25 wl_105 vdd gnd cell_6t
Xbit_r106_c25 bl_25 br_25 wl_106 vdd gnd cell_6t
Xbit_r107_c25 bl_25 br_25 wl_107 vdd gnd cell_6t
Xbit_r108_c25 bl_25 br_25 wl_108 vdd gnd cell_6t
Xbit_r109_c25 bl_25 br_25 wl_109 vdd gnd cell_6t
Xbit_r110_c25 bl_25 br_25 wl_110 vdd gnd cell_6t
Xbit_r111_c25 bl_25 br_25 wl_111 vdd gnd cell_6t
Xbit_r112_c25 bl_25 br_25 wl_112 vdd gnd cell_6t
Xbit_r113_c25 bl_25 br_25 wl_113 vdd gnd cell_6t
Xbit_r114_c25 bl_25 br_25 wl_114 vdd gnd cell_6t
Xbit_r115_c25 bl_25 br_25 wl_115 vdd gnd cell_6t
Xbit_r116_c25 bl_25 br_25 wl_116 vdd gnd cell_6t
Xbit_r117_c25 bl_25 br_25 wl_117 vdd gnd cell_6t
Xbit_r118_c25 bl_25 br_25 wl_118 vdd gnd cell_6t
Xbit_r119_c25 bl_25 br_25 wl_119 vdd gnd cell_6t
Xbit_r120_c25 bl_25 br_25 wl_120 vdd gnd cell_6t
Xbit_r121_c25 bl_25 br_25 wl_121 vdd gnd cell_6t
Xbit_r122_c25 bl_25 br_25 wl_122 vdd gnd cell_6t
Xbit_r123_c25 bl_25 br_25 wl_123 vdd gnd cell_6t
Xbit_r124_c25 bl_25 br_25 wl_124 vdd gnd cell_6t
Xbit_r125_c25 bl_25 br_25 wl_125 vdd gnd cell_6t
Xbit_r126_c25 bl_25 br_25 wl_126 vdd gnd cell_6t
Xbit_r127_c25 bl_25 br_25 wl_127 vdd gnd cell_6t
Xbit_r128_c25 bl_25 br_25 wl_128 vdd gnd cell_6t
Xbit_r129_c25 bl_25 br_25 wl_129 vdd gnd cell_6t
Xbit_r130_c25 bl_25 br_25 wl_130 vdd gnd cell_6t
Xbit_r131_c25 bl_25 br_25 wl_131 vdd gnd cell_6t
Xbit_r132_c25 bl_25 br_25 wl_132 vdd gnd cell_6t
Xbit_r133_c25 bl_25 br_25 wl_133 vdd gnd cell_6t
Xbit_r134_c25 bl_25 br_25 wl_134 vdd gnd cell_6t
Xbit_r135_c25 bl_25 br_25 wl_135 vdd gnd cell_6t
Xbit_r136_c25 bl_25 br_25 wl_136 vdd gnd cell_6t
Xbit_r137_c25 bl_25 br_25 wl_137 vdd gnd cell_6t
Xbit_r138_c25 bl_25 br_25 wl_138 vdd gnd cell_6t
Xbit_r139_c25 bl_25 br_25 wl_139 vdd gnd cell_6t
Xbit_r140_c25 bl_25 br_25 wl_140 vdd gnd cell_6t
Xbit_r141_c25 bl_25 br_25 wl_141 vdd gnd cell_6t
Xbit_r142_c25 bl_25 br_25 wl_142 vdd gnd cell_6t
Xbit_r143_c25 bl_25 br_25 wl_143 vdd gnd cell_6t
Xbit_r144_c25 bl_25 br_25 wl_144 vdd gnd cell_6t
Xbit_r145_c25 bl_25 br_25 wl_145 vdd gnd cell_6t
Xbit_r146_c25 bl_25 br_25 wl_146 vdd gnd cell_6t
Xbit_r147_c25 bl_25 br_25 wl_147 vdd gnd cell_6t
Xbit_r148_c25 bl_25 br_25 wl_148 vdd gnd cell_6t
Xbit_r149_c25 bl_25 br_25 wl_149 vdd gnd cell_6t
Xbit_r150_c25 bl_25 br_25 wl_150 vdd gnd cell_6t
Xbit_r151_c25 bl_25 br_25 wl_151 vdd gnd cell_6t
Xbit_r152_c25 bl_25 br_25 wl_152 vdd gnd cell_6t
Xbit_r153_c25 bl_25 br_25 wl_153 vdd gnd cell_6t
Xbit_r154_c25 bl_25 br_25 wl_154 vdd gnd cell_6t
Xbit_r155_c25 bl_25 br_25 wl_155 vdd gnd cell_6t
Xbit_r156_c25 bl_25 br_25 wl_156 vdd gnd cell_6t
Xbit_r157_c25 bl_25 br_25 wl_157 vdd gnd cell_6t
Xbit_r158_c25 bl_25 br_25 wl_158 vdd gnd cell_6t
Xbit_r159_c25 bl_25 br_25 wl_159 vdd gnd cell_6t
Xbit_r160_c25 bl_25 br_25 wl_160 vdd gnd cell_6t
Xbit_r161_c25 bl_25 br_25 wl_161 vdd gnd cell_6t
Xbit_r162_c25 bl_25 br_25 wl_162 vdd gnd cell_6t
Xbit_r163_c25 bl_25 br_25 wl_163 vdd gnd cell_6t
Xbit_r164_c25 bl_25 br_25 wl_164 vdd gnd cell_6t
Xbit_r165_c25 bl_25 br_25 wl_165 vdd gnd cell_6t
Xbit_r166_c25 bl_25 br_25 wl_166 vdd gnd cell_6t
Xbit_r167_c25 bl_25 br_25 wl_167 vdd gnd cell_6t
Xbit_r168_c25 bl_25 br_25 wl_168 vdd gnd cell_6t
Xbit_r169_c25 bl_25 br_25 wl_169 vdd gnd cell_6t
Xbit_r170_c25 bl_25 br_25 wl_170 vdd gnd cell_6t
Xbit_r171_c25 bl_25 br_25 wl_171 vdd gnd cell_6t
Xbit_r172_c25 bl_25 br_25 wl_172 vdd gnd cell_6t
Xbit_r173_c25 bl_25 br_25 wl_173 vdd gnd cell_6t
Xbit_r174_c25 bl_25 br_25 wl_174 vdd gnd cell_6t
Xbit_r175_c25 bl_25 br_25 wl_175 vdd gnd cell_6t
Xbit_r176_c25 bl_25 br_25 wl_176 vdd gnd cell_6t
Xbit_r177_c25 bl_25 br_25 wl_177 vdd gnd cell_6t
Xbit_r178_c25 bl_25 br_25 wl_178 vdd gnd cell_6t
Xbit_r179_c25 bl_25 br_25 wl_179 vdd gnd cell_6t
Xbit_r180_c25 bl_25 br_25 wl_180 vdd gnd cell_6t
Xbit_r181_c25 bl_25 br_25 wl_181 vdd gnd cell_6t
Xbit_r182_c25 bl_25 br_25 wl_182 vdd gnd cell_6t
Xbit_r183_c25 bl_25 br_25 wl_183 vdd gnd cell_6t
Xbit_r184_c25 bl_25 br_25 wl_184 vdd gnd cell_6t
Xbit_r185_c25 bl_25 br_25 wl_185 vdd gnd cell_6t
Xbit_r186_c25 bl_25 br_25 wl_186 vdd gnd cell_6t
Xbit_r187_c25 bl_25 br_25 wl_187 vdd gnd cell_6t
Xbit_r188_c25 bl_25 br_25 wl_188 vdd gnd cell_6t
Xbit_r189_c25 bl_25 br_25 wl_189 vdd gnd cell_6t
Xbit_r190_c25 bl_25 br_25 wl_190 vdd gnd cell_6t
Xbit_r191_c25 bl_25 br_25 wl_191 vdd gnd cell_6t
Xbit_r192_c25 bl_25 br_25 wl_192 vdd gnd cell_6t
Xbit_r193_c25 bl_25 br_25 wl_193 vdd gnd cell_6t
Xbit_r194_c25 bl_25 br_25 wl_194 vdd gnd cell_6t
Xbit_r195_c25 bl_25 br_25 wl_195 vdd gnd cell_6t
Xbit_r196_c25 bl_25 br_25 wl_196 vdd gnd cell_6t
Xbit_r197_c25 bl_25 br_25 wl_197 vdd gnd cell_6t
Xbit_r198_c25 bl_25 br_25 wl_198 vdd gnd cell_6t
Xbit_r199_c25 bl_25 br_25 wl_199 vdd gnd cell_6t
Xbit_r200_c25 bl_25 br_25 wl_200 vdd gnd cell_6t
Xbit_r201_c25 bl_25 br_25 wl_201 vdd gnd cell_6t
Xbit_r202_c25 bl_25 br_25 wl_202 vdd gnd cell_6t
Xbit_r203_c25 bl_25 br_25 wl_203 vdd gnd cell_6t
Xbit_r204_c25 bl_25 br_25 wl_204 vdd gnd cell_6t
Xbit_r205_c25 bl_25 br_25 wl_205 vdd gnd cell_6t
Xbit_r206_c25 bl_25 br_25 wl_206 vdd gnd cell_6t
Xbit_r207_c25 bl_25 br_25 wl_207 vdd gnd cell_6t
Xbit_r208_c25 bl_25 br_25 wl_208 vdd gnd cell_6t
Xbit_r209_c25 bl_25 br_25 wl_209 vdd gnd cell_6t
Xbit_r210_c25 bl_25 br_25 wl_210 vdd gnd cell_6t
Xbit_r211_c25 bl_25 br_25 wl_211 vdd gnd cell_6t
Xbit_r212_c25 bl_25 br_25 wl_212 vdd gnd cell_6t
Xbit_r213_c25 bl_25 br_25 wl_213 vdd gnd cell_6t
Xbit_r214_c25 bl_25 br_25 wl_214 vdd gnd cell_6t
Xbit_r215_c25 bl_25 br_25 wl_215 vdd gnd cell_6t
Xbit_r216_c25 bl_25 br_25 wl_216 vdd gnd cell_6t
Xbit_r217_c25 bl_25 br_25 wl_217 vdd gnd cell_6t
Xbit_r218_c25 bl_25 br_25 wl_218 vdd gnd cell_6t
Xbit_r219_c25 bl_25 br_25 wl_219 vdd gnd cell_6t
Xbit_r220_c25 bl_25 br_25 wl_220 vdd gnd cell_6t
Xbit_r221_c25 bl_25 br_25 wl_221 vdd gnd cell_6t
Xbit_r222_c25 bl_25 br_25 wl_222 vdd gnd cell_6t
Xbit_r223_c25 bl_25 br_25 wl_223 vdd gnd cell_6t
Xbit_r224_c25 bl_25 br_25 wl_224 vdd gnd cell_6t
Xbit_r225_c25 bl_25 br_25 wl_225 vdd gnd cell_6t
Xbit_r226_c25 bl_25 br_25 wl_226 vdd gnd cell_6t
Xbit_r227_c25 bl_25 br_25 wl_227 vdd gnd cell_6t
Xbit_r228_c25 bl_25 br_25 wl_228 vdd gnd cell_6t
Xbit_r229_c25 bl_25 br_25 wl_229 vdd gnd cell_6t
Xbit_r230_c25 bl_25 br_25 wl_230 vdd gnd cell_6t
Xbit_r231_c25 bl_25 br_25 wl_231 vdd gnd cell_6t
Xbit_r232_c25 bl_25 br_25 wl_232 vdd gnd cell_6t
Xbit_r233_c25 bl_25 br_25 wl_233 vdd gnd cell_6t
Xbit_r234_c25 bl_25 br_25 wl_234 vdd gnd cell_6t
Xbit_r235_c25 bl_25 br_25 wl_235 vdd gnd cell_6t
Xbit_r236_c25 bl_25 br_25 wl_236 vdd gnd cell_6t
Xbit_r237_c25 bl_25 br_25 wl_237 vdd gnd cell_6t
Xbit_r238_c25 bl_25 br_25 wl_238 vdd gnd cell_6t
Xbit_r239_c25 bl_25 br_25 wl_239 vdd gnd cell_6t
Xbit_r240_c25 bl_25 br_25 wl_240 vdd gnd cell_6t
Xbit_r241_c25 bl_25 br_25 wl_241 vdd gnd cell_6t
Xbit_r242_c25 bl_25 br_25 wl_242 vdd gnd cell_6t
Xbit_r243_c25 bl_25 br_25 wl_243 vdd gnd cell_6t
Xbit_r244_c25 bl_25 br_25 wl_244 vdd gnd cell_6t
Xbit_r245_c25 bl_25 br_25 wl_245 vdd gnd cell_6t
Xbit_r246_c25 bl_25 br_25 wl_246 vdd gnd cell_6t
Xbit_r247_c25 bl_25 br_25 wl_247 vdd gnd cell_6t
Xbit_r248_c25 bl_25 br_25 wl_248 vdd gnd cell_6t
Xbit_r249_c25 bl_25 br_25 wl_249 vdd gnd cell_6t
Xbit_r250_c25 bl_25 br_25 wl_250 vdd gnd cell_6t
Xbit_r251_c25 bl_25 br_25 wl_251 vdd gnd cell_6t
Xbit_r252_c25 bl_25 br_25 wl_252 vdd gnd cell_6t
Xbit_r253_c25 bl_25 br_25 wl_253 vdd gnd cell_6t
Xbit_r254_c25 bl_25 br_25 wl_254 vdd gnd cell_6t
Xbit_r255_c25 bl_25 br_25 wl_255 vdd gnd cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd cell_6t
Xbit_r1_c26 bl_26 br_26 wl_1 vdd gnd cell_6t
Xbit_r2_c26 bl_26 br_26 wl_2 vdd gnd cell_6t
Xbit_r3_c26 bl_26 br_26 wl_3 vdd gnd cell_6t
Xbit_r4_c26 bl_26 br_26 wl_4 vdd gnd cell_6t
Xbit_r5_c26 bl_26 br_26 wl_5 vdd gnd cell_6t
Xbit_r6_c26 bl_26 br_26 wl_6 vdd gnd cell_6t
Xbit_r7_c26 bl_26 br_26 wl_7 vdd gnd cell_6t
Xbit_r8_c26 bl_26 br_26 wl_8 vdd gnd cell_6t
Xbit_r9_c26 bl_26 br_26 wl_9 vdd gnd cell_6t
Xbit_r10_c26 bl_26 br_26 wl_10 vdd gnd cell_6t
Xbit_r11_c26 bl_26 br_26 wl_11 vdd gnd cell_6t
Xbit_r12_c26 bl_26 br_26 wl_12 vdd gnd cell_6t
Xbit_r13_c26 bl_26 br_26 wl_13 vdd gnd cell_6t
Xbit_r14_c26 bl_26 br_26 wl_14 vdd gnd cell_6t
Xbit_r15_c26 bl_26 br_26 wl_15 vdd gnd cell_6t
Xbit_r16_c26 bl_26 br_26 wl_16 vdd gnd cell_6t
Xbit_r17_c26 bl_26 br_26 wl_17 vdd gnd cell_6t
Xbit_r18_c26 bl_26 br_26 wl_18 vdd gnd cell_6t
Xbit_r19_c26 bl_26 br_26 wl_19 vdd gnd cell_6t
Xbit_r20_c26 bl_26 br_26 wl_20 vdd gnd cell_6t
Xbit_r21_c26 bl_26 br_26 wl_21 vdd gnd cell_6t
Xbit_r22_c26 bl_26 br_26 wl_22 vdd gnd cell_6t
Xbit_r23_c26 bl_26 br_26 wl_23 vdd gnd cell_6t
Xbit_r24_c26 bl_26 br_26 wl_24 vdd gnd cell_6t
Xbit_r25_c26 bl_26 br_26 wl_25 vdd gnd cell_6t
Xbit_r26_c26 bl_26 br_26 wl_26 vdd gnd cell_6t
Xbit_r27_c26 bl_26 br_26 wl_27 vdd gnd cell_6t
Xbit_r28_c26 bl_26 br_26 wl_28 vdd gnd cell_6t
Xbit_r29_c26 bl_26 br_26 wl_29 vdd gnd cell_6t
Xbit_r30_c26 bl_26 br_26 wl_30 vdd gnd cell_6t
Xbit_r31_c26 bl_26 br_26 wl_31 vdd gnd cell_6t
Xbit_r32_c26 bl_26 br_26 wl_32 vdd gnd cell_6t
Xbit_r33_c26 bl_26 br_26 wl_33 vdd gnd cell_6t
Xbit_r34_c26 bl_26 br_26 wl_34 vdd gnd cell_6t
Xbit_r35_c26 bl_26 br_26 wl_35 vdd gnd cell_6t
Xbit_r36_c26 bl_26 br_26 wl_36 vdd gnd cell_6t
Xbit_r37_c26 bl_26 br_26 wl_37 vdd gnd cell_6t
Xbit_r38_c26 bl_26 br_26 wl_38 vdd gnd cell_6t
Xbit_r39_c26 bl_26 br_26 wl_39 vdd gnd cell_6t
Xbit_r40_c26 bl_26 br_26 wl_40 vdd gnd cell_6t
Xbit_r41_c26 bl_26 br_26 wl_41 vdd gnd cell_6t
Xbit_r42_c26 bl_26 br_26 wl_42 vdd gnd cell_6t
Xbit_r43_c26 bl_26 br_26 wl_43 vdd gnd cell_6t
Xbit_r44_c26 bl_26 br_26 wl_44 vdd gnd cell_6t
Xbit_r45_c26 bl_26 br_26 wl_45 vdd gnd cell_6t
Xbit_r46_c26 bl_26 br_26 wl_46 vdd gnd cell_6t
Xbit_r47_c26 bl_26 br_26 wl_47 vdd gnd cell_6t
Xbit_r48_c26 bl_26 br_26 wl_48 vdd gnd cell_6t
Xbit_r49_c26 bl_26 br_26 wl_49 vdd gnd cell_6t
Xbit_r50_c26 bl_26 br_26 wl_50 vdd gnd cell_6t
Xbit_r51_c26 bl_26 br_26 wl_51 vdd gnd cell_6t
Xbit_r52_c26 bl_26 br_26 wl_52 vdd gnd cell_6t
Xbit_r53_c26 bl_26 br_26 wl_53 vdd gnd cell_6t
Xbit_r54_c26 bl_26 br_26 wl_54 vdd gnd cell_6t
Xbit_r55_c26 bl_26 br_26 wl_55 vdd gnd cell_6t
Xbit_r56_c26 bl_26 br_26 wl_56 vdd gnd cell_6t
Xbit_r57_c26 bl_26 br_26 wl_57 vdd gnd cell_6t
Xbit_r58_c26 bl_26 br_26 wl_58 vdd gnd cell_6t
Xbit_r59_c26 bl_26 br_26 wl_59 vdd gnd cell_6t
Xbit_r60_c26 bl_26 br_26 wl_60 vdd gnd cell_6t
Xbit_r61_c26 bl_26 br_26 wl_61 vdd gnd cell_6t
Xbit_r62_c26 bl_26 br_26 wl_62 vdd gnd cell_6t
Xbit_r63_c26 bl_26 br_26 wl_63 vdd gnd cell_6t
Xbit_r64_c26 bl_26 br_26 wl_64 vdd gnd cell_6t
Xbit_r65_c26 bl_26 br_26 wl_65 vdd gnd cell_6t
Xbit_r66_c26 bl_26 br_26 wl_66 vdd gnd cell_6t
Xbit_r67_c26 bl_26 br_26 wl_67 vdd gnd cell_6t
Xbit_r68_c26 bl_26 br_26 wl_68 vdd gnd cell_6t
Xbit_r69_c26 bl_26 br_26 wl_69 vdd gnd cell_6t
Xbit_r70_c26 bl_26 br_26 wl_70 vdd gnd cell_6t
Xbit_r71_c26 bl_26 br_26 wl_71 vdd gnd cell_6t
Xbit_r72_c26 bl_26 br_26 wl_72 vdd gnd cell_6t
Xbit_r73_c26 bl_26 br_26 wl_73 vdd gnd cell_6t
Xbit_r74_c26 bl_26 br_26 wl_74 vdd gnd cell_6t
Xbit_r75_c26 bl_26 br_26 wl_75 vdd gnd cell_6t
Xbit_r76_c26 bl_26 br_26 wl_76 vdd gnd cell_6t
Xbit_r77_c26 bl_26 br_26 wl_77 vdd gnd cell_6t
Xbit_r78_c26 bl_26 br_26 wl_78 vdd gnd cell_6t
Xbit_r79_c26 bl_26 br_26 wl_79 vdd gnd cell_6t
Xbit_r80_c26 bl_26 br_26 wl_80 vdd gnd cell_6t
Xbit_r81_c26 bl_26 br_26 wl_81 vdd gnd cell_6t
Xbit_r82_c26 bl_26 br_26 wl_82 vdd gnd cell_6t
Xbit_r83_c26 bl_26 br_26 wl_83 vdd gnd cell_6t
Xbit_r84_c26 bl_26 br_26 wl_84 vdd gnd cell_6t
Xbit_r85_c26 bl_26 br_26 wl_85 vdd gnd cell_6t
Xbit_r86_c26 bl_26 br_26 wl_86 vdd gnd cell_6t
Xbit_r87_c26 bl_26 br_26 wl_87 vdd gnd cell_6t
Xbit_r88_c26 bl_26 br_26 wl_88 vdd gnd cell_6t
Xbit_r89_c26 bl_26 br_26 wl_89 vdd gnd cell_6t
Xbit_r90_c26 bl_26 br_26 wl_90 vdd gnd cell_6t
Xbit_r91_c26 bl_26 br_26 wl_91 vdd gnd cell_6t
Xbit_r92_c26 bl_26 br_26 wl_92 vdd gnd cell_6t
Xbit_r93_c26 bl_26 br_26 wl_93 vdd gnd cell_6t
Xbit_r94_c26 bl_26 br_26 wl_94 vdd gnd cell_6t
Xbit_r95_c26 bl_26 br_26 wl_95 vdd gnd cell_6t
Xbit_r96_c26 bl_26 br_26 wl_96 vdd gnd cell_6t
Xbit_r97_c26 bl_26 br_26 wl_97 vdd gnd cell_6t
Xbit_r98_c26 bl_26 br_26 wl_98 vdd gnd cell_6t
Xbit_r99_c26 bl_26 br_26 wl_99 vdd gnd cell_6t
Xbit_r100_c26 bl_26 br_26 wl_100 vdd gnd cell_6t
Xbit_r101_c26 bl_26 br_26 wl_101 vdd gnd cell_6t
Xbit_r102_c26 bl_26 br_26 wl_102 vdd gnd cell_6t
Xbit_r103_c26 bl_26 br_26 wl_103 vdd gnd cell_6t
Xbit_r104_c26 bl_26 br_26 wl_104 vdd gnd cell_6t
Xbit_r105_c26 bl_26 br_26 wl_105 vdd gnd cell_6t
Xbit_r106_c26 bl_26 br_26 wl_106 vdd gnd cell_6t
Xbit_r107_c26 bl_26 br_26 wl_107 vdd gnd cell_6t
Xbit_r108_c26 bl_26 br_26 wl_108 vdd gnd cell_6t
Xbit_r109_c26 bl_26 br_26 wl_109 vdd gnd cell_6t
Xbit_r110_c26 bl_26 br_26 wl_110 vdd gnd cell_6t
Xbit_r111_c26 bl_26 br_26 wl_111 vdd gnd cell_6t
Xbit_r112_c26 bl_26 br_26 wl_112 vdd gnd cell_6t
Xbit_r113_c26 bl_26 br_26 wl_113 vdd gnd cell_6t
Xbit_r114_c26 bl_26 br_26 wl_114 vdd gnd cell_6t
Xbit_r115_c26 bl_26 br_26 wl_115 vdd gnd cell_6t
Xbit_r116_c26 bl_26 br_26 wl_116 vdd gnd cell_6t
Xbit_r117_c26 bl_26 br_26 wl_117 vdd gnd cell_6t
Xbit_r118_c26 bl_26 br_26 wl_118 vdd gnd cell_6t
Xbit_r119_c26 bl_26 br_26 wl_119 vdd gnd cell_6t
Xbit_r120_c26 bl_26 br_26 wl_120 vdd gnd cell_6t
Xbit_r121_c26 bl_26 br_26 wl_121 vdd gnd cell_6t
Xbit_r122_c26 bl_26 br_26 wl_122 vdd gnd cell_6t
Xbit_r123_c26 bl_26 br_26 wl_123 vdd gnd cell_6t
Xbit_r124_c26 bl_26 br_26 wl_124 vdd gnd cell_6t
Xbit_r125_c26 bl_26 br_26 wl_125 vdd gnd cell_6t
Xbit_r126_c26 bl_26 br_26 wl_126 vdd gnd cell_6t
Xbit_r127_c26 bl_26 br_26 wl_127 vdd gnd cell_6t
Xbit_r128_c26 bl_26 br_26 wl_128 vdd gnd cell_6t
Xbit_r129_c26 bl_26 br_26 wl_129 vdd gnd cell_6t
Xbit_r130_c26 bl_26 br_26 wl_130 vdd gnd cell_6t
Xbit_r131_c26 bl_26 br_26 wl_131 vdd gnd cell_6t
Xbit_r132_c26 bl_26 br_26 wl_132 vdd gnd cell_6t
Xbit_r133_c26 bl_26 br_26 wl_133 vdd gnd cell_6t
Xbit_r134_c26 bl_26 br_26 wl_134 vdd gnd cell_6t
Xbit_r135_c26 bl_26 br_26 wl_135 vdd gnd cell_6t
Xbit_r136_c26 bl_26 br_26 wl_136 vdd gnd cell_6t
Xbit_r137_c26 bl_26 br_26 wl_137 vdd gnd cell_6t
Xbit_r138_c26 bl_26 br_26 wl_138 vdd gnd cell_6t
Xbit_r139_c26 bl_26 br_26 wl_139 vdd gnd cell_6t
Xbit_r140_c26 bl_26 br_26 wl_140 vdd gnd cell_6t
Xbit_r141_c26 bl_26 br_26 wl_141 vdd gnd cell_6t
Xbit_r142_c26 bl_26 br_26 wl_142 vdd gnd cell_6t
Xbit_r143_c26 bl_26 br_26 wl_143 vdd gnd cell_6t
Xbit_r144_c26 bl_26 br_26 wl_144 vdd gnd cell_6t
Xbit_r145_c26 bl_26 br_26 wl_145 vdd gnd cell_6t
Xbit_r146_c26 bl_26 br_26 wl_146 vdd gnd cell_6t
Xbit_r147_c26 bl_26 br_26 wl_147 vdd gnd cell_6t
Xbit_r148_c26 bl_26 br_26 wl_148 vdd gnd cell_6t
Xbit_r149_c26 bl_26 br_26 wl_149 vdd gnd cell_6t
Xbit_r150_c26 bl_26 br_26 wl_150 vdd gnd cell_6t
Xbit_r151_c26 bl_26 br_26 wl_151 vdd gnd cell_6t
Xbit_r152_c26 bl_26 br_26 wl_152 vdd gnd cell_6t
Xbit_r153_c26 bl_26 br_26 wl_153 vdd gnd cell_6t
Xbit_r154_c26 bl_26 br_26 wl_154 vdd gnd cell_6t
Xbit_r155_c26 bl_26 br_26 wl_155 vdd gnd cell_6t
Xbit_r156_c26 bl_26 br_26 wl_156 vdd gnd cell_6t
Xbit_r157_c26 bl_26 br_26 wl_157 vdd gnd cell_6t
Xbit_r158_c26 bl_26 br_26 wl_158 vdd gnd cell_6t
Xbit_r159_c26 bl_26 br_26 wl_159 vdd gnd cell_6t
Xbit_r160_c26 bl_26 br_26 wl_160 vdd gnd cell_6t
Xbit_r161_c26 bl_26 br_26 wl_161 vdd gnd cell_6t
Xbit_r162_c26 bl_26 br_26 wl_162 vdd gnd cell_6t
Xbit_r163_c26 bl_26 br_26 wl_163 vdd gnd cell_6t
Xbit_r164_c26 bl_26 br_26 wl_164 vdd gnd cell_6t
Xbit_r165_c26 bl_26 br_26 wl_165 vdd gnd cell_6t
Xbit_r166_c26 bl_26 br_26 wl_166 vdd gnd cell_6t
Xbit_r167_c26 bl_26 br_26 wl_167 vdd gnd cell_6t
Xbit_r168_c26 bl_26 br_26 wl_168 vdd gnd cell_6t
Xbit_r169_c26 bl_26 br_26 wl_169 vdd gnd cell_6t
Xbit_r170_c26 bl_26 br_26 wl_170 vdd gnd cell_6t
Xbit_r171_c26 bl_26 br_26 wl_171 vdd gnd cell_6t
Xbit_r172_c26 bl_26 br_26 wl_172 vdd gnd cell_6t
Xbit_r173_c26 bl_26 br_26 wl_173 vdd gnd cell_6t
Xbit_r174_c26 bl_26 br_26 wl_174 vdd gnd cell_6t
Xbit_r175_c26 bl_26 br_26 wl_175 vdd gnd cell_6t
Xbit_r176_c26 bl_26 br_26 wl_176 vdd gnd cell_6t
Xbit_r177_c26 bl_26 br_26 wl_177 vdd gnd cell_6t
Xbit_r178_c26 bl_26 br_26 wl_178 vdd gnd cell_6t
Xbit_r179_c26 bl_26 br_26 wl_179 vdd gnd cell_6t
Xbit_r180_c26 bl_26 br_26 wl_180 vdd gnd cell_6t
Xbit_r181_c26 bl_26 br_26 wl_181 vdd gnd cell_6t
Xbit_r182_c26 bl_26 br_26 wl_182 vdd gnd cell_6t
Xbit_r183_c26 bl_26 br_26 wl_183 vdd gnd cell_6t
Xbit_r184_c26 bl_26 br_26 wl_184 vdd gnd cell_6t
Xbit_r185_c26 bl_26 br_26 wl_185 vdd gnd cell_6t
Xbit_r186_c26 bl_26 br_26 wl_186 vdd gnd cell_6t
Xbit_r187_c26 bl_26 br_26 wl_187 vdd gnd cell_6t
Xbit_r188_c26 bl_26 br_26 wl_188 vdd gnd cell_6t
Xbit_r189_c26 bl_26 br_26 wl_189 vdd gnd cell_6t
Xbit_r190_c26 bl_26 br_26 wl_190 vdd gnd cell_6t
Xbit_r191_c26 bl_26 br_26 wl_191 vdd gnd cell_6t
Xbit_r192_c26 bl_26 br_26 wl_192 vdd gnd cell_6t
Xbit_r193_c26 bl_26 br_26 wl_193 vdd gnd cell_6t
Xbit_r194_c26 bl_26 br_26 wl_194 vdd gnd cell_6t
Xbit_r195_c26 bl_26 br_26 wl_195 vdd gnd cell_6t
Xbit_r196_c26 bl_26 br_26 wl_196 vdd gnd cell_6t
Xbit_r197_c26 bl_26 br_26 wl_197 vdd gnd cell_6t
Xbit_r198_c26 bl_26 br_26 wl_198 vdd gnd cell_6t
Xbit_r199_c26 bl_26 br_26 wl_199 vdd gnd cell_6t
Xbit_r200_c26 bl_26 br_26 wl_200 vdd gnd cell_6t
Xbit_r201_c26 bl_26 br_26 wl_201 vdd gnd cell_6t
Xbit_r202_c26 bl_26 br_26 wl_202 vdd gnd cell_6t
Xbit_r203_c26 bl_26 br_26 wl_203 vdd gnd cell_6t
Xbit_r204_c26 bl_26 br_26 wl_204 vdd gnd cell_6t
Xbit_r205_c26 bl_26 br_26 wl_205 vdd gnd cell_6t
Xbit_r206_c26 bl_26 br_26 wl_206 vdd gnd cell_6t
Xbit_r207_c26 bl_26 br_26 wl_207 vdd gnd cell_6t
Xbit_r208_c26 bl_26 br_26 wl_208 vdd gnd cell_6t
Xbit_r209_c26 bl_26 br_26 wl_209 vdd gnd cell_6t
Xbit_r210_c26 bl_26 br_26 wl_210 vdd gnd cell_6t
Xbit_r211_c26 bl_26 br_26 wl_211 vdd gnd cell_6t
Xbit_r212_c26 bl_26 br_26 wl_212 vdd gnd cell_6t
Xbit_r213_c26 bl_26 br_26 wl_213 vdd gnd cell_6t
Xbit_r214_c26 bl_26 br_26 wl_214 vdd gnd cell_6t
Xbit_r215_c26 bl_26 br_26 wl_215 vdd gnd cell_6t
Xbit_r216_c26 bl_26 br_26 wl_216 vdd gnd cell_6t
Xbit_r217_c26 bl_26 br_26 wl_217 vdd gnd cell_6t
Xbit_r218_c26 bl_26 br_26 wl_218 vdd gnd cell_6t
Xbit_r219_c26 bl_26 br_26 wl_219 vdd gnd cell_6t
Xbit_r220_c26 bl_26 br_26 wl_220 vdd gnd cell_6t
Xbit_r221_c26 bl_26 br_26 wl_221 vdd gnd cell_6t
Xbit_r222_c26 bl_26 br_26 wl_222 vdd gnd cell_6t
Xbit_r223_c26 bl_26 br_26 wl_223 vdd gnd cell_6t
Xbit_r224_c26 bl_26 br_26 wl_224 vdd gnd cell_6t
Xbit_r225_c26 bl_26 br_26 wl_225 vdd gnd cell_6t
Xbit_r226_c26 bl_26 br_26 wl_226 vdd gnd cell_6t
Xbit_r227_c26 bl_26 br_26 wl_227 vdd gnd cell_6t
Xbit_r228_c26 bl_26 br_26 wl_228 vdd gnd cell_6t
Xbit_r229_c26 bl_26 br_26 wl_229 vdd gnd cell_6t
Xbit_r230_c26 bl_26 br_26 wl_230 vdd gnd cell_6t
Xbit_r231_c26 bl_26 br_26 wl_231 vdd gnd cell_6t
Xbit_r232_c26 bl_26 br_26 wl_232 vdd gnd cell_6t
Xbit_r233_c26 bl_26 br_26 wl_233 vdd gnd cell_6t
Xbit_r234_c26 bl_26 br_26 wl_234 vdd gnd cell_6t
Xbit_r235_c26 bl_26 br_26 wl_235 vdd gnd cell_6t
Xbit_r236_c26 bl_26 br_26 wl_236 vdd gnd cell_6t
Xbit_r237_c26 bl_26 br_26 wl_237 vdd gnd cell_6t
Xbit_r238_c26 bl_26 br_26 wl_238 vdd gnd cell_6t
Xbit_r239_c26 bl_26 br_26 wl_239 vdd gnd cell_6t
Xbit_r240_c26 bl_26 br_26 wl_240 vdd gnd cell_6t
Xbit_r241_c26 bl_26 br_26 wl_241 vdd gnd cell_6t
Xbit_r242_c26 bl_26 br_26 wl_242 vdd gnd cell_6t
Xbit_r243_c26 bl_26 br_26 wl_243 vdd gnd cell_6t
Xbit_r244_c26 bl_26 br_26 wl_244 vdd gnd cell_6t
Xbit_r245_c26 bl_26 br_26 wl_245 vdd gnd cell_6t
Xbit_r246_c26 bl_26 br_26 wl_246 vdd gnd cell_6t
Xbit_r247_c26 bl_26 br_26 wl_247 vdd gnd cell_6t
Xbit_r248_c26 bl_26 br_26 wl_248 vdd gnd cell_6t
Xbit_r249_c26 bl_26 br_26 wl_249 vdd gnd cell_6t
Xbit_r250_c26 bl_26 br_26 wl_250 vdd gnd cell_6t
Xbit_r251_c26 bl_26 br_26 wl_251 vdd gnd cell_6t
Xbit_r252_c26 bl_26 br_26 wl_252 vdd gnd cell_6t
Xbit_r253_c26 bl_26 br_26 wl_253 vdd gnd cell_6t
Xbit_r254_c26 bl_26 br_26 wl_254 vdd gnd cell_6t
Xbit_r255_c26 bl_26 br_26 wl_255 vdd gnd cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd cell_6t
Xbit_r1_c27 bl_27 br_27 wl_1 vdd gnd cell_6t
Xbit_r2_c27 bl_27 br_27 wl_2 vdd gnd cell_6t
Xbit_r3_c27 bl_27 br_27 wl_3 vdd gnd cell_6t
Xbit_r4_c27 bl_27 br_27 wl_4 vdd gnd cell_6t
Xbit_r5_c27 bl_27 br_27 wl_5 vdd gnd cell_6t
Xbit_r6_c27 bl_27 br_27 wl_6 vdd gnd cell_6t
Xbit_r7_c27 bl_27 br_27 wl_7 vdd gnd cell_6t
Xbit_r8_c27 bl_27 br_27 wl_8 vdd gnd cell_6t
Xbit_r9_c27 bl_27 br_27 wl_9 vdd gnd cell_6t
Xbit_r10_c27 bl_27 br_27 wl_10 vdd gnd cell_6t
Xbit_r11_c27 bl_27 br_27 wl_11 vdd gnd cell_6t
Xbit_r12_c27 bl_27 br_27 wl_12 vdd gnd cell_6t
Xbit_r13_c27 bl_27 br_27 wl_13 vdd gnd cell_6t
Xbit_r14_c27 bl_27 br_27 wl_14 vdd gnd cell_6t
Xbit_r15_c27 bl_27 br_27 wl_15 vdd gnd cell_6t
Xbit_r16_c27 bl_27 br_27 wl_16 vdd gnd cell_6t
Xbit_r17_c27 bl_27 br_27 wl_17 vdd gnd cell_6t
Xbit_r18_c27 bl_27 br_27 wl_18 vdd gnd cell_6t
Xbit_r19_c27 bl_27 br_27 wl_19 vdd gnd cell_6t
Xbit_r20_c27 bl_27 br_27 wl_20 vdd gnd cell_6t
Xbit_r21_c27 bl_27 br_27 wl_21 vdd gnd cell_6t
Xbit_r22_c27 bl_27 br_27 wl_22 vdd gnd cell_6t
Xbit_r23_c27 bl_27 br_27 wl_23 vdd gnd cell_6t
Xbit_r24_c27 bl_27 br_27 wl_24 vdd gnd cell_6t
Xbit_r25_c27 bl_27 br_27 wl_25 vdd gnd cell_6t
Xbit_r26_c27 bl_27 br_27 wl_26 vdd gnd cell_6t
Xbit_r27_c27 bl_27 br_27 wl_27 vdd gnd cell_6t
Xbit_r28_c27 bl_27 br_27 wl_28 vdd gnd cell_6t
Xbit_r29_c27 bl_27 br_27 wl_29 vdd gnd cell_6t
Xbit_r30_c27 bl_27 br_27 wl_30 vdd gnd cell_6t
Xbit_r31_c27 bl_27 br_27 wl_31 vdd gnd cell_6t
Xbit_r32_c27 bl_27 br_27 wl_32 vdd gnd cell_6t
Xbit_r33_c27 bl_27 br_27 wl_33 vdd gnd cell_6t
Xbit_r34_c27 bl_27 br_27 wl_34 vdd gnd cell_6t
Xbit_r35_c27 bl_27 br_27 wl_35 vdd gnd cell_6t
Xbit_r36_c27 bl_27 br_27 wl_36 vdd gnd cell_6t
Xbit_r37_c27 bl_27 br_27 wl_37 vdd gnd cell_6t
Xbit_r38_c27 bl_27 br_27 wl_38 vdd gnd cell_6t
Xbit_r39_c27 bl_27 br_27 wl_39 vdd gnd cell_6t
Xbit_r40_c27 bl_27 br_27 wl_40 vdd gnd cell_6t
Xbit_r41_c27 bl_27 br_27 wl_41 vdd gnd cell_6t
Xbit_r42_c27 bl_27 br_27 wl_42 vdd gnd cell_6t
Xbit_r43_c27 bl_27 br_27 wl_43 vdd gnd cell_6t
Xbit_r44_c27 bl_27 br_27 wl_44 vdd gnd cell_6t
Xbit_r45_c27 bl_27 br_27 wl_45 vdd gnd cell_6t
Xbit_r46_c27 bl_27 br_27 wl_46 vdd gnd cell_6t
Xbit_r47_c27 bl_27 br_27 wl_47 vdd gnd cell_6t
Xbit_r48_c27 bl_27 br_27 wl_48 vdd gnd cell_6t
Xbit_r49_c27 bl_27 br_27 wl_49 vdd gnd cell_6t
Xbit_r50_c27 bl_27 br_27 wl_50 vdd gnd cell_6t
Xbit_r51_c27 bl_27 br_27 wl_51 vdd gnd cell_6t
Xbit_r52_c27 bl_27 br_27 wl_52 vdd gnd cell_6t
Xbit_r53_c27 bl_27 br_27 wl_53 vdd gnd cell_6t
Xbit_r54_c27 bl_27 br_27 wl_54 vdd gnd cell_6t
Xbit_r55_c27 bl_27 br_27 wl_55 vdd gnd cell_6t
Xbit_r56_c27 bl_27 br_27 wl_56 vdd gnd cell_6t
Xbit_r57_c27 bl_27 br_27 wl_57 vdd gnd cell_6t
Xbit_r58_c27 bl_27 br_27 wl_58 vdd gnd cell_6t
Xbit_r59_c27 bl_27 br_27 wl_59 vdd gnd cell_6t
Xbit_r60_c27 bl_27 br_27 wl_60 vdd gnd cell_6t
Xbit_r61_c27 bl_27 br_27 wl_61 vdd gnd cell_6t
Xbit_r62_c27 bl_27 br_27 wl_62 vdd gnd cell_6t
Xbit_r63_c27 bl_27 br_27 wl_63 vdd gnd cell_6t
Xbit_r64_c27 bl_27 br_27 wl_64 vdd gnd cell_6t
Xbit_r65_c27 bl_27 br_27 wl_65 vdd gnd cell_6t
Xbit_r66_c27 bl_27 br_27 wl_66 vdd gnd cell_6t
Xbit_r67_c27 bl_27 br_27 wl_67 vdd gnd cell_6t
Xbit_r68_c27 bl_27 br_27 wl_68 vdd gnd cell_6t
Xbit_r69_c27 bl_27 br_27 wl_69 vdd gnd cell_6t
Xbit_r70_c27 bl_27 br_27 wl_70 vdd gnd cell_6t
Xbit_r71_c27 bl_27 br_27 wl_71 vdd gnd cell_6t
Xbit_r72_c27 bl_27 br_27 wl_72 vdd gnd cell_6t
Xbit_r73_c27 bl_27 br_27 wl_73 vdd gnd cell_6t
Xbit_r74_c27 bl_27 br_27 wl_74 vdd gnd cell_6t
Xbit_r75_c27 bl_27 br_27 wl_75 vdd gnd cell_6t
Xbit_r76_c27 bl_27 br_27 wl_76 vdd gnd cell_6t
Xbit_r77_c27 bl_27 br_27 wl_77 vdd gnd cell_6t
Xbit_r78_c27 bl_27 br_27 wl_78 vdd gnd cell_6t
Xbit_r79_c27 bl_27 br_27 wl_79 vdd gnd cell_6t
Xbit_r80_c27 bl_27 br_27 wl_80 vdd gnd cell_6t
Xbit_r81_c27 bl_27 br_27 wl_81 vdd gnd cell_6t
Xbit_r82_c27 bl_27 br_27 wl_82 vdd gnd cell_6t
Xbit_r83_c27 bl_27 br_27 wl_83 vdd gnd cell_6t
Xbit_r84_c27 bl_27 br_27 wl_84 vdd gnd cell_6t
Xbit_r85_c27 bl_27 br_27 wl_85 vdd gnd cell_6t
Xbit_r86_c27 bl_27 br_27 wl_86 vdd gnd cell_6t
Xbit_r87_c27 bl_27 br_27 wl_87 vdd gnd cell_6t
Xbit_r88_c27 bl_27 br_27 wl_88 vdd gnd cell_6t
Xbit_r89_c27 bl_27 br_27 wl_89 vdd gnd cell_6t
Xbit_r90_c27 bl_27 br_27 wl_90 vdd gnd cell_6t
Xbit_r91_c27 bl_27 br_27 wl_91 vdd gnd cell_6t
Xbit_r92_c27 bl_27 br_27 wl_92 vdd gnd cell_6t
Xbit_r93_c27 bl_27 br_27 wl_93 vdd gnd cell_6t
Xbit_r94_c27 bl_27 br_27 wl_94 vdd gnd cell_6t
Xbit_r95_c27 bl_27 br_27 wl_95 vdd gnd cell_6t
Xbit_r96_c27 bl_27 br_27 wl_96 vdd gnd cell_6t
Xbit_r97_c27 bl_27 br_27 wl_97 vdd gnd cell_6t
Xbit_r98_c27 bl_27 br_27 wl_98 vdd gnd cell_6t
Xbit_r99_c27 bl_27 br_27 wl_99 vdd gnd cell_6t
Xbit_r100_c27 bl_27 br_27 wl_100 vdd gnd cell_6t
Xbit_r101_c27 bl_27 br_27 wl_101 vdd gnd cell_6t
Xbit_r102_c27 bl_27 br_27 wl_102 vdd gnd cell_6t
Xbit_r103_c27 bl_27 br_27 wl_103 vdd gnd cell_6t
Xbit_r104_c27 bl_27 br_27 wl_104 vdd gnd cell_6t
Xbit_r105_c27 bl_27 br_27 wl_105 vdd gnd cell_6t
Xbit_r106_c27 bl_27 br_27 wl_106 vdd gnd cell_6t
Xbit_r107_c27 bl_27 br_27 wl_107 vdd gnd cell_6t
Xbit_r108_c27 bl_27 br_27 wl_108 vdd gnd cell_6t
Xbit_r109_c27 bl_27 br_27 wl_109 vdd gnd cell_6t
Xbit_r110_c27 bl_27 br_27 wl_110 vdd gnd cell_6t
Xbit_r111_c27 bl_27 br_27 wl_111 vdd gnd cell_6t
Xbit_r112_c27 bl_27 br_27 wl_112 vdd gnd cell_6t
Xbit_r113_c27 bl_27 br_27 wl_113 vdd gnd cell_6t
Xbit_r114_c27 bl_27 br_27 wl_114 vdd gnd cell_6t
Xbit_r115_c27 bl_27 br_27 wl_115 vdd gnd cell_6t
Xbit_r116_c27 bl_27 br_27 wl_116 vdd gnd cell_6t
Xbit_r117_c27 bl_27 br_27 wl_117 vdd gnd cell_6t
Xbit_r118_c27 bl_27 br_27 wl_118 vdd gnd cell_6t
Xbit_r119_c27 bl_27 br_27 wl_119 vdd gnd cell_6t
Xbit_r120_c27 bl_27 br_27 wl_120 vdd gnd cell_6t
Xbit_r121_c27 bl_27 br_27 wl_121 vdd gnd cell_6t
Xbit_r122_c27 bl_27 br_27 wl_122 vdd gnd cell_6t
Xbit_r123_c27 bl_27 br_27 wl_123 vdd gnd cell_6t
Xbit_r124_c27 bl_27 br_27 wl_124 vdd gnd cell_6t
Xbit_r125_c27 bl_27 br_27 wl_125 vdd gnd cell_6t
Xbit_r126_c27 bl_27 br_27 wl_126 vdd gnd cell_6t
Xbit_r127_c27 bl_27 br_27 wl_127 vdd gnd cell_6t
Xbit_r128_c27 bl_27 br_27 wl_128 vdd gnd cell_6t
Xbit_r129_c27 bl_27 br_27 wl_129 vdd gnd cell_6t
Xbit_r130_c27 bl_27 br_27 wl_130 vdd gnd cell_6t
Xbit_r131_c27 bl_27 br_27 wl_131 vdd gnd cell_6t
Xbit_r132_c27 bl_27 br_27 wl_132 vdd gnd cell_6t
Xbit_r133_c27 bl_27 br_27 wl_133 vdd gnd cell_6t
Xbit_r134_c27 bl_27 br_27 wl_134 vdd gnd cell_6t
Xbit_r135_c27 bl_27 br_27 wl_135 vdd gnd cell_6t
Xbit_r136_c27 bl_27 br_27 wl_136 vdd gnd cell_6t
Xbit_r137_c27 bl_27 br_27 wl_137 vdd gnd cell_6t
Xbit_r138_c27 bl_27 br_27 wl_138 vdd gnd cell_6t
Xbit_r139_c27 bl_27 br_27 wl_139 vdd gnd cell_6t
Xbit_r140_c27 bl_27 br_27 wl_140 vdd gnd cell_6t
Xbit_r141_c27 bl_27 br_27 wl_141 vdd gnd cell_6t
Xbit_r142_c27 bl_27 br_27 wl_142 vdd gnd cell_6t
Xbit_r143_c27 bl_27 br_27 wl_143 vdd gnd cell_6t
Xbit_r144_c27 bl_27 br_27 wl_144 vdd gnd cell_6t
Xbit_r145_c27 bl_27 br_27 wl_145 vdd gnd cell_6t
Xbit_r146_c27 bl_27 br_27 wl_146 vdd gnd cell_6t
Xbit_r147_c27 bl_27 br_27 wl_147 vdd gnd cell_6t
Xbit_r148_c27 bl_27 br_27 wl_148 vdd gnd cell_6t
Xbit_r149_c27 bl_27 br_27 wl_149 vdd gnd cell_6t
Xbit_r150_c27 bl_27 br_27 wl_150 vdd gnd cell_6t
Xbit_r151_c27 bl_27 br_27 wl_151 vdd gnd cell_6t
Xbit_r152_c27 bl_27 br_27 wl_152 vdd gnd cell_6t
Xbit_r153_c27 bl_27 br_27 wl_153 vdd gnd cell_6t
Xbit_r154_c27 bl_27 br_27 wl_154 vdd gnd cell_6t
Xbit_r155_c27 bl_27 br_27 wl_155 vdd gnd cell_6t
Xbit_r156_c27 bl_27 br_27 wl_156 vdd gnd cell_6t
Xbit_r157_c27 bl_27 br_27 wl_157 vdd gnd cell_6t
Xbit_r158_c27 bl_27 br_27 wl_158 vdd gnd cell_6t
Xbit_r159_c27 bl_27 br_27 wl_159 vdd gnd cell_6t
Xbit_r160_c27 bl_27 br_27 wl_160 vdd gnd cell_6t
Xbit_r161_c27 bl_27 br_27 wl_161 vdd gnd cell_6t
Xbit_r162_c27 bl_27 br_27 wl_162 vdd gnd cell_6t
Xbit_r163_c27 bl_27 br_27 wl_163 vdd gnd cell_6t
Xbit_r164_c27 bl_27 br_27 wl_164 vdd gnd cell_6t
Xbit_r165_c27 bl_27 br_27 wl_165 vdd gnd cell_6t
Xbit_r166_c27 bl_27 br_27 wl_166 vdd gnd cell_6t
Xbit_r167_c27 bl_27 br_27 wl_167 vdd gnd cell_6t
Xbit_r168_c27 bl_27 br_27 wl_168 vdd gnd cell_6t
Xbit_r169_c27 bl_27 br_27 wl_169 vdd gnd cell_6t
Xbit_r170_c27 bl_27 br_27 wl_170 vdd gnd cell_6t
Xbit_r171_c27 bl_27 br_27 wl_171 vdd gnd cell_6t
Xbit_r172_c27 bl_27 br_27 wl_172 vdd gnd cell_6t
Xbit_r173_c27 bl_27 br_27 wl_173 vdd gnd cell_6t
Xbit_r174_c27 bl_27 br_27 wl_174 vdd gnd cell_6t
Xbit_r175_c27 bl_27 br_27 wl_175 vdd gnd cell_6t
Xbit_r176_c27 bl_27 br_27 wl_176 vdd gnd cell_6t
Xbit_r177_c27 bl_27 br_27 wl_177 vdd gnd cell_6t
Xbit_r178_c27 bl_27 br_27 wl_178 vdd gnd cell_6t
Xbit_r179_c27 bl_27 br_27 wl_179 vdd gnd cell_6t
Xbit_r180_c27 bl_27 br_27 wl_180 vdd gnd cell_6t
Xbit_r181_c27 bl_27 br_27 wl_181 vdd gnd cell_6t
Xbit_r182_c27 bl_27 br_27 wl_182 vdd gnd cell_6t
Xbit_r183_c27 bl_27 br_27 wl_183 vdd gnd cell_6t
Xbit_r184_c27 bl_27 br_27 wl_184 vdd gnd cell_6t
Xbit_r185_c27 bl_27 br_27 wl_185 vdd gnd cell_6t
Xbit_r186_c27 bl_27 br_27 wl_186 vdd gnd cell_6t
Xbit_r187_c27 bl_27 br_27 wl_187 vdd gnd cell_6t
Xbit_r188_c27 bl_27 br_27 wl_188 vdd gnd cell_6t
Xbit_r189_c27 bl_27 br_27 wl_189 vdd gnd cell_6t
Xbit_r190_c27 bl_27 br_27 wl_190 vdd gnd cell_6t
Xbit_r191_c27 bl_27 br_27 wl_191 vdd gnd cell_6t
Xbit_r192_c27 bl_27 br_27 wl_192 vdd gnd cell_6t
Xbit_r193_c27 bl_27 br_27 wl_193 vdd gnd cell_6t
Xbit_r194_c27 bl_27 br_27 wl_194 vdd gnd cell_6t
Xbit_r195_c27 bl_27 br_27 wl_195 vdd gnd cell_6t
Xbit_r196_c27 bl_27 br_27 wl_196 vdd gnd cell_6t
Xbit_r197_c27 bl_27 br_27 wl_197 vdd gnd cell_6t
Xbit_r198_c27 bl_27 br_27 wl_198 vdd gnd cell_6t
Xbit_r199_c27 bl_27 br_27 wl_199 vdd gnd cell_6t
Xbit_r200_c27 bl_27 br_27 wl_200 vdd gnd cell_6t
Xbit_r201_c27 bl_27 br_27 wl_201 vdd gnd cell_6t
Xbit_r202_c27 bl_27 br_27 wl_202 vdd gnd cell_6t
Xbit_r203_c27 bl_27 br_27 wl_203 vdd gnd cell_6t
Xbit_r204_c27 bl_27 br_27 wl_204 vdd gnd cell_6t
Xbit_r205_c27 bl_27 br_27 wl_205 vdd gnd cell_6t
Xbit_r206_c27 bl_27 br_27 wl_206 vdd gnd cell_6t
Xbit_r207_c27 bl_27 br_27 wl_207 vdd gnd cell_6t
Xbit_r208_c27 bl_27 br_27 wl_208 vdd gnd cell_6t
Xbit_r209_c27 bl_27 br_27 wl_209 vdd gnd cell_6t
Xbit_r210_c27 bl_27 br_27 wl_210 vdd gnd cell_6t
Xbit_r211_c27 bl_27 br_27 wl_211 vdd gnd cell_6t
Xbit_r212_c27 bl_27 br_27 wl_212 vdd gnd cell_6t
Xbit_r213_c27 bl_27 br_27 wl_213 vdd gnd cell_6t
Xbit_r214_c27 bl_27 br_27 wl_214 vdd gnd cell_6t
Xbit_r215_c27 bl_27 br_27 wl_215 vdd gnd cell_6t
Xbit_r216_c27 bl_27 br_27 wl_216 vdd gnd cell_6t
Xbit_r217_c27 bl_27 br_27 wl_217 vdd gnd cell_6t
Xbit_r218_c27 bl_27 br_27 wl_218 vdd gnd cell_6t
Xbit_r219_c27 bl_27 br_27 wl_219 vdd gnd cell_6t
Xbit_r220_c27 bl_27 br_27 wl_220 vdd gnd cell_6t
Xbit_r221_c27 bl_27 br_27 wl_221 vdd gnd cell_6t
Xbit_r222_c27 bl_27 br_27 wl_222 vdd gnd cell_6t
Xbit_r223_c27 bl_27 br_27 wl_223 vdd gnd cell_6t
Xbit_r224_c27 bl_27 br_27 wl_224 vdd gnd cell_6t
Xbit_r225_c27 bl_27 br_27 wl_225 vdd gnd cell_6t
Xbit_r226_c27 bl_27 br_27 wl_226 vdd gnd cell_6t
Xbit_r227_c27 bl_27 br_27 wl_227 vdd gnd cell_6t
Xbit_r228_c27 bl_27 br_27 wl_228 vdd gnd cell_6t
Xbit_r229_c27 bl_27 br_27 wl_229 vdd gnd cell_6t
Xbit_r230_c27 bl_27 br_27 wl_230 vdd gnd cell_6t
Xbit_r231_c27 bl_27 br_27 wl_231 vdd gnd cell_6t
Xbit_r232_c27 bl_27 br_27 wl_232 vdd gnd cell_6t
Xbit_r233_c27 bl_27 br_27 wl_233 vdd gnd cell_6t
Xbit_r234_c27 bl_27 br_27 wl_234 vdd gnd cell_6t
Xbit_r235_c27 bl_27 br_27 wl_235 vdd gnd cell_6t
Xbit_r236_c27 bl_27 br_27 wl_236 vdd gnd cell_6t
Xbit_r237_c27 bl_27 br_27 wl_237 vdd gnd cell_6t
Xbit_r238_c27 bl_27 br_27 wl_238 vdd gnd cell_6t
Xbit_r239_c27 bl_27 br_27 wl_239 vdd gnd cell_6t
Xbit_r240_c27 bl_27 br_27 wl_240 vdd gnd cell_6t
Xbit_r241_c27 bl_27 br_27 wl_241 vdd gnd cell_6t
Xbit_r242_c27 bl_27 br_27 wl_242 vdd gnd cell_6t
Xbit_r243_c27 bl_27 br_27 wl_243 vdd gnd cell_6t
Xbit_r244_c27 bl_27 br_27 wl_244 vdd gnd cell_6t
Xbit_r245_c27 bl_27 br_27 wl_245 vdd gnd cell_6t
Xbit_r246_c27 bl_27 br_27 wl_246 vdd gnd cell_6t
Xbit_r247_c27 bl_27 br_27 wl_247 vdd gnd cell_6t
Xbit_r248_c27 bl_27 br_27 wl_248 vdd gnd cell_6t
Xbit_r249_c27 bl_27 br_27 wl_249 vdd gnd cell_6t
Xbit_r250_c27 bl_27 br_27 wl_250 vdd gnd cell_6t
Xbit_r251_c27 bl_27 br_27 wl_251 vdd gnd cell_6t
Xbit_r252_c27 bl_27 br_27 wl_252 vdd gnd cell_6t
Xbit_r253_c27 bl_27 br_27 wl_253 vdd gnd cell_6t
Xbit_r254_c27 bl_27 br_27 wl_254 vdd gnd cell_6t
Xbit_r255_c27 bl_27 br_27 wl_255 vdd gnd cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd cell_6t
Xbit_r1_c28 bl_28 br_28 wl_1 vdd gnd cell_6t
Xbit_r2_c28 bl_28 br_28 wl_2 vdd gnd cell_6t
Xbit_r3_c28 bl_28 br_28 wl_3 vdd gnd cell_6t
Xbit_r4_c28 bl_28 br_28 wl_4 vdd gnd cell_6t
Xbit_r5_c28 bl_28 br_28 wl_5 vdd gnd cell_6t
Xbit_r6_c28 bl_28 br_28 wl_6 vdd gnd cell_6t
Xbit_r7_c28 bl_28 br_28 wl_7 vdd gnd cell_6t
Xbit_r8_c28 bl_28 br_28 wl_8 vdd gnd cell_6t
Xbit_r9_c28 bl_28 br_28 wl_9 vdd gnd cell_6t
Xbit_r10_c28 bl_28 br_28 wl_10 vdd gnd cell_6t
Xbit_r11_c28 bl_28 br_28 wl_11 vdd gnd cell_6t
Xbit_r12_c28 bl_28 br_28 wl_12 vdd gnd cell_6t
Xbit_r13_c28 bl_28 br_28 wl_13 vdd gnd cell_6t
Xbit_r14_c28 bl_28 br_28 wl_14 vdd gnd cell_6t
Xbit_r15_c28 bl_28 br_28 wl_15 vdd gnd cell_6t
Xbit_r16_c28 bl_28 br_28 wl_16 vdd gnd cell_6t
Xbit_r17_c28 bl_28 br_28 wl_17 vdd gnd cell_6t
Xbit_r18_c28 bl_28 br_28 wl_18 vdd gnd cell_6t
Xbit_r19_c28 bl_28 br_28 wl_19 vdd gnd cell_6t
Xbit_r20_c28 bl_28 br_28 wl_20 vdd gnd cell_6t
Xbit_r21_c28 bl_28 br_28 wl_21 vdd gnd cell_6t
Xbit_r22_c28 bl_28 br_28 wl_22 vdd gnd cell_6t
Xbit_r23_c28 bl_28 br_28 wl_23 vdd gnd cell_6t
Xbit_r24_c28 bl_28 br_28 wl_24 vdd gnd cell_6t
Xbit_r25_c28 bl_28 br_28 wl_25 vdd gnd cell_6t
Xbit_r26_c28 bl_28 br_28 wl_26 vdd gnd cell_6t
Xbit_r27_c28 bl_28 br_28 wl_27 vdd gnd cell_6t
Xbit_r28_c28 bl_28 br_28 wl_28 vdd gnd cell_6t
Xbit_r29_c28 bl_28 br_28 wl_29 vdd gnd cell_6t
Xbit_r30_c28 bl_28 br_28 wl_30 vdd gnd cell_6t
Xbit_r31_c28 bl_28 br_28 wl_31 vdd gnd cell_6t
Xbit_r32_c28 bl_28 br_28 wl_32 vdd gnd cell_6t
Xbit_r33_c28 bl_28 br_28 wl_33 vdd gnd cell_6t
Xbit_r34_c28 bl_28 br_28 wl_34 vdd gnd cell_6t
Xbit_r35_c28 bl_28 br_28 wl_35 vdd gnd cell_6t
Xbit_r36_c28 bl_28 br_28 wl_36 vdd gnd cell_6t
Xbit_r37_c28 bl_28 br_28 wl_37 vdd gnd cell_6t
Xbit_r38_c28 bl_28 br_28 wl_38 vdd gnd cell_6t
Xbit_r39_c28 bl_28 br_28 wl_39 vdd gnd cell_6t
Xbit_r40_c28 bl_28 br_28 wl_40 vdd gnd cell_6t
Xbit_r41_c28 bl_28 br_28 wl_41 vdd gnd cell_6t
Xbit_r42_c28 bl_28 br_28 wl_42 vdd gnd cell_6t
Xbit_r43_c28 bl_28 br_28 wl_43 vdd gnd cell_6t
Xbit_r44_c28 bl_28 br_28 wl_44 vdd gnd cell_6t
Xbit_r45_c28 bl_28 br_28 wl_45 vdd gnd cell_6t
Xbit_r46_c28 bl_28 br_28 wl_46 vdd gnd cell_6t
Xbit_r47_c28 bl_28 br_28 wl_47 vdd gnd cell_6t
Xbit_r48_c28 bl_28 br_28 wl_48 vdd gnd cell_6t
Xbit_r49_c28 bl_28 br_28 wl_49 vdd gnd cell_6t
Xbit_r50_c28 bl_28 br_28 wl_50 vdd gnd cell_6t
Xbit_r51_c28 bl_28 br_28 wl_51 vdd gnd cell_6t
Xbit_r52_c28 bl_28 br_28 wl_52 vdd gnd cell_6t
Xbit_r53_c28 bl_28 br_28 wl_53 vdd gnd cell_6t
Xbit_r54_c28 bl_28 br_28 wl_54 vdd gnd cell_6t
Xbit_r55_c28 bl_28 br_28 wl_55 vdd gnd cell_6t
Xbit_r56_c28 bl_28 br_28 wl_56 vdd gnd cell_6t
Xbit_r57_c28 bl_28 br_28 wl_57 vdd gnd cell_6t
Xbit_r58_c28 bl_28 br_28 wl_58 vdd gnd cell_6t
Xbit_r59_c28 bl_28 br_28 wl_59 vdd gnd cell_6t
Xbit_r60_c28 bl_28 br_28 wl_60 vdd gnd cell_6t
Xbit_r61_c28 bl_28 br_28 wl_61 vdd gnd cell_6t
Xbit_r62_c28 bl_28 br_28 wl_62 vdd gnd cell_6t
Xbit_r63_c28 bl_28 br_28 wl_63 vdd gnd cell_6t
Xbit_r64_c28 bl_28 br_28 wl_64 vdd gnd cell_6t
Xbit_r65_c28 bl_28 br_28 wl_65 vdd gnd cell_6t
Xbit_r66_c28 bl_28 br_28 wl_66 vdd gnd cell_6t
Xbit_r67_c28 bl_28 br_28 wl_67 vdd gnd cell_6t
Xbit_r68_c28 bl_28 br_28 wl_68 vdd gnd cell_6t
Xbit_r69_c28 bl_28 br_28 wl_69 vdd gnd cell_6t
Xbit_r70_c28 bl_28 br_28 wl_70 vdd gnd cell_6t
Xbit_r71_c28 bl_28 br_28 wl_71 vdd gnd cell_6t
Xbit_r72_c28 bl_28 br_28 wl_72 vdd gnd cell_6t
Xbit_r73_c28 bl_28 br_28 wl_73 vdd gnd cell_6t
Xbit_r74_c28 bl_28 br_28 wl_74 vdd gnd cell_6t
Xbit_r75_c28 bl_28 br_28 wl_75 vdd gnd cell_6t
Xbit_r76_c28 bl_28 br_28 wl_76 vdd gnd cell_6t
Xbit_r77_c28 bl_28 br_28 wl_77 vdd gnd cell_6t
Xbit_r78_c28 bl_28 br_28 wl_78 vdd gnd cell_6t
Xbit_r79_c28 bl_28 br_28 wl_79 vdd gnd cell_6t
Xbit_r80_c28 bl_28 br_28 wl_80 vdd gnd cell_6t
Xbit_r81_c28 bl_28 br_28 wl_81 vdd gnd cell_6t
Xbit_r82_c28 bl_28 br_28 wl_82 vdd gnd cell_6t
Xbit_r83_c28 bl_28 br_28 wl_83 vdd gnd cell_6t
Xbit_r84_c28 bl_28 br_28 wl_84 vdd gnd cell_6t
Xbit_r85_c28 bl_28 br_28 wl_85 vdd gnd cell_6t
Xbit_r86_c28 bl_28 br_28 wl_86 vdd gnd cell_6t
Xbit_r87_c28 bl_28 br_28 wl_87 vdd gnd cell_6t
Xbit_r88_c28 bl_28 br_28 wl_88 vdd gnd cell_6t
Xbit_r89_c28 bl_28 br_28 wl_89 vdd gnd cell_6t
Xbit_r90_c28 bl_28 br_28 wl_90 vdd gnd cell_6t
Xbit_r91_c28 bl_28 br_28 wl_91 vdd gnd cell_6t
Xbit_r92_c28 bl_28 br_28 wl_92 vdd gnd cell_6t
Xbit_r93_c28 bl_28 br_28 wl_93 vdd gnd cell_6t
Xbit_r94_c28 bl_28 br_28 wl_94 vdd gnd cell_6t
Xbit_r95_c28 bl_28 br_28 wl_95 vdd gnd cell_6t
Xbit_r96_c28 bl_28 br_28 wl_96 vdd gnd cell_6t
Xbit_r97_c28 bl_28 br_28 wl_97 vdd gnd cell_6t
Xbit_r98_c28 bl_28 br_28 wl_98 vdd gnd cell_6t
Xbit_r99_c28 bl_28 br_28 wl_99 vdd gnd cell_6t
Xbit_r100_c28 bl_28 br_28 wl_100 vdd gnd cell_6t
Xbit_r101_c28 bl_28 br_28 wl_101 vdd gnd cell_6t
Xbit_r102_c28 bl_28 br_28 wl_102 vdd gnd cell_6t
Xbit_r103_c28 bl_28 br_28 wl_103 vdd gnd cell_6t
Xbit_r104_c28 bl_28 br_28 wl_104 vdd gnd cell_6t
Xbit_r105_c28 bl_28 br_28 wl_105 vdd gnd cell_6t
Xbit_r106_c28 bl_28 br_28 wl_106 vdd gnd cell_6t
Xbit_r107_c28 bl_28 br_28 wl_107 vdd gnd cell_6t
Xbit_r108_c28 bl_28 br_28 wl_108 vdd gnd cell_6t
Xbit_r109_c28 bl_28 br_28 wl_109 vdd gnd cell_6t
Xbit_r110_c28 bl_28 br_28 wl_110 vdd gnd cell_6t
Xbit_r111_c28 bl_28 br_28 wl_111 vdd gnd cell_6t
Xbit_r112_c28 bl_28 br_28 wl_112 vdd gnd cell_6t
Xbit_r113_c28 bl_28 br_28 wl_113 vdd gnd cell_6t
Xbit_r114_c28 bl_28 br_28 wl_114 vdd gnd cell_6t
Xbit_r115_c28 bl_28 br_28 wl_115 vdd gnd cell_6t
Xbit_r116_c28 bl_28 br_28 wl_116 vdd gnd cell_6t
Xbit_r117_c28 bl_28 br_28 wl_117 vdd gnd cell_6t
Xbit_r118_c28 bl_28 br_28 wl_118 vdd gnd cell_6t
Xbit_r119_c28 bl_28 br_28 wl_119 vdd gnd cell_6t
Xbit_r120_c28 bl_28 br_28 wl_120 vdd gnd cell_6t
Xbit_r121_c28 bl_28 br_28 wl_121 vdd gnd cell_6t
Xbit_r122_c28 bl_28 br_28 wl_122 vdd gnd cell_6t
Xbit_r123_c28 bl_28 br_28 wl_123 vdd gnd cell_6t
Xbit_r124_c28 bl_28 br_28 wl_124 vdd gnd cell_6t
Xbit_r125_c28 bl_28 br_28 wl_125 vdd gnd cell_6t
Xbit_r126_c28 bl_28 br_28 wl_126 vdd gnd cell_6t
Xbit_r127_c28 bl_28 br_28 wl_127 vdd gnd cell_6t
Xbit_r128_c28 bl_28 br_28 wl_128 vdd gnd cell_6t
Xbit_r129_c28 bl_28 br_28 wl_129 vdd gnd cell_6t
Xbit_r130_c28 bl_28 br_28 wl_130 vdd gnd cell_6t
Xbit_r131_c28 bl_28 br_28 wl_131 vdd gnd cell_6t
Xbit_r132_c28 bl_28 br_28 wl_132 vdd gnd cell_6t
Xbit_r133_c28 bl_28 br_28 wl_133 vdd gnd cell_6t
Xbit_r134_c28 bl_28 br_28 wl_134 vdd gnd cell_6t
Xbit_r135_c28 bl_28 br_28 wl_135 vdd gnd cell_6t
Xbit_r136_c28 bl_28 br_28 wl_136 vdd gnd cell_6t
Xbit_r137_c28 bl_28 br_28 wl_137 vdd gnd cell_6t
Xbit_r138_c28 bl_28 br_28 wl_138 vdd gnd cell_6t
Xbit_r139_c28 bl_28 br_28 wl_139 vdd gnd cell_6t
Xbit_r140_c28 bl_28 br_28 wl_140 vdd gnd cell_6t
Xbit_r141_c28 bl_28 br_28 wl_141 vdd gnd cell_6t
Xbit_r142_c28 bl_28 br_28 wl_142 vdd gnd cell_6t
Xbit_r143_c28 bl_28 br_28 wl_143 vdd gnd cell_6t
Xbit_r144_c28 bl_28 br_28 wl_144 vdd gnd cell_6t
Xbit_r145_c28 bl_28 br_28 wl_145 vdd gnd cell_6t
Xbit_r146_c28 bl_28 br_28 wl_146 vdd gnd cell_6t
Xbit_r147_c28 bl_28 br_28 wl_147 vdd gnd cell_6t
Xbit_r148_c28 bl_28 br_28 wl_148 vdd gnd cell_6t
Xbit_r149_c28 bl_28 br_28 wl_149 vdd gnd cell_6t
Xbit_r150_c28 bl_28 br_28 wl_150 vdd gnd cell_6t
Xbit_r151_c28 bl_28 br_28 wl_151 vdd gnd cell_6t
Xbit_r152_c28 bl_28 br_28 wl_152 vdd gnd cell_6t
Xbit_r153_c28 bl_28 br_28 wl_153 vdd gnd cell_6t
Xbit_r154_c28 bl_28 br_28 wl_154 vdd gnd cell_6t
Xbit_r155_c28 bl_28 br_28 wl_155 vdd gnd cell_6t
Xbit_r156_c28 bl_28 br_28 wl_156 vdd gnd cell_6t
Xbit_r157_c28 bl_28 br_28 wl_157 vdd gnd cell_6t
Xbit_r158_c28 bl_28 br_28 wl_158 vdd gnd cell_6t
Xbit_r159_c28 bl_28 br_28 wl_159 vdd gnd cell_6t
Xbit_r160_c28 bl_28 br_28 wl_160 vdd gnd cell_6t
Xbit_r161_c28 bl_28 br_28 wl_161 vdd gnd cell_6t
Xbit_r162_c28 bl_28 br_28 wl_162 vdd gnd cell_6t
Xbit_r163_c28 bl_28 br_28 wl_163 vdd gnd cell_6t
Xbit_r164_c28 bl_28 br_28 wl_164 vdd gnd cell_6t
Xbit_r165_c28 bl_28 br_28 wl_165 vdd gnd cell_6t
Xbit_r166_c28 bl_28 br_28 wl_166 vdd gnd cell_6t
Xbit_r167_c28 bl_28 br_28 wl_167 vdd gnd cell_6t
Xbit_r168_c28 bl_28 br_28 wl_168 vdd gnd cell_6t
Xbit_r169_c28 bl_28 br_28 wl_169 vdd gnd cell_6t
Xbit_r170_c28 bl_28 br_28 wl_170 vdd gnd cell_6t
Xbit_r171_c28 bl_28 br_28 wl_171 vdd gnd cell_6t
Xbit_r172_c28 bl_28 br_28 wl_172 vdd gnd cell_6t
Xbit_r173_c28 bl_28 br_28 wl_173 vdd gnd cell_6t
Xbit_r174_c28 bl_28 br_28 wl_174 vdd gnd cell_6t
Xbit_r175_c28 bl_28 br_28 wl_175 vdd gnd cell_6t
Xbit_r176_c28 bl_28 br_28 wl_176 vdd gnd cell_6t
Xbit_r177_c28 bl_28 br_28 wl_177 vdd gnd cell_6t
Xbit_r178_c28 bl_28 br_28 wl_178 vdd gnd cell_6t
Xbit_r179_c28 bl_28 br_28 wl_179 vdd gnd cell_6t
Xbit_r180_c28 bl_28 br_28 wl_180 vdd gnd cell_6t
Xbit_r181_c28 bl_28 br_28 wl_181 vdd gnd cell_6t
Xbit_r182_c28 bl_28 br_28 wl_182 vdd gnd cell_6t
Xbit_r183_c28 bl_28 br_28 wl_183 vdd gnd cell_6t
Xbit_r184_c28 bl_28 br_28 wl_184 vdd gnd cell_6t
Xbit_r185_c28 bl_28 br_28 wl_185 vdd gnd cell_6t
Xbit_r186_c28 bl_28 br_28 wl_186 vdd gnd cell_6t
Xbit_r187_c28 bl_28 br_28 wl_187 vdd gnd cell_6t
Xbit_r188_c28 bl_28 br_28 wl_188 vdd gnd cell_6t
Xbit_r189_c28 bl_28 br_28 wl_189 vdd gnd cell_6t
Xbit_r190_c28 bl_28 br_28 wl_190 vdd gnd cell_6t
Xbit_r191_c28 bl_28 br_28 wl_191 vdd gnd cell_6t
Xbit_r192_c28 bl_28 br_28 wl_192 vdd gnd cell_6t
Xbit_r193_c28 bl_28 br_28 wl_193 vdd gnd cell_6t
Xbit_r194_c28 bl_28 br_28 wl_194 vdd gnd cell_6t
Xbit_r195_c28 bl_28 br_28 wl_195 vdd gnd cell_6t
Xbit_r196_c28 bl_28 br_28 wl_196 vdd gnd cell_6t
Xbit_r197_c28 bl_28 br_28 wl_197 vdd gnd cell_6t
Xbit_r198_c28 bl_28 br_28 wl_198 vdd gnd cell_6t
Xbit_r199_c28 bl_28 br_28 wl_199 vdd gnd cell_6t
Xbit_r200_c28 bl_28 br_28 wl_200 vdd gnd cell_6t
Xbit_r201_c28 bl_28 br_28 wl_201 vdd gnd cell_6t
Xbit_r202_c28 bl_28 br_28 wl_202 vdd gnd cell_6t
Xbit_r203_c28 bl_28 br_28 wl_203 vdd gnd cell_6t
Xbit_r204_c28 bl_28 br_28 wl_204 vdd gnd cell_6t
Xbit_r205_c28 bl_28 br_28 wl_205 vdd gnd cell_6t
Xbit_r206_c28 bl_28 br_28 wl_206 vdd gnd cell_6t
Xbit_r207_c28 bl_28 br_28 wl_207 vdd gnd cell_6t
Xbit_r208_c28 bl_28 br_28 wl_208 vdd gnd cell_6t
Xbit_r209_c28 bl_28 br_28 wl_209 vdd gnd cell_6t
Xbit_r210_c28 bl_28 br_28 wl_210 vdd gnd cell_6t
Xbit_r211_c28 bl_28 br_28 wl_211 vdd gnd cell_6t
Xbit_r212_c28 bl_28 br_28 wl_212 vdd gnd cell_6t
Xbit_r213_c28 bl_28 br_28 wl_213 vdd gnd cell_6t
Xbit_r214_c28 bl_28 br_28 wl_214 vdd gnd cell_6t
Xbit_r215_c28 bl_28 br_28 wl_215 vdd gnd cell_6t
Xbit_r216_c28 bl_28 br_28 wl_216 vdd gnd cell_6t
Xbit_r217_c28 bl_28 br_28 wl_217 vdd gnd cell_6t
Xbit_r218_c28 bl_28 br_28 wl_218 vdd gnd cell_6t
Xbit_r219_c28 bl_28 br_28 wl_219 vdd gnd cell_6t
Xbit_r220_c28 bl_28 br_28 wl_220 vdd gnd cell_6t
Xbit_r221_c28 bl_28 br_28 wl_221 vdd gnd cell_6t
Xbit_r222_c28 bl_28 br_28 wl_222 vdd gnd cell_6t
Xbit_r223_c28 bl_28 br_28 wl_223 vdd gnd cell_6t
Xbit_r224_c28 bl_28 br_28 wl_224 vdd gnd cell_6t
Xbit_r225_c28 bl_28 br_28 wl_225 vdd gnd cell_6t
Xbit_r226_c28 bl_28 br_28 wl_226 vdd gnd cell_6t
Xbit_r227_c28 bl_28 br_28 wl_227 vdd gnd cell_6t
Xbit_r228_c28 bl_28 br_28 wl_228 vdd gnd cell_6t
Xbit_r229_c28 bl_28 br_28 wl_229 vdd gnd cell_6t
Xbit_r230_c28 bl_28 br_28 wl_230 vdd gnd cell_6t
Xbit_r231_c28 bl_28 br_28 wl_231 vdd gnd cell_6t
Xbit_r232_c28 bl_28 br_28 wl_232 vdd gnd cell_6t
Xbit_r233_c28 bl_28 br_28 wl_233 vdd gnd cell_6t
Xbit_r234_c28 bl_28 br_28 wl_234 vdd gnd cell_6t
Xbit_r235_c28 bl_28 br_28 wl_235 vdd gnd cell_6t
Xbit_r236_c28 bl_28 br_28 wl_236 vdd gnd cell_6t
Xbit_r237_c28 bl_28 br_28 wl_237 vdd gnd cell_6t
Xbit_r238_c28 bl_28 br_28 wl_238 vdd gnd cell_6t
Xbit_r239_c28 bl_28 br_28 wl_239 vdd gnd cell_6t
Xbit_r240_c28 bl_28 br_28 wl_240 vdd gnd cell_6t
Xbit_r241_c28 bl_28 br_28 wl_241 vdd gnd cell_6t
Xbit_r242_c28 bl_28 br_28 wl_242 vdd gnd cell_6t
Xbit_r243_c28 bl_28 br_28 wl_243 vdd gnd cell_6t
Xbit_r244_c28 bl_28 br_28 wl_244 vdd gnd cell_6t
Xbit_r245_c28 bl_28 br_28 wl_245 vdd gnd cell_6t
Xbit_r246_c28 bl_28 br_28 wl_246 vdd gnd cell_6t
Xbit_r247_c28 bl_28 br_28 wl_247 vdd gnd cell_6t
Xbit_r248_c28 bl_28 br_28 wl_248 vdd gnd cell_6t
Xbit_r249_c28 bl_28 br_28 wl_249 vdd gnd cell_6t
Xbit_r250_c28 bl_28 br_28 wl_250 vdd gnd cell_6t
Xbit_r251_c28 bl_28 br_28 wl_251 vdd gnd cell_6t
Xbit_r252_c28 bl_28 br_28 wl_252 vdd gnd cell_6t
Xbit_r253_c28 bl_28 br_28 wl_253 vdd gnd cell_6t
Xbit_r254_c28 bl_28 br_28 wl_254 vdd gnd cell_6t
Xbit_r255_c28 bl_28 br_28 wl_255 vdd gnd cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd cell_6t
Xbit_r1_c29 bl_29 br_29 wl_1 vdd gnd cell_6t
Xbit_r2_c29 bl_29 br_29 wl_2 vdd gnd cell_6t
Xbit_r3_c29 bl_29 br_29 wl_3 vdd gnd cell_6t
Xbit_r4_c29 bl_29 br_29 wl_4 vdd gnd cell_6t
Xbit_r5_c29 bl_29 br_29 wl_5 vdd gnd cell_6t
Xbit_r6_c29 bl_29 br_29 wl_6 vdd gnd cell_6t
Xbit_r7_c29 bl_29 br_29 wl_7 vdd gnd cell_6t
Xbit_r8_c29 bl_29 br_29 wl_8 vdd gnd cell_6t
Xbit_r9_c29 bl_29 br_29 wl_9 vdd gnd cell_6t
Xbit_r10_c29 bl_29 br_29 wl_10 vdd gnd cell_6t
Xbit_r11_c29 bl_29 br_29 wl_11 vdd gnd cell_6t
Xbit_r12_c29 bl_29 br_29 wl_12 vdd gnd cell_6t
Xbit_r13_c29 bl_29 br_29 wl_13 vdd gnd cell_6t
Xbit_r14_c29 bl_29 br_29 wl_14 vdd gnd cell_6t
Xbit_r15_c29 bl_29 br_29 wl_15 vdd gnd cell_6t
Xbit_r16_c29 bl_29 br_29 wl_16 vdd gnd cell_6t
Xbit_r17_c29 bl_29 br_29 wl_17 vdd gnd cell_6t
Xbit_r18_c29 bl_29 br_29 wl_18 vdd gnd cell_6t
Xbit_r19_c29 bl_29 br_29 wl_19 vdd gnd cell_6t
Xbit_r20_c29 bl_29 br_29 wl_20 vdd gnd cell_6t
Xbit_r21_c29 bl_29 br_29 wl_21 vdd gnd cell_6t
Xbit_r22_c29 bl_29 br_29 wl_22 vdd gnd cell_6t
Xbit_r23_c29 bl_29 br_29 wl_23 vdd gnd cell_6t
Xbit_r24_c29 bl_29 br_29 wl_24 vdd gnd cell_6t
Xbit_r25_c29 bl_29 br_29 wl_25 vdd gnd cell_6t
Xbit_r26_c29 bl_29 br_29 wl_26 vdd gnd cell_6t
Xbit_r27_c29 bl_29 br_29 wl_27 vdd gnd cell_6t
Xbit_r28_c29 bl_29 br_29 wl_28 vdd gnd cell_6t
Xbit_r29_c29 bl_29 br_29 wl_29 vdd gnd cell_6t
Xbit_r30_c29 bl_29 br_29 wl_30 vdd gnd cell_6t
Xbit_r31_c29 bl_29 br_29 wl_31 vdd gnd cell_6t
Xbit_r32_c29 bl_29 br_29 wl_32 vdd gnd cell_6t
Xbit_r33_c29 bl_29 br_29 wl_33 vdd gnd cell_6t
Xbit_r34_c29 bl_29 br_29 wl_34 vdd gnd cell_6t
Xbit_r35_c29 bl_29 br_29 wl_35 vdd gnd cell_6t
Xbit_r36_c29 bl_29 br_29 wl_36 vdd gnd cell_6t
Xbit_r37_c29 bl_29 br_29 wl_37 vdd gnd cell_6t
Xbit_r38_c29 bl_29 br_29 wl_38 vdd gnd cell_6t
Xbit_r39_c29 bl_29 br_29 wl_39 vdd gnd cell_6t
Xbit_r40_c29 bl_29 br_29 wl_40 vdd gnd cell_6t
Xbit_r41_c29 bl_29 br_29 wl_41 vdd gnd cell_6t
Xbit_r42_c29 bl_29 br_29 wl_42 vdd gnd cell_6t
Xbit_r43_c29 bl_29 br_29 wl_43 vdd gnd cell_6t
Xbit_r44_c29 bl_29 br_29 wl_44 vdd gnd cell_6t
Xbit_r45_c29 bl_29 br_29 wl_45 vdd gnd cell_6t
Xbit_r46_c29 bl_29 br_29 wl_46 vdd gnd cell_6t
Xbit_r47_c29 bl_29 br_29 wl_47 vdd gnd cell_6t
Xbit_r48_c29 bl_29 br_29 wl_48 vdd gnd cell_6t
Xbit_r49_c29 bl_29 br_29 wl_49 vdd gnd cell_6t
Xbit_r50_c29 bl_29 br_29 wl_50 vdd gnd cell_6t
Xbit_r51_c29 bl_29 br_29 wl_51 vdd gnd cell_6t
Xbit_r52_c29 bl_29 br_29 wl_52 vdd gnd cell_6t
Xbit_r53_c29 bl_29 br_29 wl_53 vdd gnd cell_6t
Xbit_r54_c29 bl_29 br_29 wl_54 vdd gnd cell_6t
Xbit_r55_c29 bl_29 br_29 wl_55 vdd gnd cell_6t
Xbit_r56_c29 bl_29 br_29 wl_56 vdd gnd cell_6t
Xbit_r57_c29 bl_29 br_29 wl_57 vdd gnd cell_6t
Xbit_r58_c29 bl_29 br_29 wl_58 vdd gnd cell_6t
Xbit_r59_c29 bl_29 br_29 wl_59 vdd gnd cell_6t
Xbit_r60_c29 bl_29 br_29 wl_60 vdd gnd cell_6t
Xbit_r61_c29 bl_29 br_29 wl_61 vdd gnd cell_6t
Xbit_r62_c29 bl_29 br_29 wl_62 vdd gnd cell_6t
Xbit_r63_c29 bl_29 br_29 wl_63 vdd gnd cell_6t
Xbit_r64_c29 bl_29 br_29 wl_64 vdd gnd cell_6t
Xbit_r65_c29 bl_29 br_29 wl_65 vdd gnd cell_6t
Xbit_r66_c29 bl_29 br_29 wl_66 vdd gnd cell_6t
Xbit_r67_c29 bl_29 br_29 wl_67 vdd gnd cell_6t
Xbit_r68_c29 bl_29 br_29 wl_68 vdd gnd cell_6t
Xbit_r69_c29 bl_29 br_29 wl_69 vdd gnd cell_6t
Xbit_r70_c29 bl_29 br_29 wl_70 vdd gnd cell_6t
Xbit_r71_c29 bl_29 br_29 wl_71 vdd gnd cell_6t
Xbit_r72_c29 bl_29 br_29 wl_72 vdd gnd cell_6t
Xbit_r73_c29 bl_29 br_29 wl_73 vdd gnd cell_6t
Xbit_r74_c29 bl_29 br_29 wl_74 vdd gnd cell_6t
Xbit_r75_c29 bl_29 br_29 wl_75 vdd gnd cell_6t
Xbit_r76_c29 bl_29 br_29 wl_76 vdd gnd cell_6t
Xbit_r77_c29 bl_29 br_29 wl_77 vdd gnd cell_6t
Xbit_r78_c29 bl_29 br_29 wl_78 vdd gnd cell_6t
Xbit_r79_c29 bl_29 br_29 wl_79 vdd gnd cell_6t
Xbit_r80_c29 bl_29 br_29 wl_80 vdd gnd cell_6t
Xbit_r81_c29 bl_29 br_29 wl_81 vdd gnd cell_6t
Xbit_r82_c29 bl_29 br_29 wl_82 vdd gnd cell_6t
Xbit_r83_c29 bl_29 br_29 wl_83 vdd gnd cell_6t
Xbit_r84_c29 bl_29 br_29 wl_84 vdd gnd cell_6t
Xbit_r85_c29 bl_29 br_29 wl_85 vdd gnd cell_6t
Xbit_r86_c29 bl_29 br_29 wl_86 vdd gnd cell_6t
Xbit_r87_c29 bl_29 br_29 wl_87 vdd gnd cell_6t
Xbit_r88_c29 bl_29 br_29 wl_88 vdd gnd cell_6t
Xbit_r89_c29 bl_29 br_29 wl_89 vdd gnd cell_6t
Xbit_r90_c29 bl_29 br_29 wl_90 vdd gnd cell_6t
Xbit_r91_c29 bl_29 br_29 wl_91 vdd gnd cell_6t
Xbit_r92_c29 bl_29 br_29 wl_92 vdd gnd cell_6t
Xbit_r93_c29 bl_29 br_29 wl_93 vdd gnd cell_6t
Xbit_r94_c29 bl_29 br_29 wl_94 vdd gnd cell_6t
Xbit_r95_c29 bl_29 br_29 wl_95 vdd gnd cell_6t
Xbit_r96_c29 bl_29 br_29 wl_96 vdd gnd cell_6t
Xbit_r97_c29 bl_29 br_29 wl_97 vdd gnd cell_6t
Xbit_r98_c29 bl_29 br_29 wl_98 vdd gnd cell_6t
Xbit_r99_c29 bl_29 br_29 wl_99 vdd gnd cell_6t
Xbit_r100_c29 bl_29 br_29 wl_100 vdd gnd cell_6t
Xbit_r101_c29 bl_29 br_29 wl_101 vdd gnd cell_6t
Xbit_r102_c29 bl_29 br_29 wl_102 vdd gnd cell_6t
Xbit_r103_c29 bl_29 br_29 wl_103 vdd gnd cell_6t
Xbit_r104_c29 bl_29 br_29 wl_104 vdd gnd cell_6t
Xbit_r105_c29 bl_29 br_29 wl_105 vdd gnd cell_6t
Xbit_r106_c29 bl_29 br_29 wl_106 vdd gnd cell_6t
Xbit_r107_c29 bl_29 br_29 wl_107 vdd gnd cell_6t
Xbit_r108_c29 bl_29 br_29 wl_108 vdd gnd cell_6t
Xbit_r109_c29 bl_29 br_29 wl_109 vdd gnd cell_6t
Xbit_r110_c29 bl_29 br_29 wl_110 vdd gnd cell_6t
Xbit_r111_c29 bl_29 br_29 wl_111 vdd gnd cell_6t
Xbit_r112_c29 bl_29 br_29 wl_112 vdd gnd cell_6t
Xbit_r113_c29 bl_29 br_29 wl_113 vdd gnd cell_6t
Xbit_r114_c29 bl_29 br_29 wl_114 vdd gnd cell_6t
Xbit_r115_c29 bl_29 br_29 wl_115 vdd gnd cell_6t
Xbit_r116_c29 bl_29 br_29 wl_116 vdd gnd cell_6t
Xbit_r117_c29 bl_29 br_29 wl_117 vdd gnd cell_6t
Xbit_r118_c29 bl_29 br_29 wl_118 vdd gnd cell_6t
Xbit_r119_c29 bl_29 br_29 wl_119 vdd gnd cell_6t
Xbit_r120_c29 bl_29 br_29 wl_120 vdd gnd cell_6t
Xbit_r121_c29 bl_29 br_29 wl_121 vdd gnd cell_6t
Xbit_r122_c29 bl_29 br_29 wl_122 vdd gnd cell_6t
Xbit_r123_c29 bl_29 br_29 wl_123 vdd gnd cell_6t
Xbit_r124_c29 bl_29 br_29 wl_124 vdd gnd cell_6t
Xbit_r125_c29 bl_29 br_29 wl_125 vdd gnd cell_6t
Xbit_r126_c29 bl_29 br_29 wl_126 vdd gnd cell_6t
Xbit_r127_c29 bl_29 br_29 wl_127 vdd gnd cell_6t
Xbit_r128_c29 bl_29 br_29 wl_128 vdd gnd cell_6t
Xbit_r129_c29 bl_29 br_29 wl_129 vdd gnd cell_6t
Xbit_r130_c29 bl_29 br_29 wl_130 vdd gnd cell_6t
Xbit_r131_c29 bl_29 br_29 wl_131 vdd gnd cell_6t
Xbit_r132_c29 bl_29 br_29 wl_132 vdd gnd cell_6t
Xbit_r133_c29 bl_29 br_29 wl_133 vdd gnd cell_6t
Xbit_r134_c29 bl_29 br_29 wl_134 vdd gnd cell_6t
Xbit_r135_c29 bl_29 br_29 wl_135 vdd gnd cell_6t
Xbit_r136_c29 bl_29 br_29 wl_136 vdd gnd cell_6t
Xbit_r137_c29 bl_29 br_29 wl_137 vdd gnd cell_6t
Xbit_r138_c29 bl_29 br_29 wl_138 vdd gnd cell_6t
Xbit_r139_c29 bl_29 br_29 wl_139 vdd gnd cell_6t
Xbit_r140_c29 bl_29 br_29 wl_140 vdd gnd cell_6t
Xbit_r141_c29 bl_29 br_29 wl_141 vdd gnd cell_6t
Xbit_r142_c29 bl_29 br_29 wl_142 vdd gnd cell_6t
Xbit_r143_c29 bl_29 br_29 wl_143 vdd gnd cell_6t
Xbit_r144_c29 bl_29 br_29 wl_144 vdd gnd cell_6t
Xbit_r145_c29 bl_29 br_29 wl_145 vdd gnd cell_6t
Xbit_r146_c29 bl_29 br_29 wl_146 vdd gnd cell_6t
Xbit_r147_c29 bl_29 br_29 wl_147 vdd gnd cell_6t
Xbit_r148_c29 bl_29 br_29 wl_148 vdd gnd cell_6t
Xbit_r149_c29 bl_29 br_29 wl_149 vdd gnd cell_6t
Xbit_r150_c29 bl_29 br_29 wl_150 vdd gnd cell_6t
Xbit_r151_c29 bl_29 br_29 wl_151 vdd gnd cell_6t
Xbit_r152_c29 bl_29 br_29 wl_152 vdd gnd cell_6t
Xbit_r153_c29 bl_29 br_29 wl_153 vdd gnd cell_6t
Xbit_r154_c29 bl_29 br_29 wl_154 vdd gnd cell_6t
Xbit_r155_c29 bl_29 br_29 wl_155 vdd gnd cell_6t
Xbit_r156_c29 bl_29 br_29 wl_156 vdd gnd cell_6t
Xbit_r157_c29 bl_29 br_29 wl_157 vdd gnd cell_6t
Xbit_r158_c29 bl_29 br_29 wl_158 vdd gnd cell_6t
Xbit_r159_c29 bl_29 br_29 wl_159 vdd gnd cell_6t
Xbit_r160_c29 bl_29 br_29 wl_160 vdd gnd cell_6t
Xbit_r161_c29 bl_29 br_29 wl_161 vdd gnd cell_6t
Xbit_r162_c29 bl_29 br_29 wl_162 vdd gnd cell_6t
Xbit_r163_c29 bl_29 br_29 wl_163 vdd gnd cell_6t
Xbit_r164_c29 bl_29 br_29 wl_164 vdd gnd cell_6t
Xbit_r165_c29 bl_29 br_29 wl_165 vdd gnd cell_6t
Xbit_r166_c29 bl_29 br_29 wl_166 vdd gnd cell_6t
Xbit_r167_c29 bl_29 br_29 wl_167 vdd gnd cell_6t
Xbit_r168_c29 bl_29 br_29 wl_168 vdd gnd cell_6t
Xbit_r169_c29 bl_29 br_29 wl_169 vdd gnd cell_6t
Xbit_r170_c29 bl_29 br_29 wl_170 vdd gnd cell_6t
Xbit_r171_c29 bl_29 br_29 wl_171 vdd gnd cell_6t
Xbit_r172_c29 bl_29 br_29 wl_172 vdd gnd cell_6t
Xbit_r173_c29 bl_29 br_29 wl_173 vdd gnd cell_6t
Xbit_r174_c29 bl_29 br_29 wl_174 vdd gnd cell_6t
Xbit_r175_c29 bl_29 br_29 wl_175 vdd gnd cell_6t
Xbit_r176_c29 bl_29 br_29 wl_176 vdd gnd cell_6t
Xbit_r177_c29 bl_29 br_29 wl_177 vdd gnd cell_6t
Xbit_r178_c29 bl_29 br_29 wl_178 vdd gnd cell_6t
Xbit_r179_c29 bl_29 br_29 wl_179 vdd gnd cell_6t
Xbit_r180_c29 bl_29 br_29 wl_180 vdd gnd cell_6t
Xbit_r181_c29 bl_29 br_29 wl_181 vdd gnd cell_6t
Xbit_r182_c29 bl_29 br_29 wl_182 vdd gnd cell_6t
Xbit_r183_c29 bl_29 br_29 wl_183 vdd gnd cell_6t
Xbit_r184_c29 bl_29 br_29 wl_184 vdd gnd cell_6t
Xbit_r185_c29 bl_29 br_29 wl_185 vdd gnd cell_6t
Xbit_r186_c29 bl_29 br_29 wl_186 vdd gnd cell_6t
Xbit_r187_c29 bl_29 br_29 wl_187 vdd gnd cell_6t
Xbit_r188_c29 bl_29 br_29 wl_188 vdd gnd cell_6t
Xbit_r189_c29 bl_29 br_29 wl_189 vdd gnd cell_6t
Xbit_r190_c29 bl_29 br_29 wl_190 vdd gnd cell_6t
Xbit_r191_c29 bl_29 br_29 wl_191 vdd gnd cell_6t
Xbit_r192_c29 bl_29 br_29 wl_192 vdd gnd cell_6t
Xbit_r193_c29 bl_29 br_29 wl_193 vdd gnd cell_6t
Xbit_r194_c29 bl_29 br_29 wl_194 vdd gnd cell_6t
Xbit_r195_c29 bl_29 br_29 wl_195 vdd gnd cell_6t
Xbit_r196_c29 bl_29 br_29 wl_196 vdd gnd cell_6t
Xbit_r197_c29 bl_29 br_29 wl_197 vdd gnd cell_6t
Xbit_r198_c29 bl_29 br_29 wl_198 vdd gnd cell_6t
Xbit_r199_c29 bl_29 br_29 wl_199 vdd gnd cell_6t
Xbit_r200_c29 bl_29 br_29 wl_200 vdd gnd cell_6t
Xbit_r201_c29 bl_29 br_29 wl_201 vdd gnd cell_6t
Xbit_r202_c29 bl_29 br_29 wl_202 vdd gnd cell_6t
Xbit_r203_c29 bl_29 br_29 wl_203 vdd gnd cell_6t
Xbit_r204_c29 bl_29 br_29 wl_204 vdd gnd cell_6t
Xbit_r205_c29 bl_29 br_29 wl_205 vdd gnd cell_6t
Xbit_r206_c29 bl_29 br_29 wl_206 vdd gnd cell_6t
Xbit_r207_c29 bl_29 br_29 wl_207 vdd gnd cell_6t
Xbit_r208_c29 bl_29 br_29 wl_208 vdd gnd cell_6t
Xbit_r209_c29 bl_29 br_29 wl_209 vdd gnd cell_6t
Xbit_r210_c29 bl_29 br_29 wl_210 vdd gnd cell_6t
Xbit_r211_c29 bl_29 br_29 wl_211 vdd gnd cell_6t
Xbit_r212_c29 bl_29 br_29 wl_212 vdd gnd cell_6t
Xbit_r213_c29 bl_29 br_29 wl_213 vdd gnd cell_6t
Xbit_r214_c29 bl_29 br_29 wl_214 vdd gnd cell_6t
Xbit_r215_c29 bl_29 br_29 wl_215 vdd gnd cell_6t
Xbit_r216_c29 bl_29 br_29 wl_216 vdd gnd cell_6t
Xbit_r217_c29 bl_29 br_29 wl_217 vdd gnd cell_6t
Xbit_r218_c29 bl_29 br_29 wl_218 vdd gnd cell_6t
Xbit_r219_c29 bl_29 br_29 wl_219 vdd gnd cell_6t
Xbit_r220_c29 bl_29 br_29 wl_220 vdd gnd cell_6t
Xbit_r221_c29 bl_29 br_29 wl_221 vdd gnd cell_6t
Xbit_r222_c29 bl_29 br_29 wl_222 vdd gnd cell_6t
Xbit_r223_c29 bl_29 br_29 wl_223 vdd gnd cell_6t
Xbit_r224_c29 bl_29 br_29 wl_224 vdd gnd cell_6t
Xbit_r225_c29 bl_29 br_29 wl_225 vdd gnd cell_6t
Xbit_r226_c29 bl_29 br_29 wl_226 vdd gnd cell_6t
Xbit_r227_c29 bl_29 br_29 wl_227 vdd gnd cell_6t
Xbit_r228_c29 bl_29 br_29 wl_228 vdd gnd cell_6t
Xbit_r229_c29 bl_29 br_29 wl_229 vdd gnd cell_6t
Xbit_r230_c29 bl_29 br_29 wl_230 vdd gnd cell_6t
Xbit_r231_c29 bl_29 br_29 wl_231 vdd gnd cell_6t
Xbit_r232_c29 bl_29 br_29 wl_232 vdd gnd cell_6t
Xbit_r233_c29 bl_29 br_29 wl_233 vdd gnd cell_6t
Xbit_r234_c29 bl_29 br_29 wl_234 vdd gnd cell_6t
Xbit_r235_c29 bl_29 br_29 wl_235 vdd gnd cell_6t
Xbit_r236_c29 bl_29 br_29 wl_236 vdd gnd cell_6t
Xbit_r237_c29 bl_29 br_29 wl_237 vdd gnd cell_6t
Xbit_r238_c29 bl_29 br_29 wl_238 vdd gnd cell_6t
Xbit_r239_c29 bl_29 br_29 wl_239 vdd gnd cell_6t
Xbit_r240_c29 bl_29 br_29 wl_240 vdd gnd cell_6t
Xbit_r241_c29 bl_29 br_29 wl_241 vdd gnd cell_6t
Xbit_r242_c29 bl_29 br_29 wl_242 vdd gnd cell_6t
Xbit_r243_c29 bl_29 br_29 wl_243 vdd gnd cell_6t
Xbit_r244_c29 bl_29 br_29 wl_244 vdd gnd cell_6t
Xbit_r245_c29 bl_29 br_29 wl_245 vdd gnd cell_6t
Xbit_r246_c29 bl_29 br_29 wl_246 vdd gnd cell_6t
Xbit_r247_c29 bl_29 br_29 wl_247 vdd gnd cell_6t
Xbit_r248_c29 bl_29 br_29 wl_248 vdd gnd cell_6t
Xbit_r249_c29 bl_29 br_29 wl_249 vdd gnd cell_6t
Xbit_r250_c29 bl_29 br_29 wl_250 vdd gnd cell_6t
Xbit_r251_c29 bl_29 br_29 wl_251 vdd gnd cell_6t
Xbit_r252_c29 bl_29 br_29 wl_252 vdd gnd cell_6t
Xbit_r253_c29 bl_29 br_29 wl_253 vdd gnd cell_6t
Xbit_r254_c29 bl_29 br_29 wl_254 vdd gnd cell_6t
Xbit_r255_c29 bl_29 br_29 wl_255 vdd gnd cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd cell_6t
Xbit_r1_c30 bl_30 br_30 wl_1 vdd gnd cell_6t
Xbit_r2_c30 bl_30 br_30 wl_2 vdd gnd cell_6t
Xbit_r3_c30 bl_30 br_30 wl_3 vdd gnd cell_6t
Xbit_r4_c30 bl_30 br_30 wl_4 vdd gnd cell_6t
Xbit_r5_c30 bl_30 br_30 wl_5 vdd gnd cell_6t
Xbit_r6_c30 bl_30 br_30 wl_6 vdd gnd cell_6t
Xbit_r7_c30 bl_30 br_30 wl_7 vdd gnd cell_6t
Xbit_r8_c30 bl_30 br_30 wl_8 vdd gnd cell_6t
Xbit_r9_c30 bl_30 br_30 wl_9 vdd gnd cell_6t
Xbit_r10_c30 bl_30 br_30 wl_10 vdd gnd cell_6t
Xbit_r11_c30 bl_30 br_30 wl_11 vdd gnd cell_6t
Xbit_r12_c30 bl_30 br_30 wl_12 vdd gnd cell_6t
Xbit_r13_c30 bl_30 br_30 wl_13 vdd gnd cell_6t
Xbit_r14_c30 bl_30 br_30 wl_14 vdd gnd cell_6t
Xbit_r15_c30 bl_30 br_30 wl_15 vdd gnd cell_6t
Xbit_r16_c30 bl_30 br_30 wl_16 vdd gnd cell_6t
Xbit_r17_c30 bl_30 br_30 wl_17 vdd gnd cell_6t
Xbit_r18_c30 bl_30 br_30 wl_18 vdd gnd cell_6t
Xbit_r19_c30 bl_30 br_30 wl_19 vdd gnd cell_6t
Xbit_r20_c30 bl_30 br_30 wl_20 vdd gnd cell_6t
Xbit_r21_c30 bl_30 br_30 wl_21 vdd gnd cell_6t
Xbit_r22_c30 bl_30 br_30 wl_22 vdd gnd cell_6t
Xbit_r23_c30 bl_30 br_30 wl_23 vdd gnd cell_6t
Xbit_r24_c30 bl_30 br_30 wl_24 vdd gnd cell_6t
Xbit_r25_c30 bl_30 br_30 wl_25 vdd gnd cell_6t
Xbit_r26_c30 bl_30 br_30 wl_26 vdd gnd cell_6t
Xbit_r27_c30 bl_30 br_30 wl_27 vdd gnd cell_6t
Xbit_r28_c30 bl_30 br_30 wl_28 vdd gnd cell_6t
Xbit_r29_c30 bl_30 br_30 wl_29 vdd gnd cell_6t
Xbit_r30_c30 bl_30 br_30 wl_30 vdd gnd cell_6t
Xbit_r31_c30 bl_30 br_30 wl_31 vdd gnd cell_6t
Xbit_r32_c30 bl_30 br_30 wl_32 vdd gnd cell_6t
Xbit_r33_c30 bl_30 br_30 wl_33 vdd gnd cell_6t
Xbit_r34_c30 bl_30 br_30 wl_34 vdd gnd cell_6t
Xbit_r35_c30 bl_30 br_30 wl_35 vdd gnd cell_6t
Xbit_r36_c30 bl_30 br_30 wl_36 vdd gnd cell_6t
Xbit_r37_c30 bl_30 br_30 wl_37 vdd gnd cell_6t
Xbit_r38_c30 bl_30 br_30 wl_38 vdd gnd cell_6t
Xbit_r39_c30 bl_30 br_30 wl_39 vdd gnd cell_6t
Xbit_r40_c30 bl_30 br_30 wl_40 vdd gnd cell_6t
Xbit_r41_c30 bl_30 br_30 wl_41 vdd gnd cell_6t
Xbit_r42_c30 bl_30 br_30 wl_42 vdd gnd cell_6t
Xbit_r43_c30 bl_30 br_30 wl_43 vdd gnd cell_6t
Xbit_r44_c30 bl_30 br_30 wl_44 vdd gnd cell_6t
Xbit_r45_c30 bl_30 br_30 wl_45 vdd gnd cell_6t
Xbit_r46_c30 bl_30 br_30 wl_46 vdd gnd cell_6t
Xbit_r47_c30 bl_30 br_30 wl_47 vdd gnd cell_6t
Xbit_r48_c30 bl_30 br_30 wl_48 vdd gnd cell_6t
Xbit_r49_c30 bl_30 br_30 wl_49 vdd gnd cell_6t
Xbit_r50_c30 bl_30 br_30 wl_50 vdd gnd cell_6t
Xbit_r51_c30 bl_30 br_30 wl_51 vdd gnd cell_6t
Xbit_r52_c30 bl_30 br_30 wl_52 vdd gnd cell_6t
Xbit_r53_c30 bl_30 br_30 wl_53 vdd gnd cell_6t
Xbit_r54_c30 bl_30 br_30 wl_54 vdd gnd cell_6t
Xbit_r55_c30 bl_30 br_30 wl_55 vdd gnd cell_6t
Xbit_r56_c30 bl_30 br_30 wl_56 vdd gnd cell_6t
Xbit_r57_c30 bl_30 br_30 wl_57 vdd gnd cell_6t
Xbit_r58_c30 bl_30 br_30 wl_58 vdd gnd cell_6t
Xbit_r59_c30 bl_30 br_30 wl_59 vdd gnd cell_6t
Xbit_r60_c30 bl_30 br_30 wl_60 vdd gnd cell_6t
Xbit_r61_c30 bl_30 br_30 wl_61 vdd gnd cell_6t
Xbit_r62_c30 bl_30 br_30 wl_62 vdd gnd cell_6t
Xbit_r63_c30 bl_30 br_30 wl_63 vdd gnd cell_6t
Xbit_r64_c30 bl_30 br_30 wl_64 vdd gnd cell_6t
Xbit_r65_c30 bl_30 br_30 wl_65 vdd gnd cell_6t
Xbit_r66_c30 bl_30 br_30 wl_66 vdd gnd cell_6t
Xbit_r67_c30 bl_30 br_30 wl_67 vdd gnd cell_6t
Xbit_r68_c30 bl_30 br_30 wl_68 vdd gnd cell_6t
Xbit_r69_c30 bl_30 br_30 wl_69 vdd gnd cell_6t
Xbit_r70_c30 bl_30 br_30 wl_70 vdd gnd cell_6t
Xbit_r71_c30 bl_30 br_30 wl_71 vdd gnd cell_6t
Xbit_r72_c30 bl_30 br_30 wl_72 vdd gnd cell_6t
Xbit_r73_c30 bl_30 br_30 wl_73 vdd gnd cell_6t
Xbit_r74_c30 bl_30 br_30 wl_74 vdd gnd cell_6t
Xbit_r75_c30 bl_30 br_30 wl_75 vdd gnd cell_6t
Xbit_r76_c30 bl_30 br_30 wl_76 vdd gnd cell_6t
Xbit_r77_c30 bl_30 br_30 wl_77 vdd gnd cell_6t
Xbit_r78_c30 bl_30 br_30 wl_78 vdd gnd cell_6t
Xbit_r79_c30 bl_30 br_30 wl_79 vdd gnd cell_6t
Xbit_r80_c30 bl_30 br_30 wl_80 vdd gnd cell_6t
Xbit_r81_c30 bl_30 br_30 wl_81 vdd gnd cell_6t
Xbit_r82_c30 bl_30 br_30 wl_82 vdd gnd cell_6t
Xbit_r83_c30 bl_30 br_30 wl_83 vdd gnd cell_6t
Xbit_r84_c30 bl_30 br_30 wl_84 vdd gnd cell_6t
Xbit_r85_c30 bl_30 br_30 wl_85 vdd gnd cell_6t
Xbit_r86_c30 bl_30 br_30 wl_86 vdd gnd cell_6t
Xbit_r87_c30 bl_30 br_30 wl_87 vdd gnd cell_6t
Xbit_r88_c30 bl_30 br_30 wl_88 vdd gnd cell_6t
Xbit_r89_c30 bl_30 br_30 wl_89 vdd gnd cell_6t
Xbit_r90_c30 bl_30 br_30 wl_90 vdd gnd cell_6t
Xbit_r91_c30 bl_30 br_30 wl_91 vdd gnd cell_6t
Xbit_r92_c30 bl_30 br_30 wl_92 vdd gnd cell_6t
Xbit_r93_c30 bl_30 br_30 wl_93 vdd gnd cell_6t
Xbit_r94_c30 bl_30 br_30 wl_94 vdd gnd cell_6t
Xbit_r95_c30 bl_30 br_30 wl_95 vdd gnd cell_6t
Xbit_r96_c30 bl_30 br_30 wl_96 vdd gnd cell_6t
Xbit_r97_c30 bl_30 br_30 wl_97 vdd gnd cell_6t
Xbit_r98_c30 bl_30 br_30 wl_98 vdd gnd cell_6t
Xbit_r99_c30 bl_30 br_30 wl_99 vdd gnd cell_6t
Xbit_r100_c30 bl_30 br_30 wl_100 vdd gnd cell_6t
Xbit_r101_c30 bl_30 br_30 wl_101 vdd gnd cell_6t
Xbit_r102_c30 bl_30 br_30 wl_102 vdd gnd cell_6t
Xbit_r103_c30 bl_30 br_30 wl_103 vdd gnd cell_6t
Xbit_r104_c30 bl_30 br_30 wl_104 vdd gnd cell_6t
Xbit_r105_c30 bl_30 br_30 wl_105 vdd gnd cell_6t
Xbit_r106_c30 bl_30 br_30 wl_106 vdd gnd cell_6t
Xbit_r107_c30 bl_30 br_30 wl_107 vdd gnd cell_6t
Xbit_r108_c30 bl_30 br_30 wl_108 vdd gnd cell_6t
Xbit_r109_c30 bl_30 br_30 wl_109 vdd gnd cell_6t
Xbit_r110_c30 bl_30 br_30 wl_110 vdd gnd cell_6t
Xbit_r111_c30 bl_30 br_30 wl_111 vdd gnd cell_6t
Xbit_r112_c30 bl_30 br_30 wl_112 vdd gnd cell_6t
Xbit_r113_c30 bl_30 br_30 wl_113 vdd gnd cell_6t
Xbit_r114_c30 bl_30 br_30 wl_114 vdd gnd cell_6t
Xbit_r115_c30 bl_30 br_30 wl_115 vdd gnd cell_6t
Xbit_r116_c30 bl_30 br_30 wl_116 vdd gnd cell_6t
Xbit_r117_c30 bl_30 br_30 wl_117 vdd gnd cell_6t
Xbit_r118_c30 bl_30 br_30 wl_118 vdd gnd cell_6t
Xbit_r119_c30 bl_30 br_30 wl_119 vdd gnd cell_6t
Xbit_r120_c30 bl_30 br_30 wl_120 vdd gnd cell_6t
Xbit_r121_c30 bl_30 br_30 wl_121 vdd gnd cell_6t
Xbit_r122_c30 bl_30 br_30 wl_122 vdd gnd cell_6t
Xbit_r123_c30 bl_30 br_30 wl_123 vdd gnd cell_6t
Xbit_r124_c30 bl_30 br_30 wl_124 vdd gnd cell_6t
Xbit_r125_c30 bl_30 br_30 wl_125 vdd gnd cell_6t
Xbit_r126_c30 bl_30 br_30 wl_126 vdd gnd cell_6t
Xbit_r127_c30 bl_30 br_30 wl_127 vdd gnd cell_6t
Xbit_r128_c30 bl_30 br_30 wl_128 vdd gnd cell_6t
Xbit_r129_c30 bl_30 br_30 wl_129 vdd gnd cell_6t
Xbit_r130_c30 bl_30 br_30 wl_130 vdd gnd cell_6t
Xbit_r131_c30 bl_30 br_30 wl_131 vdd gnd cell_6t
Xbit_r132_c30 bl_30 br_30 wl_132 vdd gnd cell_6t
Xbit_r133_c30 bl_30 br_30 wl_133 vdd gnd cell_6t
Xbit_r134_c30 bl_30 br_30 wl_134 vdd gnd cell_6t
Xbit_r135_c30 bl_30 br_30 wl_135 vdd gnd cell_6t
Xbit_r136_c30 bl_30 br_30 wl_136 vdd gnd cell_6t
Xbit_r137_c30 bl_30 br_30 wl_137 vdd gnd cell_6t
Xbit_r138_c30 bl_30 br_30 wl_138 vdd gnd cell_6t
Xbit_r139_c30 bl_30 br_30 wl_139 vdd gnd cell_6t
Xbit_r140_c30 bl_30 br_30 wl_140 vdd gnd cell_6t
Xbit_r141_c30 bl_30 br_30 wl_141 vdd gnd cell_6t
Xbit_r142_c30 bl_30 br_30 wl_142 vdd gnd cell_6t
Xbit_r143_c30 bl_30 br_30 wl_143 vdd gnd cell_6t
Xbit_r144_c30 bl_30 br_30 wl_144 vdd gnd cell_6t
Xbit_r145_c30 bl_30 br_30 wl_145 vdd gnd cell_6t
Xbit_r146_c30 bl_30 br_30 wl_146 vdd gnd cell_6t
Xbit_r147_c30 bl_30 br_30 wl_147 vdd gnd cell_6t
Xbit_r148_c30 bl_30 br_30 wl_148 vdd gnd cell_6t
Xbit_r149_c30 bl_30 br_30 wl_149 vdd gnd cell_6t
Xbit_r150_c30 bl_30 br_30 wl_150 vdd gnd cell_6t
Xbit_r151_c30 bl_30 br_30 wl_151 vdd gnd cell_6t
Xbit_r152_c30 bl_30 br_30 wl_152 vdd gnd cell_6t
Xbit_r153_c30 bl_30 br_30 wl_153 vdd gnd cell_6t
Xbit_r154_c30 bl_30 br_30 wl_154 vdd gnd cell_6t
Xbit_r155_c30 bl_30 br_30 wl_155 vdd gnd cell_6t
Xbit_r156_c30 bl_30 br_30 wl_156 vdd gnd cell_6t
Xbit_r157_c30 bl_30 br_30 wl_157 vdd gnd cell_6t
Xbit_r158_c30 bl_30 br_30 wl_158 vdd gnd cell_6t
Xbit_r159_c30 bl_30 br_30 wl_159 vdd gnd cell_6t
Xbit_r160_c30 bl_30 br_30 wl_160 vdd gnd cell_6t
Xbit_r161_c30 bl_30 br_30 wl_161 vdd gnd cell_6t
Xbit_r162_c30 bl_30 br_30 wl_162 vdd gnd cell_6t
Xbit_r163_c30 bl_30 br_30 wl_163 vdd gnd cell_6t
Xbit_r164_c30 bl_30 br_30 wl_164 vdd gnd cell_6t
Xbit_r165_c30 bl_30 br_30 wl_165 vdd gnd cell_6t
Xbit_r166_c30 bl_30 br_30 wl_166 vdd gnd cell_6t
Xbit_r167_c30 bl_30 br_30 wl_167 vdd gnd cell_6t
Xbit_r168_c30 bl_30 br_30 wl_168 vdd gnd cell_6t
Xbit_r169_c30 bl_30 br_30 wl_169 vdd gnd cell_6t
Xbit_r170_c30 bl_30 br_30 wl_170 vdd gnd cell_6t
Xbit_r171_c30 bl_30 br_30 wl_171 vdd gnd cell_6t
Xbit_r172_c30 bl_30 br_30 wl_172 vdd gnd cell_6t
Xbit_r173_c30 bl_30 br_30 wl_173 vdd gnd cell_6t
Xbit_r174_c30 bl_30 br_30 wl_174 vdd gnd cell_6t
Xbit_r175_c30 bl_30 br_30 wl_175 vdd gnd cell_6t
Xbit_r176_c30 bl_30 br_30 wl_176 vdd gnd cell_6t
Xbit_r177_c30 bl_30 br_30 wl_177 vdd gnd cell_6t
Xbit_r178_c30 bl_30 br_30 wl_178 vdd gnd cell_6t
Xbit_r179_c30 bl_30 br_30 wl_179 vdd gnd cell_6t
Xbit_r180_c30 bl_30 br_30 wl_180 vdd gnd cell_6t
Xbit_r181_c30 bl_30 br_30 wl_181 vdd gnd cell_6t
Xbit_r182_c30 bl_30 br_30 wl_182 vdd gnd cell_6t
Xbit_r183_c30 bl_30 br_30 wl_183 vdd gnd cell_6t
Xbit_r184_c30 bl_30 br_30 wl_184 vdd gnd cell_6t
Xbit_r185_c30 bl_30 br_30 wl_185 vdd gnd cell_6t
Xbit_r186_c30 bl_30 br_30 wl_186 vdd gnd cell_6t
Xbit_r187_c30 bl_30 br_30 wl_187 vdd gnd cell_6t
Xbit_r188_c30 bl_30 br_30 wl_188 vdd gnd cell_6t
Xbit_r189_c30 bl_30 br_30 wl_189 vdd gnd cell_6t
Xbit_r190_c30 bl_30 br_30 wl_190 vdd gnd cell_6t
Xbit_r191_c30 bl_30 br_30 wl_191 vdd gnd cell_6t
Xbit_r192_c30 bl_30 br_30 wl_192 vdd gnd cell_6t
Xbit_r193_c30 bl_30 br_30 wl_193 vdd gnd cell_6t
Xbit_r194_c30 bl_30 br_30 wl_194 vdd gnd cell_6t
Xbit_r195_c30 bl_30 br_30 wl_195 vdd gnd cell_6t
Xbit_r196_c30 bl_30 br_30 wl_196 vdd gnd cell_6t
Xbit_r197_c30 bl_30 br_30 wl_197 vdd gnd cell_6t
Xbit_r198_c30 bl_30 br_30 wl_198 vdd gnd cell_6t
Xbit_r199_c30 bl_30 br_30 wl_199 vdd gnd cell_6t
Xbit_r200_c30 bl_30 br_30 wl_200 vdd gnd cell_6t
Xbit_r201_c30 bl_30 br_30 wl_201 vdd gnd cell_6t
Xbit_r202_c30 bl_30 br_30 wl_202 vdd gnd cell_6t
Xbit_r203_c30 bl_30 br_30 wl_203 vdd gnd cell_6t
Xbit_r204_c30 bl_30 br_30 wl_204 vdd gnd cell_6t
Xbit_r205_c30 bl_30 br_30 wl_205 vdd gnd cell_6t
Xbit_r206_c30 bl_30 br_30 wl_206 vdd gnd cell_6t
Xbit_r207_c30 bl_30 br_30 wl_207 vdd gnd cell_6t
Xbit_r208_c30 bl_30 br_30 wl_208 vdd gnd cell_6t
Xbit_r209_c30 bl_30 br_30 wl_209 vdd gnd cell_6t
Xbit_r210_c30 bl_30 br_30 wl_210 vdd gnd cell_6t
Xbit_r211_c30 bl_30 br_30 wl_211 vdd gnd cell_6t
Xbit_r212_c30 bl_30 br_30 wl_212 vdd gnd cell_6t
Xbit_r213_c30 bl_30 br_30 wl_213 vdd gnd cell_6t
Xbit_r214_c30 bl_30 br_30 wl_214 vdd gnd cell_6t
Xbit_r215_c30 bl_30 br_30 wl_215 vdd gnd cell_6t
Xbit_r216_c30 bl_30 br_30 wl_216 vdd gnd cell_6t
Xbit_r217_c30 bl_30 br_30 wl_217 vdd gnd cell_6t
Xbit_r218_c30 bl_30 br_30 wl_218 vdd gnd cell_6t
Xbit_r219_c30 bl_30 br_30 wl_219 vdd gnd cell_6t
Xbit_r220_c30 bl_30 br_30 wl_220 vdd gnd cell_6t
Xbit_r221_c30 bl_30 br_30 wl_221 vdd gnd cell_6t
Xbit_r222_c30 bl_30 br_30 wl_222 vdd gnd cell_6t
Xbit_r223_c30 bl_30 br_30 wl_223 vdd gnd cell_6t
Xbit_r224_c30 bl_30 br_30 wl_224 vdd gnd cell_6t
Xbit_r225_c30 bl_30 br_30 wl_225 vdd gnd cell_6t
Xbit_r226_c30 bl_30 br_30 wl_226 vdd gnd cell_6t
Xbit_r227_c30 bl_30 br_30 wl_227 vdd gnd cell_6t
Xbit_r228_c30 bl_30 br_30 wl_228 vdd gnd cell_6t
Xbit_r229_c30 bl_30 br_30 wl_229 vdd gnd cell_6t
Xbit_r230_c30 bl_30 br_30 wl_230 vdd gnd cell_6t
Xbit_r231_c30 bl_30 br_30 wl_231 vdd gnd cell_6t
Xbit_r232_c30 bl_30 br_30 wl_232 vdd gnd cell_6t
Xbit_r233_c30 bl_30 br_30 wl_233 vdd gnd cell_6t
Xbit_r234_c30 bl_30 br_30 wl_234 vdd gnd cell_6t
Xbit_r235_c30 bl_30 br_30 wl_235 vdd gnd cell_6t
Xbit_r236_c30 bl_30 br_30 wl_236 vdd gnd cell_6t
Xbit_r237_c30 bl_30 br_30 wl_237 vdd gnd cell_6t
Xbit_r238_c30 bl_30 br_30 wl_238 vdd gnd cell_6t
Xbit_r239_c30 bl_30 br_30 wl_239 vdd gnd cell_6t
Xbit_r240_c30 bl_30 br_30 wl_240 vdd gnd cell_6t
Xbit_r241_c30 bl_30 br_30 wl_241 vdd gnd cell_6t
Xbit_r242_c30 bl_30 br_30 wl_242 vdd gnd cell_6t
Xbit_r243_c30 bl_30 br_30 wl_243 vdd gnd cell_6t
Xbit_r244_c30 bl_30 br_30 wl_244 vdd gnd cell_6t
Xbit_r245_c30 bl_30 br_30 wl_245 vdd gnd cell_6t
Xbit_r246_c30 bl_30 br_30 wl_246 vdd gnd cell_6t
Xbit_r247_c30 bl_30 br_30 wl_247 vdd gnd cell_6t
Xbit_r248_c30 bl_30 br_30 wl_248 vdd gnd cell_6t
Xbit_r249_c30 bl_30 br_30 wl_249 vdd gnd cell_6t
Xbit_r250_c30 bl_30 br_30 wl_250 vdd gnd cell_6t
Xbit_r251_c30 bl_30 br_30 wl_251 vdd gnd cell_6t
Xbit_r252_c30 bl_30 br_30 wl_252 vdd gnd cell_6t
Xbit_r253_c30 bl_30 br_30 wl_253 vdd gnd cell_6t
Xbit_r254_c30 bl_30 br_30 wl_254 vdd gnd cell_6t
Xbit_r255_c30 bl_30 br_30 wl_255 vdd gnd cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd cell_6t
Xbit_r1_c31 bl_31 br_31 wl_1 vdd gnd cell_6t
Xbit_r2_c31 bl_31 br_31 wl_2 vdd gnd cell_6t
Xbit_r3_c31 bl_31 br_31 wl_3 vdd gnd cell_6t
Xbit_r4_c31 bl_31 br_31 wl_4 vdd gnd cell_6t
Xbit_r5_c31 bl_31 br_31 wl_5 vdd gnd cell_6t
Xbit_r6_c31 bl_31 br_31 wl_6 vdd gnd cell_6t
Xbit_r7_c31 bl_31 br_31 wl_7 vdd gnd cell_6t
Xbit_r8_c31 bl_31 br_31 wl_8 vdd gnd cell_6t
Xbit_r9_c31 bl_31 br_31 wl_9 vdd gnd cell_6t
Xbit_r10_c31 bl_31 br_31 wl_10 vdd gnd cell_6t
Xbit_r11_c31 bl_31 br_31 wl_11 vdd gnd cell_6t
Xbit_r12_c31 bl_31 br_31 wl_12 vdd gnd cell_6t
Xbit_r13_c31 bl_31 br_31 wl_13 vdd gnd cell_6t
Xbit_r14_c31 bl_31 br_31 wl_14 vdd gnd cell_6t
Xbit_r15_c31 bl_31 br_31 wl_15 vdd gnd cell_6t
Xbit_r16_c31 bl_31 br_31 wl_16 vdd gnd cell_6t
Xbit_r17_c31 bl_31 br_31 wl_17 vdd gnd cell_6t
Xbit_r18_c31 bl_31 br_31 wl_18 vdd gnd cell_6t
Xbit_r19_c31 bl_31 br_31 wl_19 vdd gnd cell_6t
Xbit_r20_c31 bl_31 br_31 wl_20 vdd gnd cell_6t
Xbit_r21_c31 bl_31 br_31 wl_21 vdd gnd cell_6t
Xbit_r22_c31 bl_31 br_31 wl_22 vdd gnd cell_6t
Xbit_r23_c31 bl_31 br_31 wl_23 vdd gnd cell_6t
Xbit_r24_c31 bl_31 br_31 wl_24 vdd gnd cell_6t
Xbit_r25_c31 bl_31 br_31 wl_25 vdd gnd cell_6t
Xbit_r26_c31 bl_31 br_31 wl_26 vdd gnd cell_6t
Xbit_r27_c31 bl_31 br_31 wl_27 vdd gnd cell_6t
Xbit_r28_c31 bl_31 br_31 wl_28 vdd gnd cell_6t
Xbit_r29_c31 bl_31 br_31 wl_29 vdd gnd cell_6t
Xbit_r30_c31 bl_31 br_31 wl_30 vdd gnd cell_6t
Xbit_r31_c31 bl_31 br_31 wl_31 vdd gnd cell_6t
Xbit_r32_c31 bl_31 br_31 wl_32 vdd gnd cell_6t
Xbit_r33_c31 bl_31 br_31 wl_33 vdd gnd cell_6t
Xbit_r34_c31 bl_31 br_31 wl_34 vdd gnd cell_6t
Xbit_r35_c31 bl_31 br_31 wl_35 vdd gnd cell_6t
Xbit_r36_c31 bl_31 br_31 wl_36 vdd gnd cell_6t
Xbit_r37_c31 bl_31 br_31 wl_37 vdd gnd cell_6t
Xbit_r38_c31 bl_31 br_31 wl_38 vdd gnd cell_6t
Xbit_r39_c31 bl_31 br_31 wl_39 vdd gnd cell_6t
Xbit_r40_c31 bl_31 br_31 wl_40 vdd gnd cell_6t
Xbit_r41_c31 bl_31 br_31 wl_41 vdd gnd cell_6t
Xbit_r42_c31 bl_31 br_31 wl_42 vdd gnd cell_6t
Xbit_r43_c31 bl_31 br_31 wl_43 vdd gnd cell_6t
Xbit_r44_c31 bl_31 br_31 wl_44 vdd gnd cell_6t
Xbit_r45_c31 bl_31 br_31 wl_45 vdd gnd cell_6t
Xbit_r46_c31 bl_31 br_31 wl_46 vdd gnd cell_6t
Xbit_r47_c31 bl_31 br_31 wl_47 vdd gnd cell_6t
Xbit_r48_c31 bl_31 br_31 wl_48 vdd gnd cell_6t
Xbit_r49_c31 bl_31 br_31 wl_49 vdd gnd cell_6t
Xbit_r50_c31 bl_31 br_31 wl_50 vdd gnd cell_6t
Xbit_r51_c31 bl_31 br_31 wl_51 vdd gnd cell_6t
Xbit_r52_c31 bl_31 br_31 wl_52 vdd gnd cell_6t
Xbit_r53_c31 bl_31 br_31 wl_53 vdd gnd cell_6t
Xbit_r54_c31 bl_31 br_31 wl_54 vdd gnd cell_6t
Xbit_r55_c31 bl_31 br_31 wl_55 vdd gnd cell_6t
Xbit_r56_c31 bl_31 br_31 wl_56 vdd gnd cell_6t
Xbit_r57_c31 bl_31 br_31 wl_57 vdd gnd cell_6t
Xbit_r58_c31 bl_31 br_31 wl_58 vdd gnd cell_6t
Xbit_r59_c31 bl_31 br_31 wl_59 vdd gnd cell_6t
Xbit_r60_c31 bl_31 br_31 wl_60 vdd gnd cell_6t
Xbit_r61_c31 bl_31 br_31 wl_61 vdd gnd cell_6t
Xbit_r62_c31 bl_31 br_31 wl_62 vdd gnd cell_6t
Xbit_r63_c31 bl_31 br_31 wl_63 vdd gnd cell_6t
Xbit_r64_c31 bl_31 br_31 wl_64 vdd gnd cell_6t
Xbit_r65_c31 bl_31 br_31 wl_65 vdd gnd cell_6t
Xbit_r66_c31 bl_31 br_31 wl_66 vdd gnd cell_6t
Xbit_r67_c31 bl_31 br_31 wl_67 vdd gnd cell_6t
Xbit_r68_c31 bl_31 br_31 wl_68 vdd gnd cell_6t
Xbit_r69_c31 bl_31 br_31 wl_69 vdd gnd cell_6t
Xbit_r70_c31 bl_31 br_31 wl_70 vdd gnd cell_6t
Xbit_r71_c31 bl_31 br_31 wl_71 vdd gnd cell_6t
Xbit_r72_c31 bl_31 br_31 wl_72 vdd gnd cell_6t
Xbit_r73_c31 bl_31 br_31 wl_73 vdd gnd cell_6t
Xbit_r74_c31 bl_31 br_31 wl_74 vdd gnd cell_6t
Xbit_r75_c31 bl_31 br_31 wl_75 vdd gnd cell_6t
Xbit_r76_c31 bl_31 br_31 wl_76 vdd gnd cell_6t
Xbit_r77_c31 bl_31 br_31 wl_77 vdd gnd cell_6t
Xbit_r78_c31 bl_31 br_31 wl_78 vdd gnd cell_6t
Xbit_r79_c31 bl_31 br_31 wl_79 vdd gnd cell_6t
Xbit_r80_c31 bl_31 br_31 wl_80 vdd gnd cell_6t
Xbit_r81_c31 bl_31 br_31 wl_81 vdd gnd cell_6t
Xbit_r82_c31 bl_31 br_31 wl_82 vdd gnd cell_6t
Xbit_r83_c31 bl_31 br_31 wl_83 vdd gnd cell_6t
Xbit_r84_c31 bl_31 br_31 wl_84 vdd gnd cell_6t
Xbit_r85_c31 bl_31 br_31 wl_85 vdd gnd cell_6t
Xbit_r86_c31 bl_31 br_31 wl_86 vdd gnd cell_6t
Xbit_r87_c31 bl_31 br_31 wl_87 vdd gnd cell_6t
Xbit_r88_c31 bl_31 br_31 wl_88 vdd gnd cell_6t
Xbit_r89_c31 bl_31 br_31 wl_89 vdd gnd cell_6t
Xbit_r90_c31 bl_31 br_31 wl_90 vdd gnd cell_6t
Xbit_r91_c31 bl_31 br_31 wl_91 vdd gnd cell_6t
Xbit_r92_c31 bl_31 br_31 wl_92 vdd gnd cell_6t
Xbit_r93_c31 bl_31 br_31 wl_93 vdd gnd cell_6t
Xbit_r94_c31 bl_31 br_31 wl_94 vdd gnd cell_6t
Xbit_r95_c31 bl_31 br_31 wl_95 vdd gnd cell_6t
Xbit_r96_c31 bl_31 br_31 wl_96 vdd gnd cell_6t
Xbit_r97_c31 bl_31 br_31 wl_97 vdd gnd cell_6t
Xbit_r98_c31 bl_31 br_31 wl_98 vdd gnd cell_6t
Xbit_r99_c31 bl_31 br_31 wl_99 vdd gnd cell_6t
Xbit_r100_c31 bl_31 br_31 wl_100 vdd gnd cell_6t
Xbit_r101_c31 bl_31 br_31 wl_101 vdd gnd cell_6t
Xbit_r102_c31 bl_31 br_31 wl_102 vdd gnd cell_6t
Xbit_r103_c31 bl_31 br_31 wl_103 vdd gnd cell_6t
Xbit_r104_c31 bl_31 br_31 wl_104 vdd gnd cell_6t
Xbit_r105_c31 bl_31 br_31 wl_105 vdd gnd cell_6t
Xbit_r106_c31 bl_31 br_31 wl_106 vdd gnd cell_6t
Xbit_r107_c31 bl_31 br_31 wl_107 vdd gnd cell_6t
Xbit_r108_c31 bl_31 br_31 wl_108 vdd gnd cell_6t
Xbit_r109_c31 bl_31 br_31 wl_109 vdd gnd cell_6t
Xbit_r110_c31 bl_31 br_31 wl_110 vdd gnd cell_6t
Xbit_r111_c31 bl_31 br_31 wl_111 vdd gnd cell_6t
Xbit_r112_c31 bl_31 br_31 wl_112 vdd gnd cell_6t
Xbit_r113_c31 bl_31 br_31 wl_113 vdd gnd cell_6t
Xbit_r114_c31 bl_31 br_31 wl_114 vdd gnd cell_6t
Xbit_r115_c31 bl_31 br_31 wl_115 vdd gnd cell_6t
Xbit_r116_c31 bl_31 br_31 wl_116 vdd gnd cell_6t
Xbit_r117_c31 bl_31 br_31 wl_117 vdd gnd cell_6t
Xbit_r118_c31 bl_31 br_31 wl_118 vdd gnd cell_6t
Xbit_r119_c31 bl_31 br_31 wl_119 vdd gnd cell_6t
Xbit_r120_c31 bl_31 br_31 wl_120 vdd gnd cell_6t
Xbit_r121_c31 bl_31 br_31 wl_121 vdd gnd cell_6t
Xbit_r122_c31 bl_31 br_31 wl_122 vdd gnd cell_6t
Xbit_r123_c31 bl_31 br_31 wl_123 vdd gnd cell_6t
Xbit_r124_c31 bl_31 br_31 wl_124 vdd gnd cell_6t
Xbit_r125_c31 bl_31 br_31 wl_125 vdd gnd cell_6t
Xbit_r126_c31 bl_31 br_31 wl_126 vdd gnd cell_6t
Xbit_r127_c31 bl_31 br_31 wl_127 vdd gnd cell_6t
Xbit_r128_c31 bl_31 br_31 wl_128 vdd gnd cell_6t
Xbit_r129_c31 bl_31 br_31 wl_129 vdd gnd cell_6t
Xbit_r130_c31 bl_31 br_31 wl_130 vdd gnd cell_6t
Xbit_r131_c31 bl_31 br_31 wl_131 vdd gnd cell_6t
Xbit_r132_c31 bl_31 br_31 wl_132 vdd gnd cell_6t
Xbit_r133_c31 bl_31 br_31 wl_133 vdd gnd cell_6t
Xbit_r134_c31 bl_31 br_31 wl_134 vdd gnd cell_6t
Xbit_r135_c31 bl_31 br_31 wl_135 vdd gnd cell_6t
Xbit_r136_c31 bl_31 br_31 wl_136 vdd gnd cell_6t
Xbit_r137_c31 bl_31 br_31 wl_137 vdd gnd cell_6t
Xbit_r138_c31 bl_31 br_31 wl_138 vdd gnd cell_6t
Xbit_r139_c31 bl_31 br_31 wl_139 vdd gnd cell_6t
Xbit_r140_c31 bl_31 br_31 wl_140 vdd gnd cell_6t
Xbit_r141_c31 bl_31 br_31 wl_141 vdd gnd cell_6t
Xbit_r142_c31 bl_31 br_31 wl_142 vdd gnd cell_6t
Xbit_r143_c31 bl_31 br_31 wl_143 vdd gnd cell_6t
Xbit_r144_c31 bl_31 br_31 wl_144 vdd gnd cell_6t
Xbit_r145_c31 bl_31 br_31 wl_145 vdd gnd cell_6t
Xbit_r146_c31 bl_31 br_31 wl_146 vdd gnd cell_6t
Xbit_r147_c31 bl_31 br_31 wl_147 vdd gnd cell_6t
Xbit_r148_c31 bl_31 br_31 wl_148 vdd gnd cell_6t
Xbit_r149_c31 bl_31 br_31 wl_149 vdd gnd cell_6t
Xbit_r150_c31 bl_31 br_31 wl_150 vdd gnd cell_6t
Xbit_r151_c31 bl_31 br_31 wl_151 vdd gnd cell_6t
Xbit_r152_c31 bl_31 br_31 wl_152 vdd gnd cell_6t
Xbit_r153_c31 bl_31 br_31 wl_153 vdd gnd cell_6t
Xbit_r154_c31 bl_31 br_31 wl_154 vdd gnd cell_6t
Xbit_r155_c31 bl_31 br_31 wl_155 vdd gnd cell_6t
Xbit_r156_c31 bl_31 br_31 wl_156 vdd gnd cell_6t
Xbit_r157_c31 bl_31 br_31 wl_157 vdd gnd cell_6t
Xbit_r158_c31 bl_31 br_31 wl_158 vdd gnd cell_6t
Xbit_r159_c31 bl_31 br_31 wl_159 vdd gnd cell_6t
Xbit_r160_c31 bl_31 br_31 wl_160 vdd gnd cell_6t
Xbit_r161_c31 bl_31 br_31 wl_161 vdd gnd cell_6t
Xbit_r162_c31 bl_31 br_31 wl_162 vdd gnd cell_6t
Xbit_r163_c31 bl_31 br_31 wl_163 vdd gnd cell_6t
Xbit_r164_c31 bl_31 br_31 wl_164 vdd gnd cell_6t
Xbit_r165_c31 bl_31 br_31 wl_165 vdd gnd cell_6t
Xbit_r166_c31 bl_31 br_31 wl_166 vdd gnd cell_6t
Xbit_r167_c31 bl_31 br_31 wl_167 vdd gnd cell_6t
Xbit_r168_c31 bl_31 br_31 wl_168 vdd gnd cell_6t
Xbit_r169_c31 bl_31 br_31 wl_169 vdd gnd cell_6t
Xbit_r170_c31 bl_31 br_31 wl_170 vdd gnd cell_6t
Xbit_r171_c31 bl_31 br_31 wl_171 vdd gnd cell_6t
Xbit_r172_c31 bl_31 br_31 wl_172 vdd gnd cell_6t
Xbit_r173_c31 bl_31 br_31 wl_173 vdd gnd cell_6t
Xbit_r174_c31 bl_31 br_31 wl_174 vdd gnd cell_6t
Xbit_r175_c31 bl_31 br_31 wl_175 vdd gnd cell_6t
Xbit_r176_c31 bl_31 br_31 wl_176 vdd gnd cell_6t
Xbit_r177_c31 bl_31 br_31 wl_177 vdd gnd cell_6t
Xbit_r178_c31 bl_31 br_31 wl_178 vdd gnd cell_6t
Xbit_r179_c31 bl_31 br_31 wl_179 vdd gnd cell_6t
Xbit_r180_c31 bl_31 br_31 wl_180 vdd gnd cell_6t
Xbit_r181_c31 bl_31 br_31 wl_181 vdd gnd cell_6t
Xbit_r182_c31 bl_31 br_31 wl_182 vdd gnd cell_6t
Xbit_r183_c31 bl_31 br_31 wl_183 vdd gnd cell_6t
Xbit_r184_c31 bl_31 br_31 wl_184 vdd gnd cell_6t
Xbit_r185_c31 bl_31 br_31 wl_185 vdd gnd cell_6t
Xbit_r186_c31 bl_31 br_31 wl_186 vdd gnd cell_6t
Xbit_r187_c31 bl_31 br_31 wl_187 vdd gnd cell_6t
Xbit_r188_c31 bl_31 br_31 wl_188 vdd gnd cell_6t
Xbit_r189_c31 bl_31 br_31 wl_189 vdd gnd cell_6t
Xbit_r190_c31 bl_31 br_31 wl_190 vdd gnd cell_6t
Xbit_r191_c31 bl_31 br_31 wl_191 vdd gnd cell_6t
Xbit_r192_c31 bl_31 br_31 wl_192 vdd gnd cell_6t
Xbit_r193_c31 bl_31 br_31 wl_193 vdd gnd cell_6t
Xbit_r194_c31 bl_31 br_31 wl_194 vdd gnd cell_6t
Xbit_r195_c31 bl_31 br_31 wl_195 vdd gnd cell_6t
Xbit_r196_c31 bl_31 br_31 wl_196 vdd gnd cell_6t
Xbit_r197_c31 bl_31 br_31 wl_197 vdd gnd cell_6t
Xbit_r198_c31 bl_31 br_31 wl_198 vdd gnd cell_6t
Xbit_r199_c31 bl_31 br_31 wl_199 vdd gnd cell_6t
Xbit_r200_c31 bl_31 br_31 wl_200 vdd gnd cell_6t
Xbit_r201_c31 bl_31 br_31 wl_201 vdd gnd cell_6t
Xbit_r202_c31 bl_31 br_31 wl_202 vdd gnd cell_6t
Xbit_r203_c31 bl_31 br_31 wl_203 vdd gnd cell_6t
Xbit_r204_c31 bl_31 br_31 wl_204 vdd gnd cell_6t
Xbit_r205_c31 bl_31 br_31 wl_205 vdd gnd cell_6t
Xbit_r206_c31 bl_31 br_31 wl_206 vdd gnd cell_6t
Xbit_r207_c31 bl_31 br_31 wl_207 vdd gnd cell_6t
Xbit_r208_c31 bl_31 br_31 wl_208 vdd gnd cell_6t
Xbit_r209_c31 bl_31 br_31 wl_209 vdd gnd cell_6t
Xbit_r210_c31 bl_31 br_31 wl_210 vdd gnd cell_6t
Xbit_r211_c31 bl_31 br_31 wl_211 vdd gnd cell_6t
Xbit_r212_c31 bl_31 br_31 wl_212 vdd gnd cell_6t
Xbit_r213_c31 bl_31 br_31 wl_213 vdd gnd cell_6t
Xbit_r214_c31 bl_31 br_31 wl_214 vdd gnd cell_6t
Xbit_r215_c31 bl_31 br_31 wl_215 vdd gnd cell_6t
Xbit_r216_c31 bl_31 br_31 wl_216 vdd gnd cell_6t
Xbit_r217_c31 bl_31 br_31 wl_217 vdd gnd cell_6t
Xbit_r218_c31 bl_31 br_31 wl_218 vdd gnd cell_6t
Xbit_r219_c31 bl_31 br_31 wl_219 vdd gnd cell_6t
Xbit_r220_c31 bl_31 br_31 wl_220 vdd gnd cell_6t
Xbit_r221_c31 bl_31 br_31 wl_221 vdd gnd cell_6t
Xbit_r222_c31 bl_31 br_31 wl_222 vdd gnd cell_6t
Xbit_r223_c31 bl_31 br_31 wl_223 vdd gnd cell_6t
Xbit_r224_c31 bl_31 br_31 wl_224 vdd gnd cell_6t
Xbit_r225_c31 bl_31 br_31 wl_225 vdd gnd cell_6t
Xbit_r226_c31 bl_31 br_31 wl_226 vdd gnd cell_6t
Xbit_r227_c31 bl_31 br_31 wl_227 vdd gnd cell_6t
Xbit_r228_c31 bl_31 br_31 wl_228 vdd gnd cell_6t
Xbit_r229_c31 bl_31 br_31 wl_229 vdd gnd cell_6t
Xbit_r230_c31 bl_31 br_31 wl_230 vdd gnd cell_6t
Xbit_r231_c31 bl_31 br_31 wl_231 vdd gnd cell_6t
Xbit_r232_c31 bl_31 br_31 wl_232 vdd gnd cell_6t
Xbit_r233_c31 bl_31 br_31 wl_233 vdd gnd cell_6t
Xbit_r234_c31 bl_31 br_31 wl_234 vdd gnd cell_6t
Xbit_r235_c31 bl_31 br_31 wl_235 vdd gnd cell_6t
Xbit_r236_c31 bl_31 br_31 wl_236 vdd gnd cell_6t
Xbit_r237_c31 bl_31 br_31 wl_237 vdd gnd cell_6t
Xbit_r238_c31 bl_31 br_31 wl_238 vdd gnd cell_6t
Xbit_r239_c31 bl_31 br_31 wl_239 vdd gnd cell_6t
Xbit_r240_c31 bl_31 br_31 wl_240 vdd gnd cell_6t
Xbit_r241_c31 bl_31 br_31 wl_241 vdd gnd cell_6t
Xbit_r242_c31 bl_31 br_31 wl_242 vdd gnd cell_6t
Xbit_r243_c31 bl_31 br_31 wl_243 vdd gnd cell_6t
Xbit_r244_c31 bl_31 br_31 wl_244 vdd gnd cell_6t
Xbit_r245_c31 bl_31 br_31 wl_245 vdd gnd cell_6t
Xbit_r246_c31 bl_31 br_31 wl_246 vdd gnd cell_6t
Xbit_r247_c31 bl_31 br_31 wl_247 vdd gnd cell_6t
Xbit_r248_c31 bl_31 br_31 wl_248 vdd gnd cell_6t
Xbit_r249_c31 bl_31 br_31 wl_249 vdd gnd cell_6t
Xbit_r250_c31 bl_31 br_31 wl_250 vdd gnd cell_6t
Xbit_r251_c31 bl_31 br_31 wl_251 vdd gnd cell_6t
Xbit_r252_c31 bl_31 br_31 wl_252 vdd gnd cell_6t
Xbit_r253_c31 bl_31 br_31 wl_253 vdd gnd cell_6t
Xbit_r254_c31 bl_31 br_31 wl_254 vdd gnd cell_6t
Xbit_r255_c31 bl_31 br_31 wl_255 vdd gnd cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd cell_6t
Xbit_r1_c32 bl_32 br_32 wl_1 vdd gnd cell_6t
Xbit_r2_c32 bl_32 br_32 wl_2 vdd gnd cell_6t
Xbit_r3_c32 bl_32 br_32 wl_3 vdd gnd cell_6t
Xbit_r4_c32 bl_32 br_32 wl_4 vdd gnd cell_6t
Xbit_r5_c32 bl_32 br_32 wl_5 vdd gnd cell_6t
Xbit_r6_c32 bl_32 br_32 wl_6 vdd gnd cell_6t
Xbit_r7_c32 bl_32 br_32 wl_7 vdd gnd cell_6t
Xbit_r8_c32 bl_32 br_32 wl_8 vdd gnd cell_6t
Xbit_r9_c32 bl_32 br_32 wl_9 vdd gnd cell_6t
Xbit_r10_c32 bl_32 br_32 wl_10 vdd gnd cell_6t
Xbit_r11_c32 bl_32 br_32 wl_11 vdd gnd cell_6t
Xbit_r12_c32 bl_32 br_32 wl_12 vdd gnd cell_6t
Xbit_r13_c32 bl_32 br_32 wl_13 vdd gnd cell_6t
Xbit_r14_c32 bl_32 br_32 wl_14 vdd gnd cell_6t
Xbit_r15_c32 bl_32 br_32 wl_15 vdd gnd cell_6t
Xbit_r16_c32 bl_32 br_32 wl_16 vdd gnd cell_6t
Xbit_r17_c32 bl_32 br_32 wl_17 vdd gnd cell_6t
Xbit_r18_c32 bl_32 br_32 wl_18 vdd gnd cell_6t
Xbit_r19_c32 bl_32 br_32 wl_19 vdd gnd cell_6t
Xbit_r20_c32 bl_32 br_32 wl_20 vdd gnd cell_6t
Xbit_r21_c32 bl_32 br_32 wl_21 vdd gnd cell_6t
Xbit_r22_c32 bl_32 br_32 wl_22 vdd gnd cell_6t
Xbit_r23_c32 bl_32 br_32 wl_23 vdd gnd cell_6t
Xbit_r24_c32 bl_32 br_32 wl_24 vdd gnd cell_6t
Xbit_r25_c32 bl_32 br_32 wl_25 vdd gnd cell_6t
Xbit_r26_c32 bl_32 br_32 wl_26 vdd gnd cell_6t
Xbit_r27_c32 bl_32 br_32 wl_27 vdd gnd cell_6t
Xbit_r28_c32 bl_32 br_32 wl_28 vdd gnd cell_6t
Xbit_r29_c32 bl_32 br_32 wl_29 vdd gnd cell_6t
Xbit_r30_c32 bl_32 br_32 wl_30 vdd gnd cell_6t
Xbit_r31_c32 bl_32 br_32 wl_31 vdd gnd cell_6t
Xbit_r32_c32 bl_32 br_32 wl_32 vdd gnd cell_6t
Xbit_r33_c32 bl_32 br_32 wl_33 vdd gnd cell_6t
Xbit_r34_c32 bl_32 br_32 wl_34 vdd gnd cell_6t
Xbit_r35_c32 bl_32 br_32 wl_35 vdd gnd cell_6t
Xbit_r36_c32 bl_32 br_32 wl_36 vdd gnd cell_6t
Xbit_r37_c32 bl_32 br_32 wl_37 vdd gnd cell_6t
Xbit_r38_c32 bl_32 br_32 wl_38 vdd gnd cell_6t
Xbit_r39_c32 bl_32 br_32 wl_39 vdd gnd cell_6t
Xbit_r40_c32 bl_32 br_32 wl_40 vdd gnd cell_6t
Xbit_r41_c32 bl_32 br_32 wl_41 vdd gnd cell_6t
Xbit_r42_c32 bl_32 br_32 wl_42 vdd gnd cell_6t
Xbit_r43_c32 bl_32 br_32 wl_43 vdd gnd cell_6t
Xbit_r44_c32 bl_32 br_32 wl_44 vdd gnd cell_6t
Xbit_r45_c32 bl_32 br_32 wl_45 vdd gnd cell_6t
Xbit_r46_c32 bl_32 br_32 wl_46 vdd gnd cell_6t
Xbit_r47_c32 bl_32 br_32 wl_47 vdd gnd cell_6t
Xbit_r48_c32 bl_32 br_32 wl_48 vdd gnd cell_6t
Xbit_r49_c32 bl_32 br_32 wl_49 vdd gnd cell_6t
Xbit_r50_c32 bl_32 br_32 wl_50 vdd gnd cell_6t
Xbit_r51_c32 bl_32 br_32 wl_51 vdd gnd cell_6t
Xbit_r52_c32 bl_32 br_32 wl_52 vdd gnd cell_6t
Xbit_r53_c32 bl_32 br_32 wl_53 vdd gnd cell_6t
Xbit_r54_c32 bl_32 br_32 wl_54 vdd gnd cell_6t
Xbit_r55_c32 bl_32 br_32 wl_55 vdd gnd cell_6t
Xbit_r56_c32 bl_32 br_32 wl_56 vdd gnd cell_6t
Xbit_r57_c32 bl_32 br_32 wl_57 vdd gnd cell_6t
Xbit_r58_c32 bl_32 br_32 wl_58 vdd gnd cell_6t
Xbit_r59_c32 bl_32 br_32 wl_59 vdd gnd cell_6t
Xbit_r60_c32 bl_32 br_32 wl_60 vdd gnd cell_6t
Xbit_r61_c32 bl_32 br_32 wl_61 vdd gnd cell_6t
Xbit_r62_c32 bl_32 br_32 wl_62 vdd gnd cell_6t
Xbit_r63_c32 bl_32 br_32 wl_63 vdd gnd cell_6t
Xbit_r64_c32 bl_32 br_32 wl_64 vdd gnd cell_6t
Xbit_r65_c32 bl_32 br_32 wl_65 vdd gnd cell_6t
Xbit_r66_c32 bl_32 br_32 wl_66 vdd gnd cell_6t
Xbit_r67_c32 bl_32 br_32 wl_67 vdd gnd cell_6t
Xbit_r68_c32 bl_32 br_32 wl_68 vdd gnd cell_6t
Xbit_r69_c32 bl_32 br_32 wl_69 vdd gnd cell_6t
Xbit_r70_c32 bl_32 br_32 wl_70 vdd gnd cell_6t
Xbit_r71_c32 bl_32 br_32 wl_71 vdd gnd cell_6t
Xbit_r72_c32 bl_32 br_32 wl_72 vdd gnd cell_6t
Xbit_r73_c32 bl_32 br_32 wl_73 vdd gnd cell_6t
Xbit_r74_c32 bl_32 br_32 wl_74 vdd gnd cell_6t
Xbit_r75_c32 bl_32 br_32 wl_75 vdd gnd cell_6t
Xbit_r76_c32 bl_32 br_32 wl_76 vdd gnd cell_6t
Xbit_r77_c32 bl_32 br_32 wl_77 vdd gnd cell_6t
Xbit_r78_c32 bl_32 br_32 wl_78 vdd gnd cell_6t
Xbit_r79_c32 bl_32 br_32 wl_79 vdd gnd cell_6t
Xbit_r80_c32 bl_32 br_32 wl_80 vdd gnd cell_6t
Xbit_r81_c32 bl_32 br_32 wl_81 vdd gnd cell_6t
Xbit_r82_c32 bl_32 br_32 wl_82 vdd gnd cell_6t
Xbit_r83_c32 bl_32 br_32 wl_83 vdd gnd cell_6t
Xbit_r84_c32 bl_32 br_32 wl_84 vdd gnd cell_6t
Xbit_r85_c32 bl_32 br_32 wl_85 vdd gnd cell_6t
Xbit_r86_c32 bl_32 br_32 wl_86 vdd gnd cell_6t
Xbit_r87_c32 bl_32 br_32 wl_87 vdd gnd cell_6t
Xbit_r88_c32 bl_32 br_32 wl_88 vdd gnd cell_6t
Xbit_r89_c32 bl_32 br_32 wl_89 vdd gnd cell_6t
Xbit_r90_c32 bl_32 br_32 wl_90 vdd gnd cell_6t
Xbit_r91_c32 bl_32 br_32 wl_91 vdd gnd cell_6t
Xbit_r92_c32 bl_32 br_32 wl_92 vdd gnd cell_6t
Xbit_r93_c32 bl_32 br_32 wl_93 vdd gnd cell_6t
Xbit_r94_c32 bl_32 br_32 wl_94 vdd gnd cell_6t
Xbit_r95_c32 bl_32 br_32 wl_95 vdd gnd cell_6t
Xbit_r96_c32 bl_32 br_32 wl_96 vdd gnd cell_6t
Xbit_r97_c32 bl_32 br_32 wl_97 vdd gnd cell_6t
Xbit_r98_c32 bl_32 br_32 wl_98 vdd gnd cell_6t
Xbit_r99_c32 bl_32 br_32 wl_99 vdd gnd cell_6t
Xbit_r100_c32 bl_32 br_32 wl_100 vdd gnd cell_6t
Xbit_r101_c32 bl_32 br_32 wl_101 vdd gnd cell_6t
Xbit_r102_c32 bl_32 br_32 wl_102 vdd gnd cell_6t
Xbit_r103_c32 bl_32 br_32 wl_103 vdd gnd cell_6t
Xbit_r104_c32 bl_32 br_32 wl_104 vdd gnd cell_6t
Xbit_r105_c32 bl_32 br_32 wl_105 vdd gnd cell_6t
Xbit_r106_c32 bl_32 br_32 wl_106 vdd gnd cell_6t
Xbit_r107_c32 bl_32 br_32 wl_107 vdd gnd cell_6t
Xbit_r108_c32 bl_32 br_32 wl_108 vdd gnd cell_6t
Xbit_r109_c32 bl_32 br_32 wl_109 vdd gnd cell_6t
Xbit_r110_c32 bl_32 br_32 wl_110 vdd gnd cell_6t
Xbit_r111_c32 bl_32 br_32 wl_111 vdd gnd cell_6t
Xbit_r112_c32 bl_32 br_32 wl_112 vdd gnd cell_6t
Xbit_r113_c32 bl_32 br_32 wl_113 vdd gnd cell_6t
Xbit_r114_c32 bl_32 br_32 wl_114 vdd gnd cell_6t
Xbit_r115_c32 bl_32 br_32 wl_115 vdd gnd cell_6t
Xbit_r116_c32 bl_32 br_32 wl_116 vdd gnd cell_6t
Xbit_r117_c32 bl_32 br_32 wl_117 vdd gnd cell_6t
Xbit_r118_c32 bl_32 br_32 wl_118 vdd gnd cell_6t
Xbit_r119_c32 bl_32 br_32 wl_119 vdd gnd cell_6t
Xbit_r120_c32 bl_32 br_32 wl_120 vdd gnd cell_6t
Xbit_r121_c32 bl_32 br_32 wl_121 vdd gnd cell_6t
Xbit_r122_c32 bl_32 br_32 wl_122 vdd gnd cell_6t
Xbit_r123_c32 bl_32 br_32 wl_123 vdd gnd cell_6t
Xbit_r124_c32 bl_32 br_32 wl_124 vdd gnd cell_6t
Xbit_r125_c32 bl_32 br_32 wl_125 vdd gnd cell_6t
Xbit_r126_c32 bl_32 br_32 wl_126 vdd gnd cell_6t
Xbit_r127_c32 bl_32 br_32 wl_127 vdd gnd cell_6t
Xbit_r128_c32 bl_32 br_32 wl_128 vdd gnd cell_6t
Xbit_r129_c32 bl_32 br_32 wl_129 vdd gnd cell_6t
Xbit_r130_c32 bl_32 br_32 wl_130 vdd gnd cell_6t
Xbit_r131_c32 bl_32 br_32 wl_131 vdd gnd cell_6t
Xbit_r132_c32 bl_32 br_32 wl_132 vdd gnd cell_6t
Xbit_r133_c32 bl_32 br_32 wl_133 vdd gnd cell_6t
Xbit_r134_c32 bl_32 br_32 wl_134 vdd gnd cell_6t
Xbit_r135_c32 bl_32 br_32 wl_135 vdd gnd cell_6t
Xbit_r136_c32 bl_32 br_32 wl_136 vdd gnd cell_6t
Xbit_r137_c32 bl_32 br_32 wl_137 vdd gnd cell_6t
Xbit_r138_c32 bl_32 br_32 wl_138 vdd gnd cell_6t
Xbit_r139_c32 bl_32 br_32 wl_139 vdd gnd cell_6t
Xbit_r140_c32 bl_32 br_32 wl_140 vdd gnd cell_6t
Xbit_r141_c32 bl_32 br_32 wl_141 vdd gnd cell_6t
Xbit_r142_c32 bl_32 br_32 wl_142 vdd gnd cell_6t
Xbit_r143_c32 bl_32 br_32 wl_143 vdd gnd cell_6t
Xbit_r144_c32 bl_32 br_32 wl_144 vdd gnd cell_6t
Xbit_r145_c32 bl_32 br_32 wl_145 vdd gnd cell_6t
Xbit_r146_c32 bl_32 br_32 wl_146 vdd gnd cell_6t
Xbit_r147_c32 bl_32 br_32 wl_147 vdd gnd cell_6t
Xbit_r148_c32 bl_32 br_32 wl_148 vdd gnd cell_6t
Xbit_r149_c32 bl_32 br_32 wl_149 vdd gnd cell_6t
Xbit_r150_c32 bl_32 br_32 wl_150 vdd gnd cell_6t
Xbit_r151_c32 bl_32 br_32 wl_151 vdd gnd cell_6t
Xbit_r152_c32 bl_32 br_32 wl_152 vdd gnd cell_6t
Xbit_r153_c32 bl_32 br_32 wl_153 vdd gnd cell_6t
Xbit_r154_c32 bl_32 br_32 wl_154 vdd gnd cell_6t
Xbit_r155_c32 bl_32 br_32 wl_155 vdd gnd cell_6t
Xbit_r156_c32 bl_32 br_32 wl_156 vdd gnd cell_6t
Xbit_r157_c32 bl_32 br_32 wl_157 vdd gnd cell_6t
Xbit_r158_c32 bl_32 br_32 wl_158 vdd gnd cell_6t
Xbit_r159_c32 bl_32 br_32 wl_159 vdd gnd cell_6t
Xbit_r160_c32 bl_32 br_32 wl_160 vdd gnd cell_6t
Xbit_r161_c32 bl_32 br_32 wl_161 vdd gnd cell_6t
Xbit_r162_c32 bl_32 br_32 wl_162 vdd gnd cell_6t
Xbit_r163_c32 bl_32 br_32 wl_163 vdd gnd cell_6t
Xbit_r164_c32 bl_32 br_32 wl_164 vdd gnd cell_6t
Xbit_r165_c32 bl_32 br_32 wl_165 vdd gnd cell_6t
Xbit_r166_c32 bl_32 br_32 wl_166 vdd gnd cell_6t
Xbit_r167_c32 bl_32 br_32 wl_167 vdd gnd cell_6t
Xbit_r168_c32 bl_32 br_32 wl_168 vdd gnd cell_6t
Xbit_r169_c32 bl_32 br_32 wl_169 vdd gnd cell_6t
Xbit_r170_c32 bl_32 br_32 wl_170 vdd gnd cell_6t
Xbit_r171_c32 bl_32 br_32 wl_171 vdd gnd cell_6t
Xbit_r172_c32 bl_32 br_32 wl_172 vdd gnd cell_6t
Xbit_r173_c32 bl_32 br_32 wl_173 vdd gnd cell_6t
Xbit_r174_c32 bl_32 br_32 wl_174 vdd gnd cell_6t
Xbit_r175_c32 bl_32 br_32 wl_175 vdd gnd cell_6t
Xbit_r176_c32 bl_32 br_32 wl_176 vdd gnd cell_6t
Xbit_r177_c32 bl_32 br_32 wl_177 vdd gnd cell_6t
Xbit_r178_c32 bl_32 br_32 wl_178 vdd gnd cell_6t
Xbit_r179_c32 bl_32 br_32 wl_179 vdd gnd cell_6t
Xbit_r180_c32 bl_32 br_32 wl_180 vdd gnd cell_6t
Xbit_r181_c32 bl_32 br_32 wl_181 vdd gnd cell_6t
Xbit_r182_c32 bl_32 br_32 wl_182 vdd gnd cell_6t
Xbit_r183_c32 bl_32 br_32 wl_183 vdd gnd cell_6t
Xbit_r184_c32 bl_32 br_32 wl_184 vdd gnd cell_6t
Xbit_r185_c32 bl_32 br_32 wl_185 vdd gnd cell_6t
Xbit_r186_c32 bl_32 br_32 wl_186 vdd gnd cell_6t
Xbit_r187_c32 bl_32 br_32 wl_187 vdd gnd cell_6t
Xbit_r188_c32 bl_32 br_32 wl_188 vdd gnd cell_6t
Xbit_r189_c32 bl_32 br_32 wl_189 vdd gnd cell_6t
Xbit_r190_c32 bl_32 br_32 wl_190 vdd gnd cell_6t
Xbit_r191_c32 bl_32 br_32 wl_191 vdd gnd cell_6t
Xbit_r192_c32 bl_32 br_32 wl_192 vdd gnd cell_6t
Xbit_r193_c32 bl_32 br_32 wl_193 vdd gnd cell_6t
Xbit_r194_c32 bl_32 br_32 wl_194 vdd gnd cell_6t
Xbit_r195_c32 bl_32 br_32 wl_195 vdd gnd cell_6t
Xbit_r196_c32 bl_32 br_32 wl_196 vdd gnd cell_6t
Xbit_r197_c32 bl_32 br_32 wl_197 vdd gnd cell_6t
Xbit_r198_c32 bl_32 br_32 wl_198 vdd gnd cell_6t
Xbit_r199_c32 bl_32 br_32 wl_199 vdd gnd cell_6t
Xbit_r200_c32 bl_32 br_32 wl_200 vdd gnd cell_6t
Xbit_r201_c32 bl_32 br_32 wl_201 vdd gnd cell_6t
Xbit_r202_c32 bl_32 br_32 wl_202 vdd gnd cell_6t
Xbit_r203_c32 bl_32 br_32 wl_203 vdd gnd cell_6t
Xbit_r204_c32 bl_32 br_32 wl_204 vdd gnd cell_6t
Xbit_r205_c32 bl_32 br_32 wl_205 vdd gnd cell_6t
Xbit_r206_c32 bl_32 br_32 wl_206 vdd gnd cell_6t
Xbit_r207_c32 bl_32 br_32 wl_207 vdd gnd cell_6t
Xbit_r208_c32 bl_32 br_32 wl_208 vdd gnd cell_6t
Xbit_r209_c32 bl_32 br_32 wl_209 vdd gnd cell_6t
Xbit_r210_c32 bl_32 br_32 wl_210 vdd gnd cell_6t
Xbit_r211_c32 bl_32 br_32 wl_211 vdd gnd cell_6t
Xbit_r212_c32 bl_32 br_32 wl_212 vdd gnd cell_6t
Xbit_r213_c32 bl_32 br_32 wl_213 vdd gnd cell_6t
Xbit_r214_c32 bl_32 br_32 wl_214 vdd gnd cell_6t
Xbit_r215_c32 bl_32 br_32 wl_215 vdd gnd cell_6t
Xbit_r216_c32 bl_32 br_32 wl_216 vdd gnd cell_6t
Xbit_r217_c32 bl_32 br_32 wl_217 vdd gnd cell_6t
Xbit_r218_c32 bl_32 br_32 wl_218 vdd gnd cell_6t
Xbit_r219_c32 bl_32 br_32 wl_219 vdd gnd cell_6t
Xbit_r220_c32 bl_32 br_32 wl_220 vdd gnd cell_6t
Xbit_r221_c32 bl_32 br_32 wl_221 vdd gnd cell_6t
Xbit_r222_c32 bl_32 br_32 wl_222 vdd gnd cell_6t
Xbit_r223_c32 bl_32 br_32 wl_223 vdd gnd cell_6t
Xbit_r224_c32 bl_32 br_32 wl_224 vdd gnd cell_6t
Xbit_r225_c32 bl_32 br_32 wl_225 vdd gnd cell_6t
Xbit_r226_c32 bl_32 br_32 wl_226 vdd gnd cell_6t
Xbit_r227_c32 bl_32 br_32 wl_227 vdd gnd cell_6t
Xbit_r228_c32 bl_32 br_32 wl_228 vdd gnd cell_6t
Xbit_r229_c32 bl_32 br_32 wl_229 vdd gnd cell_6t
Xbit_r230_c32 bl_32 br_32 wl_230 vdd gnd cell_6t
Xbit_r231_c32 bl_32 br_32 wl_231 vdd gnd cell_6t
Xbit_r232_c32 bl_32 br_32 wl_232 vdd gnd cell_6t
Xbit_r233_c32 bl_32 br_32 wl_233 vdd gnd cell_6t
Xbit_r234_c32 bl_32 br_32 wl_234 vdd gnd cell_6t
Xbit_r235_c32 bl_32 br_32 wl_235 vdd gnd cell_6t
Xbit_r236_c32 bl_32 br_32 wl_236 vdd gnd cell_6t
Xbit_r237_c32 bl_32 br_32 wl_237 vdd gnd cell_6t
Xbit_r238_c32 bl_32 br_32 wl_238 vdd gnd cell_6t
Xbit_r239_c32 bl_32 br_32 wl_239 vdd gnd cell_6t
Xbit_r240_c32 bl_32 br_32 wl_240 vdd gnd cell_6t
Xbit_r241_c32 bl_32 br_32 wl_241 vdd gnd cell_6t
Xbit_r242_c32 bl_32 br_32 wl_242 vdd gnd cell_6t
Xbit_r243_c32 bl_32 br_32 wl_243 vdd gnd cell_6t
Xbit_r244_c32 bl_32 br_32 wl_244 vdd gnd cell_6t
Xbit_r245_c32 bl_32 br_32 wl_245 vdd gnd cell_6t
Xbit_r246_c32 bl_32 br_32 wl_246 vdd gnd cell_6t
Xbit_r247_c32 bl_32 br_32 wl_247 vdd gnd cell_6t
Xbit_r248_c32 bl_32 br_32 wl_248 vdd gnd cell_6t
Xbit_r249_c32 bl_32 br_32 wl_249 vdd gnd cell_6t
Xbit_r250_c32 bl_32 br_32 wl_250 vdd gnd cell_6t
Xbit_r251_c32 bl_32 br_32 wl_251 vdd gnd cell_6t
Xbit_r252_c32 bl_32 br_32 wl_252 vdd gnd cell_6t
Xbit_r253_c32 bl_32 br_32 wl_253 vdd gnd cell_6t
Xbit_r254_c32 bl_32 br_32 wl_254 vdd gnd cell_6t
Xbit_r255_c32 bl_32 br_32 wl_255 vdd gnd cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd cell_6t
Xbit_r1_c33 bl_33 br_33 wl_1 vdd gnd cell_6t
Xbit_r2_c33 bl_33 br_33 wl_2 vdd gnd cell_6t
Xbit_r3_c33 bl_33 br_33 wl_3 vdd gnd cell_6t
Xbit_r4_c33 bl_33 br_33 wl_4 vdd gnd cell_6t
Xbit_r5_c33 bl_33 br_33 wl_5 vdd gnd cell_6t
Xbit_r6_c33 bl_33 br_33 wl_6 vdd gnd cell_6t
Xbit_r7_c33 bl_33 br_33 wl_7 vdd gnd cell_6t
Xbit_r8_c33 bl_33 br_33 wl_8 vdd gnd cell_6t
Xbit_r9_c33 bl_33 br_33 wl_9 vdd gnd cell_6t
Xbit_r10_c33 bl_33 br_33 wl_10 vdd gnd cell_6t
Xbit_r11_c33 bl_33 br_33 wl_11 vdd gnd cell_6t
Xbit_r12_c33 bl_33 br_33 wl_12 vdd gnd cell_6t
Xbit_r13_c33 bl_33 br_33 wl_13 vdd gnd cell_6t
Xbit_r14_c33 bl_33 br_33 wl_14 vdd gnd cell_6t
Xbit_r15_c33 bl_33 br_33 wl_15 vdd gnd cell_6t
Xbit_r16_c33 bl_33 br_33 wl_16 vdd gnd cell_6t
Xbit_r17_c33 bl_33 br_33 wl_17 vdd gnd cell_6t
Xbit_r18_c33 bl_33 br_33 wl_18 vdd gnd cell_6t
Xbit_r19_c33 bl_33 br_33 wl_19 vdd gnd cell_6t
Xbit_r20_c33 bl_33 br_33 wl_20 vdd gnd cell_6t
Xbit_r21_c33 bl_33 br_33 wl_21 vdd gnd cell_6t
Xbit_r22_c33 bl_33 br_33 wl_22 vdd gnd cell_6t
Xbit_r23_c33 bl_33 br_33 wl_23 vdd gnd cell_6t
Xbit_r24_c33 bl_33 br_33 wl_24 vdd gnd cell_6t
Xbit_r25_c33 bl_33 br_33 wl_25 vdd gnd cell_6t
Xbit_r26_c33 bl_33 br_33 wl_26 vdd gnd cell_6t
Xbit_r27_c33 bl_33 br_33 wl_27 vdd gnd cell_6t
Xbit_r28_c33 bl_33 br_33 wl_28 vdd gnd cell_6t
Xbit_r29_c33 bl_33 br_33 wl_29 vdd gnd cell_6t
Xbit_r30_c33 bl_33 br_33 wl_30 vdd gnd cell_6t
Xbit_r31_c33 bl_33 br_33 wl_31 vdd gnd cell_6t
Xbit_r32_c33 bl_33 br_33 wl_32 vdd gnd cell_6t
Xbit_r33_c33 bl_33 br_33 wl_33 vdd gnd cell_6t
Xbit_r34_c33 bl_33 br_33 wl_34 vdd gnd cell_6t
Xbit_r35_c33 bl_33 br_33 wl_35 vdd gnd cell_6t
Xbit_r36_c33 bl_33 br_33 wl_36 vdd gnd cell_6t
Xbit_r37_c33 bl_33 br_33 wl_37 vdd gnd cell_6t
Xbit_r38_c33 bl_33 br_33 wl_38 vdd gnd cell_6t
Xbit_r39_c33 bl_33 br_33 wl_39 vdd gnd cell_6t
Xbit_r40_c33 bl_33 br_33 wl_40 vdd gnd cell_6t
Xbit_r41_c33 bl_33 br_33 wl_41 vdd gnd cell_6t
Xbit_r42_c33 bl_33 br_33 wl_42 vdd gnd cell_6t
Xbit_r43_c33 bl_33 br_33 wl_43 vdd gnd cell_6t
Xbit_r44_c33 bl_33 br_33 wl_44 vdd gnd cell_6t
Xbit_r45_c33 bl_33 br_33 wl_45 vdd gnd cell_6t
Xbit_r46_c33 bl_33 br_33 wl_46 vdd gnd cell_6t
Xbit_r47_c33 bl_33 br_33 wl_47 vdd gnd cell_6t
Xbit_r48_c33 bl_33 br_33 wl_48 vdd gnd cell_6t
Xbit_r49_c33 bl_33 br_33 wl_49 vdd gnd cell_6t
Xbit_r50_c33 bl_33 br_33 wl_50 vdd gnd cell_6t
Xbit_r51_c33 bl_33 br_33 wl_51 vdd gnd cell_6t
Xbit_r52_c33 bl_33 br_33 wl_52 vdd gnd cell_6t
Xbit_r53_c33 bl_33 br_33 wl_53 vdd gnd cell_6t
Xbit_r54_c33 bl_33 br_33 wl_54 vdd gnd cell_6t
Xbit_r55_c33 bl_33 br_33 wl_55 vdd gnd cell_6t
Xbit_r56_c33 bl_33 br_33 wl_56 vdd gnd cell_6t
Xbit_r57_c33 bl_33 br_33 wl_57 vdd gnd cell_6t
Xbit_r58_c33 bl_33 br_33 wl_58 vdd gnd cell_6t
Xbit_r59_c33 bl_33 br_33 wl_59 vdd gnd cell_6t
Xbit_r60_c33 bl_33 br_33 wl_60 vdd gnd cell_6t
Xbit_r61_c33 bl_33 br_33 wl_61 vdd gnd cell_6t
Xbit_r62_c33 bl_33 br_33 wl_62 vdd gnd cell_6t
Xbit_r63_c33 bl_33 br_33 wl_63 vdd gnd cell_6t
Xbit_r64_c33 bl_33 br_33 wl_64 vdd gnd cell_6t
Xbit_r65_c33 bl_33 br_33 wl_65 vdd gnd cell_6t
Xbit_r66_c33 bl_33 br_33 wl_66 vdd gnd cell_6t
Xbit_r67_c33 bl_33 br_33 wl_67 vdd gnd cell_6t
Xbit_r68_c33 bl_33 br_33 wl_68 vdd gnd cell_6t
Xbit_r69_c33 bl_33 br_33 wl_69 vdd gnd cell_6t
Xbit_r70_c33 bl_33 br_33 wl_70 vdd gnd cell_6t
Xbit_r71_c33 bl_33 br_33 wl_71 vdd gnd cell_6t
Xbit_r72_c33 bl_33 br_33 wl_72 vdd gnd cell_6t
Xbit_r73_c33 bl_33 br_33 wl_73 vdd gnd cell_6t
Xbit_r74_c33 bl_33 br_33 wl_74 vdd gnd cell_6t
Xbit_r75_c33 bl_33 br_33 wl_75 vdd gnd cell_6t
Xbit_r76_c33 bl_33 br_33 wl_76 vdd gnd cell_6t
Xbit_r77_c33 bl_33 br_33 wl_77 vdd gnd cell_6t
Xbit_r78_c33 bl_33 br_33 wl_78 vdd gnd cell_6t
Xbit_r79_c33 bl_33 br_33 wl_79 vdd gnd cell_6t
Xbit_r80_c33 bl_33 br_33 wl_80 vdd gnd cell_6t
Xbit_r81_c33 bl_33 br_33 wl_81 vdd gnd cell_6t
Xbit_r82_c33 bl_33 br_33 wl_82 vdd gnd cell_6t
Xbit_r83_c33 bl_33 br_33 wl_83 vdd gnd cell_6t
Xbit_r84_c33 bl_33 br_33 wl_84 vdd gnd cell_6t
Xbit_r85_c33 bl_33 br_33 wl_85 vdd gnd cell_6t
Xbit_r86_c33 bl_33 br_33 wl_86 vdd gnd cell_6t
Xbit_r87_c33 bl_33 br_33 wl_87 vdd gnd cell_6t
Xbit_r88_c33 bl_33 br_33 wl_88 vdd gnd cell_6t
Xbit_r89_c33 bl_33 br_33 wl_89 vdd gnd cell_6t
Xbit_r90_c33 bl_33 br_33 wl_90 vdd gnd cell_6t
Xbit_r91_c33 bl_33 br_33 wl_91 vdd gnd cell_6t
Xbit_r92_c33 bl_33 br_33 wl_92 vdd gnd cell_6t
Xbit_r93_c33 bl_33 br_33 wl_93 vdd gnd cell_6t
Xbit_r94_c33 bl_33 br_33 wl_94 vdd gnd cell_6t
Xbit_r95_c33 bl_33 br_33 wl_95 vdd gnd cell_6t
Xbit_r96_c33 bl_33 br_33 wl_96 vdd gnd cell_6t
Xbit_r97_c33 bl_33 br_33 wl_97 vdd gnd cell_6t
Xbit_r98_c33 bl_33 br_33 wl_98 vdd gnd cell_6t
Xbit_r99_c33 bl_33 br_33 wl_99 vdd gnd cell_6t
Xbit_r100_c33 bl_33 br_33 wl_100 vdd gnd cell_6t
Xbit_r101_c33 bl_33 br_33 wl_101 vdd gnd cell_6t
Xbit_r102_c33 bl_33 br_33 wl_102 vdd gnd cell_6t
Xbit_r103_c33 bl_33 br_33 wl_103 vdd gnd cell_6t
Xbit_r104_c33 bl_33 br_33 wl_104 vdd gnd cell_6t
Xbit_r105_c33 bl_33 br_33 wl_105 vdd gnd cell_6t
Xbit_r106_c33 bl_33 br_33 wl_106 vdd gnd cell_6t
Xbit_r107_c33 bl_33 br_33 wl_107 vdd gnd cell_6t
Xbit_r108_c33 bl_33 br_33 wl_108 vdd gnd cell_6t
Xbit_r109_c33 bl_33 br_33 wl_109 vdd gnd cell_6t
Xbit_r110_c33 bl_33 br_33 wl_110 vdd gnd cell_6t
Xbit_r111_c33 bl_33 br_33 wl_111 vdd gnd cell_6t
Xbit_r112_c33 bl_33 br_33 wl_112 vdd gnd cell_6t
Xbit_r113_c33 bl_33 br_33 wl_113 vdd gnd cell_6t
Xbit_r114_c33 bl_33 br_33 wl_114 vdd gnd cell_6t
Xbit_r115_c33 bl_33 br_33 wl_115 vdd gnd cell_6t
Xbit_r116_c33 bl_33 br_33 wl_116 vdd gnd cell_6t
Xbit_r117_c33 bl_33 br_33 wl_117 vdd gnd cell_6t
Xbit_r118_c33 bl_33 br_33 wl_118 vdd gnd cell_6t
Xbit_r119_c33 bl_33 br_33 wl_119 vdd gnd cell_6t
Xbit_r120_c33 bl_33 br_33 wl_120 vdd gnd cell_6t
Xbit_r121_c33 bl_33 br_33 wl_121 vdd gnd cell_6t
Xbit_r122_c33 bl_33 br_33 wl_122 vdd gnd cell_6t
Xbit_r123_c33 bl_33 br_33 wl_123 vdd gnd cell_6t
Xbit_r124_c33 bl_33 br_33 wl_124 vdd gnd cell_6t
Xbit_r125_c33 bl_33 br_33 wl_125 vdd gnd cell_6t
Xbit_r126_c33 bl_33 br_33 wl_126 vdd gnd cell_6t
Xbit_r127_c33 bl_33 br_33 wl_127 vdd gnd cell_6t
Xbit_r128_c33 bl_33 br_33 wl_128 vdd gnd cell_6t
Xbit_r129_c33 bl_33 br_33 wl_129 vdd gnd cell_6t
Xbit_r130_c33 bl_33 br_33 wl_130 vdd gnd cell_6t
Xbit_r131_c33 bl_33 br_33 wl_131 vdd gnd cell_6t
Xbit_r132_c33 bl_33 br_33 wl_132 vdd gnd cell_6t
Xbit_r133_c33 bl_33 br_33 wl_133 vdd gnd cell_6t
Xbit_r134_c33 bl_33 br_33 wl_134 vdd gnd cell_6t
Xbit_r135_c33 bl_33 br_33 wl_135 vdd gnd cell_6t
Xbit_r136_c33 bl_33 br_33 wl_136 vdd gnd cell_6t
Xbit_r137_c33 bl_33 br_33 wl_137 vdd gnd cell_6t
Xbit_r138_c33 bl_33 br_33 wl_138 vdd gnd cell_6t
Xbit_r139_c33 bl_33 br_33 wl_139 vdd gnd cell_6t
Xbit_r140_c33 bl_33 br_33 wl_140 vdd gnd cell_6t
Xbit_r141_c33 bl_33 br_33 wl_141 vdd gnd cell_6t
Xbit_r142_c33 bl_33 br_33 wl_142 vdd gnd cell_6t
Xbit_r143_c33 bl_33 br_33 wl_143 vdd gnd cell_6t
Xbit_r144_c33 bl_33 br_33 wl_144 vdd gnd cell_6t
Xbit_r145_c33 bl_33 br_33 wl_145 vdd gnd cell_6t
Xbit_r146_c33 bl_33 br_33 wl_146 vdd gnd cell_6t
Xbit_r147_c33 bl_33 br_33 wl_147 vdd gnd cell_6t
Xbit_r148_c33 bl_33 br_33 wl_148 vdd gnd cell_6t
Xbit_r149_c33 bl_33 br_33 wl_149 vdd gnd cell_6t
Xbit_r150_c33 bl_33 br_33 wl_150 vdd gnd cell_6t
Xbit_r151_c33 bl_33 br_33 wl_151 vdd gnd cell_6t
Xbit_r152_c33 bl_33 br_33 wl_152 vdd gnd cell_6t
Xbit_r153_c33 bl_33 br_33 wl_153 vdd gnd cell_6t
Xbit_r154_c33 bl_33 br_33 wl_154 vdd gnd cell_6t
Xbit_r155_c33 bl_33 br_33 wl_155 vdd gnd cell_6t
Xbit_r156_c33 bl_33 br_33 wl_156 vdd gnd cell_6t
Xbit_r157_c33 bl_33 br_33 wl_157 vdd gnd cell_6t
Xbit_r158_c33 bl_33 br_33 wl_158 vdd gnd cell_6t
Xbit_r159_c33 bl_33 br_33 wl_159 vdd gnd cell_6t
Xbit_r160_c33 bl_33 br_33 wl_160 vdd gnd cell_6t
Xbit_r161_c33 bl_33 br_33 wl_161 vdd gnd cell_6t
Xbit_r162_c33 bl_33 br_33 wl_162 vdd gnd cell_6t
Xbit_r163_c33 bl_33 br_33 wl_163 vdd gnd cell_6t
Xbit_r164_c33 bl_33 br_33 wl_164 vdd gnd cell_6t
Xbit_r165_c33 bl_33 br_33 wl_165 vdd gnd cell_6t
Xbit_r166_c33 bl_33 br_33 wl_166 vdd gnd cell_6t
Xbit_r167_c33 bl_33 br_33 wl_167 vdd gnd cell_6t
Xbit_r168_c33 bl_33 br_33 wl_168 vdd gnd cell_6t
Xbit_r169_c33 bl_33 br_33 wl_169 vdd gnd cell_6t
Xbit_r170_c33 bl_33 br_33 wl_170 vdd gnd cell_6t
Xbit_r171_c33 bl_33 br_33 wl_171 vdd gnd cell_6t
Xbit_r172_c33 bl_33 br_33 wl_172 vdd gnd cell_6t
Xbit_r173_c33 bl_33 br_33 wl_173 vdd gnd cell_6t
Xbit_r174_c33 bl_33 br_33 wl_174 vdd gnd cell_6t
Xbit_r175_c33 bl_33 br_33 wl_175 vdd gnd cell_6t
Xbit_r176_c33 bl_33 br_33 wl_176 vdd gnd cell_6t
Xbit_r177_c33 bl_33 br_33 wl_177 vdd gnd cell_6t
Xbit_r178_c33 bl_33 br_33 wl_178 vdd gnd cell_6t
Xbit_r179_c33 bl_33 br_33 wl_179 vdd gnd cell_6t
Xbit_r180_c33 bl_33 br_33 wl_180 vdd gnd cell_6t
Xbit_r181_c33 bl_33 br_33 wl_181 vdd gnd cell_6t
Xbit_r182_c33 bl_33 br_33 wl_182 vdd gnd cell_6t
Xbit_r183_c33 bl_33 br_33 wl_183 vdd gnd cell_6t
Xbit_r184_c33 bl_33 br_33 wl_184 vdd gnd cell_6t
Xbit_r185_c33 bl_33 br_33 wl_185 vdd gnd cell_6t
Xbit_r186_c33 bl_33 br_33 wl_186 vdd gnd cell_6t
Xbit_r187_c33 bl_33 br_33 wl_187 vdd gnd cell_6t
Xbit_r188_c33 bl_33 br_33 wl_188 vdd gnd cell_6t
Xbit_r189_c33 bl_33 br_33 wl_189 vdd gnd cell_6t
Xbit_r190_c33 bl_33 br_33 wl_190 vdd gnd cell_6t
Xbit_r191_c33 bl_33 br_33 wl_191 vdd gnd cell_6t
Xbit_r192_c33 bl_33 br_33 wl_192 vdd gnd cell_6t
Xbit_r193_c33 bl_33 br_33 wl_193 vdd gnd cell_6t
Xbit_r194_c33 bl_33 br_33 wl_194 vdd gnd cell_6t
Xbit_r195_c33 bl_33 br_33 wl_195 vdd gnd cell_6t
Xbit_r196_c33 bl_33 br_33 wl_196 vdd gnd cell_6t
Xbit_r197_c33 bl_33 br_33 wl_197 vdd gnd cell_6t
Xbit_r198_c33 bl_33 br_33 wl_198 vdd gnd cell_6t
Xbit_r199_c33 bl_33 br_33 wl_199 vdd gnd cell_6t
Xbit_r200_c33 bl_33 br_33 wl_200 vdd gnd cell_6t
Xbit_r201_c33 bl_33 br_33 wl_201 vdd gnd cell_6t
Xbit_r202_c33 bl_33 br_33 wl_202 vdd gnd cell_6t
Xbit_r203_c33 bl_33 br_33 wl_203 vdd gnd cell_6t
Xbit_r204_c33 bl_33 br_33 wl_204 vdd gnd cell_6t
Xbit_r205_c33 bl_33 br_33 wl_205 vdd gnd cell_6t
Xbit_r206_c33 bl_33 br_33 wl_206 vdd gnd cell_6t
Xbit_r207_c33 bl_33 br_33 wl_207 vdd gnd cell_6t
Xbit_r208_c33 bl_33 br_33 wl_208 vdd gnd cell_6t
Xbit_r209_c33 bl_33 br_33 wl_209 vdd gnd cell_6t
Xbit_r210_c33 bl_33 br_33 wl_210 vdd gnd cell_6t
Xbit_r211_c33 bl_33 br_33 wl_211 vdd gnd cell_6t
Xbit_r212_c33 bl_33 br_33 wl_212 vdd gnd cell_6t
Xbit_r213_c33 bl_33 br_33 wl_213 vdd gnd cell_6t
Xbit_r214_c33 bl_33 br_33 wl_214 vdd gnd cell_6t
Xbit_r215_c33 bl_33 br_33 wl_215 vdd gnd cell_6t
Xbit_r216_c33 bl_33 br_33 wl_216 vdd gnd cell_6t
Xbit_r217_c33 bl_33 br_33 wl_217 vdd gnd cell_6t
Xbit_r218_c33 bl_33 br_33 wl_218 vdd gnd cell_6t
Xbit_r219_c33 bl_33 br_33 wl_219 vdd gnd cell_6t
Xbit_r220_c33 bl_33 br_33 wl_220 vdd gnd cell_6t
Xbit_r221_c33 bl_33 br_33 wl_221 vdd gnd cell_6t
Xbit_r222_c33 bl_33 br_33 wl_222 vdd gnd cell_6t
Xbit_r223_c33 bl_33 br_33 wl_223 vdd gnd cell_6t
Xbit_r224_c33 bl_33 br_33 wl_224 vdd gnd cell_6t
Xbit_r225_c33 bl_33 br_33 wl_225 vdd gnd cell_6t
Xbit_r226_c33 bl_33 br_33 wl_226 vdd gnd cell_6t
Xbit_r227_c33 bl_33 br_33 wl_227 vdd gnd cell_6t
Xbit_r228_c33 bl_33 br_33 wl_228 vdd gnd cell_6t
Xbit_r229_c33 bl_33 br_33 wl_229 vdd gnd cell_6t
Xbit_r230_c33 bl_33 br_33 wl_230 vdd gnd cell_6t
Xbit_r231_c33 bl_33 br_33 wl_231 vdd gnd cell_6t
Xbit_r232_c33 bl_33 br_33 wl_232 vdd gnd cell_6t
Xbit_r233_c33 bl_33 br_33 wl_233 vdd gnd cell_6t
Xbit_r234_c33 bl_33 br_33 wl_234 vdd gnd cell_6t
Xbit_r235_c33 bl_33 br_33 wl_235 vdd gnd cell_6t
Xbit_r236_c33 bl_33 br_33 wl_236 vdd gnd cell_6t
Xbit_r237_c33 bl_33 br_33 wl_237 vdd gnd cell_6t
Xbit_r238_c33 bl_33 br_33 wl_238 vdd gnd cell_6t
Xbit_r239_c33 bl_33 br_33 wl_239 vdd gnd cell_6t
Xbit_r240_c33 bl_33 br_33 wl_240 vdd gnd cell_6t
Xbit_r241_c33 bl_33 br_33 wl_241 vdd gnd cell_6t
Xbit_r242_c33 bl_33 br_33 wl_242 vdd gnd cell_6t
Xbit_r243_c33 bl_33 br_33 wl_243 vdd gnd cell_6t
Xbit_r244_c33 bl_33 br_33 wl_244 vdd gnd cell_6t
Xbit_r245_c33 bl_33 br_33 wl_245 vdd gnd cell_6t
Xbit_r246_c33 bl_33 br_33 wl_246 vdd gnd cell_6t
Xbit_r247_c33 bl_33 br_33 wl_247 vdd gnd cell_6t
Xbit_r248_c33 bl_33 br_33 wl_248 vdd gnd cell_6t
Xbit_r249_c33 bl_33 br_33 wl_249 vdd gnd cell_6t
Xbit_r250_c33 bl_33 br_33 wl_250 vdd gnd cell_6t
Xbit_r251_c33 bl_33 br_33 wl_251 vdd gnd cell_6t
Xbit_r252_c33 bl_33 br_33 wl_252 vdd gnd cell_6t
Xbit_r253_c33 bl_33 br_33 wl_253 vdd gnd cell_6t
Xbit_r254_c33 bl_33 br_33 wl_254 vdd gnd cell_6t
Xbit_r255_c33 bl_33 br_33 wl_255 vdd gnd cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd cell_6t
Xbit_r1_c34 bl_34 br_34 wl_1 vdd gnd cell_6t
Xbit_r2_c34 bl_34 br_34 wl_2 vdd gnd cell_6t
Xbit_r3_c34 bl_34 br_34 wl_3 vdd gnd cell_6t
Xbit_r4_c34 bl_34 br_34 wl_4 vdd gnd cell_6t
Xbit_r5_c34 bl_34 br_34 wl_5 vdd gnd cell_6t
Xbit_r6_c34 bl_34 br_34 wl_6 vdd gnd cell_6t
Xbit_r7_c34 bl_34 br_34 wl_7 vdd gnd cell_6t
Xbit_r8_c34 bl_34 br_34 wl_8 vdd gnd cell_6t
Xbit_r9_c34 bl_34 br_34 wl_9 vdd gnd cell_6t
Xbit_r10_c34 bl_34 br_34 wl_10 vdd gnd cell_6t
Xbit_r11_c34 bl_34 br_34 wl_11 vdd gnd cell_6t
Xbit_r12_c34 bl_34 br_34 wl_12 vdd gnd cell_6t
Xbit_r13_c34 bl_34 br_34 wl_13 vdd gnd cell_6t
Xbit_r14_c34 bl_34 br_34 wl_14 vdd gnd cell_6t
Xbit_r15_c34 bl_34 br_34 wl_15 vdd gnd cell_6t
Xbit_r16_c34 bl_34 br_34 wl_16 vdd gnd cell_6t
Xbit_r17_c34 bl_34 br_34 wl_17 vdd gnd cell_6t
Xbit_r18_c34 bl_34 br_34 wl_18 vdd gnd cell_6t
Xbit_r19_c34 bl_34 br_34 wl_19 vdd gnd cell_6t
Xbit_r20_c34 bl_34 br_34 wl_20 vdd gnd cell_6t
Xbit_r21_c34 bl_34 br_34 wl_21 vdd gnd cell_6t
Xbit_r22_c34 bl_34 br_34 wl_22 vdd gnd cell_6t
Xbit_r23_c34 bl_34 br_34 wl_23 vdd gnd cell_6t
Xbit_r24_c34 bl_34 br_34 wl_24 vdd gnd cell_6t
Xbit_r25_c34 bl_34 br_34 wl_25 vdd gnd cell_6t
Xbit_r26_c34 bl_34 br_34 wl_26 vdd gnd cell_6t
Xbit_r27_c34 bl_34 br_34 wl_27 vdd gnd cell_6t
Xbit_r28_c34 bl_34 br_34 wl_28 vdd gnd cell_6t
Xbit_r29_c34 bl_34 br_34 wl_29 vdd gnd cell_6t
Xbit_r30_c34 bl_34 br_34 wl_30 vdd gnd cell_6t
Xbit_r31_c34 bl_34 br_34 wl_31 vdd gnd cell_6t
Xbit_r32_c34 bl_34 br_34 wl_32 vdd gnd cell_6t
Xbit_r33_c34 bl_34 br_34 wl_33 vdd gnd cell_6t
Xbit_r34_c34 bl_34 br_34 wl_34 vdd gnd cell_6t
Xbit_r35_c34 bl_34 br_34 wl_35 vdd gnd cell_6t
Xbit_r36_c34 bl_34 br_34 wl_36 vdd gnd cell_6t
Xbit_r37_c34 bl_34 br_34 wl_37 vdd gnd cell_6t
Xbit_r38_c34 bl_34 br_34 wl_38 vdd gnd cell_6t
Xbit_r39_c34 bl_34 br_34 wl_39 vdd gnd cell_6t
Xbit_r40_c34 bl_34 br_34 wl_40 vdd gnd cell_6t
Xbit_r41_c34 bl_34 br_34 wl_41 vdd gnd cell_6t
Xbit_r42_c34 bl_34 br_34 wl_42 vdd gnd cell_6t
Xbit_r43_c34 bl_34 br_34 wl_43 vdd gnd cell_6t
Xbit_r44_c34 bl_34 br_34 wl_44 vdd gnd cell_6t
Xbit_r45_c34 bl_34 br_34 wl_45 vdd gnd cell_6t
Xbit_r46_c34 bl_34 br_34 wl_46 vdd gnd cell_6t
Xbit_r47_c34 bl_34 br_34 wl_47 vdd gnd cell_6t
Xbit_r48_c34 bl_34 br_34 wl_48 vdd gnd cell_6t
Xbit_r49_c34 bl_34 br_34 wl_49 vdd gnd cell_6t
Xbit_r50_c34 bl_34 br_34 wl_50 vdd gnd cell_6t
Xbit_r51_c34 bl_34 br_34 wl_51 vdd gnd cell_6t
Xbit_r52_c34 bl_34 br_34 wl_52 vdd gnd cell_6t
Xbit_r53_c34 bl_34 br_34 wl_53 vdd gnd cell_6t
Xbit_r54_c34 bl_34 br_34 wl_54 vdd gnd cell_6t
Xbit_r55_c34 bl_34 br_34 wl_55 vdd gnd cell_6t
Xbit_r56_c34 bl_34 br_34 wl_56 vdd gnd cell_6t
Xbit_r57_c34 bl_34 br_34 wl_57 vdd gnd cell_6t
Xbit_r58_c34 bl_34 br_34 wl_58 vdd gnd cell_6t
Xbit_r59_c34 bl_34 br_34 wl_59 vdd gnd cell_6t
Xbit_r60_c34 bl_34 br_34 wl_60 vdd gnd cell_6t
Xbit_r61_c34 bl_34 br_34 wl_61 vdd gnd cell_6t
Xbit_r62_c34 bl_34 br_34 wl_62 vdd gnd cell_6t
Xbit_r63_c34 bl_34 br_34 wl_63 vdd gnd cell_6t
Xbit_r64_c34 bl_34 br_34 wl_64 vdd gnd cell_6t
Xbit_r65_c34 bl_34 br_34 wl_65 vdd gnd cell_6t
Xbit_r66_c34 bl_34 br_34 wl_66 vdd gnd cell_6t
Xbit_r67_c34 bl_34 br_34 wl_67 vdd gnd cell_6t
Xbit_r68_c34 bl_34 br_34 wl_68 vdd gnd cell_6t
Xbit_r69_c34 bl_34 br_34 wl_69 vdd gnd cell_6t
Xbit_r70_c34 bl_34 br_34 wl_70 vdd gnd cell_6t
Xbit_r71_c34 bl_34 br_34 wl_71 vdd gnd cell_6t
Xbit_r72_c34 bl_34 br_34 wl_72 vdd gnd cell_6t
Xbit_r73_c34 bl_34 br_34 wl_73 vdd gnd cell_6t
Xbit_r74_c34 bl_34 br_34 wl_74 vdd gnd cell_6t
Xbit_r75_c34 bl_34 br_34 wl_75 vdd gnd cell_6t
Xbit_r76_c34 bl_34 br_34 wl_76 vdd gnd cell_6t
Xbit_r77_c34 bl_34 br_34 wl_77 vdd gnd cell_6t
Xbit_r78_c34 bl_34 br_34 wl_78 vdd gnd cell_6t
Xbit_r79_c34 bl_34 br_34 wl_79 vdd gnd cell_6t
Xbit_r80_c34 bl_34 br_34 wl_80 vdd gnd cell_6t
Xbit_r81_c34 bl_34 br_34 wl_81 vdd gnd cell_6t
Xbit_r82_c34 bl_34 br_34 wl_82 vdd gnd cell_6t
Xbit_r83_c34 bl_34 br_34 wl_83 vdd gnd cell_6t
Xbit_r84_c34 bl_34 br_34 wl_84 vdd gnd cell_6t
Xbit_r85_c34 bl_34 br_34 wl_85 vdd gnd cell_6t
Xbit_r86_c34 bl_34 br_34 wl_86 vdd gnd cell_6t
Xbit_r87_c34 bl_34 br_34 wl_87 vdd gnd cell_6t
Xbit_r88_c34 bl_34 br_34 wl_88 vdd gnd cell_6t
Xbit_r89_c34 bl_34 br_34 wl_89 vdd gnd cell_6t
Xbit_r90_c34 bl_34 br_34 wl_90 vdd gnd cell_6t
Xbit_r91_c34 bl_34 br_34 wl_91 vdd gnd cell_6t
Xbit_r92_c34 bl_34 br_34 wl_92 vdd gnd cell_6t
Xbit_r93_c34 bl_34 br_34 wl_93 vdd gnd cell_6t
Xbit_r94_c34 bl_34 br_34 wl_94 vdd gnd cell_6t
Xbit_r95_c34 bl_34 br_34 wl_95 vdd gnd cell_6t
Xbit_r96_c34 bl_34 br_34 wl_96 vdd gnd cell_6t
Xbit_r97_c34 bl_34 br_34 wl_97 vdd gnd cell_6t
Xbit_r98_c34 bl_34 br_34 wl_98 vdd gnd cell_6t
Xbit_r99_c34 bl_34 br_34 wl_99 vdd gnd cell_6t
Xbit_r100_c34 bl_34 br_34 wl_100 vdd gnd cell_6t
Xbit_r101_c34 bl_34 br_34 wl_101 vdd gnd cell_6t
Xbit_r102_c34 bl_34 br_34 wl_102 vdd gnd cell_6t
Xbit_r103_c34 bl_34 br_34 wl_103 vdd gnd cell_6t
Xbit_r104_c34 bl_34 br_34 wl_104 vdd gnd cell_6t
Xbit_r105_c34 bl_34 br_34 wl_105 vdd gnd cell_6t
Xbit_r106_c34 bl_34 br_34 wl_106 vdd gnd cell_6t
Xbit_r107_c34 bl_34 br_34 wl_107 vdd gnd cell_6t
Xbit_r108_c34 bl_34 br_34 wl_108 vdd gnd cell_6t
Xbit_r109_c34 bl_34 br_34 wl_109 vdd gnd cell_6t
Xbit_r110_c34 bl_34 br_34 wl_110 vdd gnd cell_6t
Xbit_r111_c34 bl_34 br_34 wl_111 vdd gnd cell_6t
Xbit_r112_c34 bl_34 br_34 wl_112 vdd gnd cell_6t
Xbit_r113_c34 bl_34 br_34 wl_113 vdd gnd cell_6t
Xbit_r114_c34 bl_34 br_34 wl_114 vdd gnd cell_6t
Xbit_r115_c34 bl_34 br_34 wl_115 vdd gnd cell_6t
Xbit_r116_c34 bl_34 br_34 wl_116 vdd gnd cell_6t
Xbit_r117_c34 bl_34 br_34 wl_117 vdd gnd cell_6t
Xbit_r118_c34 bl_34 br_34 wl_118 vdd gnd cell_6t
Xbit_r119_c34 bl_34 br_34 wl_119 vdd gnd cell_6t
Xbit_r120_c34 bl_34 br_34 wl_120 vdd gnd cell_6t
Xbit_r121_c34 bl_34 br_34 wl_121 vdd gnd cell_6t
Xbit_r122_c34 bl_34 br_34 wl_122 vdd gnd cell_6t
Xbit_r123_c34 bl_34 br_34 wl_123 vdd gnd cell_6t
Xbit_r124_c34 bl_34 br_34 wl_124 vdd gnd cell_6t
Xbit_r125_c34 bl_34 br_34 wl_125 vdd gnd cell_6t
Xbit_r126_c34 bl_34 br_34 wl_126 vdd gnd cell_6t
Xbit_r127_c34 bl_34 br_34 wl_127 vdd gnd cell_6t
Xbit_r128_c34 bl_34 br_34 wl_128 vdd gnd cell_6t
Xbit_r129_c34 bl_34 br_34 wl_129 vdd gnd cell_6t
Xbit_r130_c34 bl_34 br_34 wl_130 vdd gnd cell_6t
Xbit_r131_c34 bl_34 br_34 wl_131 vdd gnd cell_6t
Xbit_r132_c34 bl_34 br_34 wl_132 vdd gnd cell_6t
Xbit_r133_c34 bl_34 br_34 wl_133 vdd gnd cell_6t
Xbit_r134_c34 bl_34 br_34 wl_134 vdd gnd cell_6t
Xbit_r135_c34 bl_34 br_34 wl_135 vdd gnd cell_6t
Xbit_r136_c34 bl_34 br_34 wl_136 vdd gnd cell_6t
Xbit_r137_c34 bl_34 br_34 wl_137 vdd gnd cell_6t
Xbit_r138_c34 bl_34 br_34 wl_138 vdd gnd cell_6t
Xbit_r139_c34 bl_34 br_34 wl_139 vdd gnd cell_6t
Xbit_r140_c34 bl_34 br_34 wl_140 vdd gnd cell_6t
Xbit_r141_c34 bl_34 br_34 wl_141 vdd gnd cell_6t
Xbit_r142_c34 bl_34 br_34 wl_142 vdd gnd cell_6t
Xbit_r143_c34 bl_34 br_34 wl_143 vdd gnd cell_6t
Xbit_r144_c34 bl_34 br_34 wl_144 vdd gnd cell_6t
Xbit_r145_c34 bl_34 br_34 wl_145 vdd gnd cell_6t
Xbit_r146_c34 bl_34 br_34 wl_146 vdd gnd cell_6t
Xbit_r147_c34 bl_34 br_34 wl_147 vdd gnd cell_6t
Xbit_r148_c34 bl_34 br_34 wl_148 vdd gnd cell_6t
Xbit_r149_c34 bl_34 br_34 wl_149 vdd gnd cell_6t
Xbit_r150_c34 bl_34 br_34 wl_150 vdd gnd cell_6t
Xbit_r151_c34 bl_34 br_34 wl_151 vdd gnd cell_6t
Xbit_r152_c34 bl_34 br_34 wl_152 vdd gnd cell_6t
Xbit_r153_c34 bl_34 br_34 wl_153 vdd gnd cell_6t
Xbit_r154_c34 bl_34 br_34 wl_154 vdd gnd cell_6t
Xbit_r155_c34 bl_34 br_34 wl_155 vdd gnd cell_6t
Xbit_r156_c34 bl_34 br_34 wl_156 vdd gnd cell_6t
Xbit_r157_c34 bl_34 br_34 wl_157 vdd gnd cell_6t
Xbit_r158_c34 bl_34 br_34 wl_158 vdd gnd cell_6t
Xbit_r159_c34 bl_34 br_34 wl_159 vdd gnd cell_6t
Xbit_r160_c34 bl_34 br_34 wl_160 vdd gnd cell_6t
Xbit_r161_c34 bl_34 br_34 wl_161 vdd gnd cell_6t
Xbit_r162_c34 bl_34 br_34 wl_162 vdd gnd cell_6t
Xbit_r163_c34 bl_34 br_34 wl_163 vdd gnd cell_6t
Xbit_r164_c34 bl_34 br_34 wl_164 vdd gnd cell_6t
Xbit_r165_c34 bl_34 br_34 wl_165 vdd gnd cell_6t
Xbit_r166_c34 bl_34 br_34 wl_166 vdd gnd cell_6t
Xbit_r167_c34 bl_34 br_34 wl_167 vdd gnd cell_6t
Xbit_r168_c34 bl_34 br_34 wl_168 vdd gnd cell_6t
Xbit_r169_c34 bl_34 br_34 wl_169 vdd gnd cell_6t
Xbit_r170_c34 bl_34 br_34 wl_170 vdd gnd cell_6t
Xbit_r171_c34 bl_34 br_34 wl_171 vdd gnd cell_6t
Xbit_r172_c34 bl_34 br_34 wl_172 vdd gnd cell_6t
Xbit_r173_c34 bl_34 br_34 wl_173 vdd gnd cell_6t
Xbit_r174_c34 bl_34 br_34 wl_174 vdd gnd cell_6t
Xbit_r175_c34 bl_34 br_34 wl_175 vdd gnd cell_6t
Xbit_r176_c34 bl_34 br_34 wl_176 vdd gnd cell_6t
Xbit_r177_c34 bl_34 br_34 wl_177 vdd gnd cell_6t
Xbit_r178_c34 bl_34 br_34 wl_178 vdd gnd cell_6t
Xbit_r179_c34 bl_34 br_34 wl_179 vdd gnd cell_6t
Xbit_r180_c34 bl_34 br_34 wl_180 vdd gnd cell_6t
Xbit_r181_c34 bl_34 br_34 wl_181 vdd gnd cell_6t
Xbit_r182_c34 bl_34 br_34 wl_182 vdd gnd cell_6t
Xbit_r183_c34 bl_34 br_34 wl_183 vdd gnd cell_6t
Xbit_r184_c34 bl_34 br_34 wl_184 vdd gnd cell_6t
Xbit_r185_c34 bl_34 br_34 wl_185 vdd gnd cell_6t
Xbit_r186_c34 bl_34 br_34 wl_186 vdd gnd cell_6t
Xbit_r187_c34 bl_34 br_34 wl_187 vdd gnd cell_6t
Xbit_r188_c34 bl_34 br_34 wl_188 vdd gnd cell_6t
Xbit_r189_c34 bl_34 br_34 wl_189 vdd gnd cell_6t
Xbit_r190_c34 bl_34 br_34 wl_190 vdd gnd cell_6t
Xbit_r191_c34 bl_34 br_34 wl_191 vdd gnd cell_6t
Xbit_r192_c34 bl_34 br_34 wl_192 vdd gnd cell_6t
Xbit_r193_c34 bl_34 br_34 wl_193 vdd gnd cell_6t
Xbit_r194_c34 bl_34 br_34 wl_194 vdd gnd cell_6t
Xbit_r195_c34 bl_34 br_34 wl_195 vdd gnd cell_6t
Xbit_r196_c34 bl_34 br_34 wl_196 vdd gnd cell_6t
Xbit_r197_c34 bl_34 br_34 wl_197 vdd gnd cell_6t
Xbit_r198_c34 bl_34 br_34 wl_198 vdd gnd cell_6t
Xbit_r199_c34 bl_34 br_34 wl_199 vdd gnd cell_6t
Xbit_r200_c34 bl_34 br_34 wl_200 vdd gnd cell_6t
Xbit_r201_c34 bl_34 br_34 wl_201 vdd gnd cell_6t
Xbit_r202_c34 bl_34 br_34 wl_202 vdd gnd cell_6t
Xbit_r203_c34 bl_34 br_34 wl_203 vdd gnd cell_6t
Xbit_r204_c34 bl_34 br_34 wl_204 vdd gnd cell_6t
Xbit_r205_c34 bl_34 br_34 wl_205 vdd gnd cell_6t
Xbit_r206_c34 bl_34 br_34 wl_206 vdd gnd cell_6t
Xbit_r207_c34 bl_34 br_34 wl_207 vdd gnd cell_6t
Xbit_r208_c34 bl_34 br_34 wl_208 vdd gnd cell_6t
Xbit_r209_c34 bl_34 br_34 wl_209 vdd gnd cell_6t
Xbit_r210_c34 bl_34 br_34 wl_210 vdd gnd cell_6t
Xbit_r211_c34 bl_34 br_34 wl_211 vdd gnd cell_6t
Xbit_r212_c34 bl_34 br_34 wl_212 vdd gnd cell_6t
Xbit_r213_c34 bl_34 br_34 wl_213 vdd gnd cell_6t
Xbit_r214_c34 bl_34 br_34 wl_214 vdd gnd cell_6t
Xbit_r215_c34 bl_34 br_34 wl_215 vdd gnd cell_6t
Xbit_r216_c34 bl_34 br_34 wl_216 vdd gnd cell_6t
Xbit_r217_c34 bl_34 br_34 wl_217 vdd gnd cell_6t
Xbit_r218_c34 bl_34 br_34 wl_218 vdd gnd cell_6t
Xbit_r219_c34 bl_34 br_34 wl_219 vdd gnd cell_6t
Xbit_r220_c34 bl_34 br_34 wl_220 vdd gnd cell_6t
Xbit_r221_c34 bl_34 br_34 wl_221 vdd gnd cell_6t
Xbit_r222_c34 bl_34 br_34 wl_222 vdd gnd cell_6t
Xbit_r223_c34 bl_34 br_34 wl_223 vdd gnd cell_6t
Xbit_r224_c34 bl_34 br_34 wl_224 vdd gnd cell_6t
Xbit_r225_c34 bl_34 br_34 wl_225 vdd gnd cell_6t
Xbit_r226_c34 bl_34 br_34 wl_226 vdd gnd cell_6t
Xbit_r227_c34 bl_34 br_34 wl_227 vdd gnd cell_6t
Xbit_r228_c34 bl_34 br_34 wl_228 vdd gnd cell_6t
Xbit_r229_c34 bl_34 br_34 wl_229 vdd gnd cell_6t
Xbit_r230_c34 bl_34 br_34 wl_230 vdd gnd cell_6t
Xbit_r231_c34 bl_34 br_34 wl_231 vdd gnd cell_6t
Xbit_r232_c34 bl_34 br_34 wl_232 vdd gnd cell_6t
Xbit_r233_c34 bl_34 br_34 wl_233 vdd gnd cell_6t
Xbit_r234_c34 bl_34 br_34 wl_234 vdd gnd cell_6t
Xbit_r235_c34 bl_34 br_34 wl_235 vdd gnd cell_6t
Xbit_r236_c34 bl_34 br_34 wl_236 vdd gnd cell_6t
Xbit_r237_c34 bl_34 br_34 wl_237 vdd gnd cell_6t
Xbit_r238_c34 bl_34 br_34 wl_238 vdd gnd cell_6t
Xbit_r239_c34 bl_34 br_34 wl_239 vdd gnd cell_6t
Xbit_r240_c34 bl_34 br_34 wl_240 vdd gnd cell_6t
Xbit_r241_c34 bl_34 br_34 wl_241 vdd gnd cell_6t
Xbit_r242_c34 bl_34 br_34 wl_242 vdd gnd cell_6t
Xbit_r243_c34 bl_34 br_34 wl_243 vdd gnd cell_6t
Xbit_r244_c34 bl_34 br_34 wl_244 vdd gnd cell_6t
Xbit_r245_c34 bl_34 br_34 wl_245 vdd gnd cell_6t
Xbit_r246_c34 bl_34 br_34 wl_246 vdd gnd cell_6t
Xbit_r247_c34 bl_34 br_34 wl_247 vdd gnd cell_6t
Xbit_r248_c34 bl_34 br_34 wl_248 vdd gnd cell_6t
Xbit_r249_c34 bl_34 br_34 wl_249 vdd gnd cell_6t
Xbit_r250_c34 bl_34 br_34 wl_250 vdd gnd cell_6t
Xbit_r251_c34 bl_34 br_34 wl_251 vdd gnd cell_6t
Xbit_r252_c34 bl_34 br_34 wl_252 vdd gnd cell_6t
Xbit_r253_c34 bl_34 br_34 wl_253 vdd gnd cell_6t
Xbit_r254_c34 bl_34 br_34 wl_254 vdd gnd cell_6t
Xbit_r255_c34 bl_34 br_34 wl_255 vdd gnd cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd cell_6t
Xbit_r1_c35 bl_35 br_35 wl_1 vdd gnd cell_6t
Xbit_r2_c35 bl_35 br_35 wl_2 vdd gnd cell_6t
Xbit_r3_c35 bl_35 br_35 wl_3 vdd gnd cell_6t
Xbit_r4_c35 bl_35 br_35 wl_4 vdd gnd cell_6t
Xbit_r5_c35 bl_35 br_35 wl_5 vdd gnd cell_6t
Xbit_r6_c35 bl_35 br_35 wl_6 vdd gnd cell_6t
Xbit_r7_c35 bl_35 br_35 wl_7 vdd gnd cell_6t
Xbit_r8_c35 bl_35 br_35 wl_8 vdd gnd cell_6t
Xbit_r9_c35 bl_35 br_35 wl_9 vdd gnd cell_6t
Xbit_r10_c35 bl_35 br_35 wl_10 vdd gnd cell_6t
Xbit_r11_c35 bl_35 br_35 wl_11 vdd gnd cell_6t
Xbit_r12_c35 bl_35 br_35 wl_12 vdd gnd cell_6t
Xbit_r13_c35 bl_35 br_35 wl_13 vdd gnd cell_6t
Xbit_r14_c35 bl_35 br_35 wl_14 vdd gnd cell_6t
Xbit_r15_c35 bl_35 br_35 wl_15 vdd gnd cell_6t
Xbit_r16_c35 bl_35 br_35 wl_16 vdd gnd cell_6t
Xbit_r17_c35 bl_35 br_35 wl_17 vdd gnd cell_6t
Xbit_r18_c35 bl_35 br_35 wl_18 vdd gnd cell_6t
Xbit_r19_c35 bl_35 br_35 wl_19 vdd gnd cell_6t
Xbit_r20_c35 bl_35 br_35 wl_20 vdd gnd cell_6t
Xbit_r21_c35 bl_35 br_35 wl_21 vdd gnd cell_6t
Xbit_r22_c35 bl_35 br_35 wl_22 vdd gnd cell_6t
Xbit_r23_c35 bl_35 br_35 wl_23 vdd gnd cell_6t
Xbit_r24_c35 bl_35 br_35 wl_24 vdd gnd cell_6t
Xbit_r25_c35 bl_35 br_35 wl_25 vdd gnd cell_6t
Xbit_r26_c35 bl_35 br_35 wl_26 vdd gnd cell_6t
Xbit_r27_c35 bl_35 br_35 wl_27 vdd gnd cell_6t
Xbit_r28_c35 bl_35 br_35 wl_28 vdd gnd cell_6t
Xbit_r29_c35 bl_35 br_35 wl_29 vdd gnd cell_6t
Xbit_r30_c35 bl_35 br_35 wl_30 vdd gnd cell_6t
Xbit_r31_c35 bl_35 br_35 wl_31 vdd gnd cell_6t
Xbit_r32_c35 bl_35 br_35 wl_32 vdd gnd cell_6t
Xbit_r33_c35 bl_35 br_35 wl_33 vdd gnd cell_6t
Xbit_r34_c35 bl_35 br_35 wl_34 vdd gnd cell_6t
Xbit_r35_c35 bl_35 br_35 wl_35 vdd gnd cell_6t
Xbit_r36_c35 bl_35 br_35 wl_36 vdd gnd cell_6t
Xbit_r37_c35 bl_35 br_35 wl_37 vdd gnd cell_6t
Xbit_r38_c35 bl_35 br_35 wl_38 vdd gnd cell_6t
Xbit_r39_c35 bl_35 br_35 wl_39 vdd gnd cell_6t
Xbit_r40_c35 bl_35 br_35 wl_40 vdd gnd cell_6t
Xbit_r41_c35 bl_35 br_35 wl_41 vdd gnd cell_6t
Xbit_r42_c35 bl_35 br_35 wl_42 vdd gnd cell_6t
Xbit_r43_c35 bl_35 br_35 wl_43 vdd gnd cell_6t
Xbit_r44_c35 bl_35 br_35 wl_44 vdd gnd cell_6t
Xbit_r45_c35 bl_35 br_35 wl_45 vdd gnd cell_6t
Xbit_r46_c35 bl_35 br_35 wl_46 vdd gnd cell_6t
Xbit_r47_c35 bl_35 br_35 wl_47 vdd gnd cell_6t
Xbit_r48_c35 bl_35 br_35 wl_48 vdd gnd cell_6t
Xbit_r49_c35 bl_35 br_35 wl_49 vdd gnd cell_6t
Xbit_r50_c35 bl_35 br_35 wl_50 vdd gnd cell_6t
Xbit_r51_c35 bl_35 br_35 wl_51 vdd gnd cell_6t
Xbit_r52_c35 bl_35 br_35 wl_52 vdd gnd cell_6t
Xbit_r53_c35 bl_35 br_35 wl_53 vdd gnd cell_6t
Xbit_r54_c35 bl_35 br_35 wl_54 vdd gnd cell_6t
Xbit_r55_c35 bl_35 br_35 wl_55 vdd gnd cell_6t
Xbit_r56_c35 bl_35 br_35 wl_56 vdd gnd cell_6t
Xbit_r57_c35 bl_35 br_35 wl_57 vdd gnd cell_6t
Xbit_r58_c35 bl_35 br_35 wl_58 vdd gnd cell_6t
Xbit_r59_c35 bl_35 br_35 wl_59 vdd gnd cell_6t
Xbit_r60_c35 bl_35 br_35 wl_60 vdd gnd cell_6t
Xbit_r61_c35 bl_35 br_35 wl_61 vdd gnd cell_6t
Xbit_r62_c35 bl_35 br_35 wl_62 vdd gnd cell_6t
Xbit_r63_c35 bl_35 br_35 wl_63 vdd gnd cell_6t
Xbit_r64_c35 bl_35 br_35 wl_64 vdd gnd cell_6t
Xbit_r65_c35 bl_35 br_35 wl_65 vdd gnd cell_6t
Xbit_r66_c35 bl_35 br_35 wl_66 vdd gnd cell_6t
Xbit_r67_c35 bl_35 br_35 wl_67 vdd gnd cell_6t
Xbit_r68_c35 bl_35 br_35 wl_68 vdd gnd cell_6t
Xbit_r69_c35 bl_35 br_35 wl_69 vdd gnd cell_6t
Xbit_r70_c35 bl_35 br_35 wl_70 vdd gnd cell_6t
Xbit_r71_c35 bl_35 br_35 wl_71 vdd gnd cell_6t
Xbit_r72_c35 bl_35 br_35 wl_72 vdd gnd cell_6t
Xbit_r73_c35 bl_35 br_35 wl_73 vdd gnd cell_6t
Xbit_r74_c35 bl_35 br_35 wl_74 vdd gnd cell_6t
Xbit_r75_c35 bl_35 br_35 wl_75 vdd gnd cell_6t
Xbit_r76_c35 bl_35 br_35 wl_76 vdd gnd cell_6t
Xbit_r77_c35 bl_35 br_35 wl_77 vdd gnd cell_6t
Xbit_r78_c35 bl_35 br_35 wl_78 vdd gnd cell_6t
Xbit_r79_c35 bl_35 br_35 wl_79 vdd gnd cell_6t
Xbit_r80_c35 bl_35 br_35 wl_80 vdd gnd cell_6t
Xbit_r81_c35 bl_35 br_35 wl_81 vdd gnd cell_6t
Xbit_r82_c35 bl_35 br_35 wl_82 vdd gnd cell_6t
Xbit_r83_c35 bl_35 br_35 wl_83 vdd gnd cell_6t
Xbit_r84_c35 bl_35 br_35 wl_84 vdd gnd cell_6t
Xbit_r85_c35 bl_35 br_35 wl_85 vdd gnd cell_6t
Xbit_r86_c35 bl_35 br_35 wl_86 vdd gnd cell_6t
Xbit_r87_c35 bl_35 br_35 wl_87 vdd gnd cell_6t
Xbit_r88_c35 bl_35 br_35 wl_88 vdd gnd cell_6t
Xbit_r89_c35 bl_35 br_35 wl_89 vdd gnd cell_6t
Xbit_r90_c35 bl_35 br_35 wl_90 vdd gnd cell_6t
Xbit_r91_c35 bl_35 br_35 wl_91 vdd gnd cell_6t
Xbit_r92_c35 bl_35 br_35 wl_92 vdd gnd cell_6t
Xbit_r93_c35 bl_35 br_35 wl_93 vdd gnd cell_6t
Xbit_r94_c35 bl_35 br_35 wl_94 vdd gnd cell_6t
Xbit_r95_c35 bl_35 br_35 wl_95 vdd gnd cell_6t
Xbit_r96_c35 bl_35 br_35 wl_96 vdd gnd cell_6t
Xbit_r97_c35 bl_35 br_35 wl_97 vdd gnd cell_6t
Xbit_r98_c35 bl_35 br_35 wl_98 vdd gnd cell_6t
Xbit_r99_c35 bl_35 br_35 wl_99 vdd gnd cell_6t
Xbit_r100_c35 bl_35 br_35 wl_100 vdd gnd cell_6t
Xbit_r101_c35 bl_35 br_35 wl_101 vdd gnd cell_6t
Xbit_r102_c35 bl_35 br_35 wl_102 vdd gnd cell_6t
Xbit_r103_c35 bl_35 br_35 wl_103 vdd gnd cell_6t
Xbit_r104_c35 bl_35 br_35 wl_104 vdd gnd cell_6t
Xbit_r105_c35 bl_35 br_35 wl_105 vdd gnd cell_6t
Xbit_r106_c35 bl_35 br_35 wl_106 vdd gnd cell_6t
Xbit_r107_c35 bl_35 br_35 wl_107 vdd gnd cell_6t
Xbit_r108_c35 bl_35 br_35 wl_108 vdd gnd cell_6t
Xbit_r109_c35 bl_35 br_35 wl_109 vdd gnd cell_6t
Xbit_r110_c35 bl_35 br_35 wl_110 vdd gnd cell_6t
Xbit_r111_c35 bl_35 br_35 wl_111 vdd gnd cell_6t
Xbit_r112_c35 bl_35 br_35 wl_112 vdd gnd cell_6t
Xbit_r113_c35 bl_35 br_35 wl_113 vdd gnd cell_6t
Xbit_r114_c35 bl_35 br_35 wl_114 vdd gnd cell_6t
Xbit_r115_c35 bl_35 br_35 wl_115 vdd gnd cell_6t
Xbit_r116_c35 bl_35 br_35 wl_116 vdd gnd cell_6t
Xbit_r117_c35 bl_35 br_35 wl_117 vdd gnd cell_6t
Xbit_r118_c35 bl_35 br_35 wl_118 vdd gnd cell_6t
Xbit_r119_c35 bl_35 br_35 wl_119 vdd gnd cell_6t
Xbit_r120_c35 bl_35 br_35 wl_120 vdd gnd cell_6t
Xbit_r121_c35 bl_35 br_35 wl_121 vdd gnd cell_6t
Xbit_r122_c35 bl_35 br_35 wl_122 vdd gnd cell_6t
Xbit_r123_c35 bl_35 br_35 wl_123 vdd gnd cell_6t
Xbit_r124_c35 bl_35 br_35 wl_124 vdd gnd cell_6t
Xbit_r125_c35 bl_35 br_35 wl_125 vdd gnd cell_6t
Xbit_r126_c35 bl_35 br_35 wl_126 vdd gnd cell_6t
Xbit_r127_c35 bl_35 br_35 wl_127 vdd gnd cell_6t
Xbit_r128_c35 bl_35 br_35 wl_128 vdd gnd cell_6t
Xbit_r129_c35 bl_35 br_35 wl_129 vdd gnd cell_6t
Xbit_r130_c35 bl_35 br_35 wl_130 vdd gnd cell_6t
Xbit_r131_c35 bl_35 br_35 wl_131 vdd gnd cell_6t
Xbit_r132_c35 bl_35 br_35 wl_132 vdd gnd cell_6t
Xbit_r133_c35 bl_35 br_35 wl_133 vdd gnd cell_6t
Xbit_r134_c35 bl_35 br_35 wl_134 vdd gnd cell_6t
Xbit_r135_c35 bl_35 br_35 wl_135 vdd gnd cell_6t
Xbit_r136_c35 bl_35 br_35 wl_136 vdd gnd cell_6t
Xbit_r137_c35 bl_35 br_35 wl_137 vdd gnd cell_6t
Xbit_r138_c35 bl_35 br_35 wl_138 vdd gnd cell_6t
Xbit_r139_c35 bl_35 br_35 wl_139 vdd gnd cell_6t
Xbit_r140_c35 bl_35 br_35 wl_140 vdd gnd cell_6t
Xbit_r141_c35 bl_35 br_35 wl_141 vdd gnd cell_6t
Xbit_r142_c35 bl_35 br_35 wl_142 vdd gnd cell_6t
Xbit_r143_c35 bl_35 br_35 wl_143 vdd gnd cell_6t
Xbit_r144_c35 bl_35 br_35 wl_144 vdd gnd cell_6t
Xbit_r145_c35 bl_35 br_35 wl_145 vdd gnd cell_6t
Xbit_r146_c35 bl_35 br_35 wl_146 vdd gnd cell_6t
Xbit_r147_c35 bl_35 br_35 wl_147 vdd gnd cell_6t
Xbit_r148_c35 bl_35 br_35 wl_148 vdd gnd cell_6t
Xbit_r149_c35 bl_35 br_35 wl_149 vdd gnd cell_6t
Xbit_r150_c35 bl_35 br_35 wl_150 vdd gnd cell_6t
Xbit_r151_c35 bl_35 br_35 wl_151 vdd gnd cell_6t
Xbit_r152_c35 bl_35 br_35 wl_152 vdd gnd cell_6t
Xbit_r153_c35 bl_35 br_35 wl_153 vdd gnd cell_6t
Xbit_r154_c35 bl_35 br_35 wl_154 vdd gnd cell_6t
Xbit_r155_c35 bl_35 br_35 wl_155 vdd gnd cell_6t
Xbit_r156_c35 bl_35 br_35 wl_156 vdd gnd cell_6t
Xbit_r157_c35 bl_35 br_35 wl_157 vdd gnd cell_6t
Xbit_r158_c35 bl_35 br_35 wl_158 vdd gnd cell_6t
Xbit_r159_c35 bl_35 br_35 wl_159 vdd gnd cell_6t
Xbit_r160_c35 bl_35 br_35 wl_160 vdd gnd cell_6t
Xbit_r161_c35 bl_35 br_35 wl_161 vdd gnd cell_6t
Xbit_r162_c35 bl_35 br_35 wl_162 vdd gnd cell_6t
Xbit_r163_c35 bl_35 br_35 wl_163 vdd gnd cell_6t
Xbit_r164_c35 bl_35 br_35 wl_164 vdd gnd cell_6t
Xbit_r165_c35 bl_35 br_35 wl_165 vdd gnd cell_6t
Xbit_r166_c35 bl_35 br_35 wl_166 vdd gnd cell_6t
Xbit_r167_c35 bl_35 br_35 wl_167 vdd gnd cell_6t
Xbit_r168_c35 bl_35 br_35 wl_168 vdd gnd cell_6t
Xbit_r169_c35 bl_35 br_35 wl_169 vdd gnd cell_6t
Xbit_r170_c35 bl_35 br_35 wl_170 vdd gnd cell_6t
Xbit_r171_c35 bl_35 br_35 wl_171 vdd gnd cell_6t
Xbit_r172_c35 bl_35 br_35 wl_172 vdd gnd cell_6t
Xbit_r173_c35 bl_35 br_35 wl_173 vdd gnd cell_6t
Xbit_r174_c35 bl_35 br_35 wl_174 vdd gnd cell_6t
Xbit_r175_c35 bl_35 br_35 wl_175 vdd gnd cell_6t
Xbit_r176_c35 bl_35 br_35 wl_176 vdd gnd cell_6t
Xbit_r177_c35 bl_35 br_35 wl_177 vdd gnd cell_6t
Xbit_r178_c35 bl_35 br_35 wl_178 vdd gnd cell_6t
Xbit_r179_c35 bl_35 br_35 wl_179 vdd gnd cell_6t
Xbit_r180_c35 bl_35 br_35 wl_180 vdd gnd cell_6t
Xbit_r181_c35 bl_35 br_35 wl_181 vdd gnd cell_6t
Xbit_r182_c35 bl_35 br_35 wl_182 vdd gnd cell_6t
Xbit_r183_c35 bl_35 br_35 wl_183 vdd gnd cell_6t
Xbit_r184_c35 bl_35 br_35 wl_184 vdd gnd cell_6t
Xbit_r185_c35 bl_35 br_35 wl_185 vdd gnd cell_6t
Xbit_r186_c35 bl_35 br_35 wl_186 vdd gnd cell_6t
Xbit_r187_c35 bl_35 br_35 wl_187 vdd gnd cell_6t
Xbit_r188_c35 bl_35 br_35 wl_188 vdd gnd cell_6t
Xbit_r189_c35 bl_35 br_35 wl_189 vdd gnd cell_6t
Xbit_r190_c35 bl_35 br_35 wl_190 vdd gnd cell_6t
Xbit_r191_c35 bl_35 br_35 wl_191 vdd gnd cell_6t
Xbit_r192_c35 bl_35 br_35 wl_192 vdd gnd cell_6t
Xbit_r193_c35 bl_35 br_35 wl_193 vdd gnd cell_6t
Xbit_r194_c35 bl_35 br_35 wl_194 vdd gnd cell_6t
Xbit_r195_c35 bl_35 br_35 wl_195 vdd gnd cell_6t
Xbit_r196_c35 bl_35 br_35 wl_196 vdd gnd cell_6t
Xbit_r197_c35 bl_35 br_35 wl_197 vdd gnd cell_6t
Xbit_r198_c35 bl_35 br_35 wl_198 vdd gnd cell_6t
Xbit_r199_c35 bl_35 br_35 wl_199 vdd gnd cell_6t
Xbit_r200_c35 bl_35 br_35 wl_200 vdd gnd cell_6t
Xbit_r201_c35 bl_35 br_35 wl_201 vdd gnd cell_6t
Xbit_r202_c35 bl_35 br_35 wl_202 vdd gnd cell_6t
Xbit_r203_c35 bl_35 br_35 wl_203 vdd gnd cell_6t
Xbit_r204_c35 bl_35 br_35 wl_204 vdd gnd cell_6t
Xbit_r205_c35 bl_35 br_35 wl_205 vdd gnd cell_6t
Xbit_r206_c35 bl_35 br_35 wl_206 vdd gnd cell_6t
Xbit_r207_c35 bl_35 br_35 wl_207 vdd gnd cell_6t
Xbit_r208_c35 bl_35 br_35 wl_208 vdd gnd cell_6t
Xbit_r209_c35 bl_35 br_35 wl_209 vdd gnd cell_6t
Xbit_r210_c35 bl_35 br_35 wl_210 vdd gnd cell_6t
Xbit_r211_c35 bl_35 br_35 wl_211 vdd gnd cell_6t
Xbit_r212_c35 bl_35 br_35 wl_212 vdd gnd cell_6t
Xbit_r213_c35 bl_35 br_35 wl_213 vdd gnd cell_6t
Xbit_r214_c35 bl_35 br_35 wl_214 vdd gnd cell_6t
Xbit_r215_c35 bl_35 br_35 wl_215 vdd gnd cell_6t
Xbit_r216_c35 bl_35 br_35 wl_216 vdd gnd cell_6t
Xbit_r217_c35 bl_35 br_35 wl_217 vdd gnd cell_6t
Xbit_r218_c35 bl_35 br_35 wl_218 vdd gnd cell_6t
Xbit_r219_c35 bl_35 br_35 wl_219 vdd gnd cell_6t
Xbit_r220_c35 bl_35 br_35 wl_220 vdd gnd cell_6t
Xbit_r221_c35 bl_35 br_35 wl_221 vdd gnd cell_6t
Xbit_r222_c35 bl_35 br_35 wl_222 vdd gnd cell_6t
Xbit_r223_c35 bl_35 br_35 wl_223 vdd gnd cell_6t
Xbit_r224_c35 bl_35 br_35 wl_224 vdd gnd cell_6t
Xbit_r225_c35 bl_35 br_35 wl_225 vdd gnd cell_6t
Xbit_r226_c35 bl_35 br_35 wl_226 vdd gnd cell_6t
Xbit_r227_c35 bl_35 br_35 wl_227 vdd gnd cell_6t
Xbit_r228_c35 bl_35 br_35 wl_228 vdd gnd cell_6t
Xbit_r229_c35 bl_35 br_35 wl_229 vdd gnd cell_6t
Xbit_r230_c35 bl_35 br_35 wl_230 vdd gnd cell_6t
Xbit_r231_c35 bl_35 br_35 wl_231 vdd gnd cell_6t
Xbit_r232_c35 bl_35 br_35 wl_232 vdd gnd cell_6t
Xbit_r233_c35 bl_35 br_35 wl_233 vdd gnd cell_6t
Xbit_r234_c35 bl_35 br_35 wl_234 vdd gnd cell_6t
Xbit_r235_c35 bl_35 br_35 wl_235 vdd gnd cell_6t
Xbit_r236_c35 bl_35 br_35 wl_236 vdd gnd cell_6t
Xbit_r237_c35 bl_35 br_35 wl_237 vdd gnd cell_6t
Xbit_r238_c35 bl_35 br_35 wl_238 vdd gnd cell_6t
Xbit_r239_c35 bl_35 br_35 wl_239 vdd gnd cell_6t
Xbit_r240_c35 bl_35 br_35 wl_240 vdd gnd cell_6t
Xbit_r241_c35 bl_35 br_35 wl_241 vdd gnd cell_6t
Xbit_r242_c35 bl_35 br_35 wl_242 vdd gnd cell_6t
Xbit_r243_c35 bl_35 br_35 wl_243 vdd gnd cell_6t
Xbit_r244_c35 bl_35 br_35 wl_244 vdd gnd cell_6t
Xbit_r245_c35 bl_35 br_35 wl_245 vdd gnd cell_6t
Xbit_r246_c35 bl_35 br_35 wl_246 vdd gnd cell_6t
Xbit_r247_c35 bl_35 br_35 wl_247 vdd gnd cell_6t
Xbit_r248_c35 bl_35 br_35 wl_248 vdd gnd cell_6t
Xbit_r249_c35 bl_35 br_35 wl_249 vdd gnd cell_6t
Xbit_r250_c35 bl_35 br_35 wl_250 vdd gnd cell_6t
Xbit_r251_c35 bl_35 br_35 wl_251 vdd gnd cell_6t
Xbit_r252_c35 bl_35 br_35 wl_252 vdd gnd cell_6t
Xbit_r253_c35 bl_35 br_35 wl_253 vdd gnd cell_6t
Xbit_r254_c35 bl_35 br_35 wl_254 vdd gnd cell_6t
Xbit_r255_c35 bl_35 br_35 wl_255 vdd gnd cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd cell_6t
Xbit_r1_c36 bl_36 br_36 wl_1 vdd gnd cell_6t
Xbit_r2_c36 bl_36 br_36 wl_2 vdd gnd cell_6t
Xbit_r3_c36 bl_36 br_36 wl_3 vdd gnd cell_6t
Xbit_r4_c36 bl_36 br_36 wl_4 vdd gnd cell_6t
Xbit_r5_c36 bl_36 br_36 wl_5 vdd gnd cell_6t
Xbit_r6_c36 bl_36 br_36 wl_6 vdd gnd cell_6t
Xbit_r7_c36 bl_36 br_36 wl_7 vdd gnd cell_6t
Xbit_r8_c36 bl_36 br_36 wl_8 vdd gnd cell_6t
Xbit_r9_c36 bl_36 br_36 wl_9 vdd gnd cell_6t
Xbit_r10_c36 bl_36 br_36 wl_10 vdd gnd cell_6t
Xbit_r11_c36 bl_36 br_36 wl_11 vdd gnd cell_6t
Xbit_r12_c36 bl_36 br_36 wl_12 vdd gnd cell_6t
Xbit_r13_c36 bl_36 br_36 wl_13 vdd gnd cell_6t
Xbit_r14_c36 bl_36 br_36 wl_14 vdd gnd cell_6t
Xbit_r15_c36 bl_36 br_36 wl_15 vdd gnd cell_6t
Xbit_r16_c36 bl_36 br_36 wl_16 vdd gnd cell_6t
Xbit_r17_c36 bl_36 br_36 wl_17 vdd gnd cell_6t
Xbit_r18_c36 bl_36 br_36 wl_18 vdd gnd cell_6t
Xbit_r19_c36 bl_36 br_36 wl_19 vdd gnd cell_6t
Xbit_r20_c36 bl_36 br_36 wl_20 vdd gnd cell_6t
Xbit_r21_c36 bl_36 br_36 wl_21 vdd gnd cell_6t
Xbit_r22_c36 bl_36 br_36 wl_22 vdd gnd cell_6t
Xbit_r23_c36 bl_36 br_36 wl_23 vdd gnd cell_6t
Xbit_r24_c36 bl_36 br_36 wl_24 vdd gnd cell_6t
Xbit_r25_c36 bl_36 br_36 wl_25 vdd gnd cell_6t
Xbit_r26_c36 bl_36 br_36 wl_26 vdd gnd cell_6t
Xbit_r27_c36 bl_36 br_36 wl_27 vdd gnd cell_6t
Xbit_r28_c36 bl_36 br_36 wl_28 vdd gnd cell_6t
Xbit_r29_c36 bl_36 br_36 wl_29 vdd gnd cell_6t
Xbit_r30_c36 bl_36 br_36 wl_30 vdd gnd cell_6t
Xbit_r31_c36 bl_36 br_36 wl_31 vdd gnd cell_6t
Xbit_r32_c36 bl_36 br_36 wl_32 vdd gnd cell_6t
Xbit_r33_c36 bl_36 br_36 wl_33 vdd gnd cell_6t
Xbit_r34_c36 bl_36 br_36 wl_34 vdd gnd cell_6t
Xbit_r35_c36 bl_36 br_36 wl_35 vdd gnd cell_6t
Xbit_r36_c36 bl_36 br_36 wl_36 vdd gnd cell_6t
Xbit_r37_c36 bl_36 br_36 wl_37 vdd gnd cell_6t
Xbit_r38_c36 bl_36 br_36 wl_38 vdd gnd cell_6t
Xbit_r39_c36 bl_36 br_36 wl_39 vdd gnd cell_6t
Xbit_r40_c36 bl_36 br_36 wl_40 vdd gnd cell_6t
Xbit_r41_c36 bl_36 br_36 wl_41 vdd gnd cell_6t
Xbit_r42_c36 bl_36 br_36 wl_42 vdd gnd cell_6t
Xbit_r43_c36 bl_36 br_36 wl_43 vdd gnd cell_6t
Xbit_r44_c36 bl_36 br_36 wl_44 vdd gnd cell_6t
Xbit_r45_c36 bl_36 br_36 wl_45 vdd gnd cell_6t
Xbit_r46_c36 bl_36 br_36 wl_46 vdd gnd cell_6t
Xbit_r47_c36 bl_36 br_36 wl_47 vdd gnd cell_6t
Xbit_r48_c36 bl_36 br_36 wl_48 vdd gnd cell_6t
Xbit_r49_c36 bl_36 br_36 wl_49 vdd gnd cell_6t
Xbit_r50_c36 bl_36 br_36 wl_50 vdd gnd cell_6t
Xbit_r51_c36 bl_36 br_36 wl_51 vdd gnd cell_6t
Xbit_r52_c36 bl_36 br_36 wl_52 vdd gnd cell_6t
Xbit_r53_c36 bl_36 br_36 wl_53 vdd gnd cell_6t
Xbit_r54_c36 bl_36 br_36 wl_54 vdd gnd cell_6t
Xbit_r55_c36 bl_36 br_36 wl_55 vdd gnd cell_6t
Xbit_r56_c36 bl_36 br_36 wl_56 vdd gnd cell_6t
Xbit_r57_c36 bl_36 br_36 wl_57 vdd gnd cell_6t
Xbit_r58_c36 bl_36 br_36 wl_58 vdd gnd cell_6t
Xbit_r59_c36 bl_36 br_36 wl_59 vdd gnd cell_6t
Xbit_r60_c36 bl_36 br_36 wl_60 vdd gnd cell_6t
Xbit_r61_c36 bl_36 br_36 wl_61 vdd gnd cell_6t
Xbit_r62_c36 bl_36 br_36 wl_62 vdd gnd cell_6t
Xbit_r63_c36 bl_36 br_36 wl_63 vdd gnd cell_6t
Xbit_r64_c36 bl_36 br_36 wl_64 vdd gnd cell_6t
Xbit_r65_c36 bl_36 br_36 wl_65 vdd gnd cell_6t
Xbit_r66_c36 bl_36 br_36 wl_66 vdd gnd cell_6t
Xbit_r67_c36 bl_36 br_36 wl_67 vdd gnd cell_6t
Xbit_r68_c36 bl_36 br_36 wl_68 vdd gnd cell_6t
Xbit_r69_c36 bl_36 br_36 wl_69 vdd gnd cell_6t
Xbit_r70_c36 bl_36 br_36 wl_70 vdd gnd cell_6t
Xbit_r71_c36 bl_36 br_36 wl_71 vdd gnd cell_6t
Xbit_r72_c36 bl_36 br_36 wl_72 vdd gnd cell_6t
Xbit_r73_c36 bl_36 br_36 wl_73 vdd gnd cell_6t
Xbit_r74_c36 bl_36 br_36 wl_74 vdd gnd cell_6t
Xbit_r75_c36 bl_36 br_36 wl_75 vdd gnd cell_6t
Xbit_r76_c36 bl_36 br_36 wl_76 vdd gnd cell_6t
Xbit_r77_c36 bl_36 br_36 wl_77 vdd gnd cell_6t
Xbit_r78_c36 bl_36 br_36 wl_78 vdd gnd cell_6t
Xbit_r79_c36 bl_36 br_36 wl_79 vdd gnd cell_6t
Xbit_r80_c36 bl_36 br_36 wl_80 vdd gnd cell_6t
Xbit_r81_c36 bl_36 br_36 wl_81 vdd gnd cell_6t
Xbit_r82_c36 bl_36 br_36 wl_82 vdd gnd cell_6t
Xbit_r83_c36 bl_36 br_36 wl_83 vdd gnd cell_6t
Xbit_r84_c36 bl_36 br_36 wl_84 vdd gnd cell_6t
Xbit_r85_c36 bl_36 br_36 wl_85 vdd gnd cell_6t
Xbit_r86_c36 bl_36 br_36 wl_86 vdd gnd cell_6t
Xbit_r87_c36 bl_36 br_36 wl_87 vdd gnd cell_6t
Xbit_r88_c36 bl_36 br_36 wl_88 vdd gnd cell_6t
Xbit_r89_c36 bl_36 br_36 wl_89 vdd gnd cell_6t
Xbit_r90_c36 bl_36 br_36 wl_90 vdd gnd cell_6t
Xbit_r91_c36 bl_36 br_36 wl_91 vdd gnd cell_6t
Xbit_r92_c36 bl_36 br_36 wl_92 vdd gnd cell_6t
Xbit_r93_c36 bl_36 br_36 wl_93 vdd gnd cell_6t
Xbit_r94_c36 bl_36 br_36 wl_94 vdd gnd cell_6t
Xbit_r95_c36 bl_36 br_36 wl_95 vdd gnd cell_6t
Xbit_r96_c36 bl_36 br_36 wl_96 vdd gnd cell_6t
Xbit_r97_c36 bl_36 br_36 wl_97 vdd gnd cell_6t
Xbit_r98_c36 bl_36 br_36 wl_98 vdd gnd cell_6t
Xbit_r99_c36 bl_36 br_36 wl_99 vdd gnd cell_6t
Xbit_r100_c36 bl_36 br_36 wl_100 vdd gnd cell_6t
Xbit_r101_c36 bl_36 br_36 wl_101 vdd gnd cell_6t
Xbit_r102_c36 bl_36 br_36 wl_102 vdd gnd cell_6t
Xbit_r103_c36 bl_36 br_36 wl_103 vdd gnd cell_6t
Xbit_r104_c36 bl_36 br_36 wl_104 vdd gnd cell_6t
Xbit_r105_c36 bl_36 br_36 wl_105 vdd gnd cell_6t
Xbit_r106_c36 bl_36 br_36 wl_106 vdd gnd cell_6t
Xbit_r107_c36 bl_36 br_36 wl_107 vdd gnd cell_6t
Xbit_r108_c36 bl_36 br_36 wl_108 vdd gnd cell_6t
Xbit_r109_c36 bl_36 br_36 wl_109 vdd gnd cell_6t
Xbit_r110_c36 bl_36 br_36 wl_110 vdd gnd cell_6t
Xbit_r111_c36 bl_36 br_36 wl_111 vdd gnd cell_6t
Xbit_r112_c36 bl_36 br_36 wl_112 vdd gnd cell_6t
Xbit_r113_c36 bl_36 br_36 wl_113 vdd gnd cell_6t
Xbit_r114_c36 bl_36 br_36 wl_114 vdd gnd cell_6t
Xbit_r115_c36 bl_36 br_36 wl_115 vdd gnd cell_6t
Xbit_r116_c36 bl_36 br_36 wl_116 vdd gnd cell_6t
Xbit_r117_c36 bl_36 br_36 wl_117 vdd gnd cell_6t
Xbit_r118_c36 bl_36 br_36 wl_118 vdd gnd cell_6t
Xbit_r119_c36 bl_36 br_36 wl_119 vdd gnd cell_6t
Xbit_r120_c36 bl_36 br_36 wl_120 vdd gnd cell_6t
Xbit_r121_c36 bl_36 br_36 wl_121 vdd gnd cell_6t
Xbit_r122_c36 bl_36 br_36 wl_122 vdd gnd cell_6t
Xbit_r123_c36 bl_36 br_36 wl_123 vdd gnd cell_6t
Xbit_r124_c36 bl_36 br_36 wl_124 vdd gnd cell_6t
Xbit_r125_c36 bl_36 br_36 wl_125 vdd gnd cell_6t
Xbit_r126_c36 bl_36 br_36 wl_126 vdd gnd cell_6t
Xbit_r127_c36 bl_36 br_36 wl_127 vdd gnd cell_6t
Xbit_r128_c36 bl_36 br_36 wl_128 vdd gnd cell_6t
Xbit_r129_c36 bl_36 br_36 wl_129 vdd gnd cell_6t
Xbit_r130_c36 bl_36 br_36 wl_130 vdd gnd cell_6t
Xbit_r131_c36 bl_36 br_36 wl_131 vdd gnd cell_6t
Xbit_r132_c36 bl_36 br_36 wl_132 vdd gnd cell_6t
Xbit_r133_c36 bl_36 br_36 wl_133 vdd gnd cell_6t
Xbit_r134_c36 bl_36 br_36 wl_134 vdd gnd cell_6t
Xbit_r135_c36 bl_36 br_36 wl_135 vdd gnd cell_6t
Xbit_r136_c36 bl_36 br_36 wl_136 vdd gnd cell_6t
Xbit_r137_c36 bl_36 br_36 wl_137 vdd gnd cell_6t
Xbit_r138_c36 bl_36 br_36 wl_138 vdd gnd cell_6t
Xbit_r139_c36 bl_36 br_36 wl_139 vdd gnd cell_6t
Xbit_r140_c36 bl_36 br_36 wl_140 vdd gnd cell_6t
Xbit_r141_c36 bl_36 br_36 wl_141 vdd gnd cell_6t
Xbit_r142_c36 bl_36 br_36 wl_142 vdd gnd cell_6t
Xbit_r143_c36 bl_36 br_36 wl_143 vdd gnd cell_6t
Xbit_r144_c36 bl_36 br_36 wl_144 vdd gnd cell_6t
Xbit_r145_c36 bl_36 br_36 wl_145 vdd gnd cell_6t
Xbit_r146_c36 bl_36 br_36 wl_146 vdd gnd cell_6t
Xbit_r147_c36 bl_36 br_36 wl_147 vdd gnd cell_6t
Xbit_r148_c36 bl_36 br_36 wl_148 vdd gnd cell_6t
Xbit_r149_c36 bl_36 br_36 wl_149 vdd gnd cell_6t
Xbit_r150_c36 bl_36 br_36 wl_150 vdd gnd cell_6t
Xbit_r151_c36 bl_36 br_36 wl_151 vdd gnd cell_6t
Xbit_r152_c36 bl_36 br_36 wl_152 vdd gnd cell_6t
Xbit_r153_c36 bl_36 br_36 wl_153 vdd gnd cell_6t
Xbit_r154_c36 bl_36 br_36 wl_154 vdd gnd cell_6t
Xbit_r155_c36 bl_36 br_36 wl_155 vdd gnd cell_6t
Xbit_r156_c36 bl_36 br_36 wl_156 vdd gnd cell_6t
Xbit_r157_c36 bl_36 br_36 wl_157 vdd gnd cell_6t
Xbit_r158_c36 bl_36 br_36 wl_158 vdd gnd cell_6t
Xbit_r159_c36 bl_36 br_36 wl_159 vdd gnd cell_6t
Xbit_r160_c36 bl_36 br_36 wl_160 vdd gnd cell_6t
Xbit_r161_c36 bl_36 br_36 wl_161 vdd gnd cell_6t
Xbit_r162_c36 bl_36 br_36 wl_162 vdd gnd cell_6t
Xbit_r163_c36 bl_36 br_36 wl_163 vdd gnd cell_6t
Xbit_r164_c36 bl_36 br_36 wl_164 vdd gnd cell_6t
Xbit_r165_c36 bl_36 br_36 wl_165 vdd gnd cell_6t
Xbit_r166_c36 bl_36 br_36 wl_166 vdd gnd cell_6t
Xbit_r167_c36 bl_36 br_36 wl_167 vdd gnd cell_6t
Xbit_r168_c36 bl_36 br_36 wl_168 vdd gnd cell_6t
Xbit_r169_c36 bl_36 br_36 wl_169 vdd gnd cell_6t
Xbit_r170_c36 bl_36 br_36 wl_170 vdd gnd cell_6t
Xbit_r171_c36 bl_36 br_36 wl_171 vdd gnd cell_6t
Xbit_r172_c36 bl_36 br_36 wl_172 vdd gnd cell_6t
Xbit_r173_c36 bl_36 br_36 wl_173 vdd gnd cell_6t
Xbit_r174_c36 bl_36 br_36 wl_174 vdd gnd cell_6t
Xbit_r175_c36 bl_36 br_36 wl_175 vdd gnd cell_6t
Xbit_r176_c36 bl_36 br_36 wl_176 vdd gnd cell_6t
Xbit_r177_c36 bl_36 br_36 wl_177 vdd gnd cell_6t
Xbit_r178_c36 bl_36 br_36 wl_178 vdd gnd cell_6t
Xbit_r179_c36 bl_36 br_36 wl_179 vdd gnd cell_6t
Xbit_r180_c36 bl_36 br_36 wl_180 vdd gnd cell_6t
Xbit_r181_c36 bl_36 br_36 wl_181 vdd gnd cell_6t
Xbit_r182_c36 bl_36 br_36 wl_182 vdd gnd cell_6t
Xbit_r183_c36 bl_36 br_36 wl_183 vdd gnd cell_6t
Xbit_r184_c36 bl_36 br_36 wl_184 vdd gnd cell_6t
Xbit_r185_c36 bl_36 br_36 wl_185 vdd gnd cell_6t
Xbit_r186_c36 bl_36 br_36 wl_186 vdd gnd cell_6t
Xbit_r187_c36 bl_36 br_36 wl_187 vdd gnd cell_6t
Xbit_r188_c36 bl_36 br_36 wl_188 vdd gnd cell_6t
Xbit_r189_c36 bl_36 br_36 wl_189 vdd gnd cell_6t
Xbit_r190_c36 bl_36 br_36 wl_190 vdd gnd cell_6t
Xbit_r191_c36 bl_36 br_36 wl_191 vdd gnd cell_6t
Xbit_r192_c36 bl_36 br_36 wl_192 vdd gnd cell_6t
Xbit_r193_c36 bl_36 br_36 wl_193 vdd gnd cell_6t
Xbit_r194_c36 bl_36 br_36 wl_194 vdd gnd cell_6t
Xbit_r195_c36 bl_36 br_36 wl_195 vdd gnd cell_6t
Xbit_r196_c36 bl_36 br_36 wl_196 vdd gnd cell_6t
Xbit_r197_c36 bl_36 br_36 wl_197 vdd gnd cell_6t
Xbit_r198_c36 bl_36 br_36 wl_198 vdd gnd cell_6t
Xbit_r199_c36 bl_36 br_36 wl_199 vdd gnd cell_6t
Xbit_r200_c36 bl_36 br_36 wl_200 vdd gnd cell_6t
Xbit_r201_c36 bl_36 br_36 wl_201 vdd gnd cell_6t
Xbit_r202_c36 bl_36 br_36 wl_202 vdd gnd cell_6t
Xbit_r203_c36 bl_36 br_36 wl_203 vdd gnd cell_6t
Xbit_r204_c36 bl_36 br_36 wl_204 vdd gnd cell_6t
Xbit_r205_c36 bl_36 br_36 wl_205 vdd gnd cell_6t
Xbit_r206_c36 bl_36 br_36 wl_206 vdd gnd cell_6t
Xbit_r207_c36 bl_36 br_36 wl_207 vdd gnd cell_6t
Xbit_r208_c36 bl_36 br_36 wl_208 vdd gnd cell_6t
Xbit_r209_c36 bl_36 br_36 wl_209 vdd gnd cell_6t
Xbit_r210_c36 bl_36 br_36 wl_210 vdd gnd cell_6t
Xbit_r211_c36 bl_36 br_36 wl_211 vdd gnd cell_6t
Xbit_r212_c36 bl_36 br_36 wl_212 vdd gnd cell_6t
Xbit_r213_c36 bl_36 br_36 wl_213 vdd gnd cell_6t
Xbit_r214_c36 bl_36 br_36 wl_214 vdd gnd cell_6t
Xbit_r215_c36 bl_36 br_36 wl_215 vdd gnd cell_6t
Xbit_r216_c36 bl_36 br_36 wl_216 vdd gnd cell_6t
Xbit_r217_c36 bl_36 br_36 wl_217 vdd gnd cell_6t
Xbit_r218_c36 bl_36 br_36 wl_218 vdd gnd cell_6t
Xbit_r219_c36 bl_36 br_36 wl_219 vdd gnd cell_6t
Xbit_r220_c36 bl_36 br_36 wl_220 vdd gnd cell_6t
Xbit_r221_c36 bl_36 br_36 wl_221 vdd gnd cell_6t
Xbit_r222_c36 bl_36 br_36 wl_222 vdd gnd cell_6t
Xbit_r223_c36 bl_36 br_36 wl_223 vdd gnd cell_6t
Xbit_r224_c36 bl_36 br_36 wl_224 vdd gnd cell_6t
Xbit_r225_c36 bl_36 br_36 wl_225 vdd gnd cell_6t
Xbit_r226_c36 bl_36 br_36 wl_226 vdd gnd cell_6t
Xbit_r227_c36 bl_36 br_36 wl_227 vdd gnd cell_6t
Xbit_r228_c36 bl_36 br_36 wl_228 vdd gnd cell_6t
Xbit_r229_c36 bl_36 br_36 wl_229 vdd gnd cell_6t
Xbit_r230_c36 bl_36 br_36 wl_230 vdd gnd cell_6t
Xbit_r231_c36 bl_36 br_36 wl_231 vdd gnd cell_6t
Xbit_r232_c36 bl_36 br_36 wl_232 vdd gnd cell_6t
Xbit_r233_c36 bl_36 br_36 wl_233 vdd gnd cell_6t
Xbit_r234_c36 bl_36 br_36 wl_234 vdd gnd cell_6t
Xbit_r235_c36 bl_36 br_36 wl_235 vdd gnd cell_6t
Xbit_r236_c36 bl_36 br_36 wl_236 vdd gnd cell_6t
Xbit_r237_c36 bl_36 br_36 wl_237 vdd gnd cell_6t
Xbit_r238_c36 bl_36 br_36 wl_238 vdd gnd cell_6t
Xbit_r239_c36 bl_36 br_36 wl_239 vdd gnd cell_6t
Xbit_r240_c36 bl_36 br_36 wl_240 vdd gnd cell_6t
Xbit_r241_c36 bl_36 br_36 wl_241 vdd gnd cell_6t
Xbit_r242_c36 bl_36 br_36 wl_242 vdd gnd cell_6t
Xbit_r243_c36 bl_36 br_36 wl_243 vdd gnd cell_6t
Xbit_r244_c36 bl_36 br_36 wl_244 vdd gnd cell_6t
Xbit_r245_c36 bl_36 br_36 wl_245 vdd gnd cell_6t
Xbit_r246_c36 bl_36 br_36 wl_246 vdd gnd cell_6t
Xbit_r247_c36 bl_36 br_36 wl_247 vdd gnd cell_6t
Xbit_r248_c36 bl_36 br_36 wl_248 vdd gnd cell_6t
Xbit_r249_c36 bl_36 br_36 wl_249 vdd gnd cell_6t
Xbit_r250_c36 bl_36 br_36 wl_250 vdd gnd cell_6t
Xbit_r251_c36 bl_36 br_36 wl_251 vdd gnd cell_6t
Xbit_r252_c36 bl_36 br_36 wl_252 vdd gnd cell_6t
Xbit_r253_c36 bl_36 br_36 wl_253 vdd gnd cell_6t
Xbit_r254_c36 bl_36 br_36 wl_254 vdd gnd cell_6t
Xbit_r255_c36 bl_36 br_36 wl_255 vdd gnd cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd cell_6t
Xbit_r1_c37 bl_37 br_37 wl_1 vdd gnd cell_6t
Xbit_r2_c37 bl_37 br_37 wl_2 vdd gnd cell_6t
Xbit_r3_c37 bl_37 br_37 wl_3 vdd gnd cell_6t
Xbit_r4_c37 bl_37 br_37 wl_4 vdd gnd cell_6t
Xbit_r5_c37 bl_37 br_37 wl_5 vdd gnd cell_6t
Xbit_r6_c37 bl_37 br_37 wl_6 vdd gnd cell_6t
Xbit_r7_c37 bl_37 br_37 wl_7 vdd gnd cell_6t
Xbit_r8_c37 bl_37 br_37 wl_8 vdd gnd cell_6t
Xbit_r9_c37 bl_37 br_37 wl_9 vdd gnd cell_6t
Xbit_r10_c37 bl_37 br_37 wl_10 vdd gnd cell_6t
Xbit_r11_c37 bl_37 br_37 wl_11 vdd gnd cell_6t
Xbit_r12_c37 bl_37 br_37 wl_12 vdd gnd cell_6t
Xbit_r13_c37 bl_37 br_37 wl_13 vdd gnd cell_6t
Xbit_r14_c37 bl_37 br_37 wl_14 vdd gnd cell_6t
Xbit_r15_c37 bl_37 br_37 wl_15 vdd gnd cell_6t
Xbit_r16_c37 bl_37 br_37 wl_16 vdd gnd cell_6t
Xbit_r17_c37 bl_37 br_37 wl_17 vdd gnd cell_6t
Xbit_r18_c37 bl_37 br_37 wl_18 vdd gnd cell_6t
Xbit_r19_c37 bl_37 br_37 wl_19 vdd gnd cell_6t
Xbit_r20_c37 bl_37 br_37 wl_20 vdd gnd cell_6t
Xbit_r21_c37 bl_37 br_37 wl_21 vdd gnd cell_6t
Xbit_r22_c37 bl_37 br_37 wl_22 vdd gnd cell_6t
Xbit_r23_c37 bl_37 br_37 wl_23 vdd gnd cell_6t
Xbit_r24_c37 bl_37 br_37 wl_24 vdd gnd cell_6t
Xbit_r25_c37 bl_37 br_37 wl_25 vdd gnd cell_6t
Xbit_r26_c37 bl_37 br_37 wl_26 vdd gnd cell_6t
Xbit_r27_c37 bl_37 br_37 wl_27 vdd gnd cell_6t
Xbit_r28_c37 bl_37 br_37 wl_28 vdd gnd cell_6t
Xbit_r29_c37 bl_37 br_37 wl_29 vdd gnd cell_6t
Xbit_r30_c37 bl_37 br_37 wl_30 vdd gnd cell_6t
Xbit_r31_c37 bl_37 br_37 wl_31 vdd gnd cell_6t
Xbit_r32_c37 bl_37 br_37 wl_32 vdd gnd cell_6t
Xbit_r33_c37 bl_37 br_37 wl_33 vdd gnd cell_6t
Xbit_r34_c37 bl_37 br_37 wl_34 vdd gnd cell_6t
Xbit_r35_c37 bl_37 br_37 wl_35 vdd gnd cell_6t
Xbit_r36_c37 bl_37 br_37 wl_36 vdd gnd cell_6t
Xbit_r37_c37 bl_37 br_37 wl_37 vdd gnd cell_6t
Xbit_r38_c37 bl_37 br_37 wl_38 vdd gnd cell_6t
Xbit_r39_c37 bl_37 br_37 wl_39 vdd gnd cell_6t
Xbit_r40_c37 bl_37 br_37 wl_40 vdd gnd cell_6t
Xbit_r41_c37 bl_37 br_37 wl_41 vdd gnd cell_6t
Xbit_r42_c37 bl_37 br_37 wl_42 vdd gnd cell_6t
Xbit_r43_c37 bl_37 br_37 wl_43 vdd gnd cell_6t
Xbit_r44_c37 bl_37 br_37 wl_44 vdd gnd cell_6t
Xbit_r45_c37 bl_37 br_37 wl_45 vdd gnd cell_6t
Xbit_r46_c37 bl_37 br_37 wl_46 vdd gnd cell_6t
Xbit_r47_c37 bl_37 br_37 wl_47 vdd gnd cell_6t
Xbit_r48_c37 bl_37 br_37 wl_48 vdd gnd cell_6t
Xbit_r49_c37 bl_37 br_37 wl_49 vdd gnd cell_6t
Xbit_r50_c37 bl_37 br_37 wl_50 vdd gnd cell_6t
Xbit_r51_c37 bl_37 br_37 wl_51 vdd gnd cell_6t
Xbit_r52_c37 bl_37 br_37 wl_52 vdd gnd cell_6t
Xbit_r53_c37 bl_37 br_37 wl_53 vdd gnd cell_6t
Xbit_r54_c37 bl_37 br_37 wl_54 vdd gnd cell_6t
Xbit_r55_c37 bl_37 br_37 wl_55 vdd gnd cell_6t
Xbit_r56_c37 bl_37 br_37 wl_56 vdd gnd cell_6t
Xbit_r57_c37 bl_37 br_37 wl_57 vdd gnd cell_6t
Xbit_r58_c37 bl_37 br_37 wl_58 vdd gnd cell_6t
Xbit_r59_c37 bl_37 br_37 wl_59 vdd gnd cell_6t
Xbit_r60_c37 bl_37 br_37 wl_60 vdd gnd cell_6t
Xbit_r61_c37 bl_37 br_37 wl_61 vdd gnd cell_6t
Xbit_r62_c37 bl_37 br_37 wl_62 vdd gnd cell_6t
Xbit_r63_c37 bl_37 br_37 wl_63 vdd gnd cell_6t
Xbit_r64_c37 bl_37 br_37 wl_64 vdd gnd cell_6t
Xbit_r65_c37 bl_37 br_37 wl_65 vdd gnd cell_6t
Xbit_r66_c37 bl_37 br_37 wl_66 vdd gnd cell_6t
Xbit_r67_c37 bl_37 br_37 wl_67 vdd gnd cell_6t
Xbit_r68_c37 bl_37 br_37 wl_68 vdd gnd cell_6t
Xbit_r69_c37 bl_37 br_37 wl_69 vdd gnd cell_6t
Xbit_r70_c37 bl_37 br_37 wl_70 vdd gnd cell_6t
Xbit_r71_c37 bl_37 br_37 wl_71 vdd gnd cell_6t
Xbit_r72_c37 bl_37 br_37 wl_72 vdd gnd cell_6t
Xbit_r73_c37 bl_37 br_37 wl_73 vdd gnd cell_6t
Xbit_r74_c37 bl_37 br_37 wl_74 vdd gnd cell_6t
Xbit_r75_c37 bl_37 br_37 wl_75 vdd gnd cell_6t
Xbit_r76_c37 bl_37 br_37 wl_76 vdd gnd cell_6t
Xbit_r77_c37 bl_37 br_37 wl_77 vdd gnd cell_6t
Xbit_r78_c37 bl_37 br_37 wl_78 vdd gnd cell_6t
Xbit_r79_c37 bl_37 br_37 wl_79 vdd gnd cell_6t
Xbit_r80_c37 bl_37 br_37 wl_80 vdd gnd cell_6t
Xbit_r81_c37 bl_37 br_37 wl_81 vdd gnd cell_6t
Xbit_r82_c37 bl_37 br_37 wl_82 vdd gnd cell_6t
Xbit_r83_c37 bl_37 br_37 wl_83 vdd gnd cell_6t
Xbit_r84_c37 bl_37 br_37 wl_84 vdd gnd cell_6t
Xbit_r85_c37 bl_37 br_37 wl_85 vdd gnd cell_6t
Xbit_r86_c37 bl_37 br_37 wl_86 vdd gnd cell_6t
Xbit_r87_c37 bl_37 br_37 wl_87 vdd gnd cell_6t
Xbit_r88_c37 bl_37 br_37 wl_88 vdd gnd cell_6t
Xbit_r89_c37 bl_37 br_37 wl_89 vdd gnd cell_6t
Xbit_r90_c37 bl_37 br_37 wl_90 vdd gnd cell_6t
Xbit_r91_c37 bl_37 br_37 wl_91 vdd gnd cell_6t
Xbit_r92_c37 bl_37 br_37 wl_92 vdd gnd cell_6t
Xbit_r93_c37 bl_37 br_37 wl_93 vdd gnd cell_6t
Xbit_r94_c37 bl_37 br_37 wl_94 vdd gnd cell_6t
Xbit_r95_c37 bl_37 br_37 wl_95 vdd gnd cell_6t
Xbit_r96_c37 bl_37 br_37 wl_96 vdd gnd cell_6t
Xbit_r97_c37 bl_37 br_37 wl_97 vdd gnd cell_6t
Xbit_r98_c37 bl_37 br_37 wl_98 vdd gnd cell_6t
Xbit_r99_c37 bl_37 br_37 wl_99 vdd gnd cell_6t
Xbit_r100_c37 bl_37 br_37 wl_100 vdd gnd cell_6t
Xbit_r101_c37 bl_37 br_37 wl_101 vdd gnd cell_6t
Xbit_r102_c37 bl_37 br_37 wl_102 vdd gnd cell_6t
Xbit_r103_c37 bl_37 br_37 wl_103 vdd gnd cell_6t
Xbit_r104_c37 bl_37 br_37 wl_104 vdd gnd cell_6t
Xbit_r105_c37 bl_37 br_37 wl_105 vdd gnd cell_6t
Xbit_r106_c37 bl_37 br_37 wl_106 vdd gnd cell_6t
Xbit_r107_c37 bl_37 br_37 wl_107 vdd gnd cell_6t
Xbit_r108_c37 bl_37 br_37 wl_108 vdd gnd cell_6t
Xbit_r109_c37 bl_37 br_37 wl_109 vdd gnd cell_6t
Xbit_r110_c37 bl_37 br_37 wl_110 vdd gnd cell_6t
Xbit_r111_c37 bl_37 br_37 wl_111 vdd gnd cell_6t
Xbit_r112_c37 bl_37 br_37 wl_112 vdd gnd cell_6t
Xbit_r113_c37 bl_37 br_37 wl_113 vdd gnd cell_6t
Xbit_r114_c37 bl_37 br_37 wl_114 vdd gnd cell_6t
Xbit_r115_c37 bl_37 br_37 wl_115 vdd gnd cell_6t
Xbit_r116_c37 bl_37 br_37 wl_116 vdd gnd cell_6t
Xbit_r117_c37 bl_37 br_37 wl_117 vdd gnd cell_6t
Xbit_r118_c37 bl_37 br_37 wl_118 vdd gnd cell_6t
Xbit_r119_c37 bl_37 br_37 wl_119 vdd gnd cell_6t
Xbit_r120_c37 bl_37 br_37 wl_120 vdd gnd cell_6t
Xbit_r121_c37 bl_37 br_37 wl_121 vdd gnd cell_6t
Xbit_r122_c37 bl_37 br_37 wl_122 vdd gnd cell_6t
Xbit_r123_c37 bl_37 br_37 wl_123 vdd gnd cell_6t
Xbit_r124_c37 bl_37 br_37 wl_124 vdd gnd cell_6t
Xbit_r125_c37 bl_37 br_37 wl_125 vdd gnd cell_6t
Xbit_r126_c37 bl_37 br_37 wl_126 vdd gnd cell_6t
Xbit_r127_c37 bl_37 br_37 wl_127 vdd gnd cell_6t
Xbit_r128_c37 bl_37 br_37 wl_128 vdd gnd cell_6t
Xbit_r129_c37 bl_37 br_37 wl_129 vdd gnd cell_6t
Xbit_r130_c37 bl_37 br_37 wl_130 vdd gnd cell_6t
Xbit_r131_c37 bl_37 br_37 wl_131 vdd gnd cell_6t
Xbit_r132_c37 bl_37 br_37 wl_132 vdd gnd cell_6t
Xbit_r133_c37 bl_37 br_37 wl_133 vdd gnd cell_6t
Xbit_r134_c37 bl_37 br_37 wl_134 vdd gnd cell_6t
Xbit_r135_c37 bl_37 br_37 wl_135 vdd gnd cell_6t
Xbit_r136_c37 bl_37 br_37 wl_136 vdd gnd cell_6t
Xbit_r137_c37 bl_37 br_37 wl_137 vdd gnd cell_6t
Xbit_r138_c37 bl_37 br_37 wl_138 vdd gnd cell_6t
Xbit_r139_c37 bl_37 br_37 wl_139 vdd gnd cell_6t
Xbit_r140_c37 bl_37 br_37 wl_140 vdd gnd cell_6t
Xbit_r141_c37 bl_37 br_37 wl_141 vdd gnd cell_6t
Xbit_r142_c37 bl_37 br_37 wl_142 vdd gnd cell_6t
Xbit_r143_c37 bl_37 br_37 wl_143 vdd gnd cell_6t
Xbit_r144_c37 bl_37 br_37 wl_144 vdd gnd cell_6t
Xbit_r145_c37 bl_37 br_37 wl_145 vdd gnd cell_6t
Xbit_r146_c37 bl_37 br_37 wl_146 vdd gnd cell_6t
Xbit_r147_c37 bl_37 br_37 wl_147 vdd gnd cell_6t
Xbit_r148_c37 bl_37 br_37 wl_148 vdd gnd cell_6t
Xbit_r149_c37 bl_37 br_37 wl_149 vdd gnd cell_6t
Xbit_r150_c37 bl_37 br_37 wl_150 vdd gnd cell_6t
Xbit_r151_c37 bl_37 br_37 wl_151 vdd gnd cell_6t
Xbit_r152_c37 bl_37 br_37 wl_152 vdd gnd cell_6t
Xbit_r153_c37 bl_37 br_37 wl_153 vdd gnd cell_6t
Xbit_r154_c37 bl_37 br_37 wl_154 vdd gnd cell_6t
Xbit_r155_c37 bl_37 br_37 wl_155 vdd gnd cell_6t
Xbit_r156_c37 bl_37 br_37 wl_156 vdd gnd cell_6t
Xbit_r157_c37 bl_37 br_37 wl_157 vdd gnd cell_6t
Xbit_r158_c37 bl_37 br_37 wl_158 vdd gnd cell_6t
Xbit_r159_c37 bl_37 br_37 wl_159 vdd gnd cell_6t
Xbit_r160_c37 bl_37 br_37 wl_160 vdd gnd cell_6t
Xbit_r161_c37 bl_37 br_37 wl_161 vdd gnd cell_6t
Xbit_r162_c37 bl_37 br_37 wl_162 vdd gnd cell_6t
Xbit_r163_c37 bl_37 br_37 wl_163 vdd gnd cell_6t
Xbit_r164_c37 bl_37 br_37 wl_164 vdd gnd cell_6t
Xbit_r165_c37 bl_37 br_37 wl_165 vdd gnd cell_6t
Xbit_r166_c37 bl_37 br_37 wl_166 vdd gnd cell_6t
Xbit_r167_c37 bl_37 br_37 wl_167 vdd gnd cell_6t
Xbit_r168_c37 bl_37 br_37 wl_168 vdd gnd cell_6t
Xbit_r169_c37 bl_37 br_37 wl_169 vdd gnd cell_6t
Xbit_r170_c37 bl_37 br_37 wl_170 vdd gnd cell_6t
Xbit_r171_c37 bl_37 br_37 wl_171 vdd gnd cell_6t
Xbit_r172_c37 bl_37 br_37 wl_172 vdd gnd cell_6t
Xbit_r173_c37 bl_37 br_37 wl_173 vdd gnd cell_6t
Xbit_r174_c37 bl_37 br_37 wl_174 vdd gnd cell_6t
Xbit_r175_c37 bl_37 br_37 wl_175 vdd gnd cell_6t
Xbit_r176_c37 bl_37 br_37 wl_176 vdd gnd cell_6t
Xbit_r177_c37 bl_37 br_37 wl_177 vdd gnd cell_6t
Xbit_r178_c37 bl_37 br_37 wl_178 vdd gnd cell_6t
Xbit_r179_c37 bl_37 br_37 wl_179 vdd gnd cell_6t
Xbit_r180_c37 bl_37 br_37 wl_180 vdd gnd cell_6t
Xbit_r181_c37 bl_37 br_37 wl_181 vdd gnd cell_6t
Xbit_r182_c37 bl_37 br_37 wl_182 vdd gnd cell_6t
Xbit_r183_c37 bl_37 br_37 wl_183 vdd gnd cell_6t
Xbit_r184_c37 bl_37 br_37 wl_184 vdd gnd cell_6t
Xbit_r185_c37 bl_37 br_37 wl_185 vdd gnd cell_6t
Xbit_r186_c37 bl_37 br_37 wl_186 vdd gnd cell_6t
Xbit_r187_c37 bl_37 br_37 wl_187 vdd gnd cell_6t
Xbit_r188_c37 bl_37 br_37 wl_188 vdd gnd cell_6t
Xbit_r189_c37 bl_37 br_37 wl_189 vdd gnd cell_6t
Xbit_r190_c37 bl_37 br_37 wl_190 vdd gnd cell_6t
Xbit_r191_c37 bl_37 br_37 wl_191 vdd gnd cell_6t
Xbit_r192_c37 bl_37 br_37 wl_192 vdd gnd cell_6t
Xbit_r193_c37 bl_37 br_37 wl_193 vdd gnd cell_6t
Xbit_r194_c37 bl_37 br_37 wl_194 vdd gnd cell_6t
Xbit_r195_c37 bl_37 br_37 wl_195 vdd gnd cell_6t
Xbit_r196_c37 bl_37 br_37 wl_196 vdd gnd cell_6t
Xbit_r197_c37 bl_37 br_37 wl_197 vdd gnd cell_6t
Xbit_r198_c37 bl_37 br_37 wl_198 vdd gnd cell_6t
Xbit_r199_c37 bl_37 br_37 wl_199 vdd gnd cell_6t
Xbit_r200_c37 bl_37 br_37 wl_200 vdd gnd cell_6t
Xbit_r201_c37 bl_37 br_37 wl_201 vdd gnd cell_6t
Xbit_r202_c37 bl_37 br_37 wl_202 vdd gnd cell_6t
Xbit_r203_c37 bl_37 br_37 wl_203 vdd gnd cell_6t
Xbit_r204_c37 bl_37 br_37 wl_204 vdd gnd cell_6t
Xbit_r205_c37 bl_37 br_37 wl_205 vdd gnd cell_6t
Xbit_r206_c37 bl_37 br_37 wl_206 vdd gnd cell_6t
Xbit_r207_c37 bl_37 br_37 wl_207 vdd gnd cell_6t
Xbit_r208_c37 bl_37 br_37 wl_208 vdd gnd cell_6t
Xbit_r209_c37 bl_37 br_37 wl_209 vdd gnd cell_6t
Xbit_r210_c37 bl_37 br_37 wl_210 vdd gnd cell_6t
Xbit_r211_c37 bl_37 br_37 wl_211 vdd gnd cell_6t
Xbit_r212_c37 bl_37 br_37 wl_212 vdd gnd cell_6t
Xbit_r213_c37 bl_37 br_37 wl_213 vdd gnd cell_6t
Xbit_r214_c37 bl_37 br_37 wl_214 vdd gnd cell_6t
Xbit_r215_c37 bl_37 br_37 wl_215 vdd gnd cell_6t
Xbit_r216_c37 bl_37 br_37 wl_216 vdd gnd cell_6t
Xbit_r217_c37 bl_37 br_37 wl_217 vdd gnd cell_6t
Xbit_r218_c37 bl_37 br_37 wl_218 vdd gnd cell_6t
Xbit_r219_c37 bl_37 br_37 wl_219 vdd gnd cell_6t
Xbit_r220_c37 bl_37 br_37 wl_220 vdd gnd cell_6t
Xbit_r221_c37 bl_37 br_37 wl_221 vdd gnd cell_6t
Xbit_r222_c37 bl_37 br_37 wl_222 vdd gnd cell_6t
Xbit_r223_c37 bl_37 br_37 wl_223 vdd gnd cell_6t
Xbit_r224_c37 bl_37 br_37 wl_224 vdd gnd cell_6t
Xbit_r225_c37 bl_37 br_37 wl_225 vdd gnd cell_6t
Xbit_r226_c37 bl_37 br_37 wl_226 vdd gnd cell_6t
Xbit_r227_c37 bl_37 br_37 wl_227 vdd gnd cell_6t
Xbit_r228_c37 bl_37 br_37 wl_228 vdd gnd cell_6t
Xbit_r229_c37 bl_37 br_37 wl_229 vdd gnd cell_6t
Xbit_r230_c37 bl_37 br_37 wl_230 vdd gnd cell_6t
Xbit_r231_c37 bl_37 br_37 wl_231 vdd gnd cell_6t
Xbit_r232_c37 bl_37 br_37 wl_232 vdd gnd cell_6t
Xbit_r233_c37 bl_37 br_37 wl_233 vdd gnd cell_6t
Xbit_r234_c37 bl_37 br_37 wl_234 vdd gnd cell_6t
Xbit_r235_c37 bl_37 br_37 wl_235 vdd gnd cell_6t
Xbit_r236_c37 bl_37 br_37 wl_236 vdd gnd cell_6t
Xbit_r237_c37 bl_37 br_37 wl_237 vdd gnd cell_6t
Xbit_r238_c37 bl_37 br_37 wl_238 vdd gnd cell_6t
Xbit_r239_c37 bl_37 br_37 wl_239 vdd gnd cell_6t
Xbit_r240_c37 bl_37 br_37 wl_240 vdd gnd cell_6t
Xbit_r241_c37 bl_37 br_37 wl_241 vdd gnd cell_6t
Xbit_r242_c37 bl_37 br_37 wl_242 vdd gnd cell_6t
Xbit_r243_c37 bl_37 br_37 wl_243 vdd gnd cell_6t
Xbit_r244_c37 bl_37 br_37 wl_244 vdd gnd cell_6t
Xbit_r245_c37 bl_37 br_37 wl_245 vdd gnd cell_6t
Xbit_r246_c37 bl_37 br_37 wl_246 vdd gnd cell_6t
Xbit_r247_c37 bl_37 br_37 wl_247 vdd gnd cell_6t
Xbit_r248_c37 bl_37 br_37 wl_248 vdd gnd cell_6t
Xbit_r249_c37 bl_37 br_37 wl_249 vdd gnd cell_6t
Xbit_r250_c37 bl_37 br_37 wl_250 vdd gnd cell_6t
Xbit_r251_c37 bl_37 br_37 wl_251 vdd gnd cell_6t
Xbit_r252_c37 bl_37 br_37 wl_252 vdd gnd cell_6t
Xbit_r253_c37 bl_37 br_37 wl_253 vdd gnd cell_6t
Xbit_r254_c37 bl_37 br_37 wl_254 vdd gnd cell_6t
Xbit_r255_c37 bl_37 br_37 wl_255 vdd gnd cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd cell_6t
Xbit_r1_c38 bl_38 br_38 wl_1 vdd gnd cell_6t
Xbit_r2_c38 bl_38 br_38 wl_2 vdd gnd cell_6t
Xbit_r3_c38 bl_38 br_38 wl_3 vdd gnd cell_6t
Xbit_r4_c38 bl_38 br_38 wl_4 vdd gnd cell_6t
Xbit_r5_c38 bl_38 br_38 wl_5 vdd gnd cell_6t
Xbit_r6_c38 bl_38 br_38 wl_6 vdd gnd cell_6t
Xbit_r7_c38 bl_38 br_38 wl_7 vdd gnd cell_6t
Xbit_r8_c38 bl_38 br_38 wl_8 vdd gnd cell_6t
Xbit_r9_c38 bl_38 br_38 wl_9 vdd gnd cell_6t
Xbit_r10_c38 bl_38 br_38 wl_10 vdd gnd cell_6t
Xbit_r11_c38 bl_38 br_38 wl_11 vdd gnd cell_6t
Xbit_r12_c38 bl_38 br_38 wl_12 vdd gnd cell_6t
Xbit_r13_c38 bl_38 br_38 wl_13 vdd gnd cell_6t
Xbit_r14_c38 bl_38 br_38 wl_14 vdd gnd cell_6t
Xbit_r15_c38 bl_38 br_38 wl_15 vdd gnd cell_6t
Xbit_r16_c38 bl_38 br_38 wl_16 vdd gnd cell_6t
Xbit_r17_c38 bl_38 br_38 wl_17 vdd gnd cell_6t
Xbit_r18_c38 bl_38 br_38 wl_18 vdd gnd cell_6t
Xbit_r19_c38 bl_38 br_38 wl_19 vdd gnd cell_6t
Xbit_r20_c38 bl_38 br_38 wl_20 vdd gnd cell_6t
Xbit_r21_c38 bl_38 br_38 wl_21 vdd gnd cell_6t
Xbit_r22_c38 bl_38 br_38 wl_22 vdd gnd cell_6t
Xbit_r23_c38 bl_38 br_38 wl_23 vdd gnd cell_6t
Xbit_r24_c38 bl_38 br_38 wl_24 vdd gnd cell_6t
Xbit_r25_c38 bl_38 br_38 wl_25 vdd gnd cell_6t
Xbit_r26_c38 bl_38 br_38 wl_26 vdd gnd cell_6t
Xbit_r27_c38 bl_38 br_38 wl_27 vdd gnd cell_6t
Xbit_r28_c38 bl_38 br_38 wl_28 vdd gnd cell_6t
Xbit_r29_c38 bl_38 br_38 wl_29 vdd gnd cell_6t
Xbit_r30_c38 bl_38 br_38 wl_30 vdd gnd cell_6t
Xbit_r31_c38 bl_38 br_38 wl_31 vdd gnd cell_6t
Xbit_r32_c38 bl_38 br_38 wl_32 vdd gnd cell_6t
Xbit_r33_c38 bl_38 br_38 wl_33 vdd gnd cell_6t
Xbit_r34_c38 bl_38 br_38 wl_34 vdd gnd cell_6t
Xbit_r35_c38 bl_38 br_38 wl_35 vdd gnd cell_6t
Xbit_r36_c38 bl_38 br_38 wl_36 vdd gnd cell_6t
Xbit_r37_c38 bl_38 br_38 wl_37 vdd gnd cell_6t
Xbit_r38_c38 bl_38 br_38 wl_38 vdd gnd cell_6t
Xbit_r39_c38 bl_38 br_38 wl_39 vdd gnd cell_6t
Xbit_r40_c38 bl_38 br_38 wl_40 vdd gnd cell_6t
Xbit_r41_c38 bl_38 br_38 wl_41 vdd gnd cell_6t
Xbit_r42_c38 bl_38 br_38 wl_42 vdd gnd cell_6t
Xbit_r43_c38 bl_38 br_38 wl_43 vdd gnd cell_6t
Xbit_r44_c38 bl_38 br_38 wl_44 vdd gnd cell_6t
Xbit_r45_c38 bl_38 br_38 wl_45 vdd gnd cell_6t
Xbit_r46_c38 bl_38 br_38 wl_46 vdd gnd cell_6t
Xbit_r47_c38 bl_38 br_38 wl_47 vdd gnd cell_6t
Xbit_r48_c38 bl_38 br_38 wl_48 vdd gnd cell_6t
Xbit_r49_c38 bl_38 br_38 wl_49 vdd gnd cell_6t
Xbit_r50_c38 bl_38 br_38 wl_50 vdd gnd cell_6t
Xbit_r51_c38 bl_38 br_38 wl_51 vdd gnd cell_6t
Xbit_r52_c38 bl_38 br_38 wl_52 vdd gnd cell_6t
Xbit_r53_c38 bl_38 br_38 wl_53 vdd gnd cell_6t
Xbit_r54_c38 bl_38 br_38 wl_54 vdd gnd cell_6t
Xbit_r55_c38 bl_38 br_38 wl_55 vdd gnd cell_6t
Xbit_r56_c38 bl_38 br_38 wl_56 vdd gnd cell_6t
Xbit_r57_c38 bl_38 br_38 wl_57 vdd gnd cell_6t
Xbit_r58_c38 bl_38 br_38 wl_58 vdd gnd cell_6t
Xbit_r59_c38 bl_38 br_38 wl_59 vdd gnd cell_6t
Xbit_r60_c38 bl_38 br_38 wl_60 vdd gnd cell_6t
Xbit_r61_c38 bl_38 br_38 wl_61 vdd gnd cell_6t
Xbit_r62_c38 bl_38 br_38 wl_62 vdd gnd cell_6t
Xbit_r63_c38 bl_38 br_38 wl_63 vdd gnd cell_6t
Xbit_r64_c38 bl_38 br_38 wl_64 vdd gnd cell_6t
Xbit_r65_c38 bl_38 br_38 wl_65 vdd gnd cell_6t
Xbit_r66_c38 bl_38 br_38 wl_66 vdd gnd cell_6t
Xbit_r67_c38 bl_38 br_38 wl_67 vdd gnd cell_6t
Xbit_r68_c38 bl_38 br_38 wl_68 vdd gnd cell_6t
Xbit_r69_c38 bl_38 br_38 wl_69 vdd gnd cell_6t
Xbit_r70_c38 bl_38 br_38 wl_70 vdd gnd cell_6t
Xbit_r71_c38 bl_38 br_38 wl_71 vdd gnd cell_6t
Xbit_r72_c38 bl_38 br_38 wl_72 vdd gnd cell_6t
Xbit_r73_c38 bl_38 br_38 wl_73 vdd gnd cell_6t
Xbit_r74_c38 bl_38 br_38 wl_74 vdd gnd cell_6t
Xbit_r75_c38 bl_38 br_38 wl_75 vdd gnd cell_6t
Xbit_r76_c38 bl_38 br_38 wl_76 vdd gnd cell_6t
Xbit_r77_c38 bl_38 br_38 wl_77 vdd gnd cell_6t
Xbit_r78_c38 bl_38 br_38 wl_78 vdd gnd cell_6t
Xbit_r79_c38 bl_38 br_38 wl_79 vdd gnd cell_6t
Xbit_r80_c38 bl_38 br_38 wl_80 vdd gnd cell_6t
Xbit_r81_c38 bl_38 br_38 wl_81 vdd gnd cell_6t
Xbit_r82_c38 bl_38 br_38 wl_82 vdd gnd cell_6t
Xbit_r83_c38 bl_38 br_38 wl_83 vdd gnd cell_6t
Xbit_r84_c38 bl_38 br_38 wl_84 vdd gnd cell_6t
Xbit_r85_c38 bl_38 br_38 wl_85 vdd gnd cell_6t
Xbit_r86_c38 bl_38 br_38 wl_86 vdd gnd cell_6t
Xbit_r87_c38 bl_38 br_38 wl_87 vdd gnd cell_6t
Xbit_r88_c38 bl_38 br_38 wl_88 vdd gnd cell_6t
Xbit_r89_c38 bl_38 br_38 wl_89 vdd gnd cell_6t
Xbit_r90_c38 bl_38 br_38 wl_90 vdd gnd cell_6t
Xbit_r91_c38 bl_38 br_38 wl_91 vdd gnd cell_6t
Xbit_r92_c38 bl_38 br_38 wl_92 vdd gnd cell_6t
Xbit_r93_c38 bl_38 br_38 wl_93 vdd gnd cell_6t
Xbit_r94_c38 bl_38 br_38 wl_94 vdd gnd cell_6t
Xbit_r95_c38 bl_38 br_38 wl_95 vdd gnd cell_6t
Xbit_r96_c38 bl_38 br_38 wl_96 vdd gnd cell_6t
Xbit_r97_c38 bl_38 br_38 wl_97 vdd gnd cell_6t
Xbit_r98_c38 bl_38 br_38 wl_98 vdd gnd cell_6t
Xbit_r99_c38 bl_38 br_38 wl_99 vdd gnd cell_6t
Xbit_r100_c38 bl_38 br_38 wl_100 vdd gnd cell_6t
Xbit_r101_c38 bl_38 br_38 wl_101 vdd gnd cell_6t
Xbit_r102_c38 bl_38 br_38 wl_102 vdd gnd cell_6t
Xbit_r103_c38 bl_38 br_38 wl_103 vdd gnd cell_6t
Xbit_r104_c38 bl_38 br_38 wl_104 vdd gnd cell_6t
Xbit_r105_c38 bl_38 br_38 wl_105 vdd gnd cell_6t
Xbit_r106_c38 bl_38 br_38 wl_106 vdd gnd cell_6t
Xbit_r107_c38 bl_38 br_38 wl_107 vdd gnd cell_6t
Xbit_r108_c38 bl_38 br_38 wl_108 vdd gnd cell_6t
Xbit_r109_c38 bl_38 br_38 wl_109 vdd gnd cell_6t
Xbit_r110_c38 bl_38 br_38 wl_110 vdd gnd cell_6t
Xbit_r111_c38 bl_38 br_38 wl_111 vdd gnd cell_6t
Xbit_r112_c38 bl_38 br_38 wl_112 vdd gnd cell_6t
Xbit_r113_c38 bl_38 br_38 wl_113 vdd gnd cell_6t
Xbit_r114_c38 bl_38 br_38 wl_114 vdd gnd cell_6t
Xbit_r115_c38 bl_38 br_38 wl_115 vdd gnd cell_6t
Xbit_r116_c38 bl_38 br_38 wl_116 vdd gnd cell_6t
Xbit_r117_c38 bl_38 br_38 wl_117 vdd gnd cell_6t
Xbit_r118_c38 bl_38 br_38 wl_118 vdd gnd cell_6t
Xbit_r119_c38 bl_38 br_38 wl_119 vdd gnd cell_6t
Xbit_r120_c38 bl_38 br_38 wl_120 vdd gnd cell_6t
Xbit_r121_c38 bl_38 br_38 wl_121 vdd gnd cell_6t
Xbit_r122_c38 bl_38 br_38 wl_122 vdd gnd cell_6t
Xbit_r123_c38 bl_38 br_38 wl_123 vdd gnd cell_6t
Xbit_r124_c38 bl_38 br_38 wl_124 vdd gnd cell_6t
Xbit_r125_c38 bl_38 br_38 wl_125 vdd gnd cell_6t
Xbit_r126_c38 bl_38 br_38 wl_126 vdd gnd cell_6t
Xbit_r127_c38 bl_38 br_38 wl_127 vdd gnd cell_6t
Xbit_r128_c38 bl_38 br_38 wl_128 vdd gnd cell_6t
Xbit_r129_c38 bl_38 br_38 wl_129 vdd gnd cell_6t
Xbit_r130_c38 bl_38 br_38 wl_130 vdd gnd cell_6t
Xbit_r131_c38 bl_38 br_38 wl_131 vdd gnd cell_6t
Xbit_r132_c38 bl_38 br_38 wl_132 vdd gnd cell_6t
Xbit_r133_c38 bl_38 br_38 wl_133 vdd gnd cell_6t
Xbit_r134_c38 bl_38 br_38 wl_134 vdd gnd cell_6t
Xbit_r135_c38 bl_38 br_38 wl_135 vdd gnd cell_6t
Xbit_r136_c38 bl_38 br_38 wl_136 vdd gnd cell_6t
Xbit_r137_c38 bl_38 br_38 wl_137 vdd gnd cell_6t
Xbit_r138_c38 bl_38 br_38 wl_138 vdd gnd cell_6t
Xbit_r139_c38 bl_38 br_38 wl_139 vdd gnd cell_6t
Xbit_r140_c38 bl_38 br_38 wl_140 vdd gnd cell_6t
Xbit_r141_c38 bl_38 br_38 wl_141 vdd gnd cell_6t
Xbit_r142_c38 bl_38 br_38 wl_142 vdd gnd cell_6t
Xbit_r143_c38 bl_38 br_38 wl_143 vdd gnd cell_6t
Xbit_r144_c38 bl_38 br_38 wl_144 vdd gnd cell_6t
Xbit_r145_c38 bl_38 br_38 wl_145 vdd gnd cell_6t
Xbit_r146_c38 bl_38 br_38 wl_146 vdd gnd cell_6t
Xbit_r147_c38 bl_38 br_38 wl_147 vdd gnd cell_6t
Xbit_r148_c38 bl_38 br_38 wl_148 vdd gnd cell_6t
Xbit_r149_c38 bl_38 br_38 wl_149 vdd gnd cell_6t
Xbit_r150_c38 bl_38 br_38 wl_150 vdd gnd cell_6t
Xbit_r151_c38 bl_38 br_38 wl_151 vdd gnd cell_6t
Xbit_r152_c38 bl_38 br_38 wl_152 vdd gnd cell_6t
Xbit_r153_c38 bl_38 br_38 wl_153 vdd gnd cell_6t
Xbit_r154_c38 bl_38 br_38 wl_154 vdd gnd cell_6t
Xbit_r155_c38 bl_38 br_38 wl_155 vdd gnd cell_6t
Xbit_r156_c38 bl_38 br_38 wl_156 vdd gnd cell_6t
Xbit_r157_c38 bl_38 br_38 wl_157 vdd gnd cell_6t
Xbit_r158_c38 bl_38 br_38 wl_158 vdd gnd cell_6t
Xbit_r159_c38 bl_38 br_38 wl_159 vdd gnd cell_6t
Xbit_r160_c38 bl_38 br_38 wl_160 vdd gnd cell_6t
Xbit_r161_c38 bl_38 br_38 wl_161 vdd gnd cell_6t
Xbit_r162_c38 bl_38 br_38 wl_162 vdd gnd cell_6t
Xbit_r163_c38 bl_38 br_38 wl_163 vdd gnd cell_6t
Xbit_r164_c38 bl_38 br_38 wl_164 vdd gnd cell_6t
Xbit_r165_c38 bl_38 br_38 wl_165 vdd gnd cell_6t
Xbit_r166_c38 bl_38 br_38 wl_166 vdd gnd cell_6t
Xbit_r167_c38 bl_38 br_38 wl_167 vdd gnd cell_6t
Xbit_r168_c38 bl_38 br_38 wl_168 vdd gnd cell_6t
Xbit_r169_c38 bl_38 br_38 wl_169 vdd gnd cell_6t
Xbit_r170_c38 bl_38 br_38 wl_170 vdd gnd cell_6t
Xbit_r171_c38 bl_38 br_38 wl_171 vdd gnd cell_6t
Xbit_r172_c38 bl_38 br_38 wl_172 vdd gnd cell_6t
Xbit_r173_c38 bl_38 br_38 wl_173 vdd gnd cell_6t
Xbit_r174_c38 bl_38 br_38 wl_174 vdd gnd cell_6t
Xbit_r175_c38 bl_38 br_38 wl_175 vdd gnd cell_6t
Xbit_r176_c38 bl_38 br_38 wl_176 vdd gnd cell_6t
Xbit_r177_c38 bl_38 br_38 wl_177 vdd gnd cell_6t
Xbit_r178_c38 bl_38 br_38 wl_178 vdd gnd cell_6t
Xbit_r179_c38 bl_38 br_38 wl_179 vdd gnd cell_6t
Xbit_r180_c38 bl_38 br_38 wl_180 vdd gnd cell_6t
Xbit_r181_c38 bl_38 br_38 wl_181 vdd gnd cell_6t
Xbit_r182_c38 bl_38 br_38 wl_182 vdd gnd cell_6t
Xbit_r183_c38 bl_38 br_38 wl_183 vdd gnd cell_6t
Xbit_r184_c38 bl_38 br_38 wl_184 vdd gnd cell_6t
Xbit_r185_c38 bl_38 br_38 wl_185 vdd gnd cell_6t
Xbit_r186_c38 bl_38 br_38 wl_186 vdd gnd cell_6t
Xbit_r187_c38 bl_38 br_38 wl_187 vdd gnd cell_6t
Xbit_r188_c38 bl_38 br_38 wl_188 vdd gnd cell_6t
Xbit_r189_c38 bl_38 br_38 wl_189 vdd gnd cell_6t
Xbit_r190_c38 bl_38 br_38 wl_190 vdd gnd cell_6t
Xbit_r191_c38 bl_38 br_38 wl_191 vdd gnd cell_6t
Xbit_r192_c38 bl_38 br_38 wl_192 vdd gnd cell_6t
Xbit_r193_c38 bl_38 br_38 wl_193 vdd gnd cell_6t
Xbit_r194_c38 bl_38 br_38 wl_194 vdd gnd cell_6t
Xbit_r195_c38 bl_38 br_38 wl_195 vdd gnd cell_6t
Xbit_r196_c38 bl_38 br_38 wl_196 vdd gnd cell_6t
Xbit_r197_c38 bl_38 br_38 wl_197 vdd gnd cell_6t
Xbit_r198_c38 bl_38 br_38 wl_198 vdd gnd cell_6t
Xbit_r199_c38 bl_38 br_38 wl_199 vdd gnd cell_6t
Xbit_r200_c38 bl_38 br_38 wl_200 vdd gnd cell_6t
Xbit_r201_c38 bl_38 br_38 wl_201 vdd gnd cell_6t
Xbit_r202_c38 bl_38 br_38 wl_202 vdd gnd cell_6t
Xbit_r203_c38 bl_38 br_38 wl_203 vdd gnd cell_6t
Xbit_r204_c38 bl_38 br_38 wl_204 vdd gnd cell_6t
Xbit_r205_c38 bl_38 br_38 wl_205 vdd gnd cell_6t
Xbit_r206_c38 bl_38 br_38 wl_206 vdd gnd cell_6t
Xbit_r207_c38 bl_38 br_38 wl_207 vdd gnd cell_6t
Xbit_r208_c38 bl_38 br_38 wl_208 vdd gnd cell_6t
Xbit_r209_c38 bl_38 br_38 wl_209 vdd gnd cell_6t
Xbit_r210_c38 bl_38 br_38 wl_210 vdd gnd cell_6t
Xbit_r211_c38 bl_38 br_38 wl_211 vdd gnd cell_6t
Xbit_r212_c38 bl_38 br_38 wl_212 vdd gnd cell_6t
Xbit_r213_c38 bl_38 br_38 wl_213 vdd gnd cell_6t
Xbit_r214_c38 bl_38 br_38 wl_214 vdd gnd cell_6t
Xbit_r215_c38 bl_38 br_38 wl_215 vdd gnd cell_6t
Xbit_r216_c38 bl_38 br_38 wl_216 vdd gnd cell_6t
Xbit_r217_c38 bl_38 br_38 wl_217 vdd gnd cell_6t
Xbit_r218_c38 bl_38 br_38 wl_218 vdd gnd cell_6t
Xbit_r219_c38 bl_38 br_38 wl_219 vdd gnd cell_6t
Xbit_r220_c38 bl_38 br_38 wl_220 vdd gnd cell_6t
Xbit_r221_c38 bl_38 br_38 wl_221 vdd gnd cell_6t
Xbit_r222_c38 bl_38 br_38 wl_222 vdd gnd cell_6t
Xbit_r223_c38 bl_38 br_38 wl_223 vdd gnd cell_6t
Xbit_r224_c38 bl_38 br_38 wl_224 vdd gnd cell_6t
Xbit_r225_c38 bl_38 br_38 wl_225 vdd gnd cell_6t
Xbit_r226_c38 bl_38 br_38 wl_226 vdd gnd cell_6t
Xbit_r227_c38 bl_38 br_38 wl_227 vdd gnd cell_6t
Xbit_r228_c38 bl_38 br_38 wl_228 vdd gnd cell_6t
Xbit_r229_c38 bl_38 br_38 wl_229 vdd gnd cell_6t
Xbit_r230_c38 bl_38 br_38 wl_230 vdd gnd cell_6t
Xbit_r231_c38 bl_38 br_38 wl_231 vdd gnd cell_6t
Xbit_r232_c38 bl_38 br_38 wl_232 vdd gnd cell_6t
Xbit_r233_c38 bl_38 br_38 wl_233 vdd gnd cell_6t
Xbit_r234_c38 bl_38 br_38 wl_234 vdd gnd cell_6t
Xbit_r235_c38 bl_38 br_38 wl_235 vdd gnd cell_6t
Xbit_r236_c38 bl_38 br_38 wl_236 vdd gnd cell_6t
Xbit_r237_c38 bl_38 br_38 wl_237 vdd gnd cell_6t
Xbit_r238_c38 bl_38 br_38 wl_238 vdd gnd cell_6t
Xbit_r239_c38 bl_38 br_38 wl_239 vdd gnd cell_6t
Xbit_r240_c38 bl_38 br_38 wl_240 vdd gnd cell_6t
Xbit_r241_c38 bl_38 br_38 wl_241 vdd gnd cell_6t
Xbit_r242_c38 bl_38 br_38 wl_242 vdd gnd cell_6t
Xbit_r243_c38 bl_38 br_38 wl_243 vdd gnd cell_6t
Xbit_r244_c38 bl_38 br_38 wl_244 vdd gnd cell_6t
Xbit_r245_c38 bl_38 br_38 wl_245 vdd gnd cell_6t
Xbit_r246_c38 bl_38 br_38 wl_246 vdd gnd cell_6t
Xbit_r247_c38 bl_38 br_38 wl_247 vdd gnd cell_6t
Xbit_r248_c38 bl_38 br_38 wl_248 vdd gnd cell_6t
Xbit_r249_c38 bl_38 br_38 wl_249 vdd gnd cell_6t
Xbit_r250_c38 bl_38 br_38 wl_250 vdd gnd cell_6t
Xbit_r251_c38 bl_38 br_38 wl_251 vdd gnd cell_6t
Xbit_r252_c38 bl_38 br_38 wl_252 vdd gnd cell_6t
Xbit_r253_c38 bl_38 br_38 wl_253 vdd gnd cell_6t
Xbit_r254_c38 bl_38 br_38 wl_254 vdd gnd cell_6t
Xbit_r255_c38 bl_38 br_38 wl_255 vdd gnd cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd cell_6t
Xbit_r1_c39 bl_39 br_39 wl_1 vdd gnd cell_6t
Xbit_r2_c39 bl_39 br_39 wl_2 vdd gnd cell_6t
Xbit_r3_c39 bl_39 br_39 wl_3 vdd gnd cell_6t
Xbit_r4_c39 bl_39 br_39 wl_4 vdd gnd cell_6t
Xbit_r5_c39 bl_39 br_39 wl_5 vdd gnd cell_6t
Xbit_r6_c39 bl_39 br_39 wl_6 vdd gnd cell_6t
Xbit_r7_c39 bl_39 br_39 wl_7 vdd gnd cell_6t
Xbit_r8_c39 bl_39 br_39 wl_8 vdd gnd cell_6t
Xbit_r9_c39 bl_39 br_39 wl_9 vdd gnd cell_6t
Xbit_r10_c39 bl_39 br_39 wl_10 vdd gnd cell_6t
Xbit_r11_c39 bl_39 br_39 wl_11 vdd gnd cell_6t
Xbit_r12_c39 bl_39 br_39 wl_12 vdd gnd cell_6t
Xbit_r13_c39 bl_39 br_39 wl_13 vdd gnd cell_6t
Xbit_r14_c39 bl_39 br_39 wl_14 vdd gnd cell_6t
Xbit_r15_c39 bl_39 br_39 wl_15 vdd gnd cell_6t
Xbit_r16_c39 bl_39 br_39 wl_16 vdd gnd cell_6t
Xbit_r17_c39 bl_39 br_39 wl_17 vdd gnd cell_6t
Xbit_r18_c39 bl_39 br_39 wl_18 vdd gnd cell_6t
Xbit_r19_c39 bl_39 br_39 wl_19 vdd gnd cell_6t
Xbit_r20_c39 bl_39 br_39 wl_20 vdd gnd cell_6t
Xbit_r21_c39 bl_39 br_39 wl_21 vdd gnd cell_6t
Xbit_r22_c39 bl_39 br_39 wl_22 vdd gnd cell_6t
Xbit_r23_c39 bl_39 br_39 wl_23 vdd gnd cell_6t
Xbit_r24_c39 bl_39 br_39 wl_24 vdd gnd cell_6t
Xbit_r25_c39 bl_39 br_39 wl_25 vdd gnd cell_6t
Xbit_r26_c39 bl_39 br_39 wl_26 vdd gnd cell_6t
Xbit_r27_c39 bl_39 br_39 wl_27 vdd gnd cell_6t
Xbit_r28_c39 bl_39 br_39 wl_28 vdd gnd cell_6t
Xbit_r29_c39 bl_39 br_39 wl_29 vdd gnd cell_6t
Xbit_r30_c39 bl_39 br_39 wl_30 vdd gnd cell_6t
Xbit_r31_c39 bl_39 br_39 wl_31 vdd gnd cell_6t
Xbit_r32_c39 bl_39 br_39 wl_32 vdd gnd cell_6t
Xbit_r33_c39 bl_39 br_39 wl_33 vdd gnd cell_6t
Xbit_r34_c39 bl_39 br_39 wl_34 vdd gnd cell_6t
Xbit_r35_c39 bl_39 br_39 wl_35 vdd gnd cell_6t
Xbit_r36_c39 bl_39 br_39 wl_36 vdd gnd cell_6t
Xbit_r37_c39 bl_39 br_39 wl_37 vdd gnd cell_6t
Xbit_r38_c39 bl_39 br_39 wl_38 vdd gnd cell_6t
Xbit_r39_c39 bl_39 br_39 wl_39 vdd gnd cell_6t
Xbit_r40_c39 bl_39 br_39 wl_40 vdd gnd cell_6t
Xbit_r41_c39 bl_39 br_39 wl_41 vdd gnd cell_6t
Xbit_r42_c39 bl_39 br_39 wl_42 vdd gnd cell_6t
Xbit_r43_c39 bl_39 br_39 wl_43 vdd gnd cell_6t
Xbit_r44_c39 bl_39 br_39 wl_44 vdd gnd cell_6t
Xbit_r45_c39 bl_39 br_39 wl_45 vdd gnd cell_6t
Xbit_r46_c39 bl_39 br_39 wl_46 vdd gnd cell_6t
Xbit_r47_c39 bl_39 br_39 wl_47 vdd gnd cell_6t
Xbit_r48_c39 bl_39 br_39 wl_48 vdd gnd cell_6t
Xbit_r49_c39 bl_39 br_39 wl_49 vdd gnd cell_6t
Xbit_r50_c39 bl_39 br_39 wl_50 vdd gnd cell_6t
Xbit_r51_c39 bl_39 br_39 wl_51 vdd gnd cell_6t
Xbit_r52_c39 bl_39 br_39 wl_52 vdd gnd cell_6t
Xbit_r53_c39 bl_39 br_39 wl_53 vdd gnd cell_6t
Xbit_r54_c39 bl_39 br_39 wl_54 vdd gnd cell_6t
Xbit_r55_c39 bl_39 br_39 wl_55 vdd gnd cell_6t
Xbit_r56_c39 bl_39 br_39 wl_56 vdd gnd cell_6t
Xbit_r57_c39 bl_39 br_39 wl_57 vdd gnd cell_6t
Xbit_r58_c39 bl_39 br_39 wl_58 vdd gnd cell_6t
Xbit_r59_c39 bl_39 br_39 wl_59 vdd gnd cell_6t
Xbit_r60_c39 bl_39 br_39 wl_60 vdd gnd cell_6t
Xbit_r61_c39 bl_39 br_39 wl_61 vdd gnd cell_6t
Xbit_r62_c39 bl_39 br_39 wl_62 vdd gnd cell_6t
Xbit_r63_c39 bl_39 br_39 wl_63 vdd gnd cell_6t
Xbit_r64_c39 bl_39 br_39 wl_64 vdd gnd cell_6t
Xbit_r65_c39 bl_39 br_39 wl_65 vdd gnd cell_6t
Xbit_r66_c39 bl_39 br_39 wl_66 vdd gnd cell_6t
Xbit_r67_c39 bl_39 br_39 wl_67 vdd gnd cell_6t
Xbit_r68_c39 bl_39 br_39 wl_68 vdd gnd cell_6t
Xbit_r69_c39 bl_39 br_39 wl_69 vdd gnd cell_6t
Xbit_r70_c39 bl_39 br_39 wl_70 vdd gnd cell_6t
Xbit_r71_c39 bl_39 br_39 wl_71 vdd gnd cell_6t
Xbit_r72_c39 bl_39 br_39 wl_72 vdd gnd cell_6t
Xbit_r73_c39 bl_39 br_39 wl_73 vdd gnd cell_6t
Xbit_r74_c39 bl_39 br_39 wl_74 vdd gnd cell_6t
Xbit_r75_c39 bl_39 br_39 wl_75 vdd gnd cell_6t
Xbit_r76_c39 bl_39 br_39 wl_76 vdd gnd cell_6t
Xbit_r77_c39 bl_39 br_39 wl_77 vdd gnd cell_6t
Xbit_r78_c39 bl_39 br_39 wl_78 vdd gnd cell_6t
Xbit_r79_c39 bl_39 br_39 wl_79 vdd gnd cell_6t
Xbit_r80_c39 bl_39 br_39 wl_80 vdd gnd cell_6t
Xbit_r81_c39 bl_39 br_39 wl_81 vdd gnd cell_6t
Xbit_r82_c39 bl_39 br_39 wl_82 vdd gnd cell_6t
Xbit_r83_c39 bl_39 br_39 wl_83 vdd gnd cell_6t
Xbit_r84_c39 bl_39 br_39 wl_84 vdd gnd cell_6t
Xbit_r85_c39 bl_39 br_39 wl_85 vdd gnd cell_6t
Xbit_r86_c39 bl_39 br_39 wl_86 vdd gnd cell_6t
Xbit_r87_c39 bl_39 br_39 wl_87 vdd gnd cell_6t
Xbit_r88_c39 bl_39 br_39 wl_88 vdd gnd cell_6t
Xbit_r89_c39 bl_39 br_39 wl_89 vdd gnd cell_6t
Xbit_r90_c39 bl_39 br_39 wl_90 vdd gnd cell_6t
Xbit_r91_c39 bl_39 br_39 wl_91 vdd gnd cell_6t
Xbit_r92_c39 bl_39 br_39 wl_92 vdd gnd cell_6t
Xbit_r93_c39 bl_39 br_39 wl_93 vdd gnd cell_6t
Xbit_r94_c39 bl_39 br_39 wl_94 vdd gnd cell_6t
Xbit_r95_c39 bl_39 br_39 wl_95 vdd gnd cell_6t
Xbit_r96_c39 bl_39 br_39 wl_96 vdd gnd cell_6t
Xbit_r97_c39 bl_39 br_39 wl_97 vdd gnd cell_6t
Xbit_r98_c39 bl_39 br_39 wl_98 vdd gnd cell_6t
Xbit_r99_c39 bl_39 br_39 wl_99 vdd gnd cell_6t
Xbit_r100_c39 bl_39 br_39 wl_100 vdd gnd cell_6t
Xbit_r101_c39 bl_39 br_39 wl_101 vdd gnd cell_6t
Xbit_r102_c39 bl_39 br_39 wl_102 vdd gnd cell_6t
Xbit_r103_c39 bl_39 br_39 wl_103 vdd gnd cell_6t
Xbit_r104_c39 bl_39 br_39 wl_104 vdd gnd cell_6t
Xbit_r105_c39 bl_39 br_39 wl_105 vdd gnd cell_6t
Xbit_r106_c39 bl_39 br_39 wl_106 vdd gnd cell_6t
Xbit_r107_c39 bl_39 br_39 wl_107 vdd gnd cell_6t
Xbit_r108_c39 bl_39 br_39 wl_108 vdd gnd cell_6t
Xbit_r109_c39 bl_39 br_39 wl_109 vdd gnd cell_6t
Xbit_r110_c39 bl_39 br_39 wl_110 vdd gnd cell_6t
Xbit_r111_c39 bl_39 br_39 wl_111 vdd gnd cell_6t
Xbit_r112_c39 bl_39 br_39 wl_112 vdd gnd cell_6t
Xbit_r113_c39 bl_39 br_39 wl_113 vdd gnd cell_6t
Xbit_r114_c39 bl_39 br_39 wl_114 vdd gnd cell_6t
Xbit_r115_c39 bl_39 br_39 wl_115 vdd gnd cell_6t
Xbit_r116_c39 bl_39 br_39 wl_116 vdd gnd cell_6t
Xbit_r117_c39 bl_39 br_39 wl_117 vdd gnd cell_6t
Xbit_r118_c39 bl_39 br_39 wl_118 vdd gnd cell_6t
Xbit_r119_c39 bl_39 br_39 wl_119 vdd gnd cell_6t
Xbit_r120_c39 bl_39 br_39 wl_120 vdd gnd cell_6t
Xbit_r121_c39 bl_39 br_39 wl_121 vdd gnd cell_6t
Xbit_r122_c39 bl_39 br_39 wl_122 vdd gnd cell_6t
Xbit_r123_c39 bl_39 br_39 wl_123 vdd gnd cell_6t
Xbit_r124_c39 bl_39 br_39 wl_124 vdd gnd cell_6t
Xbit_r125_c39 bl_39 br_39 wl_125 vdd gnd cell_6t
Xbit_r126_c39 bl_39 br_39 wl_126 vdd gnd cell_6t
Xbit_r127_c39 bl_39 br_39 wl_127 vdd gnd cell_6t
Xbit_r128_c39 bl_39 br_39 wl_128 vdd gnd cell_6t
Xbit_r129_c39 bl_39 br_39 wl_129 vdd gnd cell_6t
Xbit_r130_c39 bl_39 br_39 wl_130 vdd gnd cell_6t
Xbit_r131_c39 bl_39 br_39 wl_131 vdd gnd cell_6t
Xbit_r132_c39 bl_39 br_39 wl_132 vdd gnd cell_6t
Xbit_r133_c39 bl_39 br_39 wl_133 vdd gnd cell_6t
Xbit_r134_c39 bl_39 br_39 wl_134 vdd gnd cell_6t
Xbit_r135_c39 bl_39 br_39 wl_135 vdd gnd cell_6t
Xbit_r136_c39 bl_39 br_39 wl_136 vdd gnd cell_6t
Xbit_r137_c39 bl_39 br_39 wl_137 vdd gnd cell_6t
Xbit_r138_c39 bl_39 br_39 wl_138 vdd gnd cell_6t
Xbit_r139_c39 bl_39 br_39 wl_139 vdd gnd cell_6t
Xbit_r140_c39 bl_39 br_39 wl_140 vdd gnd cell_6t
Xbit_r141_c39 bl_39 br_39 wl_141 vdd gnd cell_6t
Xbit_r142_c39 bl_39 br_39 wl_142 vdd gnd cell_6t
Xbit_r143_c39 bl_39 br_39 wl_143 vdd gnd cell_6t
Xbit_r144_c39 bl_39 br_39 wl_144 vdd gnd cell_6t
Xbit_r145_c39 bl_39 br_39 wl_145 vdd gnd cell_6t
Xbit_r146_c39 bl_39 br_39 wl_146 vdd gnd cell_6t
Xbit_r147_c39 bl_39 br_39 wl_147 vdd gnd cell_6t
Xbit_r148_c39 bl_39 br_39 wl_148 vdd gnd cell_6t
Xbit_r149_c39 bl_39 br_39 wl_149 vdd gnd cell_6t
Xbit_r150_c39 bl_39 br_39 wl_150 vdd gnd cell_6t
Xbit_r151_c39 bl_39 br_39 wl_151 vdd gnd cell_6t
Xbit_r152_c39 bl_39 br_39 wl_152 vdd gnd cell_6t
Xbit_r153_c39 bl_39 br_39 wl_153 vdd gnd cell_6t
Xbit_r154_c39 bl_39 br_39 wl_154 vdd gnd cell_6t
Xbit_r155_c39 bl_39 br_39 wl_155 vdd gnd cell_6t
Xbit_r156_c39 bl_39 br_39 wl_156 vdd gnd cell_6t
Xbit_r157_c39 bl_39 br_39 wl_157 vdd gnd cell_6t
Xbit_r158_c39 bl_39 br_39 wl_158 vdd gnd cell_6t
Xbit_r159_c39 bl_39 br_39 wl_159 vdd gnd cell_6t
Xbit_r160_c39 bl_39 br_39 wl_160 vdd gnd cell_6t
Xbit_r161_c39 bl_39 br_39 wl_161 vdd gnd cell_6t
Xbit_r162_c39 bl_39 br_39 wl_162 vdd gnd cell_6t
Xbit_r163_c39 bl_39 br_39 wl_163 vdd gnd cell_6t
Xbit_r164_c39 bl_39 br_39 wl_164 vdd gnd cell_6t
Xbit_r165_c39 bl_39 br_39 wl_165 vdd gnd cell_6t
Xbit_r166_c39 bl_39 br_39 wl_166 vdd gnd cell_6t
Xbit_r167_c39 bl_39 br_39 wl_167 vdd gnd cell_6t
Xbit_r168_c39 bl_39 br_39 wl_168 vdd gnd cell_6t
Xbit_r169_c39 bl_39 br_39 wl_169 vdd gnd cell_6t
Xbit_r170_c39 bl_39 br_39 wl_170 vdd gnd cell_6t
Xbit_r171_c39 bl_39 br_39 wl_171 vdd gnd cell_6t
Xbit_r172_c39 bl_39 br_39 wl_172 vdd gnd cell_6t
Xbit_r173_c39 bl_39 br_39 wl_173 vdd gnd cell_6t
Xbit_r174_c39 bl_39 br_39 wl_174 vdd gnd cell_6t
Xbit_r175_c39 bl_39 br_39 wl_175 vdd gnd cell_6t
Xbit_r176_c39 bl_39 br_39 wl_176 vdd gnd cell_6t
Xbit_r177_c39 bl_39 br_39 wl_177 vdd gnd cell_6t
Xbit_r178_c39 bl_39 br_39 wl_178 vdd gnd cell_6t
Xbit_r179_c39 bl_39 br_39 wl_179 vdd gnd cell_6t
Xbit_r180_c39 bl_39 br_39 wl_180 vdd gnd cell_6t
Xbit_r181_c39 bl_39 br_39 wl_181 vdd gnd cell_6t
Xbit_r182_c39 bl_39 br_39 wl_182 vdd gnd cell_6t
Xbit_r183_c39 bl_39 br_39 wl_183 vdd gnd cell_6t
Xbit_r184_c39 bl_39 br_39 wl_184 vdd gnd cell_6t
Xbit_r185_c39 bl_39 br_39 wl_185 vdd gnd cell_6t
Xbit_r186_c39 bl_39 br_39 wl_186 vdd gnd cell_6t
Xbit_r187_c39 bl_39 br_39 wl_187 vdd gnd cell_6t
Xbit_r188_c39 bl_39 br_39 wl_188 vdd gnd cell_6t
Xbit_r189_c39 bl_39 br_39 wl_189 vdd gnd cell_6t
Xbit_r190_c39 bl_39 br_39 wl_190 vdd gnd cell_6t
Xbit_r191_c39 bl_39 br_39 wl_191 vdd gnd cell_6t
Xbit_r192_c39 bl_39 br_39 wl_192 vdd gnd cell_6t
Xbit_r193_c39 bl_39 br_39 wl_193 vdd gnd cell_6t
Xbit_r194_c39 bl_39 br_39 wl_194 vdd gnd cell_6t
Xbit_r195_c39 bl_39 br_39 wl_195 vdd gnd cell_6t
Xbit_r196_c39 bl_39 br_39 wl_196 vdd gnd cell_6t
Xbit_r197_c39 bl_39 br_39 wl_197 vdd gnd cell_6t
Xbit_r198_c39 bl_39 br_39 wl_198 vdd gnd cell_6t
Xbit_r199_c39 bl_39 br_39 wl_199 vdd gnd cell_6t
Xbit_r200_c39 bl_39 br_39 wl_200 vdd gnd cell_6t
Xbit_r201_c39 bl_39 br_39 wl_201 vdd gnd cell_6t
Xbit_r202_c39 bl_39 br_39 wl_202 vdd gnd cell_6t
Xbit_r203_c39 bl_39 br_39 wl_203 vdd gnd cell_6t
Xbit_r204_c39 bl_39 br_39 wl_204 vdd gnd cell_6t
Xbit_r205_c39 bl_39 br_39 wl_205 vdd gnd cell_6t
Xbit_r206_c39 bl_39 br_39 wl_206 vdd gnd cell_6t
Xbit_r207_c39 bl_39 br_39 wl_207 vdd gnd cell_6t
Xbit_r208_c39 bl_39 br_39 wl_208 vdd gnd cell_6t
Xbit_r209_c39 bl_39 br_39 wl_209 vdd gnd cell_6t
Xbit_r210_c39 bl_39 br_39 wl_210 vdd gnd cell_6t
Xbit_r211_c39 bl_39 br_39 wl_211 vdd gnd cell_6t
Xbit_r212_c39 bl_39 br_39 wl_212 vdd gnd cell_6t
Xbit_r213_c39 bl_39 br_39 wl_213 vdd gnd cell_6t
Xbit_r214_c39 bl_39 br_39 wl_214 vdd gnd cell_6t
Xbit_r215_c39 bl_39 br_39 wl_215 vdd gnd cell_6t
Xbit_r216_c39 bl_39 br_39 wl_216 vdd gnd cell_6t
Xbit_r217_c39 bl_39 br_39 wl_217 vdd gnd cell_6t
Xbit_r218_c39 bl_39 br_39 wl_218 vdd gnd cell_6t
Xbit_r219_c39 bl_39 br_39 wl_219 vdd gnd cell_6t
Xbit_r220_c39 bl_39 br_39 wl_220 vdd gnd cell_6t
Xbit_r221_c39 bl_39 br_39 wl_221 vdd gnd cell_6t
Xbit_r222_c39 bl_39 br_39 wl_222 vdd gnd cell_6t
Xbit_r223_c39 bl_39 br_39 wl_223 vdd gnd cell_6t
Xbit_r224_c39 bl_39 br_39 wl_224 vdd gnd cell_6t
Xbit_r225_c39 bl_39 br_39 wl_225 vdd gnd cell_6t
Xbit_r226_c39 bl_39 br_39 wl_226 vdd gnd cell_6t
Xbit_r227_c39 bl_39 br_39 wl_227 vdd gnd cell_6t
Xbit_r228_c39 bl_39 br_39 wl_228 vdd gnd cell_6t
Xbit_r229_c39 bl_39 br_39 wl_229 vdd gnd cell_6t
Xbit_r230_c39 bl_39 br_39 wl_230 vdd gnd cell_6t
Xbit_r231_c39 bl_39 br_39 wl_231 vdd gnd cell_6t
Xbit_r232_c39 bl_39 br_39 wl_232 vdd gnd cell_6t
Xbit_r233_c39 bl_39 br_39 wl_233 vdd gnd cell_6t
Xbit_r234_c39 bl_39 br_39 wl_234 vdd gnd cell_6t
Xbit_r235_c39 bl_39 br_39 wl_235 vdd gnd cell_6t
Xbit_r236_c39 bl_39 br_39 wl_236 vdd gnd cell_6t
Xbit_r237_c39 bl_39 br_39 wl_237 vdd gnd cell_6t
Xbit_r238_c39 bl_39 br_39 wl_238 vdd gnd cell_6t
Xbit_r239_c39 bl_39 br_39 wl_239 vdd gnd cell_6t
Xbit_r240_c39 bl_39 br_39 wl_240 vdd gnd cell_6t
Xbit_r241_c39 bl_39 br_39 wl_241 vdd gnd cell_6t
Xbit_r242_c39 bl_39 br_39 wl_242 vdd gnd cell_6t
Xbit_r243_c39 bl_39 br_39 wl_243 vdd gnd cell_6t
Xbit_r244_c39 bl_39 br_39 wl_244 vdd gnd cell_6t
Xbit_r245_c39 bl_39 br_39 wl_245 vdd gnd cell_6t
Xbit_r246_c39 bl_39 br_39 wl_246 vdd gnd cell_6t
Xbit_r247_c39 bl_39 br_39 wl_247 vdd gnd cell_6t
Xbit_r248_c39 bl_39 br_39 wl_248 vdd gnd cell_6t
Xbit_r249_c39 bl_39 br_39 wl_249 vdd gnd cell_6t
Xbit_r250_c39 bl_39 br_39 wl_250 vdd gnd cell_6t
Xbit_r251_c39 bl_39 br_39 wl_251 vdd gnd cell_6t
Xbit_r252_c39 bl_39 br_39 wl_252 vdd gnd cell_6t
Xbit_r253_c39 bl_39 br_39 wl_253 vdd gnd cell_6t
Xbit_r254_c39 bl_39 br_39 wl_254 vdd gnd cell_6t
Xbit_r255_c39 bl_39 br_39 wl_255 vdd gnd cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd cell_6t
Xbit_r1_c40 bl_40 br_40 wl_1 vdd gnd cell_6t
Xbit_r2_c40 bl_40 br_40 wl_2 vdd gnd cell_6t
Xbit_r3_c40 bl_40 br_40 wl_3 vdd gnd cell_6t
Xbit_r4_c40 bl_40 br_40 wl_4 vdd gnd cell_6t
Xbit_r5_c40 bl_40 br_40 wl_5 vdd gnd cell_6t
Xbit_r6_c40 bl_40 br_40 wl_6 vdd gnd cell_6t
Xbit_r7_c40 bl_40 br_40 wl_7 vdd gnd cell_6t
Xbit_r8_c40 bl_40 br_40 wl_8 vdd gnd cell_6t
Xbit_r9_c40 bl_40 br_40 wl_9 vdd gnd cell_6t
Xbit_r10_c40 bl_40 br_40 wl_10 vdd gnd cell_6t
Xbit_r11_c40 bl_40 br_40 wl_11 vdd gnd cell_6t
Xbit_r12_c40 bl_40 br_40 wl_12 vdd gnd cell_6t
Xbit_r13_c40 bl_40 br_40 wl_13 vdd gnd cell_6t
Xbit_r14_c40 bl_40 br_40 wl_14 vdd gnd cell_6t
Xbit_r15_c40 bl_40 br_40 wl_15 vdd gnd cell_6t
Xbit_r16_c40 bl_40 br_40 wl_16 vdd gnd cell_6t
Xbit_r17_c40 bl_40 br_40 wl_17 vdd gnd cell_6t
Xbit_r18_c40 bl_40 br_40 wl_18 vdd gnd cell_6t
Xbit_r19_c40 bl_40 br_40 wl_19 vdd gnd cell_6t
Xbit_r20_c40 bl_40 br_40 wl_20 vdd gnd cell_6t
Xbit_r21_c40 bl_40 br_40 wl_21 vdd gnd cell_6t
Xbit_r22_c40 bl_40 br_40 wl_22 vdd gnd cell_6t
Xbit_r23_c40 bl_40 br_40 wl_23 vdd gnd cell_6t
Xbit_r24_c40 bl_40 br_40 wl_24 vdd gnd cell_6t
Xbit_r25_c40 bl_40 br_40 wl_25 vdd gnd cell_6t
Xbit_r26_c40 bl_40 br_40 wl_26 vdd gnd cell_6t
Xbit_r27_c40 bl_40 br_40 wl_27 vdd gnd cell_6t
Xbit_r28_c40 bl_40 br_40 wl_28 vdd gnd cell_6t
Xbit_r29_c40 bl_40 br_40 wl_29 vdd gnd cell_6t
Xbit_r30_c40 bl_40 br_40 wl_30 vdd gnd cell_6t
Xbit_r31_c40 bl_40 br_40 wl_31 vdd gnd cell_6t
Xbit_r32_c40 bl_40 br_40 wl_32 vdd gnd cell_6t
Xbit_r33_c40 bl_40 br_40 wl_33 vdd gnd cell_6t
Xbit_r34_c40 bl_40 br_40 wl_34 vdd gnd cell_6t
Xbit_r35_c40 bl_40 br_40 wl_35 vdd gnd cell_6t
Xbit_r36_c40 bl_40 br_40 wl_36 vdd gnd cell_6t
Xbit_r37_c40 bl_40 br_40 wl_37 vdd gnd cell_6t
Xbit_r38_c40 bl_40 br_40 wl_38 vdd gnd cell_6t
Xbit_r39_c40 bl_40 br_40 wl_39 vdd gnd cell_6t
Xbit_r40_c40 bl_40 br_40 wl_40 vdd gnd cell_6t
Xbit_r41_c40 bl_40 br_40 wl_41 vdd gnd cell_6t
Xbit_r42_c40 bl_40 br_40 wl_42 vdd gnd cell_6t
Xbit_r43_c40 bl_40 br_40 wl_43 vdd gnd cell_6t
Xbit_r44_c40 bl_40 br_40 wl_44 vdd gnd cell_6t
Xbit_r45_c40 bl_40 br_40 wl_45 vdd gnd cell_6t
Xbit_r46_c40 bl_40 br_40 wl_46 vdd gnd cell_6t
Xbit_r47_c40 bl_40 br_40 wl_47 vdd gnd cell_6t
Xbit_r48_c40 bl_40 br_40 wl_48 vdd gnd cell_6t
Xbit_r49_c40 bl_40 br_40 wl_49 vdd gnd cell_6t
Xbit_r50_c40 bl_40 br_40 wl_50 vdd gnd cell_6t
Xbit_r51_c40 bl_40 br_40 wl_51 vdd gnd cell_6t
Xbit_r52_c40 bl_40 br_40 wl_52 vdd gnd cell_6t
Xbit_r53_c40 bl_40 br_40 wl_53 vdd gnd cell_6t
Xbit_r54_c40 bl_40 br_40 wl_54 vdd gnd cell_6t
Xbit_r55_c40 bl_40 br_40 wl_55 vdd gnd cell_6t
Xbit_r56_c40 bl_40 br_40 wl_56 vdd gnd cell_6t
Xbit_r57_c40 bl_40 br_40 wl_57 vdd gnd cell_6t
Xbit_r58_c40 bl_40 br_40 wl_58 vdd gnd cell_6t
Xbit_r59_c40 bl_40 br_40 wl_59 vdd gnd cell_6t
Xbit_r60_c40 bl_40 br_40 wl_60 vdd gnd cell_6t
Xbit_r61_c40 bl_40 br_40 wl_61 vdd gnd cell_6t
Xbit_r62_c40 bl_40 br_40 wl_62 vdd gnd cell_6t
Xbit_r63_c40 bl_40 br_40 wl_63 vdd gnd cell_6t
Xbit_r64_c40 bl_40 br_40 wl_64 vdd gnd cell_6t
Xbit_r65_c40 bl_40 br_40 wl_65 vdd gnd cell_6t
Xbit_r66_c40 bl_40 br_40 wl_66 vdd gnd cell_6t
Xbit_r67_c40 bl_40 br_40 wl_67 vdd gnd cell_6t
Xbit_r68_c40 bl_40 br_40 wl_68 vdd gnd cell_6t
Xbit_r69_c40 bl_40 br_40 wl_69 vdd gnd cell_6t
Xbit_r70_c40 bl_40 br_40 wl_70 vdd gnd cell_6t
Xbit_r71_c40 bl_40 br_40 wl_71 vdd gnd cell_6t
Xbit_r72_c40 bl_40 br_40 wl_72 vdd gnd cell_6t
Xbit_r73_c40 bl_40 br_40 wl_73 vdd gnd cell_6t
Xbit_r74_c40 bl_40 br_40 wl_74 vdd gnd cell_6t
Xbit_r75_c40 bl_40 br_40 wl_75 vdd gnd cell_6t
Xbit_r76_c40 bl_40 br_40 wl_76 vdd gnd cell_6t
Xbit_r77_c40 bl_40 br_40 wl_77 vdd gnd cell_6t
Xbit_r78_c40 bl_40 br_40 wl_78 vdd gnd cell_6t
Xbit_r79_c40 bl_40 br_40 wl_79 vdd gnd cell_6t
Xbit_r80_c40 bl_40 br_40 wl_80 vdd gnd cell_6t
Xbit_r81_c40 bl_40 br_40 wl_81 vdd gnd cell_6t
Xbit_r82_c40 bl_40 br_40 wl_82 vdd gnd cell_6t
Xbit_r83_c40 bl_40 br_40 wl_83 vdd gnd cell_6t
Xbit_r84_c40 bl_40 br_40 wl_84 vdd gnd cell_6t
Xbit_r85_c40 bl_40 br_40 wl_85 vdd gnd cell_6t
Xbit_r86_c40 bl_40 br_40 wl_86 vdd gnd cell_6t
Xbit_r87_c40 bl_40 br_40 wl_87 vdd gnd cell_6t
Xbit_r88_c40 bl_40 br_40 wl_88 vdd gnd cell_6t
Xbit_r89_c40 bl_40 br_40 wl_89 vdd gnd cell_6t
Xbit_r90_c40 bl_40 br_40 wl_90 vdd gnd cell_6t
Xbit_r91_c40 bl_40 br_40 wl_91 vdd gnd cell_6t
Xbit_r92_c40 bl_40 br_40 wl_92 vdd gnd cell_6t
Xbit_r93_c40 bl_40 br_40 wl_93 vdd gnd cell_6t
Xbit_r94_c40 bl_40 br_40 wl_94 vdd gnd cell_6t
Xbit_r95_c40 bl_40 br_40 wl_95 vdd gnd cell_6t
Xbit_r96_c40 bl_40 br_40 wl_96 vdd gnd cell_6t
Xbit_r97_c40 bl_40 br_40 wl_97 vdd gnd cell_6t
Xbit_r98_c40 bl_40 br_40 wl_98 vdd gnd cell_6t
Xbit_r99_c40 bl_40 br_40 wl_99 vdd gnd cell_6t
Xbit_r100_c40 bl_40 br_40 wl_100 vdd gnd cell_6t
Xbit_r101_c40 bl_40 br_40 wl_101 vdd gnd cell_6t
Xbit_r102_c40 bl_40 br_40 wl_102 vdd gnd cell_6t
Xbit_r103_c40 bl_40 br_40 wl_103 vdd gnd cell_6t
Xbit_r104_c40 bl_40 br_40 wl_104 vdd gnd cell_6t
Xbit_r105_c40 bl_40 br_40 wl_105 vdd gnd cell_6t
Xbit_r106_c40 bl_40 br_40 wl_106 vdd gnd cell_6t
Xbit_r107_c40 bl_40 br_40 wl_107 vdd gnd cell_6t
Xbit_r108_c40 bl_40 br_40 wl_108 vdd gnd cell_6t
Xbit_r109_c40 bl_40 br_40 wl_109 vdd gnd cell_6t
Xbit_r110_c40 bl_40 br_40 wl_110 vdd gnd cell_6t
Xbit_r111_c40 bl_40 br_40 wl_111 vdd gnd cell_6t
Xbit_r112_c40 bl_40 br_40 wl_112 vdd gnd cell_6t
Xbit_r113_c40 bl_40 br_40 wl_113 vdd gnd cell_6t
Xbit_r114_c40 bl_40 br_40 wl_114 vdd gnd cell_6t
Xbit_r115_c40 bl_40 br_40 wl_115 vdd gnd cell_6t
Xbit_r116_c40 bl_40 br_40 wl_116 vdd gnd cell_6t
Xbit_r117_c40 bl_40 br_40 wl_117 vdd gnd cell_6t
Xbit_r118_c40 bl_40 br_40 wl_118 vdd gnd cell_6t
Xbit_r119_c40 bl_40 br_40 wl_119 vdd gnd cell_6t
Xbit_r120_c40 bl_40 br_40 wl_120 vdd gnd cell_6t
Xbit_r121_c40 bl_40 br_40 wl_121 vdd gnd cell_6t
Xbit_r122_c40 bl_40 br_40 wl_122 vdd gnd cell_6t
Xbit_r123_c40 bl_40 br_40 wl_123 vdd gnd cell_6t
Xbit_r124_c40 bl_40 br_40 wl_124 vdd gnd cell_6t
Xbit_r125_c40 bl_40 br_40 wl_125 vdd gnd cell_6t
Xbit_r126_c40 bl_40 br_40 wl_126 vdd gnd cell_6t
Xbit_r127_c40 bl_40 br_40 wl_127 vdd gnd cell_6t
Xbit_r128_c40 bl_40 br_40 wl_128 vdd gnd cell_6t
Xbit_r129_c40 bl_40 br_40 wl_129 vdd gnd cell_6t
Xbit_r130_c40 bl_40 br_40 wl_130 vdd gnd cell_6t
Xbit_r131_c40 bl_40 br_40 wl_131 vdd gnd cell_6t
Xbit_r132_c40 bl_40 br_40 wl_132 vdd gnd cell_6t
Xbit_r133_c40 bl_40 br_40 wl_133 vdd gnd cell_6t
Xbit_r134_c40 bl_40 br_40 wl_134 vdd gnd cell_6t
Xbit_r135_c40 bl_40 br_40 wl_135 vdd gnd cell_6t
Xbit_r136_c40 bl_40 br_40 wl_136 vdd gnd cell_6t
Xbit_r137_c40 bl_40 br_40 wl_137 vdd gnd cell_6t
Xbit_r138_c40 bl_40 br_40 wl_138 vdd gnd cell_6t
Xbit_r139_c40 bl_40 br_40 wl_139 vdd gnd cell_6t
Xbit_r140_c40 bl_40 br_40 wl_140 vdd gnd cell_6t
Xbit_r141_c40 bl_40 br_40 wl_141 vdd gnd cell_6t
Xbit_r142_c40 bl_40 br_40 wl_142 vdd gnd cell_6t
Xbit_r143_c40 bl_40 br_40 wl_143 vdd gnd cell_6t
Xbit_r144_c40 bl_40 br_40 wl_144 vdd gnd cell_6t
Xbit_r145_c40 bl_40 br_40 wl_145 vdd gnd cell_6t
Xbit_r146_c40 bl_40 br_40 wl_146 vdd gnd cell_6t
Xbit_r147_c40 bl_40 br_40 wl_147 vdd gnd cell_6t
Xbit_r148_c40 bl_40 br_40 wl_148 vdd gnd cell_6t
Xbit_r149_c40 bl_40 br_40 wl_149 vdd gnd cell_6t
Xbit_r150_c40 bl_40 br_40 wl_150 vdd gnd cell_6t
Xbit_r151_c40 bl_40 br_40 wl_151 vdd gnd cell_6t
Xbit_r152_c40 bl_40 br_40 wl_152 vdd gnd cell_6t
Xbit_r153_c40 bl_40 br_40 wl_153 vdd gnd cell_6t
Xbit_r154_c40 bl_40 br_40 wl_154 vdd gnd cell_6t
Xbit_r155_c40 bl_40 br_40 wl_155 vdd gnd cell_6t
Xbit_r156_c40 bl_40 br_40 wl_156 vdd gnd cell_6t
Xbit_r157_c40 bl_40 br_40 wl_157 vdd gnd cell_6t
Xbit_r158_c40 bl_40 br_40 wl_158 vdd gnd cell_6t
Xbit_r159_c40 bl_40 br_40 wl_159 vdd gnd cell_6t
Xbit_r160_c40 bl_40 br_40 wl_160 vdd gnd cell_6t
Xbit_r161_c40 bl_40 br_40 wl_161 vdd gnd cell_6t
Xbit_r162_c40 bl_40 br_40 wl_162 vdd gnd cell_6t
Xbit_r163_c40 bl_40 br_40 wl_163 vdd gnd cell_6t
Xbit_r164_c40 bl_40 br_40 wl_164 vdd gnd cell_6t
Xbit_r165_c40 bl_40 br_40 wl_165 vdd gnd cell_6t
Xbit_r166_c40 bl_40 br_40 wl_166 vdd gnd cell_6t
Xbit_r167_c40 bl_40 br_40 wl_167 vdd gnd cell_6t
Xbit_r168_c40 bl_40 br_40 wl_168 vdd gnd cell_6t
Xbit_r169_c40 bl_40 br_40 wl_169 vdd gnd cell_6t
Xbit_r170_c40 bl_40 br_40 wl_170 vdd gnd cell_6t
Xbit_r171_c40 bl_40 br_40 wl_171 vdd gnd cell_6t
Xbit_r172_c40 bl_40 br_40 wl_172 vdd gnd cell_6t
Xbit_r173_c40 bl_40 br_40 wl_173 vdd gnd cell_6t
Xbit_r174_c40 bl_40 br_40 wl_174 vdd gnd cell_6t
Xbit_r175_c40 bl_40 br_40 wl_175 vdd gnd cell_6t
Xbit_r176_c40 bl_40 br_40 wl_176 vdd gnd cell_6t
Xbit_r177_c40 bl_40 br_40 wl_177 vdd gnd cell_6t
Xbit_r178_c40 bl_40 br_40 wl_178 vdd gnd cell_6t
Xbit_r179_c40 bl_40 br_40 wl_179 vdd gnd cell_6t
Xbit_r180_c40 bl_40 br_40 wl_180 vdd gnd cell_6t
Xbit_r181_c40 bl_40 br_40 wl_181 vdd gnd cell_6t
Xbit_r182_c40 bl_40 br_40 wl_182 vdd gnd cell_6t
Xbit_r183_c40 bl_40 br_40 wl_183 vdd gnd cell_6t
Xbit_r184_c40 bl_40 br_40 wl_184 vdd gnd cell_6t
Xbit_r185_c40 bl_40 br_40 wl_185 vdd gnd cell_6t
Xbit_r186_c40 bl_40 br_40 wl_186 vdd gnd cell_6t
Xbit_r187_c40 bl_40 br_40 wl_187 vdd gnd cell_6t
Xbit_r188_c40 bl_40 br_40 wl_188 vdd gnd cell_6t
Xbit_r189_c40 bl_40 br_40 wl_189 vdd gnd cell_6t
Xbit_r190_c40 bl_40 br_40 wl_190 vdd gnd cell_6t
Xbit_r191_c40 bl_40 br_40 wl_191 vdd gnd cell_6t
Xbit_r192_c40 bl_40 br_40 wl_192 vdd gnd cell_6t
Xbit_r193_c40 bl_40 br_40 wl_193 vdd gnd cell_6t
Xbit_r194_c40 bl_40 br_40 wl_194 vdd gnd cell_6t
Xbit_r195_c40 bl_40 br_40 wl_195 vdd gnd cell_6t
Xbit_r196_c40 bl_40 br_40 wl_196 vdd gnd cell_6t
Xbit_r197_c40 bl_40 br_40 wl_197 vdd gnd cell_6t
Xbit_r198_c40 bl_40 br_40 wl_198 vdd gnd cell_6t
Xbit_r199_c40 bl_40 br_40 wl_199 vdd gnd cell_6t
Xbit_r200_c40 bl_40 br_40 wl_200 vdd gnd cell_6t
Xbit_r201_c40 bl_40 br_40 wl_201 vdd gnd cell_6t
Xbit_r202_c40 bl_40 br_40 wl_202 vdd gnd cell_6t
Xbit_r203_c40 bl_40 br_40 wl_203 vdd gnd cell_6t
Xbit_r204_c40 bl_40 br_40 wl_204 vdd gnd cell_6t
Xbit_r205_c40 bl_40 br_40 wl_205 vdd gnd cell_6t
Xbit_r206_c40 bl_40 br_40 wl_206 vdd gnd cell_6t
Xbit_r207_c40 bl_40 br_40 wl_207 vdd gnd cell_6t
Xbit_r208_c40 bl_40 br_40 wl_208 vdd gnd cell_6t
Xbit_r209_c40 bl_40 br_40 wl_209 vdd gnd cell_6t
Xbit_r210_c40 bl_40 br_40 wl_210 vdd gnd cell_6t
Xbit_r211_c40 bl_40 br_40 wl_211 vdd gnd cell_6t
Xbit_r212_c40 bl_40 br_40 wl_212 vdd gnd cell_6t
Xbit_r213_c40 bl_40 br_40 wl_213 vdd gnd cell_6t
Xbit_r214_c40 bl_40 br_40 wl_214 vdd gnd cell_6t
Xbit_r215_c40 bl_40 br_40 wl_215 vdd gnd cell_6t
Xbit_r216_c40 bl_40 br_40 wl_216 vdd gnd cell_6t
Xbit_r217_c40 bl_40 br_40 wl_217 vdd gnd cell_6t
Xbit_r218_c40 bl_40 br_40 wl_218 vdd gnd cell_6t
Xbit_r219_c40 bl_40 br_40 wl_219 vdd gnd cell_6t
Xbit_r220_c40 bl_40 br_40 wl_220 vdd gnd cell_6t
Xbit_r221_c40 bl_40 br_40 wl_221 vdd gnd cell_6t
Xbit_r222_c40 bl_40 br_40 wl_222 vdd gnd cell_6t
Xbit_r223_c40 bl_40 br_40 wl_223 vdd gnd cell_6t
Xbit_r224_c40 bl_40 br_40 wl_224 vdd gnd cell_6t
Xbit_r225_c40 bl_40 br_40 wl_225 vdd gnd cell_6t
Xbit_r226_c40 bl_40 br_40 wl_226 vdd gnd cell_6t
Xbit_r227_c40 bl_40 br_40 wl_227 vdd gnd cell_6t
Xbit_r228_c40 bl_40 br_40 wl_228 vdd gnd cell_6t
Xbit_r229_c40 bl_40 br_40 wl_229 vdd gnd cell_6t
Xbit_r230_c40 bl_40 br_40 wl_230 vdd gnd cell_6t
Xbit_r231_c40 bl_40 br_40 wl_231 vdd gnd cell_6t
Xbit_r232_c40 bl_40 br_40 wl_232 vdd gnd cell_6t
Xbit_r233_c40 bl_40 br_40 wl_233 vdd gnd cell_6t
Xbit_r234_c40 bl_40 br_40 wl_234 vdd gnd cell_6t
Xbit_r235_c40 bl_40 br_40 wl_235 vdd gnd cell_6t
Xbit_r236_c40 bl_40 br_40 wl_236 vdd gnd cell_6t
Xbit_r237_c40 bl_40 br_40 wl_237 vdd gnd cell_6t
Xbit_r238_c40 bl_40 br_40 wl_238 vdd gnd cell_6t
Xbit_r239_c40 bl_40 br_40 wl_239 vdd gnd cell_6t
Xbit_r240_c40 bl_40 br_40 wl_240 vdd gnd cell_6t
Xbit_r241_c40 bl_40 br_40 wl_241 vdd gnd cell_6t
Xbit_r242_c40 bl_40 br_40 wl_242 vdd gnd cell_6t
Xbit_r243_c40 bl_40 br_40 wl_243 vdd gnd cell_6t
Xbit_r244_c40 bl_40 br_40 wl_244 vdd gnd cell_6t
Xbit_r245_c40 bl_40 br_40 wl_245 vdd gnd cell_6t
Xbit_r246_c40 bl_40 br_40 wl_246 vdd gnd cell_6t
Xbit_r247_c40 bl_40 br_40 wl_247 vdd gnd cell_6t
Xbit_r248_c40 bl_40 br_40 wl_248 vdd gnd cell_6t
Xbit_r249_c40 bl_40 br_40 wl_249 vdd gnd cell_6t
Xbit_r250_c40 bl_40 br_40 wl_250 vdd gnd cell_6t
Xbit_r251_c40 bl_40 br_40 wl_251 vdd gnd cell_6t
Xbit_r252_c40 bl_40 br_40 wl_252 vdd gnd cell_6t
Xbit_r253_c40 bl_40 br_40 wl_253 vdd gnd cell_6t
Xbit_r254_c40 bl_40 br_40 wl_254 vdd gnd cell_6t
Xbit_r255_c40 bl_40 br_40 wl_255 vdd gnd cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd cell_6t
Xbit_r1_c41 bl_41 br_41 wl_1 vdd gnd cell_6t
Xbit_r2_c41 bl_41 br_41 wl_2 vdd gnd cell_6t
Xbit_r3_c41 bl_41 br_41 wl_3 vdd gnd cell_6t
Xbit_r4_c41 bl_41 br_41 wl_4 vdd gnd cell_6t
Xbit_r5_c41 bl_41 br_41 wl_5 vdd gnd cell_6t
Xbit_r6_c41 bl_41 br_41 wl_6 vdd gnd cell_6t
Xbit_r7_c41 bl_41 br_41 wl_7 vdd gnd cell_6t
Xbit_r8_c41 bl_41 br_41 wl_8 vdd gnd cell_6t
Xbit_r9_c41 bl_41 br_41 wl_9 vdd gnd cell_6t
Xbit_r10_c41 bl_41 br_41 wl_10 vdd gnd cell_6t
Xbit_r11_c41 bl_41 br_41 wl_11 vdd gnd cell_6t
Xbit_r12_c41 bl_41 br_41 wl_12 vdd gnd cell_6t
Xbit_r13_c41 bl_41 br_41 wl_13 vdd gnd cell_6t
Xbit_r14_c41 bl_41 br_41 wl_14 vdd gnd cell_6t
Xbit_r15_c41 bl_41 br_41 wl_15 vdd gnd cell_6t
Xbit_r16_c41 bl_41 br_41 wl_16 vdd gnd cell_6t
Xbit_r17_c41 bl_41 br_41 wl_17 vdd gnd cell_6t
Xbit_r18_c41 bl_41 br_41 wl_18 vdd gnd cell_6t
Xbit_r19_c41 bl_41 br_41 wl_19 vdd gnd cell_6t
Xbit_r20_c41 bl_41 br_41 wl_20 vdd gnd cell_6t
Xbit_r21_c41 bl_41 br_41 wl_21 vdd gnd cell_6t
Xbit_r22_c41 bl_41 br_41 wl_22 vdd gnd cell_6t
Xbit_r23_c41 bl_41 br_41 wl_23 vdd gnd cell_6t
Xbit_r24_c41 bl_41 br_41 wl_24 vdd gnd cell_6t
Xbit_r25_c41 bl_41 br_41 wl_25 vdd gnd cell_6t
Xbit_r26_c41 bl_41 br_41 wl_26 vdd gnd cell_6t
Xbit_r27_c41 bl_41 br_41 wl_27 vdd gnd cell_6t
Xbit_r28_c41 bl_41 br_41 wl_28 vdd gnd cell_6t
Xbit_r29_c41 bl_41 br_41 wl_29 vdd gnd cell_6t
Xbit_r30_c41 bl_41 br_41 wl_30 vdd gnd cell_6t
Xbit_r31_c41 bl_41 br_41 wl_31 vdd gnd cell_6t
Xbit_r32_c41 bl_41 br_41 wl_32 vdd gnd cell_6t
Xbit_r33_c41 bl_41 br_41 wl_33 vdd gnd cell_6t
Xbit_r34_c41 bl_41 br_41 wl_34 vdd gnd cell_6t
Xbit_r35_c41 bl_41 br_41 wl_35 vdd gnd cell_6t
Xbit_r36_c41 bl_41 br_41 wl_36 vdd gnd cell_6t
Xbit_r37_c41 bl_41 br_41 wl_37 vdd gnd cell_6t
Xbit_r38_c41 bl_41 br_41 wl_38 vdd gnd cell_6t
Xbit_r39_c41 bl_41 br_41 wl_39 vdd gnd cell_6t
Xbit_r40_c41 bl_41 br_41 wl_40 vdd gnd cell_6t
Xbit_r41_c41 bl_41 br_41 wl_41 vdd gnd cell_6t
Xbit_r42_c41 bl_41 br_41 wl_42 vdd gnd cell_6t
Xbit_r43_c41 bl_41 br_41 wl_43 vdd gnd cell_6t
Xbit_r44_c41 bl_41 br_41 wl_44 vdd gnd cell_6t
Xbit_r45_c41 bl_41 br_41 wl_45 vdd gnd cell_6t
Xbit_r46_c41 bl_41 br_41 wl_46 vdd gnd cell_6t
Xbit_r47_c41 bl_41 br_41 wl_47 vdd gnd cell_6t
Xbit_r48_c41 bl_41 br_41 wl_48 vdd gnd cell_6t
Xbit_r49_c41 bl_41 br_41 wl_49 vdd gnd cell_6t
Xbit_r50_c41 bl_41 br_41 wl_50 vdd gnd cell_6t
Xbit_r51_c41 bl_41 br_41 wl_51 vdd gnd cell_6t
Xbit_r52_c41 bl_41 br_41 wl_52 vdd gnd cell_6t
Xbit_r53_c41 bl_41 br_41 wl_53 vdd gnd cell_6t
Xbit_r54_c41 bl_41 br_41 wl_54 vdd gnd cell_6t
Xbit_r55_c41 bl_41 br_41 wl_55 vdd gnd cell_6t
Xbit_r56_c41 bl_41 br_41 wl_56 vdd gnd cell_6t
Xbit_r57_c41 bl_41 br_41 wl_57 vdd gnd cell_6t
Xbit_r58_c41 bl_41 br_41 wl_58 vdd gnd cell_6t
Xbit_r59_c41 bl_41 br_41 wl_59 vdd gnd cell_6t
Xbit_r60_c41 bl_41 br_41 wl_60 vdd gnd cell_6t
Xbit_r61_c41 bl_41 br_41 wl_61 vdd gnd cell_6t
Xbit_r62_c41 bl_41 br_41 wl_62 vdd gnd cell_6t
Xbit_r63_c41 bl_41 br_41 wl_63 vdd gnd cell_6t
Xbit_r64_c41 bl_41 br_41 wl_64 vdd gnd cell_6t
Xbit_r65_c41 bl_41 br_41 wl_65 vdd gnd cell_6t
Xbit_r66_c41 bl_41 br_41 wl_66 vdd gnd cell_6t
Xbit_r67_c41 bl_41 br_41 wl_67 vdd gnd cell_6t
Xbit_r68_c41 bl_41 br_41 wl_68 vdd gnd cell_6t
Xbit_r69_c41 bl_41 br_41 wl_69 vdd gnd cell_6t
Xbit_r70_c41 bl_41 br_41 wl_70 vdd gnd cell_6t
Xbit_r71_c41 bl_41 br_41 wl_71 vdd gnd cell_6t
Xbit_r72_c41 bl_41 br_41 wl_72 vdd gnd cell_6t
Xbit_r73_c41 bl_41 br_41 wl_73 vdd gnd cell_6t
Xbit_r74_c41 bl_41 br_41 wl_74 vdd gnd cell_6t
Xbit_r75_c41 bl_41 br_41 wl_75 vdd gnd cell_6t
Xbit_r76_c41 bl_41 br_41 wl_76 vdd gnd cell_6t
Xbit_r77_c41 bl_41 br_41 wl_77 vdd gnd cell_6t
Xbit_r78_c41 bl_41 br_41 wl_78 vdd gnd cell_6t
Xbit_r79_c41 bl_41 br_41 wl_79 vdd gnd cell_6t
Xbit_r80_c41 bl_41 br_41 wl_80 vdd gnd cell_6t
Xbit_r81_c41 bl_41 br_41 wl_81 vdd gnd cell_6t
Xbit_r82_c41 bl_41 br_41 wl_82 vdd gnd cell_6t
Xbit_r83_c41 bl_41 br_41 wl_83 vdd gnd cell_6t
Xbit_r84_c41 bl_41 br_41 wl_84 vdd gnd cell_6t
Xbit_r85_c41 bl_41 br_41 wl_85 vdd gnd cell_6t
Xbit_r86_c41 bl_41 br_41 wl_86 vdd gnd cell_6t
Xbit_r87_c41 bl_41 br_41 wl_87 vdd gnd cell_6t
Xbit_r88_c41 bl_41 br_41 wl_88 vdd gnd cell_6t
Xbit_r89_c41 bl_41 br_41 wl_89 vdd gnd cell_6t
Xbit_r90_c41 bl_41 br_41 wl_90 vdd gnd cell_6t
Xbit_r91_c41 bl_41 br_41 wl_91 vdd gnd cell_6t
Xbit_r92_c41 bl_41 br_41 wl_92 vdd gnd cell_6t
Xbit_r93_c41 bl_41 br_41 wl_93 vdd gnd cell_6t
Xbit_r94_c41 bl_41 br_41 wl_94 vdd gnd cell_6t
Xbit_r95_c41 bl_41 br_41 wl_95 vdd gnd cell_6t
Xbit_r96_c41 bl_41 br_41 wl_96 vdd gnd cell_6t
Xbit_r97_c41 bl_41 br_41 wl_97 vdd gnd cell_6t
Xbit_r98_c41 bl_41 br_41 wl_98 vdd gnd cell_6t
Xbit_r99_c41 bl_41 br_41 wl_99 vdd gnd cell_6t
Xbit_r100_c41 bl_41 br_41 wl_100 vdd gnd cell_6t
Xbit_r101_c41 bl_41 br_41 wl_101 vdd gnd cell_6t
Xbit_r102_c41 bl_41 br_41 wl_102 vdd gnd cell_6t
Xbit_r103_c41 bl_41 br_41 wl_103 vdd gnd cell_6t
Xbit_r104_c41 bl_41 br_41 wl_104 vdd gnd cell_6t
Xbit_r105_c41 bl_41 br_41 wl_105 vdd gnd cell_6t
Xbit_r106_c41 bl_41 br_41 wl_106 vdd gnd cell_6t
Xbit_r107_c41 bl_41 br_41 wl_107 vdd gnd cell_6t
Xbit_r108_c41 bl_41 br_41 wl_108 vdd gnd cell_6t
Xbit_r109_c41 bl_41 br_41 wl_109 vdd gnd cell_6t
Xbit_r110_c41 bl_41 br_41 wl_110 vdd gnd cell_6t
Xbit_r111_c41 bl_41 br_41 wl_111 vdd gnd cell_6t
Xbit_r112_c41 bl_41 br_41 wl_112 vdd gnd cell_6t
Xbit_r113_c41 bl_41 br_41 wl_113 vdd gnd cell_6t
Xbit_r114_c41 bl_41 br_41 wl_114 vdd gnd cell_6t
Xbit_r115_c41 bl_41 br_41 wl_115 vdd gnd cell_6t
Xbit_r116_c41 bl_41 br_41 wl_116 vdd gnd cell_6t
Xbit_r117_c41 bl_41 br_41 wl_117 vdd gnd cell_6t
Xbit_r118_c41 bl_41 br_41 wl_118 vdd gnd cell_6t
Xbit_r119_c41 bl_41 br_41 wl_119 vdd gnd cell_6t
Xbit_r120_c41 bl_41 br_41 wl_120 vdd gnd cell_6t
Xbit_r121_c41 bl_41 br_41 wl_121 vdd gnd cell_6t
Xbit_r122_c41 bl_41 br_41 wl_122 vdd gnd cell_6t
Xbit_r123_c41 bl_41 br_41 wl_123 vdd gnd cell_6t
Xbit_r124_c41 bl_41 br_41 wl_124 vdd gnd cell_6t
Xbit_r125_c41 bl_41 br_41 wl_125 vdd gnd cell_6t
Xbit_r126_c41 bl_41 br_41 wl_126 vdd gnd cell_6t
Xbit_r127_c41 bl_41 br_41 wl_127 vdd gnd cell_6t
Xbit_r128_c41 bl_41 br_41 wl_128 vdd gnd cell_6t
Xbit_r129_c41 bl_41 br_41 wl_129 vdd gnd cell_6t
Xbit_r130_c41 bl_41 br_41 wl_130 vdd gnd cell_6t
Xbit_r131_c41 bl_41 br_41 wl_131 vdd gnd cell_6t
Xbit_r132_c41 bl_41 br_41 wl_132 vdd gnd cell_6t
Xbit_r133_c41 bl_41 br_41 wl_133 vdd gnd cell_6t
Xbit_r134_c41 bl_41 br_41 wl_134 vdd gnd cell_6t
Xbit_r135_c41 bl_41 br_41 wl_135 vdd gnd cell_6t
Xbit_r136_c41 bl_41 br_41 wl_136 vdd gnd cell_6t
Xbit_r137_c41 bl_41 br_41 wl_137 vdd gnd cell_6t
Xbit_r138_c41 bl_41 br_41 wl_138 vdd gnd cell_6t
Xbit_r139_c41 bl_41 br_41 wl_139 vdd gnd cell_6t
Xbit_r140_c41 bl_41 br_41 wl_140 vdd gnd cell_6t
Xbit_r141_c41 bl_41 br_41 wl_141 vdd gnd cell_6t
Xbit_r142_c41 bl_41 br_41 wl_142 vdd gnd cell_6t
Xbit_r143_c41 bl_41 br_41 wl_143 vdd gnd cell_6t
Xbit_r144_c41 bl_41 br_41 wl_144 vdd gnd cell_6t
Xbit_r145_c41 bl_41 br_41 wl_145 vdd gnd cell_6t
Xbit_r146_c41 bl_41 br_41 wl_146 vdd gnd cell_6t
Xbit_r147_c41 bl_41 br_41 wl_147 vdd gnd cell_6t
Xbit_r148_c41 bl_41 br_41 wl_148 vdd gnd cell_6t
Xbit_r149_c41 bl_41 br_41 wl_149 vdd gnd cell_6t
Xbit_r150_c41 bl_41 br_41 wl_150 vdd gnd cell_6t
Xbit_r151_c41 bl_41 br_41 wl_151 vdd gnd cell_6t
Xbit_r152_c41 bl_41 br_41 wl_152 vdd gnd cell_6t
Xbit_r153_c41 bl_41 br_41 wl_153 vdd gnd cell_6t
Xbit_r154_c41 bl_41 br_41 wl_154 vdd gnd cell_6t
Xbit_r155_c41 bl_41 br_41 wl_155 vdd gnd cell_6t
Xbit_r156_c41 bl_41 br_41 wl_156 vdd gnd cell_6t
Xbit_r157_c41 bl_41 br_41 wl_157 vdd gnd cell_6t
Xbit_r158_c41 bl_41 br_41 wl_158 vdd gnd cell_6t
Xbit_r159_c41 bl_41 br_41 wl_159 vdd gnd cell_6t
Xbit_r160_c41 bl_41 br_41 wl_160 vdd gnd cell_6t
Xbit_r161_c41 bl_41 br_41 wl_161 vdd gnd cell_6t
Xbit_r162_c41 bl_41 br_41 wl_162 vdd gnd cell_6t
Xbit_r163_c41 bl_41 br_41 wl_163 vdd gnd cell_6t
Xbit_r164_c41 bl_41 br_41 wl_164 vdd gnd cell_6t
Xbit_r165_c41 bl_41 br_41 wl_165 vdd gnd cell_6t
Xbit_r166_c41 bl_41 br_41 wl_166 vdd gnd cell_6t
Xbit_r167_c41 bl_41 br_41 wl_167 vdd gnd cell_6t
Xbit_r168_c41 bl_41 br_41 wl_168 vdd gnd cell_6t
Xbit_r169_c41 bl_41 br_41 wl_169 vdd gnd cell_6t
Xbit_r170_c41 bl_41 br_41 wl_170 vdd gnd cell_6t
Xbit_r171_c41 bl_41 br_41 wl_171 vdd gnd cell_6t
Xbit_r172_c41 bl_41 br_41 wl_172 vdd gnd cell_6t
Xbit_r173_c41 bl_41 br_41 wl_173 vdd gnd cell_6t
Xbit_r174_c41 bl_41 br_41 wl_174 vdd gnd cell_6t
Xbit_r175_c41 bl_41 br_41 wl_175 vdd gnd cell_6t
Xbit_r176_c41 bl_41 br_41 wl_176 vdd gnd cell_6t
Xbit_r177_c41 bl_41 br_41 wl_177 vdd gnd cell_6t
Xbit_r178_c41 bl_41 br_41 wl_178 vdd gnd cell_6t
Xbit_r179_c41 bl_41 br_41 wl_179 vdd gnd cell_6t
Xbit_r180_c41 bl_41 br_41 wl_180 vdd gnd cell_6t
Xbit_r181_c41 bl_41 br_41 wl_181 vdd gnd cell_6t
Xbit_r182_c41 bl_41 br_41 wl_182 vdd gnd cell_6t
Xbit_r183_c41 bl_41 br_41 wl_183 vdd gnd cell_6t
Xbit_r184_c41 bl_41 br_41 wl_184 vdd gnd cell_6t
Xbit_r185_c41 bl_41 br_41 wl_185 vdd gnd cell_6t
Xbit_r186_c41 bl_41 br_41 wl_186 vdd gnd cell_6t
Xbit_r187_c41 bl_41 br_41 wl_187 vdd gnd cell_6t
Xbit_r188_c41 bl_41 br_41 wl_188 vdd gnd cell_6t
Xbit_r189_c41 bl_41 br_41 wl_189 vdd gnd cell_6t
Xbit_r190_c41 bl_41 br_41 wl_190 vdd gnd cell_6t
Xbit_r191_c41 bl_41 br_41 wl_191 vdd gnd cell_6t
Xbit_r192_c41 bl_41 br_41 wl_192 vdd gnd cell_6t
Xbit_r193_c41 bl_41 br_41 wl_193 vdd gnd cell_6t
Xbit_r194_c41 bl_41 br_41 wl_194 vdd gnd cell_6t
Xbit_r195_c41 bl_41 br_41 wl_195 vdd gnd cell_6t
Xbit_r196_c41 bl_41 br_41 wl_196 vdd gnd cell_6t
Xbit_r197_c41 bl_41 br_41 wl_197 vdd gnd cell_6t
Xbit_r198_c41 bl_41 br_41 wl_198 vdd gnd cell_6t
Xbit_r199_c41 bl_41 br_41 wl_199 vdd gnd cell_6t
Xbit_r200_c41 bl_41 br_41 wl_200 vdd gnd cell_6t
Xbit_r201_c41 bl_41 br_41 wl_201 vdd gnd cell_6t
Xbit_r202_c41 bl_41 br_41 wl_202 vdd gnd cell_6t
Xbit_r203_c41 bl_41 br_41 wl_203 vdd gnd cell_6t
Xbit_r204_c41 bl_41 br_41 wl_204 vdd gnd cell_6t
Xbit_r205_c41 bl_41 br_41 wl_205 vdd gnd cell_6t
Xbit_r206_c41 bl_41 br_41 wl_206 vdd gnd cell_6t
Xbit_r207_c41 bl_41 br_41 wl_207 vdd gnd cell_6t
Xbit_r208_c41 bl_41 br_41 wl_208 vdd gnd cell_6t
Xbit_r209_c41 bl_41 br_41 wl_209 vdd gnd cell_6t
Xbit_r210_c41 bl_41 br_41 wl_210 vdd gnd cell_6t
Xbit_r211_c41 bl_41 br_41 wl_211 vdd gnd cell_6t
Xbit_r212_c41 bl_41 br_41 wl_212 vdd gnd cell_6t
Xbit_r213_c41 bl_41 br_41 wl_213 vdd gnd cell_6t
Xbit_r214_c41 bl_41 br_41 wl_214 vdd gnd cell_6t
Xbit_r215_c41 bl_41 br_41 wl_215 vdd gnd cell_6t
Xbit_r216_c41 bl_41 br_41 wl_216 vdd gnd cell_6t
Xbit_r217_c41 bl_41 br_41 wl_217 vdd gnd cell_6t
Xbit_r218_c41 bl_41 br_41 wl_218 vdd gnd cell_6t
Xbit_r219_c41 bl_41 br_41 wl_219 vdd gnd cell_6t
Xbit_r220_c41 bl_41 br_41 wl_220 vdd gnd cell_6t
Xbit_r221_c41 bl_41 br_41 wl_221 vdd gnd cell_6t
Xbit_r222_c41 bl_41 br_41 wl_222 vdd gnd cell_6t
Xbit_r223_c41 bl_41 br_41 wl_223 vdd gnd cell_6t
Xbit_r224_c41 bl_41 br_41 wl_224 vdd gnd cell_6t
Xbit_r225_c41 bl_41 br_41 wl_225 vdd gnd cell_6t
Xbit_r226_c41 bl_41 br_41 wl_226 vdd gnd cell_6t
Xbit_r227_c41 bl_41 br_41 wl_227 vdd gnd cell_6t
Xbit_r228_c41 bl_41 br_41 wl_228 vdd gnd cell_6t
Xbit_r229_c41 bl_41 br_41 wl_229 vdd gnd cell_6t
Xbit_r230_c41 bl_41 br_41 wl_230 vdd gnd cell_6t
Xbit_r231_c41 bl_41 br_41 wl_231 vdd gnd cell_6t
Xbit_r232_c41 bl_41 br_41 wl_232 vdd gnd cell_6t
Xbit_r233_c41 bl_41 br_41 wl_233 vdd gnd cell_6t
Xbit_r234_c41 bl_41 br_41 wl_234 vdd gnd cell_6t
Xbit_r235_c41 bl_41 br_41 wl_235 vdd gnd cell_6t
Xbit_r236_c41 bl_41 br_41 wl_236 vdd gnd cell_6t
Xbit_r237_c41 bl_41 br_41 wl_237 vdd gnd cell_6t
Xbit_r238_c41 bl_41 br_41 wl_238 vdd gnd cell_6t
Xbit_r239_c41 bl_41 br_41 wl_239 vdd gnd cell_6t
Xbit_r240_c41 bl_41 br_41 wl_240 vdd gnd cell_6t
Xbit_r241_c41 bl_41 br_41 wl_241 vdd gnd cell_6t
Xbit_r242_c41 bl_41 br_41 wl_242 vdd gnd cell_6t
Xbit_r243_c41 bl_41 br_41 wl_243 vdd gnd cell_6t
Xbit_r244_c41 bl_41 br_41 wl_244 vdd gnd cell_6t
Xbit_r245_c41 bl_41 br_41 wl_245 vdd gnd cell_6t
Xbit_r246_c41 bl_41 br_41 wl_246 vdd gnd cell_6t
Xbit_r247_c41 bl_41 br_41 wl_247 vdd gnd cell_6t
Xbit_r248_c41 bl_41 br_41 wl_248 vdd gnd cell_6t
Xbit_r249_c41 bl_41 br_41 wl_249 vdd gnd cell_6t
Xbit_r250_c41 bl_41 br_41 wl_250 vdd gnd cell_6t
Xbit_r251_c41 bl_41 br_41 wl_251 vdd gnd cell_6t
Xbit_r252_c41 bl_41 br_41 wl_252 vdd gnd cell_6t
Xbit_r253_c41 bl_41 br_41 wl_253 vdd gnd cell_6t
Xbit_r254_c41 bl_41 br_41 wl_254 vdd gnd cell_6t
Xbit_r255_c41 bl_41 br_41 wl_255 vdd gnd cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd cell_6t
Xbit_r1_c42 bl_42 br_42 wl_1 vdd gnd cell_6t
Xbit_r2_c42 bl_42 br_42 wl_2 vdd gnd cell_6t
Xbit_r3_c42 bl_42 br_42 wl_3 vdd gnd cell_6t
Xbit_r4_c42 bl_42 br_42 wl_4 vdd gnd cell_6t
Xbit_r5_c42 bl_42 br_42 wl_5 vdd gnd cell_6t
Xbit_r6_c42 bl_42 br_42 wl_6 vdd gnd cell_6t
Xbit_r7_c42 bl_42 br_42 wl_7 vdd gnd cell_6t
Xbit_r8_c42 bl_42 br_42 wl_8 vdd gnd cell_6t
Xbit_r9_c42 bl_42 br_42 wl_9 vdd gnd cell_6t
Xbit_r10_c42 bl_42 br_42 wl_10 vdd gnd cell_6t
Xbit_r11_c42 bl_42 br_42 wl_11 vdd gnd cell_6t
Xbit_r12_c42 bl_42 br_42 wl_12 vdd gnd cell_6t
Xbit_r13_c42 bl_42 br_42 wl_13 vdd gnd cell_6t
Xbit_r14_c42 bl_42 br_42 wl_14 vdd gnd cell_6t
Xbit_r15_c42 bl_42 br_42 wl_15 vdd gnd cell_6t
Xbit_r16_c42 bl_42 br_42 wl_16 vdd gnd cell_6t
Xbit_r17_c42 bl_42 br_42 wl_17 vdd gnd cell_6t
Xbit_r18_c42 bl_42 br_42 wl_18 vdd gnd cell_6t
Xbit_r19_c42 bl_42 br_42 wl_19 vdd gnd cell_6t
Xbit_r20_c42 bl_42 br_42 wl_20 vdd gnd cell_6t
Xbit_r21_c42 bl_42 br_42 wl_21 vdd gnd cell_6t
Xbit_r22_c42 bl_42 br_42 wl_22 vdd gnd cell_6t
Xbit_r23_c42 bl_42 br_42 wl_23 vdd gnd cell_6t
Xbit_r24_c42 bl_42 br_42 wl_24 vdd gnd cell_6t
Xbit_r25_c42 bl_42 br_42 wl_25 vdd gnd cell_6t
Xbit_r26_c42 bl_42 br_42 wl_26 vdd gnd cell_6t
Xbit_r27_c42 bl_42 br_42 wl_27 vdd gnd cell_6t
Xbit_r28_c42 bl_42 br_42 wl_28 vdd gnd cell_6t
Xbit_r29_c42 bl_42 br_42 wl_29 vdd gnd cell_6t
Xbit_r30_c42 bl_42 br_42 wl_30 vdd gnd cell_6t
Xbit_r31_c42 bl_42 br_42 wl_31 vdd gnd cell_6t
Xbit_r32_c42 bl_42 br_42 wl_32 vdd gnd cell_6t
Xbit_r33_c42 bl_42 br_42 wl_33 vdd gnd cell_6t
Xbit_r34_c42 bl_42 br_42 wl_34 vdd gnd cell_6t
Xbit_r35_c42 bl_42 br_42 wl_35 vdd gnd cell_6t
Xbit_r36_c42 bl_42 br_42 wl_36 vdd gnd cell_6t
Xbit_r37_c42 bl_42 br_42 wl_37 vdd gnd cell_6t
Xbit_r38_c42 bl_42 br_42 wl_38 vdd gnd cell_6t
Xbit_r39_c42 bl_42 br_42 wl_39 vdd gnd cell_6t
Xbit_r40_c42 bl_42 br_42 wl_40 vdd gnd cell_6t
Xbit_r41_c42 bl_42 br_42 wl_41 vdd gnd cell_6t
Xbit_r42_c42 bl_42 br_42 wl_42 vdd gnd cell_6t
Xbit_r43_c42 bl_42 br_42 wl_43 vdd gnd cell_6t
Xbit_r44_c42 bl_42 br_42 wl_44 vdd gnd cell_6t
Xbit_r45_c42 bl_42 br_42 wl_45 vdd gnd cell_6t
Xbit_r46_c42 bl_42 br_42 wl_46 vdd gnd cell_6t
Xbit_r47_c42 bl_42 br_42 wl_47 vdd gnd cell_6t
Xbit_r48_c42 bl_42 br_42 wl_48 vdd gnd cell_6t
Xbit_r49_c42 bl_42 br_42 wl_49 vdd gnd cell_6t
Xbit_r50_c42 bl_42 br_42 wl_50 vdd gnd cell_6t
Xbit_r51_c42 bl_42 br_42 wl_51 vdd gnd cell_6t
Xbit_r52_c42 bl_42 br_42 wl_52 vdd gnd cell_6t
Xbit_r53_c42 bl_42 br_42 wl_53 vdd gnd cell_6t
Xbit_r54_c42 bl_42 br_42 wl_54 vdd gnd cell_6t
Xbit_r55_c42 bl_42 br_42 wl_55 vdd gnd cell_6t
Xbit_r56_c42 bl_42 br_42 wl_56 vdd gnd cell_6t
Xbit_r57_c42 bl_42 br_42 wl_57 vdd gnd cell_6t
Xbit_r58_c42 bl_42 br_42 wl_58 vdd gnd cell_6t
Xbit_r59_c42 bl_42 br_42 wl_59 vdd gnd cell_6t
Xbit_r60_c42 bl_42 br_42 wl_60 vdd gnd cell_6t
Xbit_r61_c42 bl_42 br_42 wl_61 vdd gnd cell_6t
Xbit_r62_c42 bl_42 br_42 wl_62 vdd gnd cell_6t
Xbit_r63_c42 bl_42 br_42 wl_63 vdd gnd cell_6t
Xbit_r64_c42 bl_42 br_42 wl_64 vdd gnd cell_6t
Xbit_r65_c42 bl_42 br_42 wl_65 vdd gnd cell_6t
Xbit_r66_c42 bl_42 br_42 wl_66 vdd gnd cell_6t
Xbit_r67_c42 bl_42 br_42 wl_67 vdd gnd cell_6t
Xbit_r68_c42 bl_42 br_42 wl_68 vdd gnd cell_6t
Xbit_r69_c42 bl_42 br_42 wl_69 vdd gnd cell_6t
Xbit_r70_c42 bl_42 br_42 wl_70 vdd gnd cell_6t
Xbit_r71_c42 bl_42 br_42 wl_71 vdd gnd cell_6t
Xbit_r72_c42 bl_42 br_42 wl_72 vdd gnd cell_6t
Xbit_r73_c42 bl_42 br_42 wl_73 vdd gnd cell_6t
Xbit_r74_c42 bl_42 br_42 wl_74 vdd gnd cell_6t
Xbit_r75_c42 bl_42 br_42 wl_75 vdd gnd cell_6t
Xbit_r76_c42 bl_42 br_42 wl_76 vdd gnd cell_6t
Xbit_r77_c42 bl_42 br_42 wl_77 vdd gnd cell_6t
Xbit_r78_c42 bl_42 br_42 wl_78 vdd gnd cell_6t
Xbit_r79_c42 bl_42 br_42 wl_79 vdd gnd cell_6t
Xbit_r80_c42 bl_42 br_42 wl_80 vdd gnd cell_6t
Xbit_r81_c42 bl_42 br_42 wl_81 vdd gnd cell_6t
Xbit_r82_c42 bl_42 br_42 wl_82 vdd gnd cell_6t
Xbit_r83_c42 bl_42 br_42 wl_83 vdd gnd cell_6t
Xbit_r84_c42 bl_42 br_42 wl_84 vdd gnd cell_6t
Xbit_r85_c42 bl_42 br_42 wl_85 vdd gnd cell_6t
Xbit_r86_c42 bl_42 br_42 wl_86 vdd gnd cell_6t
Xbit_r87_c42 bl_42 br_42 wl_87 vdd gnd cell_6t
Xbit_r88_c42 bl_42 br_42 wl_88 vdd gnd cell_6t
Xbit_r89_c42 bl_42 br_42 wl_89 vdd gnd cell_6t
Xbit_r90_c42 bl_42 br_42 wl_90 vdd gnd cell_6t
Xbit_r91_c42 bl_42 br_42 wl_91 vdd gnd cell_6t
Xbit_r92_c42 bl_42 br_42 wl_92 vdd gnd cell_6t
Xbit_r93_c42 bl_42 br_42 wl_93 vdd gnd cell_6t
Xbit_r94_c42 bl_42 br_42 wl_94 vdd gnd cell_6t
Xbit_r95_c42 bl_42 br_42 wl_95 vdd gnd cell_6t
Xbit_r96_c42 bl_42 br_42 wl_96 vdd gnd cell_6t
Xbit_r97_c42 bl_42 br_42 wl_97 vdd gnd cell_6t
Xbit_r98_c42 bl_42 br_42 wl_98 vdd gnd cell_6t
Xbit_r99_c42 bl_42 br_42 wl_99 vdd gnd cell_6t
Xbit_r100_c42 bl_42 br_42 wl_100 vdd gnd cell_6t
Xbit_r101_c42 bl_42 br_42 wl_101 vdd gnd cell_6t
Xbit_r102_c42 bl_42 br_42 wl_102 vdd gnd cell_6t
Xbit_r103_c42 bl_42 br_42 wl_103 vdd gnd cell_6t
Xbit_r104_c42 bl_42 br_42 wl_104 vdd gnd cell_6t
Xbit_r105_c42 bl_42 br_42 wl_105 vdd gnd cell_6t
Xbit_r106_c42 bl_42 br_42 wl_106 vdd gnd cell_6t
Xbit_r107_c42 bl_42 br_42 wl_107 vdd gnd cell_6t
Xbit_r108_c42 bl_42 br_42 wl_108 vdd gnd cell_6t
Xbit_r109_c42 bl_42 br_42 wl_109 vdd gnd cell_6t
Xbit_r110_c42 bl_42 br_42 wl_110 vdd gnd cell_6t
Xbit_r111_c42 bl_42 br_42 wl_111 vdd gnd cell_6t
Xbit_r112_c42 bl_42 br_42 wl_112 vdd gnd cell_6t
Xbit_r113_c42 bl_42 br_42 wl_113 vdd gnd cell_6t
Xbit_r114_c42 bl_42 br_42 wl_114 vdd gnd cell_6t
Xbit_r115_c42 bl_42 br_42 wl_115 vdd gnd cell_6t
Xbit_r116_c42 bl_42 br_42 wl_116 vdd gnd cell_6t
Xbit_r117_c42 bl_42 br_42 wl_117 vdd gnd cell_6t
Xbit_r118_c42 bl_42 br_42 wl_118 vdd gnd cell_6t
Xbit_r119_c42 bl_42 br_42 wl_119 vdd gnd cell_6t
Xbit_r120_c42 bl_42 br_42 wl_120 vdd gnd cell_6t
Xbit_r121_c42 bl_42 br_42 wl_121 vdd gnd cell_6t
Xbit_r122_c42 bl_42 br_42 wl_122 vdd gnd cell_6t
Xbit_r123_c42 bl_42 br_42 wl_123 vdd gnd cell_6t
Xbit_r124_c42 bl_42 br_42 wl_124 vdd gnd cell_6t
Xbit_r125_c42 bl_42 br_42 wl_125 vdd gnd cell_6t
Xbit_r126_c42 bl_42 br_42 wl_126 vdd gnd cell_6t
Xbit_r127_c42 bl_42 br_42 wl_127 vdd gnd cell_6t
Xbit_r128_c42 bl_42 br_42 wl_128 vdd gnd cell_6t
Xbit_r129_c42 bl_42 br_42 wl_129 vdd gnd cell_6t
Xbit_r130_c42 bl_42 br_42 wl_130 vdd gnd cell_6t
Xbit_r131_c42 bl_42 br_42 wl_131 vdd gnd cell_6t
Xbit_r132_c42 bl_42 br_42 wl_132 vdd gnd cell_6t
Xbit_r133_c42 bl_42 br_42 wl_133 vdd gnd cell_6t
Xbit_r134_c42 bl_42 br_42 wl_134 vdd gnd cell_6t
Xbit_r135_c42 bl_42 br_42 wl_135 vdd gnd cell_6t
Xbit_r136_c42 bl_42 br_42 wl_136 vdd gnd cell_6t
Xbit_r137_c42 bl_42 br_42 wl_137 vdd gnd cell_6t
Xbit_r138_c42 bl_42 br_42 wl_138 vdd gnd cell_6t
Xbit_r139_c42 bl_42 br_42 wl_139 vdd gnd cell_6t
Xbit_r140_c42 bl_42 br_42 wl_140 vdd gnd cell_6t
Xbit_r141_c42 bl_42 br_42 wl_141 vdd gnd cell_6t
Xbit_r142_c42 bl_42 br_42 wl_142 vdd gnd cell_6t
Xbit_r143_c42 bl_42 br_42 wl_143 vdd gnd cell_6t
Xbit_r144_c42 bl_42 br_42 wl_144 vdd gnd cell_6t
Xbit_r145_c42 bl_42 br_42 wl_145 vdd gnd cell_6t
Xbit_r146_c42 bl_42 br_42 wl_146 vdd gnd cell_6t
Xbit_r147_c42 bl_42 br_42 wl_147 vdd gnd cell_6t
Xbit_r148_c42 bl_42 br_42 wl_148 vdd gnd cell_6t
Xbit_r149_c42 bl_42 br_42 wl_149 vdd gnd cell_6t
Xbit_r150_c42 bl_42 br_42 wl_150 vdd gnd cell_6t
Xbit_r151_c42 bl_42 br_42 wl_151 vdd gnd cell_6t
Xbit_r152_c42 bl_42 br_42 wl_152 vdd gnd cell_6t
Xbit_r153_c42 bl_42 br_42 wl_153 vdd gnd cell_6t
Xbit_r154_c42 bl_42 br_42 wl_154 vdd gnd cell_6t
Xbit_r155_c42 bl_42 br_42 wl_155 vdd gnd cell_6t
Xbit_r156_c42 bl_42 br_42 wl_156 vdd gnd cell_6t
Xbit_r157_c42 bl_42 br_42 wl_157 vdd gnd cell_6t
Xbit_r158_c42 bl_42 br_42 wl_158 vdd gnd cell_6t
Xbit_r159_c42 bl_42 br_42 wl_159 vdd gnd cell_6t
Xbit_r160_c42 bl_42 br_42 wl_160 vdd gnd cell_6t
Xbit_r161_c42 bl_42 br_42 wl_161 vdd gnd cell_6t
Xbit_r162_c42 bl_42 br_42 wl_162 vdd gnd cell_6t
Xbit_r163_c42 bl_42 br_42 wl_163 vdd gnd cell_6t
Xbit_r164_c42 bl_42 br_42 wl_164 vdd gnd cell_6t
Xbit_r165_c42 bl_42 br_42 wl_165 vdd gnd cell_6t
Xbit_r166_c42 bl_42 br_42 wl_166 vdd gnd cell_6t
Xbit_r167_c42 bl_42 br_42 wl_167 vdd gnd cell_6t
Xbit_r168_c42 bl_42 br_42 wl_168 vdd gnd cell_6t
Xbit_r169_c42 bl_42 br_42 wl_169 vdd gnd cell_6t
Xbit_r170_c42 bl_42 br_42 wl_170 vdd gnd cell_6t
Xbit_r171_c42 bl_42 br_42 wl_171 vdd gnd cell_6t
Xbit_r172_c42 bl_42 br_42 wl_172 vdd gnd cell_6t
Xbit_r173_c42 bl_42 br_42 wl_173 vdd gnd cell_6t
Xbit_r174_c42 bl_42 br_42 wl_174 vdd gnd cell_6t
Xbit_r175_c42 bl_42 br_42 wl_175 vdd gnd cell_6t
Xbit_r176_c42 bl_42 br_42 wl_176 vdd gnd cell_6t
Xbit_r177_c42 bl_42 br_42 wl_177 vdd gnd cell_6t
Xbit_r178_c42 bl_42 br_42 wl_178 vdd gnd cell_6t
Xbit_r179_c42 bl_42 br_42 wl_179 vdd gnd cell_6t
Xbit_r180_c42 bl_42 br_42 wl_180 vdd gnd cell_6t
Xbit_r181_c42 bl_42 br_42 wl_181 vdd gnd cell_6t
Xbit_r182_c42 bl_42 br_42 wl_182 vdd gnd cell_6t
Xbit_r183_c42 bl_42 br_42 wl_183 vdd gnd cell_6t
Xbit_r184_c42 bl_42 br_42 wl_184 vdd gnd cell_6t
Xbit_r185_c42 bl_42 br_42 wl_185 vdd gnd cell_6t
Xbit_r186_c42 bl_42 br_42 wl_186 vdd gnd cell_6t
Xbit_r187_c42 bl_42 br_42 wl_187 vdd gnd cell_6t
Xbit_r188_c42 bl_42 br_42 wl_188 vdd gnd cell_6t
Xbit_r189_c42 bl_42 br_42 wl_189 vdd gnd cell_6t
Xbit_r190_c42 bl_42 br_42 wl_190 vdd gnd cell_6t
Xbit_r191_c42 bl_42 br_42 wl_191 vdd gnd cell_6t
Xbit_r192_c42 bl_42 br_42 wl_192 vdd gnd cell_6t
Xbit_r193_c42 bl_42 br_42 wl_193 vdd gnd cell_6t
Xbit_r194_c42 bl_42 br_42 wl_194 vdd gnd cell_6t
Xbit_r195_c42 bl_42 br_42 wl_195 vdd gnd cell_6t
Xbit_r196_c42 bl_42 br_42 wl_196 vdd gnd cell_6t
Xbit_r197_c42 bl_42 br_42 wl_197 vdd gnd cell_6t
Xbit_r198_c42 bl_42 br_42 wl_198 vdd gnd cell_6t
Xbit_r199_c42 bl_42 br_42 wl_199 vdd gnd cell_6t
Xbit_r200_c42 bl_42 br_42 wl_200 vdd gnd cell_6t
Xbit_r201_c42 bl_42 br_42 wl_201 vdd gnd cell_6t
Xbit_r202_c42 bl_42 br_42 wl_202 vdd gnd cell_6t
Xbit_r203_c42 bl_42 br_42 wl_203 vdd gnd cell_6t
Xbit_r204_c42 bl_42 br_42 wl_204 vdd gnd cell_6t
Xbit_r205_c42 bl_42 br_42 wl_205 vdd gnd cell_6t
Xbit_r206_c42 bl_42 br_42 wl_206 vdd gnd cell_6t
Xbit_r207_c42 bl_42 br_42 wl_207 vdd gnd cell_6t
Xbit_r208_c42 bl_42 br_42 wl_208 vdd gnd cell_6t
Xbit_r209_c42 bl_42 br_42 wl_209 vdd gnd cell_6t
Xbit_r210_c42 bl_42 br_42 wl_210 vdd gnd cell_6t
Xbit_r211_c42 bl_42 br_42 wl_211 vdd gnd cell_6t
Xbit_r212_c42 bl_42 br_42 wl_212 vdd gnd cell_6t
Xbit_r213_c42 bl_42 br_42 wl_213 vdd gnd cell_6t
Xbit_r214_c42 bl_42 br_42 wl_214 vdd gnd cell_6t
Xbit_r215_c42 bl_42 br_42 wl_215 vdd gnd cell_6t
Xbit_r216_c42 bl_42 br_42 wl_216 vdd gnd cell_6t
Xbit_r217_c42 bl_42 br_42 wl_217 vdd gnd cell_6t
Xbit_r218_c42 bl_42 br_42 wl_218 vdd gnd cell_6t
Xbit_r219_c42 bl_42 br_42 wl_219 vdd gnd cell_6t
Xbit_r220_c42 bl_42 br_42 wl_220 vdd gnd cell_6t
Xbit_r221_c42 bl_42 br_42 wl_221 vdd gnd cell_6t
Xbit_r222_c42 bl_42 br_42 wl_222 vdd gnd cell_6t
Xbit_r223_c42 bl_42 br_42 wl_223 vdd gnd cell_6t
Xbit_r224_c42 bl_42 br_42 wl_224 vdd gnd cell_6t
Xbit_r225_c42 bl_42 br_42 wl_225 vdd gnd cell_6t
Xbit_r226_c42 bl_42 br_42 wl_226 vdd gnd cell_6t
Xbit_r227_c42 bl_42 br_42 wl_227 vdd gnd cell_6t
Xbit_r228_c42 bl_42 br_42 wl_228 vdd gnd cell_6t
Xbit_r229_c42 bl_42 br_42 wl_229 vdd gnd cell_6t
Xbit_r230_c42 bl_42 br_42 wl_230 vdd gnd cell_6t
Xbit_r231_c42 bl_42 br_42 wl_231 vdd gnd cell_6t
Xbit_r232_c42 bl_42 br_42 wl_232 vdd gnd cell_6t
Xbit_r233_c42 bl_42 br_42 wl_233 vdd gnd cell_6t
Xbit_r234_c42 bl_42 br_42 wl_234 vdd gnd cell_6t
Xbit_r235_c42 bl_42 br_42 wl_235 vdd gnd cell_6t
Xbit_r236_c42 bl_42 br_42 wl_236 vdd gnd cell_6t
Xbit_r237_c42 bl_42 br_42 wl_237 vdd gnd cell_6t
Xbit_r238_c42 bl_42 br_42 wl_238 vdd gnd cell_6t
Xbit_r239_c42 bl_42 br_42 wl_239 vdd gnd cell_6t
Xbit_r240_c42 bl_42 br_42 wl_240 vdd gnd cell_6t
Xbit_r241_c42 bl_42 br_42 wl_241 vdd gnd cell_6t
Xbit_r242_c42 bl_42 br_42 wl_242 vdd gnd cell_6t
Xbit_r243_c42 bl_42 br_42 wl_243 vdd gnd cell_6t
Xbit_r244_c42 bl_42 br_42 wl_244 vdd gnd cell_6t
Xbit_r245_c42 bl_42 br_42 wl_245 vdd gnd cell_6t
Xbit_r246_c42 bl_42 br_42 wl_246 vdd gnd cell_6t
Xbit_r247_c42 bl_42 br_42 wl_247 vdd gnd cell_6t
Xbit_r248_c42 bl_42 br_42 wl_248 vdd gnd cell_6t
Xbit_r249_c42 bl_42 br_42 wl_249 vdd gnd cell_6t
Xbit_r250_c42 bl_42 br_42 wl_250 vdd gnd cell_6t
Xbit_r251_c42 bl_42 br_42 wl_251 vdd gnd cell_6t
Xbit_r252_c42 bl_42 br_42 wl_252 vdd gnd cell_6t
Xbit_r253_c42 bl_42 br_42 wl_253 vdd gnd cell_6t
Xbit_r254_c42 bl_42 br_42 wl_254 vdd gnd cell_6t
Xbit_r255_c42 bl_42 br_42 wl_255 vdd gnd cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd cell_6t
Xbit_r1_c43 bl_43 br_43 wl_1 vdd gnd cell_6t
Xbit_r2_c43 bl_43 br_43 wl_2 vdd gnd cell_6t
Xbit_r3_c43 bl_43 br_43 wl_3 vdd gnd cell_6t
Xbit_r4_c43 bl_43 br_43 wl_4 vdd gnd cell_6t
Xbit_r5_c43 bl_43 br_43 wl_5 vdd gnd cell_6t
Xbit_r6_c43 bl_43 br_43 wl_6 vdd gnd cell_6t
Xbit_r7_c43 bl_43 br_43 wl_7 vdd gnd cell_6t
Xbit_r8_c43 bl_43 br_43 wl_8 vdd gnd cell_6t
Xbit_r9_c43 bl_43 br_43 wl_9 vdd gnd cell_6t
Xbit_r10_c43 bl_43 br_43 wl_10 vdd gnd cell_6t
Xbit_r11_c43 bl_43 br_43 wl_11 vdd gnd cell_6t
Xbit_r12_c43 bl_43 br_43 wl_12 vdd gnd cell_6t
Xbit_r13_c43 bl_43 br_43 wl_13 vdd gnd cell_6t
Xbit_r14_c43 bl_43 br_43 wl_14 vdd gnd cell_6t
Xbit_r15_c43 bl_43 br_43 wl_15 vdd gnd cell_6t
Xbit_r16_c43 bl_43 br_43 wl_16 vdd gnd cell_6t
Xbit_r17_c43 bl_43 br_43 wl_17 vdd gnd cell_6t
Xbit_r18_c43 bl_43 br_43 wl_18 vdd gnd cell_6t
Xbit_r19_c43 bl_43 br_43 wl_19 vdd gnd cell_6t
Xbit_r20_c43 bl_43 br_43 wl_20 vdd gnd cell_6t
Xbit_r21_c43 bl_43 br_43 wl_21 vdd gnd cell_6t
Xbit_r22_c43 bl_43 br_43 wl_22 vdd gnd cell_6t
Xbit_r23_c43 bl_43 br_43 wl_23 vdd gnd cell_6t
Xbit_r24_c43 bl_43 br_43 wl_24 vdd gnd cell_6t
Xbit_r25_c43 bl_43 br_43 wl_25 vdd gnd cell_6t
Xbit_r26_c43 bl_43 br_43 wl_26 vdd gnd cell_6t
Xbit_r27_c43 bl_43 br_43 wl_27 vdd gnd cell_6t
Xbit_r28_c43 bl_43 br_43 wl_28 vdd gnd cell_6t
Xbit_r29_c43 bl_43 br_43 wl_29 vdd gnd cell_6t
Xbit_r30_c43 bl_43 br_43 wl_30 vdd gnd cell_6t
Xbit_r31_c43 bl_43 br_43 wl_31 vdd gnd cell_6t
Xbit_r32_c43 bl_43 br_43 wl_32 vdd gnd cell_6t
Xbit_r33_c43 bl_43 br_43 wl_33 vdd gnd cell_6t
Xbit_r34_c43 bl_43 br_43 wl_34 vdd gnd cell_6t
Xbit_r35_c43 bl_43 br_43 wl_35 vdd gnd cell_6t
Xbit_r36_c43 bl_43 br_43 wl_36 vdd gnd cell_6t
Xbit_r37_c43 bl_43 br_43 wl_37 vdd gnd cell_6t
Xbit_r38_c43 bl_43 br_43 wl_38 vdd gnd cell_6t
Xbit_r39_c43 bl_43 br_43 wl_39 vdd gnd cell_6t
Xbit_r40_c43 bl_43 br_43 wl_40 vdd gnd cell_6t
Xbit_r41_c43 bl_43 br_43 wl_41 vdd gnd cell_6t
Xbit_r42_c43 bl_43 br_43 wl_42 vdd gnd cell_6t
Xbit_r43_c43 bl_43 br_43 wl_43 vdd gnd cell_6t
Xbit_r44_c43 bl_43 br_43 wl_44 vdd gnd cell_6t
Xbit_r45_c43 bl_43 br_43 wl_45 vdd gnd cell_6t
Xbit_r46_c43 bl_43 br_43 wl_46 vdd gnd cell_6t
Xbit_r47_c43 bl_43 br_43 wl_47 vdd gnd cell_6t
Xbit_r48_c43 bl_43 br_43 wl_48 vdd gnd cell_6t
Xbit_r49_c43 bl_43 br_43 wl_49 vdd gnd cell_6t
Xbit_r50_c43 bl_43 br_43 wl_50 vdd gnd cell_6t
Xbit_r51_c43 bl_43 br_43 wl_51 vdd gnd cell_6t
Xbit_r52_c43 bl_43 br_43 wl_52 vdd gnd cell_6t
Xbit_r53_c43 bl_43 br_43 wl_53 vdd gnd cell_6t
Xbit_r54_c43 bl_43 br_43 wl_54 vdd gnd cell_6t
Xbit_r55_c43 bl_43 br_43 wl_55 vdd gnd cell_6t
Xbit_r56_c43 bl_43 br_43 wl_56 vdd gnd cell_6t
Xbit_r57_c43 bl_43 br_43 wl_57 vdd gnd cell_6t
Xbit_r58_c43 bl_43 br_43 wl_58 vdd gnd cell_6t
Xbit_r59_c43 bl_43 br_43 wl_59 vdd gnd cell_6t
Xbit_r60_c43 bl_43 br_43 wl_60 vdd gnd cell_6t
Xbit_r61_c43 bl_43 br_43 wl_61 vdd gnd cell_6t
Xbit_r62_c43 bl_43 br_43 wl_62 vdd gnd cell_6t
Xbit_r63_c43 bl_43 br_43 wl_63 vdd gnd cell_6t
Xbit_r64_c43 bl_43 br_43 wl_64 vdd gnd cell_6t
Xbit_r65_c43 bl_43 br_43 wl_65 vdd gnd cell_6t
Xbit_r66_c43 bl_43 br_43 wl_66 vdd gnd cell_6t
Xbit_r67_c43 bl_43 br_43 wl_67 vdd gnd cell_6t
Xbit_r68_c43 bl_43 br_43 wl_68 vdd gnd cell_6t
Xbit_r69_c43 bl_43 br_43 wl_69 vdd gnd cell_6t
Xbit_r70_c43 bl_43 br_43 wl_70 vdd gnd cell_6t
Xbit_r71_c43 bl_43 br_43 wl_71 vdd gnd cell_6t
Xbit_r72_c43 bl_43 br_43 wl_72 vdd gnd cell_6t
Xbit_r73_c43 bl_43 br_43 wl_73 vdd gnd cell_6t
Xbit_r74_c43 bl_43 br_43 wl_74 vdd gnd cell_6t
Xbit_r75_c43 bl_43 br_43 wl_75 vdd gnd cell_6t
Xbit_r76_c43 bl_43 br_43 wl_76 vdd gnd cell_6t
Xbit_r77_c43 bl_43 br_43 wl_77 vdd gnd cell_6t
Xbit_r78_c43 bl_43 br_43 wl_78 vdd gnd cell_6t
Xbit_r79_c43 bl_43 br_43 wl_79 vdd gnd cell_6t
Xbit_r80_c43 bl_43 br_43 wl_80 vdd gnd cell_6t
Xbit_r81_c43 bl_43 br_43 wl_81 vdd gnd cell_6t
Xbit_r82_c43 bl_43 br_43 wl_82 vdd gnd cell_6t
Xbit_r83_c43 bl_43 br_43 wl_83 vdd gnd cell_6t
Xbit_r84_c43 bl_43 br_43 wl_84 vdd gnd cell_6t
Xbit_r85_c43 bl_43 br_43 wl_85 vdd gnd cell_6t
Xbit_r86_c43 bl_43 br_43 wl_86 vdd gnd cell_6t
Xbit_r87_c43 bl_43 br_43 wl_87 vdd gnd cell_6t
Xbit_r88_c43 bl_43 br_43 wl_88 vdd gnd cell_6t
Xbit_r89_c43 bl_43 br_43 wl_89 vdd gnd cell_6t
Xbit_r90_c43 bl_43 br_43 wl_90 vdd gnd cell_6t
Xbit_r91_c43 bl_43 br_43 wl_91 vdd gnd cell_6t
Xbit_r92_c43 bl_43 br_43 wl_92 vdd gnd cell_6t
Xbit_r93_c43 bl_43 br_43 wl_93 vdd gnd cell_6t
Xbit_r94_c43 bl_43 br_43 wl_94 vdd gnd cell_6t
Xbit_r95_c43 bl_43 br_43 wl_95 vdd gnd cell_6t
Xbit_r96_c43 bl_43 br_43 wl_96 vdd gnd cell_6t
Xbit_r97_c43 bl_43 br_43 wl_97 vdd gnd cell_6t
Xbit_r98_c43 bl_43 br_43 wl_98 vdd gnd cell_6t
Xbit_r99_c43 bl_43 br_43 wl_99 vdd gnd cell_6t
Xbit_r100_c43 bl_43 br_43 wl_100 vdd gnd cell_6t
Xbit_r101_c43 bl_43 br_43 wl_101 vdd gnd cell_6t
Xbit_r102_c43 bl_43 br_43 wl_102 vdd gnd cell_6t
Xbit_r103_c43 bl_43 br_43 wl_103 vdd gnd cell_6t
Xbit_r104_c43 bl_43 br_43 wl_104 vdd gnd cell_6t
Xbit_r105_c43 bl_43 br_43 wl_105 vdd gnd cell_6t
Xbit_r106_c43 bl_43 br_43 wl_106 vdd gnd cell_6t
Xbit_r107_c43 bl_43 br_43 wl_107 vdd gnd cell_6t
Xbit_r108_c43 bl_43 br_43 wl_108 vdd gnd cell_6t
Xbit_r109_c43 bl_43 br_43 wl_109 vdd gnd cell_6t
Xbit_r110_c43 bl_43 br_43 wl_110 vdd gnd cell_6t
Xbit_r111_c43 bl_43 br_43 wl_111 vdd gnd cell_6t
Xbit_r112_c43 bl_43 br_43 wl_112 vdd gnd cell_6t
Xbit_r113_c43 bl_43 br_43 wl_113 vdd gnd cell_6t
Xbit_r114_c43 bl_43 br_43 wl_114 vdd gnd cell_6t
Xbit_r115_c43 bl_43 br_43 wl_115 vdd gnd cell_6t
Xbit_r116_c43 bl_43 br_43 wl_116 vdd gnd cell_6t
Xbit_r117_c43 bl_43 br_43 wl_117 vdd gnd cell_6t
Xbit_r118_c43 bl_43 br_43 wl_118 vdd gnd cell_6t
Xbit_r119_c43 bl_43 br_43 wl_119 vdd gnd cell_6t
Xbit_r120_c43 bl_43 br_43 wl_120 vdd gnd cell_6t
Xbit_r121_c43 bl_43 br_43 wl_121 vdd gnd cell_6t
Xbit_r122_c43 bl_43 br_43 wl_122 vdd gnd cell_6t
Xbit_r123_c43 bl_43 br_43 wl_123 vdd gnd cell_6t
Xbit_r124_c43 bl_43 br_43 wl_124 vdd gnd cell_6t
Xbit_r125_c43 bl_43 br_43 wl_125 vdd gnd cell_6t
Xbit_r126_c43 bl_43 br_43 wl_126 vdd gnd cell_6t
Xbit_r127_c43 bl_43 br_43 wl_127 vdd gnd cell_6t
Xbit_r128_c43 bl_43 br_43 wl_128 vdd gnd cell_6t
Xbit_r129_c43 bl_43 br_43 wl_129 vdd gnd cell_6t
Xbit_r130_c43 bl_43 br_43 wl_130 vdd gnd cell_6t
Xbit_r131_c43 bl_43 br_43 wl_131 vdd gnd cell_6t
Xbit_r132_c43 bl_43 br_43 wl_132 vdd gnd cell_6t
Xbit_r133_c43 bl_43 br_43 wl_133 vdd gnd cell_6t
Xbit_r134_c43 bl_43 br_43 wl_134 vdd gnd cell_6t
Xbit_r135_c43 bl_43 br_43 wl_135 vdd gnd cell_6t
Xbit_r136_c43 bl_43 br_43 wl_136 vdd gnd cell_6t
Xbit_r137_c43 bl_43 br_43 wl_137 vdd gnd cell_6t
Xbit_r138_c43 bl_43 br_43 wl_138 vdd gnd cell_6t
Xbit_r139_c43 bl_43 br_43 wl_139 vdd gnd cell_6t
Xbit_r140_c43 bl_43 br_43 wl_140 vdd gnd cell_6t
Xbit_r141_c43 bl_43 br_43 wl_141 vdd gnd cell_6t
Xbit_r142_c43 bl_43 br_43 wl_142 vdd gnd cell_6t
Xbit_r143_c43 bl_43 br_43 wl_143 vdd gnd cell_6t
Xbit_r144_c43 bl_43 br_43 wl_144 vdd gnd cell_6t
Xbit_r145_c43 bl_43 br_43 wl_145 vdd gnd cell_6t
Xbit_r146_c43 bl_43 br_43 wl_146 vdd gnd cell_6t
Xbit_r147_c43 bl_43 br_43 wl_147 vdd gnd cell_6t
Xbit_r148_c43 bl_43 br_43 wl_148 vdd gnd cell_6t
Xbit_r149_c43 bl_43 br_43 wl_149 vdd gnd cell_6t
Xbit_r150_c43 bl_43 br_43 wl_150 vdd gnd cell_6t
Xbit_r151_c43 bl_43 br_43 wl_151 vdd gnd cell_6t
Xbit_r152_c43 bl_43 br_43 wl_152 vdd gnd cell_6t
Xbit_r153_c43 bl_43 br_43 wl_153 vdd gnd cell_6t
Xbit_r154_c43 bl_43 br_43 wl_154 vdd gnd cell_6t
Xbit_r155_c43 bl_43 br_43 wl_155 vdd gnd cell_6t
Xbit_r156_c43 bl_43 br_43 wl_156 vdd gnd cell_6t
Xbit_r157_c43 bl_43 br_43 wl_157 vdd gnd cell_6t
Xbit_r158_c43 bl_43 br_43 wl_158 vdd gnd cell_6t
Xbit_r159_c43 bl_43 br_43 wl_159 vdd gnd cell_6t
Xbit_r160_c43 bl_43 br_43 wl_160 vdd gnd cell_6t
Xbit_r161_c43 bl_43 br_43 wl_161 vdd gnd cell_6t
Xbit_r162_c43 bl_43 br_43 wl_162 vdd gnd cell_6t
Xbit_r163_c43 bl_43 br_43 wl_163 vdd gnd cell_6t
Xbit_r164_c43 bl_43 br_43 wl_164 vdd gnd cell_6t
Xbit_r165_c43 bl_43 br_43 wl_165 vdd gnd cell_6t
Xbit_r166_c43 bl_43 br_43 wl_166 vdd gnd cell_6t
Xbit_r167_c43 bl_43 br_43 wl_167 vdd gnd cell_6t
Xbit_r168_c43 bl_43 br_43 wl_168 vdd gnd cell_6t
Xbit_r169_c43 bl_43 br_43 wl_169 vdd gnd cell_6t
Xbit_r170_c43 bl_43 br_43 wl_170 vdd gnd cell_6t
Xbit_r171_c43 bl_43 br_43 wl_171 vdd gnd cell_6t
Xbit_r172_c43 bl_43 br_43 wl_172 vdd gnd cell_6t
Xbit_r173_c43 bl_43 br_43 wl_173 vdd gnd cell_6t
Xbit_r174_c43 bl_43 br_43 wl_174 vdd gnd cell_6t
Xbit_r175_c43 bl_43 br_43 wl_175 vdd gnd cell_6t
Xbit_r176_c43 bl_43 br_43 wl_176 vdd gnd cell_6t
Xbit_r177_c43 bl_43 br_43 wl_177 vdd gnd cell_6t
Xbit_r178_c43 bl_43 br_43 wl_178 vdd gnd cell_6t
Xbit_r179_c43 bl_43 br_43 wl_179 vdd gnd cell_6t
Xbit_r180_c43 bl_43 br_43 wl_180 vdd gnd cell_6t
Xbit_r181_c43 bl_43 br_43 wl_181 vdd gnd cell_6t
Xbit_r182_c43 bl_43 br_43 wl_182 vdd gnd cell_6t
Xbit_r183_c43 bl_43 br_43 wl_183 vdd gnd cell_6t
Xbit_r184_c43 bl_43 br_43 wl_184 vdd gnd cell_6t
Xbit_r185_c43 bl_43 br_43 wl_185 vdd gnd cell_6t
Xbit_r186_c43 bl_43 br_43 wl_186 vdd gnd cell_6t
Xbit_r187_c43 bl_43 br_43 wl_187 vdd gnd cell_6t
Xbit_r188_c43 bl_43 br_43 wl_188 vdd gnd cell_6t
Xbit_r189_c43 bl_43 br_43 wl_189 vdd gnd cell_6t
Xbit_r190_c43 bl_43 br_43 wl_190 vdd gnd cell_6t
Xbit_r191_c43 bl_43 br_43 wl_191 vdd gnd cell_6t
Xbit_r192_c43 bl_43 br_43 wl_192 vdd gnd cell_6t
Xbit_r193_c43 bl_43 br_43 wl_193 vdd gnd cell_6t
Xbit_r194_c43 bl_43 br_43 wl_194 vdd gnd cell_6t
Xbit_r195_c43 bl_43 br_43 wl_195 vdd gnd cell_6t
Xbit_r196_c43 bl_43 br_43 wl_196 vdd gnd cell_6t
Xbit_r197_c43 bl_43 br_43 wl_197 vdd gnd cell_6t
Xbit_r198_c43 bl_43 br_43 wl_198 vdd gnd cell_6t
Xbit_r199_c43 bl_43 br_43 wl_199 vdd gnd cell_6t
Xbit_r200_c43 bl_43 br_43 wl_200 vdd gnd cell_6t
Xbit_r201_c43 bl_43 br_43 wl_201 vdd gnd cell_6t
Xbit_r202_c43 bl_43 br_43 wl_202 vdd gnd cell_6t
Xbit_r203_c43 bl_43 br_43 wl_203 vdd gnd cell_6t
Xbit_r204_c43 bl_43 br_43 wl_204 vdd gnd cell_6t
Xbit_r205_c43 bl_43 br_43 wl_205 vdd gnd cell_6t
Xbit_r206_c43 bl_43 br_43 wl_206 vdd gnd cell_6t
Xbit_r207_c43 bl_43 br_43 wl_207 vdd gnd cell_6t
Xbit_r208_c43 bl_43 br_43 wl_208 vdd gnd cell_6t
Xbit_r209_c43 bl_43 br_43 wl_209 vdd gnd cell_6t
Xbit_r210_c43 bl_43 br_43 wl_210 vdd gnd cell_6t
Xbit_r211_c43 bl_43 br_43 wl_211 vdd gnd cell_6t
Xbit_r212_c43 bl_43 br_43 wl_212 vdd gnd cell_6t
Xbit_r213_c43 bl_43 br_43 wl_213 vdd gnd cell_6t
Xbit_r214_c43 bl_43 br_43 wl_214 vdd gnd cell_6t
Xbit_r215_c43 bl_43 br_43 wl_215 vdd gnd cell_6t
Xbit_r216_c43 bl_43 br_43 wl_216 vdd gnd cell_6t
Xbit_r217_c43 bl_43 br_43 wl_217 vdd gnd cell_6t
Xbit_r218_c43 bl_43 br_43 wl_218 vdd gnd cell_6t
Xbit_r219_c43 bl_43 br_43 wl_219 vdd gnd cell_6t
Xbit_r220_c43 bl_43 br_43 wl_220 vdd gnd cell_6t
Xbit_r221_c43 bl_43 br_43 wl_221 vdd gnd cell_6t
Xbit_r222_c43 bl_43 br_43 wl_222 vdd gnd cell_6t
Xbit_r223_c43 bl_43 br_43 wl_223 vdd gnd cell_6t
Xbit_r224_c43 bl_43 br_43 wl_224 vdd gnd cell_6t
Xbit_r225_c43 bl_43 br_43 wl_225 vdd gnd cell_6t
Xbit_r226_c43 bl_43 br_43 wl_226 vdd gnd cell_6t
Xbit_r227_c43 bl_43 br_43 wl_227 vdd gnd cell_6t
Xbit_r228_c43 bl_43 br_43 wl_228 vdd gnd cell_6t
Xbit_r229_c43 bl_43 br_43 wl_229 vdd gnd cell_6t
Xbit_r230_c43 bl_43 br_43 wl_230 vdd gnd cell_6t
Xbit_r231_c43 bl_43 br_43 wl_231 vdd gnd cell_6t
Xbit_r232_c43 bl_43 br_43 wl_232 vdd gnd cell_6t
Xbit_r233_c43 bl_43 br_43 wl_233 vdd gnd cell_6t
Xbit_r234_c43 bl_43 br_43 wl_234 vdd gnd cell_6t
Xbit_r235_c43 bl_43 br_43 wl_235 vdd gnd cell_6t
Xbit_r236_c43 bl_43 br_43 wl_236 vdd gnd cell_6t
Xbit_r237_c43 bl_43 br_43 wl_237 vdd gnd cell_6t
Xbit_r238_c43 bl_43 br_43 wl_238 vdd gnd cell_6t
Xbit_r239_c43 bl_43 br_43 wl_239 vdd gnd cell_6t
Xbit_r240_c43 bl_43 br_43 wl_240 vdd gnd cell_6t
Xbit_r241_c43 bl_43 br_43 wl_241 vdd gnd cell_6t
Xbit_r242_c43 bl_43 br_43 wl_242 vdd gnd cell_6t
Xbit_r243_c43 bl_43 br_43 wl_243 vdd gnd cell_6t
Xbit_r244_c43 bl_43 br_43 wl_244 vdd gnd cell_6t
Xbit_r245_c43 bl_43 br_43 wl_245 vdd gnd cell_6t
Xbit_r246_c43 bl_43 br_43 wl_246 vdd gnd cell_6t
Xbit_r247_c43 bl_43 br_43 wl_247 vdd gnd cell_6t
Xbit_r248_c43 bl_43 br_43 wl_248 vdd gnd cell_6t
Xbit_r249_c43 bl_43 br_43 wl_249 vdd gnd cell_6t
Xbit_r250_c43 bl_43 br_43 wl_250 vdd gnd cell_6t
Xbit_r251_c43 bl_43 br_43 wl_251 vdd gnd cell_6t
Xbit_r252_c43 bl_43 br_43 wl_252 vdd gnd cell_6t
Xbit_r253_c43 bl_43 br_43 wl_253 vdd gnd cell_6t
Xbit_r254_c43 bl_43 br_43 wl_254 vdd gnd cell_6t
Xbit_r255_c43 bl_43 br_43 wl_255 vdd gnd cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd cell_6t
Xbit_r1_c44 bl_44 br_44 wl_1 vdd gnd cell_6t
Xbit_r2_c44 bl_44 br_44 wl_2 vdd gnd cell_6t
Xbit_r3_c44 bl_44 br_44 wl_3 vdd gnd cell_6t
Xbit_r4_c44 bl_44 br_44 wl_4 vdd gnd cell_6t
Xbit_r5_c44 bl_44 br_44 wl_5 vdd gnd cell_6t
Xbit_r6_c44 bl_44 br_44 wl_6 vdd gnd cell_6t
Xbit_r7_c44 bl_44 br_44 wl_7 vdd gnd cell_6t
Xbit_r8_c44 bl_44 br_44 wl_8 vdd gnd cell_6t
Xbit_r9_c44 bl_44 br_44 wl_9 vdd gnd cell_6t
Xbit_r10_c44 bl_44 br_44 wl_10 vdd gnd cell_6t
Xbit_r11_c44 bl_44 br_44 wl_11 vdd gnd cell_6t
Xbit_r12_c44 bl_44 br_44 wl_12 vdd gnd cell_6t
Xbit_r13_c44 bl_44 br_44 wl_13 vdd gnd cell_6t
Xbit_r14_c44 bl_44 br_44 wl_14 vdd gnd cell_6t
Xbit_r15_c44 bl_44 br_44 wl_15 vdd gnd cell_6t
Xbit_r16_c44 bl_44 br_44 wl_16 vdd gnd cell_6t
Xbit_r17_c44 bl_44 br_44 wl_17 vdd gnd cell_6t
Xbit_r18_c44 bl_44 br_44 wl_18 vdd gnd cell_6t
Xbit_r19_c44 bl_44 br_44 wl_19 vdd gnd cell_6t
Xbit_r20_c44 bl_44 br_44 wl_20 vdd gnd cell_6t
Xbit_r21_c44 bl_44 br_44 wl_21 vdd gnd cell_6t
Xbit_r22_c44 bl_44 br_44 wl_22 vdd gnd cell_6t
Xbit_r23_c44 bl_44 br_44 wl_23 vdd gnd cell_6t
Xbit_r24_c44 bl_44 br_44 wl_24 vdd gnd cell_6t
Xbit_r25_c44 bl_44 br_44 wl_25 vdd gnd cell_6t
Xbit_r26_c44 bl_44 br_44 wl_26 vdd gnd cell_6t
Xbit_r27_c44 bl_44 br_44 wl_27 vdd gnd cell_6t
Xbit_r28_c44 bl_44 br_44 wl_28 vdd gnd cell_6t
Xbit_r29_c44 bl_44 br_44 wl_29 vdd gnd cell_6t
Xbit_r30_c44 bl_44 br_44 wl_30 vdd gnd cell_6t
Xbit_r31_c44 bl_44 br_44 wl_31 vdd gnd cell_6t
Xbit_r32_c44 bl_44 br_44 wl_32 vdd gnd cell_6t
Xbit_r33_c44 bl_44 br_44 wl_33 vdd gnd cell_6t
Xbit_r34_c44 bl_44 br_44 wl_34 vdd gnd cell_6t
Xbit_r35_c44 bl_44 br_44 wl_35 vdd gnd cell_6t
Xbit_r36_c44 bl_44 br_44 wl_36 vdd gnd cell_6t
Xbit_r37_c44 bl_44 br_44 wl_37 vdd gnd cell_6t
Xbit_r38_c44 bl_44 br_44 wl_38 vdd gnd cell_6t
Xbit_r39_c44 bl_44 br_44 wl_39 vdd gnd cell_6t
Xbit_r40_c44 bl_44 br_44 wl_40 vdd gnd cell_6t
Xbit_r41_c44 bl_44 br_44 wl_41 vdd gnd cell_6t
Xbit_r42_c44 bl_44 br_44 wl_42 vdd gnd cell_6t
Xbit_r43_c44 bl_44 br_44 wl_43 vdd gnd cell_6t
Xbit_r44_c44 bl_44 br_44 wl_44 vdd gnd cell_6t
Xbit_r45_c44 bl_44 br_44 wl_45 vdd gnd cell_6t
Xbit_r46_c44 bl_44 br_44 wl_46 vdd gnd cell_6t
Xbit_r47_c44 bl_44 br_44 wl_47 vdd gnd cell_6t
Xbit_r48_c44 bl_44 br_44 wl_48 vdd gnd cell_6t
Xbit_r49_c44 bl_44 br_44 wl_49 vdd gnd cell_6t
Xbit_r50_c44 bl_44 br_44 wl_50 vdd gnd cell_6t
Xbit_r51_c44 bl_44 br_44 wl_51 vdd gnd cell_6t
Xbit_r52_c44 bl_44 br_44 wl_52 vdd gnd cell_6t
Xbit_r53_c44 bl_44 br_44 wl_53 vdd gnd cell_6t
Xbit_r54_c44 bl_44 br_44 wl_54 vdd gnd cell_6t
Xbit_r55_c44 bl_44 br_44 wl_55 vdd gnd cell_6t
Xbit_r56_c44 bl_44 br_44 wl_56 vdd gnd cell_6t
Xbit_r57_c44 bl_44 br_44 wl_57 vdd gnd cell_6t
Xbit_r58_c44 bl_44 br_44 wl_58 vdd gnd cell_6t
Xbit_r59_c44 bl_44 br_44 wl_59 vdd gnd cell_6t
Xbit_r60_c44 bl_44 br_44 wl_60 vdd gnd cell_6t
Xbit_r61_c44 bl_44 br_44 wl_61 vdd gnd cell_6t
Xbit_r62_c44 bl_44 br_44 wl_62 vdd gnd cell_6t
Xbit_r63_c44 bl_44 br_44 wl_63 vdd gnd cell_6t
Xbit_r64_c44 bl_44 br_44 wl_64 vdd gnd cell_6t
Xbit_r65_c44 bl_44 br_44 wl_65 vdd gnd cell_6t
Xbit_r66_c44 bl_44 br_44 wl_66 vdd gnd cell_6t
Xbit_r67_c44 bl_44 br_44 wl_67 vdd gnd cell_6t
Xbit_r68_c44 bl_44 br_44 wl_68 vdd gnd cell_6t
Xbit_r69_c44 bl_44 br_44 wl_69 vdd gnd cell_6t
Xbit_r70_c44 bl_44 br_44 wl_70 vdd gnd cell_6t
Xbit_r71_c44 bl_44 br_44 wl_71 vdd gnd cell_6t
Xbit_r72_c44 bl_44 br_44 wl_72 vdd gnd cell_6t
Xbit_r73_c44 bl_44 br_44 wl_73 vdd gnd cell_6t
Xbit_r74_c44 bl_44 br_44 wl_74 vdd gnd cell_6t
Xbit_r75_c44 bl_44 br_44 wl_75 vdd gnd cell_6t
Xbit_r76_c44 bl_44 br_44 wl_76 vdd gnd cell_6t
Xbit_r77_c44 bl_44 br_44 wl_77 vdd gnd cell_6t
Xbit_r78_c44 bl_44 br_44 wl_78 vdd gnd cell_6t
Xbit_r79_c44 bl_44 br_44 wl_79 vdd gnd cell_6t
Xbit_r80_c44 bl_44 br_44 wl_80 vdd gnd cell_6t
Xbit_r81_c44 bl_44 br_44 wl_81 vdd gnd cell_6t
Xbit_r82_c44 bl_44 br_44 wl_82 vdd gnd cell_6t
Xbit_r83_c44 bl_44 br_44 wl_83 vdd gnd cell_6t
Xbit_r84_c44 bl_44 br_44 wl_84 vdd gnd cell_6t
Xbit_r85_c44 bl_44 br_44 wl_85 vdd gnd cell_6t
Xbit_r86_c44 bl_44 br_44 wl_86 vdd gnd cell_6t
Xbit_r87_c44 bl_44 br_44 wl_87 vdd gnd cell_6t
Xbit_r88_c44 bl_44 br_44 wl_88 vdd gnd cell_6t
Xbit_r89_c44 bl_44 br_44 wl_89 vdd gnd cell_6t
Xbit_r90_c44 bl_44 br_44 wl_90 vdd gnd cell_6t
Xbit_r91_c44 bl_44 br_44 wl_91 vdd gnd cell_6t
Xbit_r92_c44 bl_44 br_44 wl_92 vdd gnd cell_6t
Xbit_r93_c44 bl_44 br_44 wl_93 vdd gnd cell_6t
Xbit_r94_c44 bl_44 br_44 wl_94 vdd gnd cell_6t
Xbit_r95_c44 bl_44 br_44 wl_95 vdd gnd cell_6t
Xbit_r96_c44 bl_44 br_44 wl_96 vdd gnd cell_6t
Xbit_r97_c44 bl_44 br_44 wl_97 vdd gnd cell_6t
Xbit_r98_c44 bl_44 br_44 wl_98 vdd gnd cell_6t
Xbit_r99_c44 bl_44 br_44 wl_99 vdd gnd cell_6t
Xbit_r100_c44 bl_44 br_44 wl_100 vdd gnd cell_6t
Xbit_r101_c44 bl_44 br_44 wl_101 vdd gnd cell_6t
Xbit_r102_c44 bl_44 br_44 wl_102 vdd gnd cell_6t
Xbit_r103_c44 bl_44 br_44 wl_103 vdd gnd cell_6t
Xbit_r104_c44 bl_44 br_44 wl_104 vdd gnd cell_6t
Xbit_r105_c44 bl_44 br_44 wl_105 vdd gnd cell_6t
Xbit_r106_c44 bl_44 br_44 wl_106 vdd gnd cell_6t
Xbit_r107_c44 bl_44 br_44 wl_107 vdd gnd cell_6t
Xbit_r108_c44 bl_44 br_44 wl_108 vdd gnd cell_6t
Xbit_r109_c44 bl_44 br_44 wl_109 vdd gnd cell_6t
Xbit_r110_c44 bl_44 br_44 wl_110 vdd gnd cell_6t
Xbit_r111_c44 bl_44 br_44 wl_111 vdd gnd cell_6t
Xbit_r112_c44 bl_44 br_44 wl_112 vdd gnd cell_6t
Xbit_r113_c44 bl_44 br_44 wl_113 vdd gnd cell_6t
Xbit_r114_c44 bl_44 br_44 wl_114 vdd gnd cell_6t
Xbit_r115_c44 bl_44 br_44 wl_115 vdd gnd cell_6t
Xbit_r116_c44 bl_44 br_44 wl_116 vdd gnd cell_6t
Xbit_r117_c44 bl_44 br_44 wl_117 vdd gnd cell_6t
Xbit_r118_c44 bl_44 br_44 wl_118 vdd gnd cell_6t
Xbit_r119_c44 bl_44 br_44 wl_119 vdd gnd cell_6t
Xbit_r120_c44 bl_44 br_44 wl_120 vdd gnd cell_6t
Xbit_r121_c44 bl_44 br_44 wl_121 vdd gnd cell_6t
Xbit_r122_c44 bl_44 br_44 wl_122 vdd gnd cell_6t
Xbit_r123_c44 bl_44 br_44 wl_123 vdd gnd cell_6t
Xbit_r124_c44 bl_44 br_44 wl_124 vdd gnd cell_6t
Xbit_r125_c44 bl_44 br_44 wl_125 vdd gnd cell_6t
Xbit_r126_c44 bl_44 br_44 wl_126 vdd gnd cell_6t
Xbit_r127_c44 bl_44 br_44 wl_127 vdd gnd cell_6t
Xbit_r128_c44 bl_44 br_44 wl_128 vdd gnd cell_6t
Xbit_r129_c44 bl_44 br_44 wl_129 vdd gnd cell_6t
Xbit_r130_c44 bl_44 br_44 wl_130 vdd gnd cell_6t
Xbit_r131_c44 bl_44 br_44 wl_131 vdd gnd cell_6t
Xbit_r132_c44 bl_44 br_44 wl_132 vdd gnd cell_6t
Xbit_r133_c44 bl_44 br_44 wl_133 vdd gnd cell_6t
Xbit_r134_c44 bl_44 br_44 wl_134 vdd gnd cell_6t
Xbit_r135_c44 bl_44 br_44 wl_135 vdd gnd cell_6t
Xbit_r136_c44 bl_44 br_44 wl_136 vdd gnd cell_6t
Xbit_r137_c44 bl_44 br_44 wl_137 vdd gnd cell_6t
Xbit_r138_c44 bl_44 br_44 wl_138 vdd gnd cell_6t
Xbit_r139_c44 bl_44 br_44 wl_139 vdd gnd cell_6t
Xbit_r140_c44 bl_44 br_44 wl_140 vdd gnd cell_6t
Xbit_r141_c44 bl_44 br_44 wl_141 vdd gnd cell_6t
Xbit_r142_c44 bl_44 br_44 wl_142 vdd gnd cell_6t
Xbit_r143_c44 bl_44 br_44 wl_143 vdd gnd cell_6t
Xbit_r144_c44 bl_44 br_44 wl_144 vdd gnd cell_6t
Xbit_r145_c44 bl_44 br_44 wl_145 vdd gnd cell_6t
Xbit_r146_c44 bl_44 br_44 wl_146 vdd gnd cell_6t
Xbit_r147_c44 bl_44 br_44 wl_147 vdd gnd cell_6t
Xbit_r148_c44 bl_44 br_44 wl_148 vdd gnd cell_6t
Xbit_r149_c44 bl_44 br_44 wl_149 vdd gnd cell_6t
Xbit_r150_c44 bl_44 br_44 wl_150 vdd gnd cell_6t
Xbit_r151_c44 bl_44 br_44 wl_151 vdd gnd cell_6t
Xbit_r152_c44 bl_44 br_44 wl_152 vdd gnd cell_6t
Xbit_r153_c44 bl_44 br_44 wl_153 vdd gnd cell_6t
Xbit_r154_c44 bl_44 br_44 wl_154 vdd gnd cell_6t
Xbit_r155_c44 bl_44 br_44 wl_155 vdd gnd cell_6t
Xbit_r156_c44 bl_44 br_44 wl_156 vdd gnd cell_6t
Xbit_r157_c44 bl_44 br_44 wl_157 vdd gnd cell_6t
Xbit_r158_c44 bl_44 br_44 wl_158 vdd gnd cell_6t
Xbit_r159_c44 bl_44 br_44 wl_159 vdd gnd cell_6t
Xbit_r160_c44 bl_44 br_44 wl_160 vdd gnd cell_6t
Xbit_r161_c44 bl_44 br_44 wl_161 vdd gnd cell_6t
Xbit_r162_c44 bl_44 br_44 wl_162 vdd gnd cell_6t
Xbit_r163_c44 bl_44 br_44 wl_163 vdd gnd cell_6t
Xbit_r164_c44 bl_44 br_44 wl_164 vdd gnd cell_6t
Xbit_r165_c44 bl_44 br_44 wl_165 vdd gnd cell_6t
Xbit_r166_c44 bl_44 br_44 wl_166 vdd gnd cell_6t
Xbit_r167_c44 bl_44 br_44 wl_167 vdd gnd cell_6t
Xbit_r168_c44 bl_44 br_44 wl_168 vdd gnd cell_6t
Xbit_r169_c44 bl_44 br_44 wl_169 vdd gnd cell_6t
Xbit_r170_c44 bl_44 br_44 wl_170 vdd gnd cell_6t
Xbit_r171_c44 bl_44 br_44 wl_171 vdd gnd cell_6t
Xbit_r172_c44 bl_44 br_44 wl_172 vdd gnd cell_6t
Xbit_r173_c44 bl_44 br_44 wl_173 vdd gnd cell_6t
Xbit_r174_c44 bl_44 br_44 wl_174 vdd gnd cell_6t
Xbit_r175_c44 bl_44 br_44 wl_175 vdd gnd cell_6t
Xbit_r176_c44 bl_44 br_44 wl_176 vdd gnd cell_6t
Xbit_r177_c44 bl_44 br_44 wl_177 vdd gnd cell_6t
Xbit_r178_c44 bl_44 br_44 wl_178 vdd gnd cell_6t
Xbit_r179_c44 bl_44 br_44 wl_179 vdd gnd cell_6t
Xbit_r180_c44 bl_44 br_44 wl_180 vdd gnd cell_6t
Xbit_r181_c44 bl_44 br_44 wl_181 vdd gnd cell_6t
Xbit_r182_c44 bl_44 br_44 wl_182 vdd gnd cell_6t
Xbit_r183_c44 bl_44 br_44 wl_183 vdd gnd cell_6t
Xbit_r184_c44 bl_44 br_44 wl_184 vdd gnd cell_6t
Xbit_r185_c44 bl_44 br_44 wl_185 vdd gnd cell_6t
Xbit_r186_c44 bl_44 br_44 wl_186 vdd gnd cell_6t
Xbit_r187_c44 bl_44 br_44 wl_187 vdd gnd cell_6t
Xbit_r188_c44 bl_44 br_44 wl_188 vdd gnd cell_6t
Xbit_r189_c44 bl_44 br_44 wl_189 vdd gnd cell_6t
Xbit_r190_c44 bl_44 br_44 wl_190 vdd gnd cell_6t
Xbit_r191_c44 bl_44 br_44 wl_191 vdd gnd cell_6t
Xbit_r192_c44 bl_44 br_44 wl_192 vdd gnd cell_6t
Xbit_r193_c44 bl_44 br_44 wl_193 vdd gnd cell_6t
Xbit_r194_c44 bl_44 br_44 wl_194 vdd gnd cell_6t
Xbit_r195_c44 bl_44 br_44 wl_195 vdd gnd cell_6t
Xbit_r196_c44 bl_44 br_44 wl_196 vdd gnd cell_6t
Xbit_r197_c44 bl_44 br_44 wl_197 vdd gnd cell_6t
Xbit_r198_c44 bl_44 br_44 wl_198 vdd gnd cell_6t
Xbit_r199_c44 bl_44 br_44 wl_199 vdd gnd cell_6t
Xbit_r200_c44 bl_44 br_44 wl_200 vdd gnd cell_6t
Xbit_r201_c44 bl_44 br_44 wl_201 vdd gnd cell_6t
Xbit_r202_c44 bl_44 br_44 wl_202 vdd gnd cell_6t
Xbit_r203_c44 bl_44 br_44 wl_203 vdd gnd cell_6t
Xbit_r204_c44 bl_44 br_44 wl_204 vdd gnd cell_6t
Xbit_r205_c44 bl_44 br_44 wl_205 vdd gnd cell_6t
Xbit_r206_c44 bl_44 br_44 wl_206 vdd gnd cell_6t
Xbit_r207_c44 bl_44 br_44 wl_207 vdd gnd cell_6t
Xbit_r208_c44 bl_44 br_44 wl_208 vdd gnd cell_6t
Xbit_r209_c44 bl_44 br_44 wl_209 vdd gnd cell_6t
Xbit_r210_c44 bl_44 br_44 wl_210 vdd gnd cell_6t
Xbit_r211_c44 bl_44 br_44 wl_211 vdd gnd cell_6t
Xbit_r212_c44 bl_44 br_44 wl_212 vdd gnd cell_6t
Xbit_r213_c44 bl_44 br_44 wl_213 vdd gnd cell_6t
Xbit_r214_c44 bl_44 br_44 wl_214 vdd gnd cell_6t
Xbit_r215_c44 bl_44 br_44 wl_215 vdd gnd cell_6t
Xbit_r216_c44 bl_44 br_44 wl_216 vdd gnd cell_6t
Xbit_r217_c44 bl_44 br_44 wl_217 vdd gnd cell_6t
Xbit_r218_c44 bl_44 br_44 wl_218 vdd gnd cell_6t
Xbit_r219_c44 bl_44 br_44 wl_219 vdd gnd cell_6t
Xbit_r220_c44 bl_44 br_44 wl_220 vdd gnd cell_6t
Xbit_r221_c44 bl_44 br_44 wl_221 vdd gnd cell_6t
Xbit_r222_c44 bl_44 br_44 wl_222 vdd gnd cell_6t
Xbit_r223_c44 bl_44 br_44 wl_223 vdd gnd cell_6t
Xbit_r224_c44 bl_44 br_44 wl_224 vdd gnd cell_6t
Xbit_r225_c44 bl_44 br_44 wl_225 vdd gnd cell_6t
Xbit_r226_c44 bl_44 br_44 wl_226 vdd gnd cell_6t
Xbit_r227_c44 bl_44 br_44 wl_227 vdd gnd cell_6t
Xbit_r228_c44 bl_44 br_44 wl_228 vdd gnd cell_6t
Xbit_r229_c44 bl_44 br_44 wl_229 vdd gnd cell_6t
Xbit_r230_c44 bl_44 br_44 wl_230 vdd gnd cell_6t
Xbit_r231_c44 bl_44 br_44 wl_231 vdd gnd cell_6t
Xbit_r232_c44 bl_44 br_44 wl_232 vdd gnd cell_6t
Xbit_r233_c44 bl_44 br_44 wl_233 vdd gnd cell_6t
Xbit_r234_c44 bl_44 br_44 wl_234 vdd gnd cell_6t
Xbit_r235_c44 bl_44 br_44 wl_235 vdd gnd cell_6t
Xbit_r236_c44 bl_44 br_44 wl_236 vdd gnd cell_6t
Xbit_r237_c44 bl_44 br_44 wl_237 vdd gnd cell_6t
Xbit_r238_c44 bl_44 br_44 wl_238 vdd gnd cell_6t
Xbit_r239_c44 bl_44 br_44 wl_239 vdd gnd cell_6t
Xbit_r240_c44 bl_44 br_44 wl_240 vdd gnd cell_6t
Xbit_r241_c44 bl_44 br_44 wl_241 vdd gnd cell_6t
Xbit_r242_c44 bl_44 br_44 wl_242 vdd gnd cell_6t
Xbit_r243_c44 bl_44 br_44 wl_243 vdd gnd cell_6t
Xbit_r244_c44 bl_44 br_44 wl_244 vdd gnd cell_6t
Xbit_r245_c44 bl_44 br_44 wl_245 vdd gnd cell_6t
Xbit_r246_c44 bl_44 br_44 wl_246 vdd gnd cell_6t
Xbit_r247_c44 bl_44 br_44 wl_247 vdd gnd cell_6t
Xbit_r248_c44 bl_44 br_44 wl_248 vdd gnd cell_6t
Xbit_r249_c44 bl_44 br_44 wl_249 vdd gnd cell_6t
Xbit_r250_c44 bl_44 br_44 wl_250 vdd gnd cell_6t
Xbit_r251_c44 bl_44 br_44 wl_251 vdd gnd cell_6t
Xbit_r252_c44 bl_44 br_44 wl_252 vdd gnd cell_6t
Xbit_r253_c44 bl_44 br_44 wl_253 vdd gnd cell_6t
Xbit_r254_c44 bl_44 br_44 wl_254 vdd gnd cell_6t
Xbit_r255_c44 bl_44 br_44 wl_255 vdd gnd cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd cell_6t
Xbit_r1_c45 bl_45 br_45 wl_1 vdd gnd cell_6t
Xbit_r2_c45 bl_45 br_45 wl_2 vdd gnd cell_6t
Xbit_r3_c45 bl_45 br_45 wl_3 vdd gnd cell_6t
Xbit_r4_c45 bl_45 br_45 wl_4 vdd gnd cell_6t
Xbit_r5_c45 bl_45 br_45 wl_5 vdd gnd cell_6t
Xbit_r6_c45 bl_45 br_45 wl_6 vdd gnd cell_6t
Xbit_r7_c45 bl_45 br_45 wl_7 vdd gnd cell_6t
Xbit_r8_c45 bl_45 br_45 wl_8 vdd gnd cell_6t
Xbit_r9_c45 bl_45 br_45 wl_9 vdd gnd cell_6t
Xbit_r10_c45 bl_45 br_45 wl_10 vdd gnd cell_6t
Xbit_r11_c45 bl_45 br_45 wl_11 vdd gnd cell_6t
Xbit_r12_c45 bl_45 br_45 wl_12 vdd gnd cell_6t
Xbit_r13_c45 bl_45 br_45 wl_13 vdd gnd cell_6t
Xbit_r14_c45 bl_45 br_45 wl_14 vdd gnd cell_6t
Xbit_r15_c45 bl_45 br_45 wl_15 vdd gnd cell_6t
Xbit_r16_c45 bl_45 br_45 wl_16 vdd gnd cell_6t
Xbit_r17_c45 bl_45 br_45 wl_17 vdd gnd cell_6t
Xbit_r18_c45 bl_45 br_45 wl_18 vdd gnd cell_6t
Xbit_r19_c45 bl_45 br_45 wl_19 vdd gnd cell_6t
Xbit_r20_c45 bl_45 br_45 wl_20 vdd gnd cell_6t
Xbit_r21_c45 bl_45 br_45 wl_21 vdd gnd cell_6t
Xbit_r22_c45 bl_45 br_45 wl_22 vdd gnd cell_6t
Xbit_r23_c45 bl_45 br_45 wl_23 vdd gnd cell_6t
Xbit_r24_c45 bl_45 br_45 wl_24 vdd gnd cell_6t
Xbit_r25_c45 bl_45 br_45 wl_25 vdd gnd cell_6t
Xbit_r26_c45 bl_45 br_45 wl_26 vdd gnd cell_6t
Xbit_r27_c45 bl_45 br_45 wl_27 vdd gnd cell_6t
Xbit_r28_c45 bl_45 br_45 wl_28 vdd gnd cell_6t
Xbit_r29_c45 bl_45 br_45 wl_29 vdd gnd cell_6t
Xbit_r30_c45 bl_45 br_45 wl_30 vdd gnd cell_6t
Xbit_r31_c45 bl_45 br_45 wl_31 vdd gnd cell_6t
Xbit_r32_c45 bl_45 br_45 wl_32 vdd gnd cell_6t
Xbit_r33_c45 bl_45 br_45 wl_33 vdd gnd cell_6t
Xbit_r34_c45 bl_45 br_45 wl_34 vdd gnd cell_6t
Xbit_r35_c45 bl_45 br_45 wl_35 vdd gnd cell_6t
Xbit_r36_c45 bl_45 br_45 wl_36 vdd gnd cell_6t
Xbit_r37_c45 bl_45 br_45 wl_37 vdd gnd cell_6t
Xbit_r38_c45 bl_45 br_45 wl_38 vdd gnd cell_6t
Xbit_r39_c45 bl_45 br_45 wl_39 vdd gnd cell_6t
Xbit_r40_c45 bl_45 br_45 wl_40 vdd gnd cell_6t
Xbit_r41_c45 bl_45 br_45 wl_41 vdd gnd cell_6t
Xbit_r42_c45 bl_45 br_45 wl_42 vdd gnd cell_6t
Xbit_r43_c45 bl_45 br_45 wl_43 vdd gnd cell_6t
Xbit_r44_c45 bl_45 br_45 wl_44 vdd gnd cell_6t
Xbit_r45_c45 bl_45 br_45 wl_45 vdd gnd cell_6t
Xbit_r46_c45 bl_45 br_45 wl_46 vdd gnd cell_6t
Xbit_r47_c45 bl_45 br_45 wl_47 vdd gnd cell_6t
Xbit_r48_c45 bl_45 br_45 wl_48 vdd gnd cell_6t
Xbit_r49_c45 bl_45 br_45 wl_49 vdd gnd cell_6t
Xbit_r50_c45 bl_45 br_45 wl_50 vdd gnd cell_6t
Xbit_r51_c45 bl_45 br_45 wl_51 vdd gnd cell_6t
Xbit_r52_c45 bl_45 br_45 wl_52 vdd gnd cell_6t
Xbit_r53_c45 bl_45 br_45 wl_53 vdd gnd cell_6t
Xbit_r54_c45 bl_45 br_45 wl_54 vdd gnd cell_6t
Xbit_r55_c45 bl_45 br_45 wl_55 vdd gnd cell_6t
Xbit_r56_c45 bl_45 br_45 wl_56 vdd gnd cell_6t
Xbit_r57_c45 bl_45 br_45 wl_57 vdd gnd cell_6t
Xbit_r58_c45 bl_45 br_45 wl_58 vdd gnd cell_6t
Xbit_r59_c45 bl_45 br_45 wl_59 vdd gnd cell_6t
Xbit_r60_c45 bl_45 br_45 wl_60 vdd gnd cell_6t
Xbit_r61_c45 bl_45 br_45 wl_61 vdd gnd cell_6t
Xbit_r62_c45 bl_45 br_45 wl_62 vdd gnd cell_6t
Xbit_r63_c45 bl_45 br_45 wl_63 vdd gnd cell_6t
Xbit_r64_c45 bl_45 br_45 wl_64 vdd gnd cell_6t
Xbit_r65_c45 bl_45 br_45 wl_65 vdd gnd cell_6t
Xbit_r66_c45 bl_45 br_45 wl_66 vdd gnd cell_6t
Xbit_r67_c45 bl_45 br_45 wl_67 vdd gnd cell_6t
Xbit_r68_c45 bl_45 br_45 wl_68 vdd gnd cell_6t
Xbit_r69_c45 bl_45 br_45 wl_69 vdd gnd cell_6t
Xbit_r70_c45 bl_45 br_45 wl_70 vdd gnd cell_6t
Xbit_r71_c45 bl_45 br_45 wl_71 vdd gnd cell_6t
Xbit_r72_c45 bl_45 br_45 wl_72 vdd gnd cell_6t
Xbit_r73_c45 bl_45 br_45 wl_73 vdd gnd cell_6t
Xbit_r74_c45 bl_45 br_45 wl_74 vdd gnd cell_6t
Xbit_r75_c45 bl_45 br_45 wl_75 vdd gnd cell_6t
Xbit_r76_c45 bl_45 br_45 wl_76 vdd gnd cell_6t
Xbit_r77_c45 bl_45 br_45 wl_77 vdd gnd cell_6t
Xbit_r78_c45 bl_45 br_45 wl_78 vdd gnd cell_6t
Xbit_r79_c45 bl_45 br_45 wl_79 vdd gnd cell_6t
Xbit_r80_c45 bl_45 br_45 wl_80 vdd gnd cell_6t
Xbit_r81_c45 bl_45 br_45 wl_81 vdd gnd cell_6t
Xbit_r82_c45 bl_45 br_45 wl_82 vdd gnd cell_6t
Xbit_r83_c45 bl_45 br_45 wl_83 vdd gnd cell_6t
Xbit_r84_c45 bl_45 br_45 wl_84 vdd gnd cell_6t
Xbit_r85_c45 bl_45 br_45 wl_85 vdd gnd cell_6t
Xbit_r86_c45 bl_45 br_45 wl_86 vdd gnd cell_6t
Xbit_r87_c45 bl_45 br_45 wl_87 vdd gnd cell_6t
Xbit_r88_c45 bl_45 br_45 wl_88 vdd gnd cell_6t
Xbit_r89_c45 bl_45 br_45 wl_89 vdd gnd cell_6t
Xbit_r90_c45 bl_45 br_45 wl_90 vdd gnd cell_6t
Xbit_r91_c45 bl_45 br_45 wl_91 vdd gnd cell_6t
Xbit_r92_c45 bl_45 br_45 wl_92 vdd gnd cell_6t
Xbit_r93_c45 bl_45 br_45 wl_93 vdd gnd cell_6t
Xbit_r94_c45 bl_45 br_45 wl_94 vdd gnd cell_6t
Xbit_r95_c45 bl_45 br_45 wl_95 vdd gnd cell_6t
Xbit_r96_c45 bl_45 br_45 wl_96 vdd gnd cell_6t
Xbit_r97_c45 bl_45 br_45 wl_97 vdd gnd cell_6t
Xbit_r98_c45 bl_45 br_45 wl_98 vdd gnd cell_6t
Xbit_r99_c45 bl_45 br_45 wl_99 vdd gnd cell_6t
Xbit_r100_c45 bl_45 br_45 wl_100 vdd gnd cell_6t
Xbit_r101_c45 bl_45 br_45 wl_101 vdd gnd cell_6t
Xbit_r102_c45 bl_45 br_45 wl_102 vdd gnd cell_6t
Xbit_r103_c45 bl_45 br_45 wl_103 vdd gnd cell_6t
Xbit_r104_c45 bl_45 br_45 wl_104 vdd gnd cell_6t
Xbit_r105_c45 bl_45 br_45 wl_105 vdd gnd cell_6t
Xbit_r106_c45 bl_45 br_45 wl_106 vdd gnd cell_6t
Xbit_r107_c45 bl_45 br_45 wl_107 vdd gnd cell_6t
Xbit_r108_c45 bl_45 br_45 wl_108 vdd gnd cell_6t
Xbit_r109_c45 bl_45 br_45 wl_109 vdd gnd cell_6t
Xbit_r110_c45 bl_45 br_45 wl_110 vdd gnd cell_6t
Xbit_r111_c45 bl_45 br_45 wl_111 vdd gnd cell_6t
Xbit_r112_c45 bl_45 br_45 wl_112 vdd gnd cell_6t
Xbit_r113_c45 bl_45 br_45 wl_113 vdd gnd cell_6t
Xbit_r114_c45 bl_45 br_45 wl_114 vdd gnd cell_6t
Xbit_r115_c45 bl_45 br_45 wl_115 vdd gnd cell_6t
Xbit_r116_c45 bl_45 br_45 wl_116 vdd gnd cell_6t
Xbit_r117_c45 bl_45 br_45 wl_117 vdd gnd cell_6t
Xbit_r118_c45 bl_45 br_45 wl_118 vdd gnd cell_6t
Xbit_r119_c45 bl_45 br_45 wl_119 vdd gnd cell_6t
Xbit_r120_c45 bl_45 br_45 wl_120 vdd gnd cell_6t
Xbit_r121_c45 bl_45 br_45 wl_121 vdd gnd cell_6t
Xbit_r122_c45 bl_45 br_45 wl_122 vdd gnd cell_6t
Xbit_r123_c45 bl_45 br_45 wl_123 vdd gnd cell_6t
Xbit_r124_c45 bl_45 br_45 wl_124 vdd gnd cell_6t
Xbit_r125_c45 bl_45 br_45 wl_125 vdd gnd cell_6t
Xbit_r126_c45 bl_45 br_45 wl_126 vdd gnd cell_6t
Xbit_r127_c45 bl_45 br_45 wl_127 vdd gnd cell_6t
Xbit_r128_c45 bl_45 br_45 wl_128 vdd gnd cell_6t
Xbit_r129_c45 bl_45 br_45 wl_129 vdd gnd cell_6t
Xbit_r130_c45 bl_45 br_45 wl_130 vdd gnd cell_6t
Xbit_r131_c45 bl_45 br_45 wl_131 vdd gnd cell_6t
Xbit_r132_c45 bl_45 br_45 wl_132 vdd gnd cell_6t
Xbit_r133_c45 bl_45 br_45 wl_133 vdd gnd cell_6t
Xbit_r134_c45 bl_45 br_45 wl_134 vdd gnd cell_6t
Xbit_r135_c45 bl_45 br_45 wl_135 vdd gnd cell_6t
Xbit_r136_c45 bl_45 br_45 wl_136 vdd gnd cell_6t
Xbit_r137_c45 bl_45 br_45 wl_137 vdd gnd cell_6t
Xbit_r138_c45 bl_45 br_45 wl_138 vdd gnd cell_6t
Xbit_r139_c45 bl_45 br_45 wl_139 vdd gnd cell_6t
Xbit_r140_c45 bl_45 br_45 wl_140 vdd gnd cell_6t
Xbit_r141_c45 bl_45 br_45 wl_141 vdd gnd cell_6t
Xbit_r142_c45 bl_45 br_45 wl_142 vdd gnd cell_6t
Xbit_r143_c45 bl_45 br_45 wl_143 vdd gnd cell_6t
Xbit_r144_c45 bl_45 br_45 wl_144 vdd gnd cell_6t
Xbit_r145_c45 bl_45 br_45 wl_145 vdd gnd cell_6t
Xbit_r146_c45 bl_45 br_45 wl_146 vdd gnd cell_6t
Xbit_r147_c45 bl_45 br_45 wl_147 vdd gnd cell_6t
Xbit_r148_c45 bl_45 br_45 wl_148 vdd gnd cell_6t
Xbit_r149_c45 bl_45 br_45 wl_149 vdd gnd cell_6t
Xbit_r150_c45 bl_45 br_45 wl_150 vdd gnd cell_6t
Xbit_r151_c45 bl_45 br_45 wl_151 vdd gnd cell_6t
Xbit_r152_c45 bl_45 br_45 wl_152 vdd gnd cell_6t
Xbit_r153_c45 bl_45 br_45 wl_153 vdd gnd cell_6t
Xbit_r154_c45 bl_45 br_45 wl_154 vdd gnd cell_6t
Xbit_r155_c45 bl_45 br_45 wl_155 vdd gnd cell_6t
Xbit_r156_c45 bl_45 br_45 wl_156 vdd gnd cell_6t
Xbit_r157_c45 bl_45 br_45 wl_157 vdd gnd cell_6t
Xbit_r158_c45 bl_45 br_45 wl_158 vdd gnd cell_6t
Xbit_r159_c45 bl_45 br_45 wl_159 vdd gnd cell_6t
Xbit_r160_c45 bl_45 br_45 wl_160 vdd gnd cell_6t
Xbit_r161_c45 bl_45 br_45 wl_161 vdd gnd cell_6t
Xbit_r162_c45 bl_45 br_45 wl_162 vdd gnd cell_6t
Xbit_r163_c45 bl_45 br_45 wl_163 vdd gnd cell_6t
Xbit_r164_c45 bl_45 br_45 wl_164 vdd gnd cell_6t
Xbit_r165_c45 bl_45 br_45 wl_165 vdd gnd cell_6t
Xbit_r166_c45 bl_45 br_45 wl_166 vdd gnd cell_6t
Xbit_r167_c45 bl_45 br_45 wl_167 vdd gnd cell_6t
Xbit_r168_c45 bl_45 br_45 wl_168 vdd gnd cell_6t
Xbit_r169_c45 bl_45 br_45 wl_169 vdd gnd cell_6t
Xbit_r170_c45 bl_45 br_45 wl_170 vdd gnd cell_6t
Xbit_r171_c45 bl_45 br_45 wl_171 vdd gnd cell_6t
Xbit_r172_c45 bl_45 br_45 wl_172 vdd gnd cell_6t
Xbit_r173_c45 bl_45 br_45 wl_173 vdd gnd cell_6t
Xbit_r174_c45 bl_45 br_45 wl_174 vdd gnd cell_6t
Xbit_r175_c45 bl_45 br_45 wl_175 vdd gnd cell_6t
Xbit_r176_c45 bl_45 br_45 wl_176 vdd gnd cell_6t
Xbit_r177_c45 bl_45 br_45 wl_177 vdd gnd cell_6t
Xbit_r178_c45 bl_45 br_45 wl_178 vdd gnd cell_6t
Xbit_r179_c45 bl_45 br_45 wl_179 vdd gnd cell_6t
Xbit_r180_c45 bl_45 br_45 wl_180 vdd gnd cell_6t
Xbit_r181_c45 bl_45 br_45 wl_181 vdd gnd cell_6t
Xbit_r182_c45 bl_45 br_45 wl_182 vdd gnd cell_6t
Xbit_r183_c45 bl_45 br_45 wl_183 vdd gnd cell_6t
Xbit_r184_c45 bl_45 br_45 wl_184 vdd gnd cell_6t
Xbit_r185_c45 bl_45 br_45 wl_185 vdd gnd cell_6t
Xbit_r186_c45 bl_45 br_45 wl_186 vdd gnd cell_6t
Xbit_r187_c45 bl_45 br_45 wl_187 vdd gnd cell_6t
Xbit_r188_c45 bl_45 br_45 wl_188 vdd gnd cell_6t
Xbit_r189_c45 bl_45 br_45 wl_189 vdd gnd cell_6t
Xbit_r190_c45 bl_45 br_45 wl_190 vdd gnd cell_6t
Xbit_r191_c45 bl_45 br_45 wl_191 vdd gnd cell_6t
Xbit_r192_c45 bl_45 br_45 wl_192 vdd gnd cell_6t
Xbit_r193_c45 bl_45 br_45 wl_193 vdd gnd cell_6t
Xbit_r194_c45 bl_45 br_45 wl_194 vdd gnd cell_6t
Xbit_r195_c45 bl_45 br_45 wl_195 vdd gnd cell_6t
Xbit_r196_c45 bl_45 br_45 wl_196 vdd gnd cell_6t
Xbit_r197_c45 bl_45 br_45 wl_197 vdd gnd cell_6t
Xbit_r198_c45 bl_45 br_45 wl_198 vdd gnd cell_6t
Xbit_r199_c45 bl_45 br_45 wl_199 vdd gnd cell_6t
Xbit_r200_c45 bl_45 br_45 wl_200 vdd gnd cell_6t
Xbit_r201_c45 bl_45 br_45 wl_201 vdd gnd cell_6t
Xbit_r202_c45 bl_45 br_45 wl_202 vdd gnd cell_6t
Xbit_r203_c45 bl_45 br_45 wl_203 vdd gnd cell_6t
Xbit_r204_c45 bl_45 br_45 wl_204 vdd gnd cell_6t
Xbit_r205_c45 bl_45 br_45 wl_205 vdd gnd cell_6t
Xbit_r206_c45 bl_45 br_45 wl_206 vdd gnd cell_6t
Xbit_r207_c45 bl_45 br_45 wl_207 vdd gnd cell_6t
Xbit_r208_c45 bl_45 br_45 wl_208 vdd gnd cell_6t
Xbit_r209_c45 bl_45 br_45 wl_209 vdd gnd cell_6t
Xbit_r210_c45 bl_45 br_45 wl_210 vdd gnd cell_6t
Xbit_r211_c45 bl_45 br_45 wl_211 vdd gnd cell_6t
Xbit_r212_c45 bl_45 br_45 wl_212 vdd gnd cell_6t
Xbit_r213_c45 bl_45 br_45 wl_213 vdd gnd cell_6t
Xbit_r214_c45 bl_45 br_45 wl_214 vdd gnd cell_6t
Xbit_r215_c45 bl_45 br_45 wl_215 vdd gnd cell_6t
Xbit_r216_c45 bl_45 br_45 wl_216 vdd gnd cell_6t
Xbit_r217_c45 bl_45 br_45 wl_217 vdd gnd cell_6t
Xbit_r218_c45 bl_45 br_45 wl_218 vdd gnd cell_6t
Xbit_r219_c45 bl_45 br_45 wl_219 vdd gnd cell_6t
Xbit_r220_c45 bl_45 br_45 wl_220 vdd gnd cell_6t
Xbit_r221_c45 bl_45 br_45 wl_221 vdd gnd cell_6t
Xbit_r222_c45 bl_45 br_45 wl_222 vdd gnd cell_6t
Xbit_r223_c45 bl_45 br_45 wl_223 vdd gnd cell_6t
Xbit_r224_c45 bl_45 br_45 wl_224 vdd gnd cell_6t
Xbit_r225_c45 bl_45 br_45 wl_225 vdd gnd cell_6t
Xbit_r226_c45 bl_45 br_45 wl_226 vdd gnd cell_6t
Xbit_r227_c45 bl_45 br_45 wl_227 vdd gnd cell_6t
Xbit_r228_c45 bl_45 br_45 wl_228 vdd gnd cell_6t
Xbit_r229_c45 bl_45 br_45 wl_229 vdd gnd cell_6t
Xbit_r230_c45 bl_45 br_45 wl_230 vdd gnd cell_6t
Xbit_r231_c45 bl_45 br_45 wl_231 vdd gnd cell_6t
Xbit_r232_c45 bl_45 br_45 wl_232 vdd gnd cell_6t
Xbit_r233_c45 bl_45 br_45 wl_233 vdd gnd cell_6t
Xbit_r234_c45 bl_45 br_45 wl_234 vdd gnd cell_6t
Xbit_r235_c45 bl_45 br_45 wl_235 vdd gnd cell_6t
Xbit_r236_c45 bl_45 br_45 wl_236 vdd gnd cell_6t
Xbit_r237_c45 bl_45 br_45 wl_237 vdd gnd cell_6t
Xbit_r238_c45 bl_45 br_45 wl_238 vdd gnd cell_6t
Xbit_r239_c45 bl_45 br_45 wl_239 vdd gnd cell_6t
Xbit_r240_c45 bl_45 br_45 wl_240 vdd gnd cell_6t
Xbit_r241_c45 bl_45 br_45 wl_241 vdd gnd cell_6t
Xbit_r242_c45 bl_45 br_45 wl_242 vdd gnd cell_6t
Xbit_r243_c45 bl_45 br_45 wl_243 vdd gnd cell_6t
Xbit_r244_c45 bl_45 br_45 wl_244 vdd gnd cell_6t
Xbit_r245_c45 bl_45 br_45 wl_245 vdd gnd cell_6t
Xbit_r246_c45 bl_45 br_45 wl_246 vdd gnd cell_6t
Xbit_r247_c45 bl_45 br_45 wl_247 vdd gnd cell_6t
Xbit_r248_c45 bl_45 br_45 wl_248 vdd gnd cell_6t
Xbit_r249_c45 bl_45 br_45 wl_249 vdd gnd cell_6t
Xbit_r250_c45 bl_45 br_45 wl_250 vdd gnd cell_6t
Xbit_r251_c45 bl_45 br_45 wl_251 vdd gnd cell_6t
Xbit_r252_c45 bl_45 br_45 wl_252 vdd gnd cell_6t
Xbit_r253_c45 bl_45 br_45 wl_253 vdd gnd cell_6t
Xbit_r254_c45 bl_45 br_45 wl_254 vdd gnd cell_6t
Xbit_r255_c45 bl_45 br_45 wl_255 vdd gnd cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd cell_6t
Xbit_r1_c46 bl_46 br_46 wl_1 vdd gnd cell_6t
Xbit_r2_c46 bl_46 br_46 wl_2 vdd gnd cell_6t
Xbit_r3_c46 bl_46 br_46 wl_3 vdd gnd cell_6t
Xbit_r4_c46 bl_46 br_46 wl_4 vdd gnd cell_6t
Xbit_r5_c46 bl_46 br_46 wl_5 vdd gnd cell_6t
Xbit_r6_c46 bl_46 br_46 wl_6 vdd gnd cell_6t
Xbit_r7_c46 bl_46 br_46 wl_7 vdd gnd cell_6t
Xbit_r8_c46 bl_46 br_46 wl_8 vdd gnd cell_6t
Xbit_r9_c46 bl_46 br_46 wl_9 vdd gnd cell_6t
Xbit_r10_c46 bl_46 br_46 wl_10 vdd gnd cell_6t
Xbit_r11_c46 bl_46 br_46 wl_11 vdd gnd cell_6t
Xbit_r12_c46 bl_46 br_46 wl_12 vdd gnd cell_6t
Xbit_r13_c46 bl_46 br_46 wl_13 vdd gnd cell_6t
Xbit_r14_c46 bl_46 br_46 wl_14 vdd gnd cell_6t
Xbit_r15_c46 bl_46 br_46 wl_15 vdd gnd cell_6t
Xbit_r16_c46 bl_46 br_46 wl_16 vdd gnd cell_6t
Xbit_r17_c46 bl_46 br_46 wl_17 vdd gnd cell_6t
Xbit_r18_c46 bl_46 br_46 wl_18 vdd gnd cell_6t
Xbit_r19_c46 bl_46 br_46 wl_19 vdd gnd cell_6t
Xbit_r20_c46 bl_46 br_46 wl_20 vdd gnd cell_6t
Xbit_r21_c46 bl_46 br_46 wl_21 vdd gnd cell_6t
Xbit_r22_c46 bl_46 br_46 wl_22 vdd gnd cell_6t
Xbit_r23_c46 bl_46 br_46 wl_23 vdd gnd cell_6t
Xbit_r24_c46 bl_46 br_46 wl_24 vdd gnd cell_6t
Xbit_r25_c46 bl_46 br_46 wl_25 vdd gnd cell_6t
Xbit_r26_c46 bl_46 br_46 wl_26 vdd gnd cell_6t
Xbit_r27_c46 bl_46 br_46 wl_27 vdd gnd cell_6t
Xbit_r28_c46 bl_46 br_46 wl_28 vdd gnd cell_6t
Xbit_r29_c46 bl_46 br_46 wl_29 vdd gnd cell_6t
Xbit_r30_c46 bl_46 br_46 wl_30 vdd gnd cell_6t
Xbit_r31_c46 bl_46 br_46 wl_31 vdd gnd cell_6t
Xbit_r32_c46 bl_46 br_46 wl_32 vdd gnd cell_6t
Xbit_r33_c46 bl_46 br_46 wl_33 vdd gnd cell_6t
Xbit_r34_c46 bl_46 br_46 wl_34 vdd gnd cell_6t
Xbit_r35_c46 bl_46 br_46 wl_35 vdd gnd cell_6t
Xbit_r36_c46 bl_46 br_46 wl_36 vdd gnd cell_6t
Xbit_r37_c46 bl_46 br_46 wl_37 vdd gnd cell_6t
Xbit_r38_c46 bl_46 br_46 wl_38 vdd gnd cell_6t
Xbit_r39_c46 bl_46 br_46 wl_39 vdd gnd cell_6t
Xbit_r40_c46 bl_46 br_46 wl_40 vdd gnd cell_6t
Xbit_r41_c46 bl_46 br_46 wl_41 vdd gnd cell_6t
Xbit_r42_c46 bl_46 br_46 wl_42 vdd gnd cell_6t
Xbit_r43_c46 bl_46 br_46 wl_43 vdd gnd cell_6t
Xbit_r44_c46 bl_46 br_46 wl_44 vdd gnd cell_6t
Xbit_r45_c46 bl_46 br_46 wl_45 vdd gnd cell_6t
Xbit_r46_c46 bl_46 br_46 wl_46 vdd gnd cell_6t
Xbit_r47_c46 bl_46 br_46 wl_47 vdd gnd cell_6t
Xbit_r48_c46 bl_46 br_46 wl_48 vdd gnd cell_6t
Xbit_r49_c46 bl_46 br_46 wl_49 vdd gnd cell_6t
Xbit_r50_c46 bl_46 br_46 wl_50 vdd gnd cell_6t
Xbit_r51_c46 bl_46 br_46 wl_51 vdd gnd cell_6t
Xbit_r52_c46 bl_46 br_46 wl_52 vdd gnd cell_6t
Xbit_r53_c46 bl_46 br_46 wl_53 vdd gnd cell_6t
Xbit_r54_c46 bl_46 br_46 wl_54 vdd gnd cell_6t
Xbit_r55_c46 bl_46 br_46 wl_55 vdd gnd cell_6t
Xbit_r56_c46 bl_46 br_46 wl_56 vdd gnd cell_6t
Xbit_r57_c46 bl_46 br_46 wl_57 vdd gnd cell_6t
Xbit_r58_c46 bl_46 br_46 wl_58 vdd gnd cell_6t
Xbit_r59_c46 bl_46 br_46 wl_59 vdd gnd cell_6t
Xbit_r60_c46 bl_46 br_46 wl_60 vdd gnd cell_6t
Xbit_r61_c46 bl_46 br_46 wl_61 vdd gnd cell_6t
Xbit_r62_c46 bl_46 br_46 wl_62 vdd gnd cell_6t
Xbit_r63_c46 bl_46 br_46 wl_63 vdd gnd cell_6t
Xbit_r64_c46 bl_46 br_46 wl_64 vdd gnd cell_6t
Xbit_r65_c46 bl_46 br_46 wl_65 vdd gnd cell_6t
Xbit_r66_c46 bl_46 br_46 wl_66 vdd gnd cell_6t
Xbit_r67_c46 bl_46 br_46 wl_67 vdd gnd cell_6t
Xbit_r68_c46 bl_46 br_46 wl_68 vdd gnd cell_6t
Xbit_r69_c46 bl_46 br_46 wl_69 vdd gnd cell_6t
Xbit_r70_c46 bl_46 br_46 wl_70 vdd gnd cell_6t
Xbit_r71_c46 bl_46 br_46 wl_71 vdd gnd cell_6t
Xbit_r72_c46 bl_46 br_46 wl_72 vdd gnd cell_6t
Xbit_r73_c46 bl_46 br_46 wl_73 vdd gnd cell_6t
Xbit_r74_c46 bl_46 br_46 wl_74 vdd gnd cell_6t
Xbit_r75_c46 bl_46 br_46 wl_75 vdd gnd cell_6t
Xbit_r76_c46 bl_46 br_46 wl_76 vdd gnd cell_6t
Xbit_r77_c46 bl_46 br_46 wl_77 vdd gnd cell_6t
Xbit_r78_c46 bl_46 br_46 wl_78 vdd gnd cell_6t
Xbit_r79_c46 bl_46 br_46 wl_79 vdd gnd cell_6t
Xbit_r80_c46 bl_46 br_46 wl_80 vdd gnd cell_6t
Xbit_r81_c46 bl_46 br_46 wl_81 vdd gnd cell_6t
Xbit_r82_c46 bl_46 br_46 wl_82 vdd gnd cell_6t
Xbit_r83_c46 bl_46 br_46 wl_83 vdd gnd cell_6t
Xbit_r84_c46 bl_46 br_46 wl_84 vdd gnd cell_6t
Xbit_r85_c46 bl_46 br_46 wl_85 vdd gnd cell_6t
Xbit_r86_c46 bl_46 br_46 wl_86 vdd gnd cell_6t
Xbit_r87_c46 bl_46 br_46 wl_87 vdd gnd cell_6t
Xbit_r88_c46 bl_46 br_46 wl_88 vdd gnd cell_6t
Xbit_r89_c46 bl_46 br_46 wl_89 vdd gnd cell_6t
Xbit_r90_c46 bl_46 br_46 wl_90 vdd gnd cell_6t
Xbit_r91_c46 bl_46 br_46 wl_91 vdd gnd cell_6t
Xbit_r92_c46 bl_46 br_46 wl_92 vdd gnd cell_6t
Xbit_r93_c46 bl_46 br_46 wl_93 vdd gnd cell_6t
Xbit_r94_c46 bl_46 br_46 wl_94 vdd gnd cell_6t
Xbit_r95_c46 bl_46 br_46 wl_95 vdd gnd cell_6t
Xbit_r96_c46 bl_46 br_46 wl_96 vdd gnd cell_6t
Xbit_r97_c46 bl_46 br_46 wl_97 vdd gnd cell_6t
Xbit_r98_c46 bl_46 br_46 wl_98 vdd gnd cell_6t
Xbit_r99_c46 bl_46 br_46 wl_99 vdd gnd cell_6t
Xbit_r100_c46 bl_46 br_46 wl_100 vdd gnd cell_6t
Xbit_r101_c46 bl_46 br_46 wl_101 vdd gnd cell_6t
Xbit_r102_c46 bl_46 br_46 wl_102 vdd gnd cell_6t
Xbit_r103_c46 bl_46 br_46 wl_103 vdd gnd cell_6t
Xbit_r104_c46 bl_46 br_46 wl_104 vdd gnd cell_6t
Xbit_r105_c46 bl_46 br_46 wl_105 vdd gnd cell_6t
Xbit_r106_c46 bl_46 br_46 wl_106 vdd gnd cell_6t
Xbit_r107_c46 bl_46 br_46 wl_107 vdd gnd cell_6t
Xbit_r108_c46 bl_46 br_46 wl_108 vdd gnd cell_6t
Xbit_r109_c46 bl_46 br_46 wl_109 vdd gnd cell_6t
Xbit_r110_c46 bl_46 br_46 wl_110 vdd gnd cell_6t
Xbit_r111_c46 bl_46 br_46 wl_111 vdd gnd cell_6t
Xbit_r112_c46 bl_46 br_46 wl_112 vdd gnd cell_6t
Xbit_r113_c46 bl_46 br_46 wl_113 vdd gnd cell_6t
Xbit_r114_c46 bl_46 br_46 wl_114 vdd gnd cell_6t
Xbit_r115_c46 bl_46 br_46 wl_115 vdd gnd cell_6t
Xbit_r116_c46 bl_46 br_46 wl_116 vdd gnd cell_6t
Xbit_r117_c46 bl_46 br_46 wl_117 vdd gnd cell_6t
Xbit_r118_c46 bl_46 br_46 wl_118 vdd gnd cell_6t
Xbit_r119_c46 bl_46 br_46 wl_119 vdd gnd cell_6t
Xbit_r120_c46 bl_46 br_46 wl_120 vdd gnd cell_6t
Xbit_r121_c46 bl_46 br_46 wl_121 vdd gnd cell_6t
Xbit_r122_c46 bl_46 br_46 wl_122 vdd gnd cell_6t
Xbit_r123_c46 bl_46 br_46 wl_123 vdd gnd cell_6t
Xbit_r124_c46 bl_46 br_46 wl_124 vdd gnd cell_6t
Xbit_r125_c46 bl_46 br_46 wl_125 vdd gnd cell_6t
Xbit_r126_c46 bl_46 br_46 wl_126 vdd gnd cell_6t
Xbit_r127_c46 bl_46 br_46 wl_127 vdd gnd cell_6t
Xbit_r128_c46 bl_46 br_46 wl_128 vdd gnd cell_6t
Xbit_r129_c46 bl_46 br_46 wl_129 vdd gnd cell_6t
Xbit_r130_c46 bl_46 br_46 wl_130 vdd gnd cell_6t
Xbit_r131_c46 bl_46 br_46 wl_131 vdd gnd cell_6t
Xbit_r132_c46 bl_46 br_46 wl_132 vdd gnd cell_6t
Xbit_r133_c46 bl_46 br_46 wl_133 vdd gnd cell_6t
Xbit_r134_c46 bl_46 br_46 wl_134 vdd gnd cell_6t
Xbit_r135_c46 bl_46 br_46 wl_135 vdd gnd cell_6t
Xbit_r136_c46 bl_46 br_46 wl_136 vdd gnd cell_6t
Xbit_r137_c46 bl_46 br_46 wl_137 vdd gnd cell_6t
Xbit_r138_c46 bl_46 br_46 wl_138 vdd gnd cell_6t
Xbit_r139_c46 bl_46 br_46 wl_139 vdd gnd cell_6t
Xbit_r140_c46 bl_46 br_46 wl_140 vdd gnd cell_6t
Xbit_r141_c46 bl_46 br_46 wl_141 vdd gnd cell_6t
Xbit_r142_c46 bl_46 br_46 wl_142 vdd gnd cell_6t
Xbit_r143_c46 bl_46 br_46 wl_143 vdd gnd cell_6t
Xbit_r144_c46 bl_46 br_46 wl_144 vdd gnd cell_6t
Xbit_r145_c46 bl_46 br_46 wl_145 vdd gnd cell_6t
Xbit_r146_c46 bl_46 br_46 wl_146 vdd gnd cell_6t
Xbit_r147_c46 bl_46 br_46 wl_147 vdd gnd cell_6t
Xbit_r148_c46 bl_46 br_46 wl_148 vdd gnd cell_6t
Xbit_r149_c46 bl_46 br_46 wl_149 vdd gnd cell_6t
Xbit_r150_c46 bl_46 br_46 wl_150 vdd gnd cell_6t
Xbit_r151_c46 bl_46 br_46 wl_151 vdd gnd cell_6t
Xbit_r152_c46 bl_46 br_46 wl_152 vdd gnd cell_6t
Xbit_r153_c46 bl_46 br_46 wl_153 vdd gnd cell_6t
Xbit_r154_c46 bl_46 br_46 wl_154 vdd gnd cell_6t
Xbit_r155_c46 bl_46 br_46 wl_155 vdd gnd cell_6t
Xbit_r156_c46 bl_46 br_46 wl_156 vdd gnd cell_6t
Xbit_r157_c46 bl_46 br_46 wl_157 vdd gnd cell_6t
Xbit_r158_c46 bl_46 br_46 wl_158 vdd gnd cell_6t
Xbit_r159_c46 bl_46 br_46 wl_159 vdd gnd cell_6t
Xbit_r160_c46 bl_46 br_46 wl_160 vdd gnd cell_6t
Xbit_r161_c46 bl_46 br_46 wl_161 vdd gnd cell_6t
Xbit_r162_c46 bl_46 br_46 wl_162 vdd gnd cell_6t
Xbit_r163_c46 bl_46 br_46 wl_163 vdd gnd cell_6t
Xbit_r164_c46 bl_46 br_46 wl_164 vdd gnd cell_6t
Xbit_r165_c46 bl_46 br_46 wl_165 vdd gnd cell_6t
Xbit_r166_c46 bl_46 br_46 wl_166 vdd gnd cell_6t
Xbit_r167_c46 bl_46 br_46 wl_167 vdd gnd cell_6t
Xbit_r168_c46 bl_46 br_46 wl_168 vdd gnd cell_6t
Xbit_r169_c46 bl_46 br_46 wl_169 vdd gnd cell_6t
Xbit_r170_c46 bl_46 br_46 wl_170 vdd gnd cell_6t
Xbit_r171_c46 bl_46 br_46 wl_171 vdd gnd cell_6t
Xbit_r172_c46 bl_46 br_46 wl_172 vdd gnd cell_6t
Xbit_r173_c46 bl_46 br_46 wl_173 vdd gnd cell_6t
Xbit_r174_c46 bl_46 br_46 wl_174 vdd gnd cell_6t
Xbit_r175_c46 bl_46 br_46 wl_175 vdd gnd cell_6t
Xbit_r176_c46 bl_46 br_46 wl_176 vdd gnd cell_6t
Xbit_r177_c46 bl_46 br_46 wl_177 vdd gnd cell_6t
Xbit_r178_c46 bl_46 br_46 wl_178 vdd gnd cell_6t
Xbit_r179_c46 bl_46 br_46 wl_179 vdd gnd cell_6t
Xbit_r180_c46 bl_46 br_46 wl_180 vdd gnd cell_6t
Xbit_r181_c46 bl_46 br_46 wl_181 vdd gnd cell_6t
Xbit_r182_c46 bl_46 br_46 wl_182 vdd gnd cell_6t
Xbit_r183_c46 bl_46 br_46 wl_183 vdd gnd cell_6t
Xbit_r184_c46 bl_46 br_46 wl_184 vdd gnd cell_6t
Xbit_r185_c46 bl_46 br_46 wl_185 vdd gnd cell_6t
Xbit_r186_c46 bl_46 br_46 wl_186 vdd gnd cell_6t
Xbit_r187_c46 bl_46 br_46 wl_187 vdd gnd cell_6t
Xbit_r188_c46 bl_46 br_46 wl_188 vdd gnd cell_6t
Xbit_r189_c46 bl_46 br_46 wl_189 vdd gnd cell_6t
Xbit_r190_c46 bl_46 br_46 wl_190 vdd gnd cell_6t
Xbit_r191_c46 bl_46 br_46 wl_191 vdd gnd cell_6t
Xbit_r192_c46 bl_46 br_46 wl_192 vdd gnd cell_6t
Xbit_r193_c46 bl_46 br_46 wl_193 vdd gnd cell_6t
Xbit_r194_c46 bl_46 br_46 wl_194 vdd gnd cell_6t
Xbit_r195_c46 bl_46 br_46 wl_195 vdd gnd cell_6t
Xbit_r196_c46 bl_46 br_46 wl_196 vdd gnd cell_6t
Xbit_r197_c46 bl_46 br_46 wl_197 vdd gnd cell_6t
Xbit_r198_c46 bl_46 br_46 wl_198 vdd gnd cell_6t
Xbit_r199_c46 bl_46 br_46 wl_199 vdd gnd cell_6t
Xbit_r200_c46 bl_46 br_46 wl_200 vdd gnd cell_6t
Xbit_r201_c46 bl_46 br_46 wl_201 vdd gnd cell_6t
Xbit_r202_c46 bl_46 br_46 wl_202 vdd gnd cell_6t
Xbit_r203_c46 bl_46 br_46 wl_203 vdd gnd cell_6t
Xbit_r204_c46 bl_46 br_46 wl_204 vdd gnd cell_6t
Xbit_r205_c46 bl_46 br_46 wl_205 vdd gnd cell_6t
Xbit_r206_c46 bl_46 br_46 wl_206 vdd gnd cell_6t
Xbit_r207_c46 bl_46 br_46 wl_207 vdd gnd cell_6t
Xbit_r208_c46 bl_46 br_46 wl_208 vdd gnd cell_6t
Xbit_r209_c46 bl_46 br_46 wl_209 vdd gnd cell_6t
Xbit_r210_c46 bl_46 br_46 wl_210 vdd gnd cell_6t
Xbit_r211_c46 bl_46 br_46 wl_211 vdd gnd cell_6t
Xbit_r212_c46 bl_46 br_46 wl_212 vdd gnd cell_6t
Xbit_r213_c46 bl_46 br_46 wl_213 vdd gnd cell_6t
Xbit_r214_c46 bl_46 br_46 wl_214 vdd gnd cell_6t
Xbit_r215_c46 bl_46 br_46 wl_215 vdd gnd cell_6t
Xbit_r216_c46 bl_46 br_46 wl_216 vdd gnd cell_6t
Xbit_r217_c46 bl_46 br_46 wl_217 vdd gnd cell_6t
Xbit_r218_c46 bl_46 br_46 wl_218 vdd gnd cell_6t
Xbit_r219_c46 bl_46 br_46 wl_219 vdd gnd cell_6t
Xbit_r220_c46 bl_46 br_46 wl_220 vdd gnd cell_6t
Xbit_r221_c46 bl_46 br_46 wl_221 vdd gnd cell_6t
Xbit_r222_c46 bl_46 br_46 wl_222 vdd gnd cell_6t
Xbit_r223_c46 bl_46 br_46 wl_223 vdd gnd cell_6t
Xbit_r224_c46 bl_46 br_46 wl_224 vdd gnd cell_6t
Xbit_r225_c46 bl_46 br_46 wl_225 vdd gnd cell_6t
Xbit_r226_c46 bl_46 br_46 wl_226 vdd gnd cell_6t
Xbit_r227_c46 bl_46 br_46 wl_227 vdd gnd cell_6t
Xbit_r228_c46 bl_46 br_46 wl_228 vdd gnd cell_6t
Xbit_r229_c46 bl_46 br_46 wl_229 vdd gnd cell_6t
Xbit_r230_c46 bl_46 br_46 wl_230 vdd gnd cell_6t
Xbit_r231_c46 bl_46 br_46 wl_231 vdd gnd cell_6t
Xbit_r232_c46 bl_46 br_46 wl_232 vdd gnd cell_6t
Xbit_r233_c46 bl_46 br_46 wl_233 vdd gnd cell_6t
Xbit_r234_c46 bl_46 br_46 wl_234 vdd gnd cell_6t
Xbit_r235_c46 bl_46 br_46 wl_235 vdd gnd cell_6t
Xbit_r236_c46 bl_46 br_46 wl_236 vdd gnd cell_6t
Xbit_r237_c46 bl_46 br_46 wl_237 vdd gnd cell_6t
Xbit_r238_c46 bl_46 br_46 wl_238 vdd gnd cell_6t
Xbit_r239_c46 bl_46 br_46 wl_239 vdd gnd cell_6t
Xbit_r240_c46 bl_46 br_46 wl_240 vdd gnd cell_6t
Xbit_r241_c46 bl_46 br_46 wl_241 vdd gnd cell_6t
Xbit_r242_c46 bl_46 br_46 wl_242 vdd gnd cell_6t
Xbit_r243_c46 bl_46 br_46 wl_243 vdd gnd cell_6t
Xbit_r244_c46 bl_46 br_46 wl_244 vdd gnd cell_6t
Xbit_r245_c46 bl_46 br_46 wl_245 vdd gnd cell_6t
Xbit_r246_c46 bl_46 br_46 wl_246 vdd gnd cell_6t
Xbit_r247_c46 bl_46 br_46 wl_247 vdd gnd cell_6t
Xbit_r248_c46 bl_46 br_46 wl_248 vdd gnd cell_6t
Xbit_r249_c46 bl_46 br_46 wl_249 vdd gnd cell_6t
Xbit_r250_c46 bl_46 br_46 wl_250 vdd gnd cell_6t
Xbit_r251_c46 bl_46 br_46 wl_251 vdd gnd cell_6t
Xbit_r252_c46 bl_46 br_46 wl_252 vdd gnd cell_6t
Xbit_r253_c46 bl_46 br_46 wl_253 vdd gnd cell_6t
Xbit_r254_c46 bl_46 br_46 wl_254 vdd gnd cell_6t
Xbit_r255_c46 bl_46 br_46 wl_255 vdd gnd cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd cell_6t
Xbit_r1_c47 bl_47 br_47 wl_1 vdd gnd cell_6t
Xbit_r2_c47 bl_47 br_47 wl_2 vdd gnd cell_6t
Xbit_r3_c47 bl_47 br_47 wl_3 vdd gnd cell_6t
Xbit_r4_c47 bl_47 br_47 wl_4 vdd gnd cell_6t
Xbit_r5_c47 bl_47 br_47 wl_5 vdd gnd cell_6t
Xbit_r6_c47 bl_47 br_47 wl_6 vdd gnd cell_6t
Xbit_r7_c47 bl_47 br_47 wl_7 vdd gnd cell_6t
Xbit_r8_c47 bl_47 br_47 wl_8 vdd gnd cell_6t
Xbit_r9_c47 bl_47 br_47 wl_9 vdd gnd cell_6t
Xbit_r10_c47 bl_47 br_47 wl_10 vdd gnd cell_6t
Xbit_r11_c47 bl_47 br_47 wl_11 vdd gnd cell_6t
Xbit_r12_c47 bl_47 br_47 wl_12 vdd gnd cell_6t
Xbit_r13_c47 bl_47 br_47 wl_13 vdd gnd cell_6t
Xbit_r14_c47 bl_47 br_47 wl_14 vdd gnd cell_6t
Xbit_r15_c47 bl_47 br_47 wl_15 vdd gnd cell_6t
Xbit_r16_c47 bl_47 br_47 wl_16 vdd gnd cell_6t
Xbit_r17_c47 bl_47 br_47 wl_17 vdd gnd cell_6t
Xbit_r18_c47 bl_47 br_47 wl_18 vdd gnd cell_6t
Xbit_r19_c47 bl_47 br_47 wl_19 vdd gnd cell_6t
Xbit_r20_c47 bl_47 br_47 wl_20 vdd gnd cell_6t
Xbit_r21_c47 bl_47 br_47 wl_21 vdd gnd cell_6t
Xbit_r22_c47 bl_47 br_47 wl_22 vdd gnd cell_6t
Xbit_r23_c47 bl_47 br_47 wl_23 vdd gnd cell_6t
Xbit_r24_c47 bl_47 br_47 wl_24 vdd gnd cell_6t
Xbit_r25_c47 bl_47 br_47 wl_25 vdd gnd cell_6t
Xbit_r26_c47 bl_47 br_47 wl_26 vdd gnd cell_6t
Xbit_r27_c47 bl_47 br_47 wl_27 vdd gnd cell_6t
Xbit_r28_c47 bl_47 br_47 wl_28 vdd gnd cell_6t
Xbit_r29_c47 bl_47 br_47 wl_29 vdd gnd cell_6t
Xbit_r30_c47 bl_47 br_47 wl_30 vdd gnd cell_6t
Xbit_r31_c47 bl_47 br_47 wl_31 vdd gnd cell_6t
Xbit_r32_c47 bl_47 br_47 wl_32 vdd gnd cell_6t
Xbit_r33_c47 bl_47 br_47 wl_33 vdd gnd cell_6t
Xbit_r34_c47 bl_47 br_47 wl_34 vdd gnd cell_6t
Xbit_r35_c47 bl_47 br_47 wl_35 vdd gnd cell_6t
Xbit_r36_c47 bl_47 br_47 wl_36 vdd gnd cell_6t
Xbit_r37_c47 bl_47 br_47 wl_37 vdd gnd cell_6t
Xbit_r38_c47 bl_47 br_47 wl_38 vdd gnd cell_6t
Xbit_r39_c47 bl_47 br_47 wl_39 vdd gnd cell_6t
Xbit_r40_c47 bl_47 br_47 wl_40 vdd gnd cell_6t
Xbit_r41_c47 bl_47 br_47 wl_41 vdd gnd cell_6t
Xbit_r42_c47 bl_47 br_47 wl_42 vdd gnd cell_6t
Xbit_r43_c47 bl_47 br_47 wl_43 vdd gnd cell_6t
Xbit_r44_c47 bl_47 br_47 wl_44 vdd gnd cell_6t
Xbit_r45_c47 bl_47 br_47 wl_45 vdd gnd cell_6t
Xbit_r46_c47 bl_47 br_47 wl_46 vdd gnd cell_6t
Xbit_r47_c47 bl_47 br_47 wl_47 vdd gnd cell_6t
Xbit_r48_c47 bl_47 br_47 wl_48 vdd gnd cell_6t
Xbit_r49_c47 bl_47 br_47 wl_49 vdd gnd cell_6t
Xbit_r50_c47 bl_47 br_47 wl_50 vdd gnd cell_6t
Xbit_r51_c47 bl_47 br_47 wl_51 vdd gnd cell_6t
Xbit_r52_c47 bl_47 br_47 wl_52 vdd gnd cell_6t
Xbit_r53_c47 bl_47 br_47 wl_53 vdd gnd cell_6t
Xbit_r54_c47 bl_47 br_47 wl_54 vdd gnd cell_6t
Xbit_r55_c47 bl_47 br_47 wl_55 vdd gnd cell_6t
Xbit_r56_c47 bl_47 br_47 wl_56 vdd gnd cell_6t
Xbit_r57_c47 bl_47 br_47 wl_57 vdd gnd cell_6t
Xbit_r58_c47 bl_47 br_47 wl_58 vdd gnd cell_6t
Xbit_r59_c47 bl_47 br_47 wl_59 vdd gnd cell_6t
Xbit_r60_c47 bl_47 br_47 wl_60 vdd gnd cell_6t
Xbit_r61_c47 bl_47 br_47 wl_61 vdd gnd cell_6t
Xbit_r62_c47 bl_47 br_47 wl_62 vdd gnd cell_6t
Xbit_r63_c47 bl_47 br_47 wl_63 vdd gnd cell_6t
Xbit_r64_c47 bl_47 br_47 wl_64 vdd gnd cell_6t
Xbit_r65_c47 bl_47 br_47 wl_65 vdd gnd cell_6t
Xbit_r66_c47 bl_47 br_47 wl_66 vdd gnd cell_6t
Xbit_r67_c47 bl_47 br_47 wl_67 vdd gnd cell_6t
Xbit_r68_c47 bl_47 br_47 wl_68 vdd gnd cell_6t
Xbit_r69_c47 bl_47 br_47 wl_69 vdd gnd cell_6t
Xbit_r70_c47 bl_47 br_47 wl_70 vdd gnd cell_6t
Xbit_r71_c47 bl_47 br_47 wl_71 vdd gnd cell_6t
Xbit_r72_c47 bl_47 br_47 wl_72 vdd gnd cell_6t
Xbit_r73_c47 bl_47 br_47 wl_73 vdd gnd cell_6t
Xbit_r74_c47 bl_47 br_47 wl_74 vdd gnd cell_6t
Xbit_r75_c47 bl_47 br_47 wl_75 vdd gnd cell_6t
Xbit_r76_c47 bl_47 br_47 wl_76 vdd gnd cell_6t
Xbit_r77_c47 bl_47 br_47 wl_77 vdd gnd cell_6t
Xbit_r78_c47 bl_47 br_47 wl_78 vdd gnd cell_6t
Xbit_r79_c47 bl_47 br_47 wl_79 vdd gnd cell_6t
Xbit_r80_c47 bl_47 br_47 wl_80 vdd gnd cell_6t
Xbit_r81_c47 bl_47 br_47 wl_81 vdd gnd cell_6t
Xbit_r82_c47 bl_47 br_47 wl_82 vdd gnd cell_6t
Xbit_r83_c47 bl_47 br_47 wl_83 vdd gnd cell_6t
Xbit_r84_c47 bl_47 br_47 wl_84 vdd gnd cell_6t
Xbit_r85_c47 bl_47 br_47 wl_85 vdd gnd cell_6t
Xbit_r86_c47 bl_47 br_47 wl_86 vdd gnd cell_6t
Xbit_r87_c47 bl_47 br_47 wl_87 vdd gnd cell_6t
Xbit_r88_c47 bl_47 br_47 wl_88 vdd gnd cell_6t
Xbit_r89_c47 bl_47 br_47 wl_89 vdd gnd cell_6t
Xbit_r90_c47 bl_47 br_47 wl_90 vdd gnd cell_6t
Xbit_r91_c47 bl_47 br_47 wl_91 vdd gnd cell_6t
Xbit_r92_c47 bl_47 br_47 wl_92 vdd gnd cell_6t
Xbit_r93_c47 bl_47 br_47 wl_93 vdd gnd cell_6t
Xbit_r94_c47 bl_47 br_47 wl_94 vdd gnd cell_6t
Xbit_r95_c47 bl_47 br_47 wl_95 vdd gnd cell_6t
Xbit_r96_c47 bl_47 br_47 wl_96 vdd gnd cell_6t
Xbit_r97_c47 bl_47 br_47 wl_97 vdd gnd cell_6t
Xbit_r98_c47 bl_47 br_47 wl_98 vdd gnd cell_6t
Xbit_r99_c47 bl_47 br_47 wl_99 vdd gnd cell_6t
Xbit_r100_c47 bl_47 br_47 wl_100 vdd gnd cell_6t
Xbit_r101_c47 bl_47 br_47 wl_101 vdd gnd cell_6t
Xbit_r102_c47 bl_47 br_47 wl_102 vdd gnd cell_6t
Xbit_r103_c47 bl_47 br_47 wl_103 vdd gnd cell_6t
Xbit_r104_c47 bl_47 br_47 wl_104 vdd gnd cell_6t
Xbit_r105_c47 bl_47 br_47 wl_105 vdd gnd cell_6t
Xbit_r106_c47 bl_47 br_47 wl_106 vdd gnd cell_6t
Xbit_r107_c47 bl_47 br_47 wl_107 vdd gnd cell_6t
Xbit_r108_c47 bl_47 br_47 wl_108 vdd gnd cell_6t
Xbit_r109_c47 bl_47 br_47 wl_109 vdd gnd cell_6t
Xbit_r110_c47 bl_47 br_47 wl_110 vdd gnd cell_6t
Xbit_r111_c47 bl_47 br_47 wl_111 vdd gnd cell_6t
Xbit_r112_c47 bl_47 br_47 wl_112 vdd gnd cell_6t
Xbit_r113_c47 bl_47 br_47 wl_113 vdd gnd cell_6t
Xbit_r114_c47 bl_47 br_47 wl_114 vdd gnd cell_6t
Xbit_r115_c47 bl_47 br_47 wl_115 vdd gnd cell_6t
Xbit_r116_c47 bl_47 br_47 wl_116 vdd gnd cell_6t
Xbit_r117_c47 bl_47 br_47 wl_117 vdd gnd cell_6t
Xbit_r118_c47 bl_47 br_47 wl_118 vdd gnd cell_6t
Xbit_r119_c47 bl_47 br_47 wl_119 vdd gnd cell_6t
Xbit_r120_c47 bl_47 br_47 wl_120 vdd gnd cell_6t
Xbit_r121_c47 bl_47 br_47 wl_121 vdd gnd cell_6t
Xbit_r122_c47 bl_47 br_47 wl_122 vdd gnd cell_6t
Xbit_r123_c47 bl_47 br_47 wl_123 vdd gnd cell_6t
Xbit_r124_c47 bl_47 br_47 wl_124 vdd gnd cell_6t
Xbit_r125_c47 bl_47 br_47 wl_125 vdd gnd cell_6t
Xbit_r126_c47 bl_47 br_47 wl_126 vdd gnd cell_6t
Xbit_r127_c47 bl_47 br_47 wl_127 vdd gnd cell_6t
Xbit_r128_c47 bl_47 br_47 wl_128 vdd gnd cell_6t
Xbit_r129_c47 bl_47 br_47 wl_129 vdd gnd cell_6t
Xbit_r130_c47 bl_47 br_47 wl_130 vdd gnd cell_6t
Xbit_r131_c47 bl_47 br_47 wl_131 vdd gnd cell_6t
Xbit_r132_c47 bl_47 br_47 wl_132 vdd gnd cell_6t
Xbit_r133_c47 bl_47 br_47 wl_133 vdd gnd cell_6t
Xbit_r134_c47 bl_47 br_47 wl_134 vdd gnd cell_6t
Xbit_r135_c47 bl_47 br_47 wl_135 vdd gnd cell_6t
Xbit_r136_c47 bl_47 br_47 wl_136 vdd gnd cell_6t
Xbit_r137_c47 bl_47 br_47 wl_137 vdd gnd cell_6t
Xbit_r138_c47 bl_47 br_47 wl_138 vdd gnd cell_6t
Xbit_r139_c47 bl_47 br_47 wl_139 vdd gnd cell_6t
Xbit_r140_c47 bl_47 br_47 wl_140 vdd gnd cell_6t
Xbit_r141_c47 bl_47 br_47 wl_141 vdd gnd cell_6t
Xbit_r142_c47 bl_47 br_47 wl_142 vdd gnd cell_6t
Xbit_r143_c47 bl_47 br_47 wl_143 vdd gnd cell_6t
Xbit_r144_c47 bl_47 br_47 wl_144 vdd gnd cell_6t
Xbit_r145_c47 bl_47 br_47 wl_145 vdd gnd cell_6t
Xbit_r146_c47 bl_47 br_47 wl_146 vdd gnd cell_6t
Xbit_r147_c47 bl_47 br_47 wl_147 vdd gnd cell_6t
Xbit_r148_c47 bl_47 br_47 wl_148 vdd gnd cell_6t
Xbit_r149_c47 bl_47 br_47 wl_149 vdd gnd cell_6t
Xbit_r150_c47 bl_47 br_47 wl_150 vdd gnd cell_6t
Xbit_r151_c47 bl_47 br_47 wl_151 vdd gnd cell_6t
Xbit_r152_c47 bl_47 br_47 wl_152 vdd gnd cell_6t
Xbit_r153_c47 bl_47 br_47 wl_153 vdd gnd cell_6t
Xbit_r154_c47 bl_47 br_47 wl_154 vdd gnd cell_6t
Xbit_r155_c47 bl_47 br_47 wl_155 vdd gnd cell_6t
Xbit_r156_c47 bl_47 br_47 wl_156 vdd gnd cell_6t
Xbit_r157_c47 bl_47 br_47 wl_157 vdd gnd cell_6t
Xbit_r158_c47 bl_47 br_47 wl_158 vdd gnd cell_6t
Xbit_r159_c47 bl_47 br_47 wl_159 vdd gnd cell_6t
Xbit_r160_c47 bl_47 br_47 wl_160 vdd gnd cell_6t
Xbit_r161_c47 bl_47 br_47 wl_161 vdd gnd cell_6t
Xbit_r162_c47 bl_47 br_47 wl_162 vdd gnd cell_6t
Xbit_r163_c47 bl_47 br_47 wl_163 vdd gnd cell_6t
Xbit_r164_c47 bl_47 br_47 wl_164 vdd gnd cell_6t
Xbit_r165_c47 bl_47 br_47 wl_165 vdd gnd cell_6t
Xbit_r166_c47 bl_47 br_47 wl_166 vdd gnd cell_6t
Xbit_r167_c47 bl_47 br_47 wl_167 vdd gnd cell_6t
Xbit_r168_c47 bl_47 br_47 wl_168 vdd gnd cell_6t
Xbit_r169_c47 bl_47 br_47 wl_169 vdd gnd cell_6t
Xbit_r170_c47 bl_47 br_47 wl_170 vdd gnd cell_6t
Xbit_r171_c47 bl_47 br_47 wl_171 vdd gnd cell_6t
Xbit_r172_c47 bl_47 br_47 wl_172 vdd gnd cell_6t
Xbit_r173_c47 bl_47 br_47 wl_173 vdd gnd cell_6t
Xbit_r174_c47 bl_47 br_47 wl_174 vdd gnd cell_6t
Xbit_r175_c47 bl_47 br_47 wl_175 vdd gnd cell_6t
Xbit_r176_c47 bl_47 br_47 wl_176 vdd gnd cell_6t
Xbit_r177_c47 bl_47 br_47 wl_177 vdd gnd cell_6t
Xbit_r178_c47 bl_47 br_47 wl_178 vdd gnd cell_6t
Xbit_r179_c47 bl_47 br_47 wl_179 vdd gnd cell_6t
Xbit_r180_c47 bl_47 br_47 wl_180 vdd gnd cell_6t
Xbit_r181_c47 bl_47 br_47 wl_181 vdd gnd cell_6t
Xbit_r182_c47 bl_47 br_47 wl_182 vdd gnd cell_6t
Xbit_r183_c47 bl_47 br_47 wl_183 vdd gnd cell_6t
Xbit_r184_c47 bl_47 br_47 wl_184 vdd gnd cell_6t
Xbit_r185_c47 bl_47 br_47 wl_185 vdd gnd cell_6t
Xbit_r186_c47 bl_47 br_47 wl_186 vdd gnd cell_6t
Xbit_r187_c47 bl_47 br_47 wl_187 vdd gnd cell_6t
Xbit_r188_c47 bl_47 br_47 wl_188 vdd gnd cell_6t
Xbit_r189_c47 bl_47 br_47 wl_189 vdd gnd cell_6t
Xbit_r190_c47 bl_47 br_47 wl_190 vdd gnd cell_6t
Xbit_r191_c47 bl_47 br_47 wl_191 vdd gnd cell_6t
Xbit_r192_c47 bl_47 br_47 wl_192 vdd gnd cell_6t
Xbit_r193_c47 bl_47 br_47 wl_193 vdd gnd cell_6t
Xbit_r194_c47 bl_47 br_47 wl_194 vdd gnd cell_6t
Xbit_r195_c47 bl_47 br_47 wl_195 vdd gnd cell_6t
Xbit_r196_c47 bl_47 br_47 wl_196 vdd gnd cell_6t
Xbit_r197_c47 bl_47 br_47 wl_197 vdd gnd cell_6t
Xbit_r198_c47 bl_47 br_47 wl_198 vdd gnd cell_6t
Xbit_r199_c47 bl_47 br_47 wl_199 vdd gnd cell_6t
Xbit_r200_c47 bl_47 br_47 wl_200 vdd gnd cell_6t
Xbit_r201_c47 bl_47 br_47 wl_201 vdd gnd cell_6t
Xbit_r202_c47 bl_47 br_47 wl_202 vdd gnd cell_6t
Xbit_r203_c47 bl_47 br_47 wl_203 vdd gnd cell_6t
Xbit_r204_c47 bl_47 br_47 wl_204 vdd gnd cell_6t
Xbit_r205_c47 bl_47 br_47 wl_205 vdd gnd cell_6t
Xbit_r206_c47 bl_47 br_47 wl_206 vdd gnd cell_6t
Xbit_r207_c47 bl_47 br_47 wl_207 vdd gnd cell_6t
Xbit_r208_c47 bl_47 br_47 wl_208 vdd gnd cell_6t
Xbit_r209_c47 bl_47 br_47 wl_209 vdd gnd cell_6t
Xbit_r210_c47 bl_47 br_47 wl_210 vdd gnd cell_6t
Xbit_r211_c47 bl_47 br_47 wl_211 vdd gnd cell_6t
Xbit_r212_c47 bl_47 br_47 wl_212 vdd gnd cell_6t
Xbit_r213_c47 bl_47 br_47 wl_213 vdd gnd cell_6t
Xbit_r214_c47 bl_47 br_47 wl_214 vdd gnd cell_6t
Xbit_r215_c47 bl_47 br_47 wl_215 vdd gnd cell_6t
Xbit_r216_c47 bl_47 br_47 wl_216 vdd gnd cell_6t
Xbit_r217_c47 bl_47 br_47 wl_217 vdd gnd cell_6t
Xbit_r218_c47 bl_47 br_47 wl_218 vdd gnd cell_6t
Xbit_r219_c47 bl_47 br_47 wl_219 vdd gnd cell_6t
Xbit_r220_c47 bl_47 br_47 wl_220 vdd gnd cell_6t
Xbit_r221_c47 bl_47 br_47 wl_221 vdd gnd cell_6t
Xbit_r222_c47 bl_47 br_47 wl_222 vdd gnd cell_6t
Xbit_r223_c47 bl_47 br_47 wl_223 vdd gnd cell_6t
Xbit_r224_c47 bl_47 br_47 wl_224 vdd gnd cell_6t
Xbit_r225_c47 bl_47 br_47 wl_225 vdd gnd cell_6t
Xbit_r226_c47 bl_47 br_47 wl_226 vdd gnd cell_6t
Xbit_r227_c47 bl_47 br_47 wl_227 vdd gnd cell_6t
Xbit_r228_c47 bl_47 br_47 wl_228 vdd gnd cell_6t
Xbit_r229_c47 bl_47 br_47 wl_229 vdd gnd cell_6t
Xbit_r230_c47 bl_47 br_47 wl_230 vdd gnd cell_6t
Xbit_r231_c47 bl_47 br_47 wl_231 vdd gnd cell_6t
Xbit_r232_c47 bl_47 br_47 wl_232 vdd gnd cell_6t
Xbit_r233_c47 bl_47 br_47 wl_233 vdd gnd cell_6t
Xbit_r234_c47 bl_47 br_47 wl_234 vdd gnd cell_6t
Xbit_r235_c47 bl_47 br_47 wl_235 vdd gnd cell_6t
Xbit_r236_c47 bl_47 br_47 wl_236 vdd gnd cell_6t
Xbit_r237_c47 bl_47 br_47 wl_237 vdd gnd cell_6t
Xbit_r238_c47 bl_47 br_47 wl_238 vdd gnd cell_6t
Xbit_r239_c47 bl_47 br_47 wl_239 vdd gnd cell_6t
Xbit_r240_c47 bl_47 br_47 wl_240 vdd gnd cell_6t
Xbit_r241_c47 bl_47 br_47 wl_241 vdd gnd cell_6t
Xbit_r242_c47 bl_47 br_47 wl_242 vdd gnd cell_6t
Xbit_r243_c47 bl_47 br_47 wl_243 vdd gnd cell_6t
Xbit_r244_c47 bl_47 br_47 wl_244 vdd gnd cell_6t
Xbit_r245_c47 bl_47 br_47 wl_245 vdd gnd cell_6t
Xbit_r246_c47 bl_47 br_47 wl_246 vdd gnd cell_6t
Xbit_r247_c47 bl_47 br_47 wl_247 vdd gnd cell_6t
Xbit_r248_c47 bl_47 br_47 wl_248 vdd gnd cell_6t
Xbit_r249_c47 bl_47 br_47 wl_249 vdd gnd cell_6t
Xbit_r250_c47 bl_47 br_47 wl_250 vdd gnd cell_6t
Xbit_r251_c47 bl_47 br_47 wl_251 vdd gnd cell_6t
Xbit_r252_c47 bl_47 br_47 wl_252 vdd gnd cell_6t
Xbit_r253_c47 bl_47 br_47 wl_253 vdd gnd cell_6t
Xbit_r254_c47 bl_47 br_47 wl_254 vdd gnd cell_6t
Xbit_r255_c47 bl_47 br_47 wl_255 vdd gnd cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd cell_6t
Xbit_r1_c48 bl_48 br_48 wl_1 vdd gnd cell_6t
Xbit_r2_c48 bl_48 br_48 wl_2 vdd gnd cell_6t
Xbit_r3_c48 bl_48 br_48 wl_3 vdd gnd cell_6t
Xbit_r4_c48 bl_48 br_48 wl_4 vdd gnd cell_6t
Xbit_r5_c48 bl_48 br_48 wl_5 vdd gnd cell_6t
Xbit_r6_c48 bl_48 br_48 wl_6 vdd gnd cell_6t
Xbit_r7_c48 bl_48 br_48 wl_7 vdd gnd cell_6t
Xbit_r8_c48 bl_48 br_48 wl_8 vdd gnd cell_6t
Xbit_r9_c48 bl_48 br_48 wl_9 vdd gnd cell_6t
Xbit_r10_c48 bl_48 br_48 wl_10 vdd gnd cell_6t
Xbit_r11_c48 bl_48 br_48 wl_11 vdd gnd cell_6t
Xbit_r12_c48 bl_48 br_48 wl_12 vdd gnd cell_6t
Xbit_r13_c48 bl_48 br_48 wl_13 vdd gnd cell_6t
Xbit_r14_c48 bl_48 br_48 wl_14 vdd gnd cell_6t
Xbit_r15_c48 bl_48 br_48 wl_15 vdd gnd cell_6t
Xbit_r16_c48 bl_48 br_48 wl_16 vdd gnd cell_6t
Xbit_r17_c48 bl_48 br_48 wl_17 vdd gnd cell_6t
Xbit_r18_c48 bl_48 br_48 wl_18 vdd gnd cell_6t
Xbit_r19_c48 bl_48 br_48 wl_19 vdd gnd cell_6t
Xbit_r20_c48 bl_48 br_48 wl_20 vdd gnd cell_6t
Xbit_r21_c48 bl_48 br_48 wl_21 vdd gnd cell_6t
Xbit_r22_c48 bl_48 br_48 wl_22 vdd gnd cell_6t
Xbit_r23_c48 bl_48 br_48 wl_23 vdd gnd cell_6t
Xbit_r24_c48 bl_48 br_48 wl_24 vdd gnd cell_6t
Xbit_r25_c48 bl_48 br_48 wl_25 vdd gnd cell_6t
Xbit_r26_c48 bl_48 br_48 wl_26 vdd gnd cell_6t
Xbit_r27_c48 bl_48 br_48 wl_27 vdd gnd cell_6t
Xbit_r28_c48 bl_48 br_48 wl_28 vdd gnd cell_6t
Xbit_r29_c48 bl_48 br_48 wl_29 vdd gnd cell_6t
Xbit_r30_c48 bl_48 br_48 wl_30 vdd gnd cell_6t
Xbit_r31_c48 bl_48 br_48 wl_31 vdd gnd cell_6t
Xbit_r32_c48 bl_48 br_48 wl_32 vdd gnd cell_6t
Xbit_r33_c48 bl_48 br_48 wl_33 vdd gnd cell_6t
Xbit_r34_c48 bl_48 br_48 wl_34 vdd gnd cell_6t
Xbit_r35_c48 bl_48 br_48 wl_35 vdd gnd cell_6t
Xbit_r36_c48 bl_48 br_48 wl_36 vdd gnd cell_6t
Xbit_r37_c48 bl_48 br_48 wl_37 vdd gnd cell_6t
Xbit_r38_c48 bl_48 br_48 wl_38 vdd gnd cell_6t
Xbit_r39_c48 bl_48 br_48 wl_39 vdd gnd cell_6t
Xbit_r40_c48 bl_48 br_48 wl_40 vdd gnd cell_6t
Xbit_r41_c48 bl_48 br_48 wl_41 vdd gnd cell_6t
Xbit_r42_c48 bl_48 br_48 wl_42 vdd gnd cell_6t
Xbit_r43_c48 bl_48 br_48 wl_43 vdd gnd cell_6t
Xbit_r44_c48 bl_48 br_48 wl_44 vdd gnd cell_6t
Xbit_r45_c48 bl_48 br_48 wl_45 vdd gnd cell_6t
Xbit_r46_c48 bl_48 br_48 wl_46 vdd gnd cell_6t
Xbit_r47_c48 bl_48 br_48 wl_47 vdd gnd cell_6t
Xbit_r48_c48 bl_48 br_48 wl_48 vdd gnd cell_6t
Xbit_r49_c48 bl_48 br_48 wl_49 vdd gnd cell_6t
Xbit_r50_c48 bl_48 br_48 wl_50 vdd gnd cell_6t
Xbit_r51_c48 bl_48 br_48 wl_51 vdd gnd cell_6t
Xbit_r52_c48 bl_48 br_48 wl_52 vdd gnd cell_6t
Xbit_r53_c48 bl_48 br_48 wl_53 vdd gnd cell_6t
Xbit_r54_c48 bl_48 br_48 wl_54 vdd gnd cell_6t
Xbit_r55_c48 bl_48 br_48 wl_55 vdd gnd cell_6t
Xbit_r56_c48 bl_48 br_48 wl_56 vdd gnd cell_6t
Xbit_r57_c48 bl_48 br_48 wl_57 vdd gnd cell_6t
Xbit_r58_c48 bl_48 br_48 wl_58 vdd gnd cell_6t
Xbit_r59_c48 bl_48 br_48 wl_59 vdd gnd cell_6t
Xbit_r60_c48 bl_48 br_48 wl_60 vdd gnd cell_6t
Xbit_r61_c48 bl_48 br_48 wl_61 vdd gnd cell_6t
Xbit_r62_c48 bl_48 br_48 wl_62 vdd gnd cell_6t
Xbit_r63_c48 bl_48 br_48 wl_63 vdd gnd cell_6t
Xbit_r64_c48 bl_48 br_48 wl_64 vdd gnd cell_6t
Xbit_r65_c48 bl_48 br_48 wl_65 vdd gnd cell_6t
Xbit_r66_c48 bl_48 br_48 wl_66 vdd gnd cell_6t
Xbit_r67_c48 bl_48 br_48 wl_67 vdd gnd cell_6t
Xbit_r68_c48 bl_48 br_48 wl_68 vdd gnd cell_6t
Xbit_r69_c48 bl_48 br_48 wl_69 vdd gnd cell_6t
Xbit_r70_c48 bl_48 br_48 wl_70 vdd gnd cell_6t
Xbit_r71_c48 bl_48 br_48 wl_71 vdd gnd cell_6t
Xbit_r72_c48 bl_48 br_48 wl_72 vdd gnd cell_6t
Xbit_r73_c48 bl_48 br_48 wl_73 vdd gnd cell_6t
Xbit_r74_c48 bl_48 br_48 wl_74 vdd gnd cell_6t
Xbit_r75_c48 bl_48 br_48 wl_75 vdd gnd cell_6t
Xbit_r76_c48 bl_48 br_48 wl_76 vdd gnd cell_6t
Xbit_r77_c48 bl_48 br_48 wl_77 vdd gnd cell_6t
Xbit_r78_c48 bl_48 br_48 wl_78 vdd gnd cell_6t
Xbit_r79_c48 bl_48 br_48 wl_79 vdd gnd cell_6t
Xbit_r80_c48 bl_48 br_48 wl_80 vdd gnd cell_6t
Xbit_r81_c48 bl_48 br_48 wl_81 vdd gnd cell_6t
Xbit_r82_c48 bl_48 br_48 wl_82 vdd gnd cell_6t
Xbit_r83_c48 bl_48 br_48 wl_83 vdd gnd cell_6t
Xbit_r84_c48 bl_48 br_48 wl_84 vdd gnd cell_6t
Xbit_r85_c48 bl_48 br_48 wl_85 vdd gnd cell_6t
Xbit_r86_c48 bl_48 br_48 wl_86 vdd gnd cell_6t
Xbit_r87_c48 bl_48 br_48 wl_87 vdd gnd cell_6t
Xbit_r88_c48 bl_48 br_48 wl_88 vdd gnd cell_6t
Xbit_r89_c48 bl_48 br_48 wl_89 vdd gnd cell_6t
Xbit_r90_c48 bl_48 br_48 wl_90 vdd gnd cell_6t
Xbit_r91_c48 bl_48 br_48 wl_91 vdd gnd cell_6t
Xbit_r92_c48 bl_48 br_48 wl_92 vdd gnd cell_6t
Xbit_r93_c48 bl_48 br_48 wl_93 vdd gnd cell_6t
Xbit_r94_c48 bl_48 br_48 wl_94 vdd gnd cell_6t
Xbit_r95_c48 bl_48 br_48 wl_95 vdd gnd cell_6t
Xbit_r96_c48 bl_48 br_48 wl_96 vdd gnd cell_6t
Xbit_r97_c48 bl_48 br_48 wl_97 vdd gnd cell_6t
Xbit_r98_c48 bl_48 br_48 wl_98 vdd gnd cell_6t
Xbit_r99_c48 bl_48 br_48 wl_99 vdd gnd cell_6t
Xbit_r100_c48 bl_48 br_48 wl_100 vdd gnd cell_6t
Xbit_r101_c48 bl_48 br_48 wl_101 vdd gnd cell_6t
Xbit_r102_c48 bl_48 br_48 wl_102 vdd gnd cell_6t
Xbit_r103_c48 bl_48 br_48 wl_103 vdd gnd cell_6t
Xbit_r104_c48 bl_48 br_48 wl_104 vdd gnd cell_6t
Xbit_r105_c48 bl_48 br_48 wl_105 vdd gnd cell_6t
Xbit_r106_c48 bl_48 br_48 wl_106 vdd gnd cell_6t
Xbit_r107_c48 bl_48 br_48 wl_107 vdd gnd cell_6t
Xbit_r108_c48 bl_48 br_48 wl_108 vdd gnd cell_6t
Xbit_r109_c48 bl_48 br_48 wl_109 vdd gnd cell_6t
Xbit_r110_c48 bl_48 br_48 wl_110 vdd gnd cell_6t
Xbit_r111_c48 bl_48 br_48 wl_111 vdd gnd cell_6t
Xbit_r112_c48 bl_48 br_48 wl_112 vdd gnd cell_6t
Xbit_r113_c48 bl_48 br_48 wl_113 vdd gnd cell_6t
Xbit_r114_c48 bl_48 br_48 wl_114 vdd gnd cell_6t
Xbit_r115_c48 bl_48 br_48 wl_115 vdd gnd cell_6t
Xbit_r116_c48 bl_48 br_48 wl_116 vdd gnd cell_6t
Xbit_r117_c48 bl_48 br_48 wl_117 vdd gnd cell_6t
Xbit_r118_c48 bl_48 br_48 wl_118 vdd gnd cell_6t
Xbit_r119_c48 bl_48 br_48 wl_119 vdd gnd cell_6t
Xbit_r120_c48 bl_48 br_48 wl_120 vdd gnd cell_6t
Xbit_r121_c48 bl_48 br_48 wl_121 vdd gnd cell_6t
Xbit_r122_c48 bl_48 br_48 wl_122 vdd gnd cell_6t
Xbit_r123_c48 bl_48 br_48 wl_123 vdd gnd cell_6t
Xbit_r124_c48 bl_48 br_48 wl_124 vdd gnd cell_6t
Xbit_r125_c48 bl_48 br_48 wl_125 vdd gnd cell_6t
Xbit_r126_c48 bl_48 br_48 wl_126 vdd gnd cell_6t
Xbit_r127_c48 bl_48 br_48 wl_127 vdd gnd cell_6t
Xbit_r128_c48 bl_48 br_48 wl_128 vdd gnd cell_6t
Xbit_r129_c48 bl_48 br_48 wl_129 vdd gnd cell_6t
Xbit_r130_c48 bl_48 br_48 wl_130 vdd gnd cell_6t
Xbit_r131_c48 bl_48 br_48 wl_131 vdd gnd cell_6t
Xbit_r132_c48 bl_48 br_48 wl_132 vdd gnd cell_6t
Xbit_r133_c48 bl_48 br_48 wl_133 vdd gnd cell_6t
Xbit_r134_c48 bl_48 br_48 wl_134 vdd gnd cell_6t
Xbit_r135_c48 bl_48 br_48 wl_135 vdd gnd cell_6t
Xbit_r136_c48 bl_48 br_48 wl_136 vdd gnd cell_6t
Xbit_r137_c48 bl_48 br_48 wl_137 vdd gnd cell_6t
Xbit_r138_c48 bl_48 br_48 wl_138 vdd gnd cell_6t
Xbit_r139_c48 bl_48 br_48 wl_139 vdd gnd cell_6t
Xbit_r140_c48 bl_48 br_48 wl_140 vdd gnd cell_6t
Xbit_r141_c48 bl_48 br_48 wl_141 vdd gnd cell_6t
Xbit_r142_c48 bl_48 br_48 wl_142 vdd gnd cell_6t
Xbit_r143_c48 bl_48 br_48 wl_143 vdd gnd cell_6t
Xbit_r144_c48 bl_48 br_48 wl_144 vdd gnd cell_6t
Xbit_r145_c48 bl_48 br_48 wl_145 vdd gnd cell_6t
Xbit_r146_c48 bl_48 br_48 wl_146 vdd gnd cell_6t
Xbit_r147_c48 bl_48 br_48 wl_147 vdd gnd cell_6t
Xbit_r148_c48 bl_48 br_48 wl_148 vdd gnd cell_6t
Xbit_r149_c48 bl_48 br_48 wl_149 vdd gnd cell_6t
Xbit_r150_c48 bl_48 br_48 wl_150 vdd gnd cell_6t
Xbit_r151_c48 bl_48 br_48 wl_151 vdd gnd cell_6t
Xbit_r152_c48 bl_48 br_48 wl_152 vdd gnd cell_6t
Xbit_r153_c48 bl_48 br_48 wl_153 vdd gnd cell_6t
Xbit_r154_c48 bl_48 br_48 wl_154 vdd gnd cell_6t
Xbit_r155_c48 bl_48 br_48 wl_155 vdd gnd cell_6t
Xbit_r156_c48 bl_48 br_48 wl_156 vdd gnd cell_6t
Xbit_r157_c48 bl_48 br_48 wl_157 vdd gnd cell_6t
Xbit_r158_c48 bl_48 br_48 wl_158 vdd gnd cell_6t
Xbit_r159_c48 bl_48 br_48 wl_159 vdd gnd cell_6t
Xbit_r160_c48 bl_48 br_48 wl_160 vdd gnd cell_6t
Xbit_r161_c48 bl_48 br_48 wl_161 vdd gnd cell_6t
Xbit_r162_c48 bl_48 br_48 wl_162 vdd gnd cell_6t
Xbit_r163_c48 bl_48 br_48 wl_163 vdd gnd cell_6t
Xbit_r164_c48 bl_48 br_48 wl_164 vdd gnd cell_6t
Xbit_r165_c48 bl_48 br_48 wl_165 vdd gnd cell_6t
Xbit_r166_c48 bl_48 br_48 wl_166 vdd gnd cell_6t
Xbit_r167_c48 bl_48 br_48 wl_167 vdd gnd cell_6t
Xbit_r168_c48 bl_48 br_48 wl_168 vdd gnd cell_6t
Xbit_r169_c48 bl_48 br_48 wl_169 vdd gnd cell_6t
Xbit_r170_c48 bl_48 br_48 wl_170 vdd gnd cell_6t
Xbit_r171_c48 bl_48 br_48 wl_171 vdd gnd cell_6t
Xbit_r172_c48 bl_48 br_48 wl_172 vdd gnd cell_6t
Xbit_r173_c48 bl_48 br_48 wl_173 vdd gnd cell_6t
Xbit_r174_c48 bl_48 br_48 wl_174 vdd gnd cell_6t
Xbit_r175_c48 bl_48 br_48 wl_175 vdd gnd cell_6t
Xbit_r176_c48 bl_48 br_48 wl_176 vdd gnd cell_6t
Xbit_r177_c48 bl_48 br_48 wl_177 vdd gnd cell_6t
Xbit_r178_c48 bl_48 br_48 wl_178 vdd gnd cell_6t
Xbit_r179_c48 bl_48 br_48 wl_179 vdd gnd cell_6t
Xbit_r180_c48 bl_48 br_48 wl_180 vdd gnd cell_6t
Xbit_r181_c48 bl_48 br_48 wl_181 vdd gnd cell_6t
Xbit_r182_c48 bl_48 br_48 wl_182 vdd gnd cell_6t
Xbit_r183_c48 bl_48 br_48 wl_183 vdd gnd cell_6t
Xbit_r184_c48 bl_48 br_48 wl_184 vdd gnd cell_6t
Xbit_r185_c48 bl_48 br_48 wl_185 vdd gnd cell_6t
Xbit_r186_c48 bl_48 br_48 wl_186 vdd gnd cell_6t
Xbit_r187_c48 bl_48 br_48 wl_187 vdd gnd cell_6t
Xbit_r188_c48 bl_48 br_48 wl_188 vdd gnd cell_6t
Xbit_r189_c48 bl_48 br_48 wl_189 vdd gnd cell_6t
Xbit_r190_c48 bl_48 br_48 wl_190 vdd gnd cell_6t
Xbit_r191_c48 bl_48 br_48 wl_191 vdd gnd cell_6t
Xbit_r192_c48 bl_48 br_48 wl_192 vdd gnd cell_6t
Xbit_r193_c48 bl_48 br_48 wl_193 vdd gnd cell_6t
Xbit_r194_c48 bl_48 br_48 wl_194 vdd gnd cell_6t
Xbit_r195_c48 bl_48 br_48 wl_195 vdd gnd cell_6t
Xbit_r196_c48 bl_48 br_48 wl_196 vdd gnd cell_6t
Xbit_r197_c48 bl_48 br_48 wl_197 vdd gnd cell_6t
Xbit_r198_c48 bl_48 br_48 wl_198 vdd gnd cell_6t
Xbit_r199_c48 bl_48 br_48 wl_199 vdd gnd cell_6t
Xbit_r200_c48 bl_48 br_48 wl_200 vdd gnd cell_6t
Xbit_r201_c48 bl_48 br_48 wl_201 vdd gnd cell_6t
Xbit_r202_c48 bl_48 br_48 wl_202 vdd gnd cell_6t
Xbit_r203_c48 bl_48 br_48 wl_203 vdd gnd cell_6t
Xbit_r204_c48 bl_48 br_48 wl_204 vdd gnd cell_6t
Xbit_r205_c48 bl_48 br_48 wl_205 vdd gnd cell_6t
Xbit_r206_c48 bl_48 br_48 wl_206 vdd gnd cell_6t
Xbit_r207_c48 bl_48 br_48 wl_207 vdd gnd cell_6t
Xbit_r208_c48 bl_48 br_48 wl_208 vdd gnd cell_6t
Xbit_r209_c48 bl_48 br_48 wl_209 vdd gnd cell_6t
Xbit_r210_c48 bl_48 br_48 wl_210 vdd gnd cell_6t
Xbit_r211_c48 bl_48 br_48 wl_211 vdd gnd cell_6t
Xbit_r212_c48 bl_48 br_48 wl_212 vdd gnd cell_6t
Xbit_r213_c48 bl_48 br_48 wl_213 vdd gnd cell_6t
Xbit_r214_c48 bl_48 br_48 wl_214 vdd gnd cell_6t
Xbit_r215_c48 bl_48 br_48 wl_215 vdd gnd cell_6t
Xbit_r216_c48 bl_48 br_48 wl_216 vdd gnd cell_6t
Xbit_r217_c48 bl_48 br_48 wl_217 vdd gnd cell_6t
Xbit_r218_c48 bl_48 br_48 wl_218 vdd gnd cell_6t
Xbit_r219_c48 bl_48 br_48 wl_219 vdd gnd cell_6t
Xbit_r220_c48 bl_48 br_48 wl_220 vdd gnd cell_6t
Xbit_r221_c48 bl_48 br_48 wl_221 vdd gnd cell_6t
Xbit_r222_c48 bl_48 br_48 wl_222 vdd gnd cell_6t
Xbit_r223_c48 bl_48 br_48 wl_223 vdd gnd cell_6t
Xbit_r224_c48 bl_48 br_48 wl_224 vdd gnd cell_6t
Xbit_r225_c48 bl_48 br_48 wl_225 vdd gnd cell_6t
Xbit_r226_c48 bl_48 br_48 wl_226 vdd gnd cell_6t
Xbit_r227_c48 bl_48 br_48 wl_227 vdd gnd cell_6t
Xbit_r228_c48 bl_48 br_48 wl_228 vdd gnd cell_6t
Xbit_r229_c48 bl_48 br_48 wl_229 vdd gnd cell_6t
Xbit_r230_c48 bl_48 br_48 wl_230 vdd gnd cell_6t
Xbit_r231_c48 bl_48 br_48 wl_231 vdd gnd cell_6t
Xbit_r232_c48 bl_48 br_48 wl_232 vdd gnd cell_6t
Xbit_r233_c48 bl_48 br_48 wl_233 vdd gnd cell_6t
Xbit_r234_c48 bl_48 br_48 wl_234 vdd gnd cell_6t
Xbit_r235_c48 bl_48 br_48 wl_235 vdd gnd cell_6t
Xbit_r236_c48 bl_48 br_48 wl_236 vdd gnd cell_6t
Xbit_r237_c48 bl_48 br_48 wl_237 vdd gnd cell_6t
Xbit_r238_c48 bl_48 br_48 wl_238 vdd gnd cell_6t
Xbit_r239_c48 bl_48 br_48 wl_239 vdd gnd cell_6t
Xbit_r240_c48 bl_48 br_48 wl_240 vdd gnd cell_6t
Xbit_r241_c48 bl_48 br_48 wl_241 vdd gnd cell_6t
Xbit_r242_c48 bl_48 br_48 wl_242 vdd gnd cell_6t
Xbit_r243_c48 bl_48 br_48 wl_243 vdd gnd cell_6t
Xbit_r244_c48 bl_48 br_48 wl_244 vdd gnd cell_6t
Xbit_r245_c48 bl_48 br_48 wl_245 vdd gnd cell_6t
Xbit_r246_c48 bl_48 br_48 wl_246 vdd gnd cell_6t
Xbit_r247_c48 bl_48 br_48 wl_247 vdd gnd cell_6t
Xbit_r248_c48 bl_48 br_48 wl_248 vdd gnd cell_6t
Xbit_r249_c48 bl_48 br_48 wl_249 vdd gnd cell_6t
Xbit_r250_c48 bl_48 br_48 wl_250 vdd gnd cell_6t
Xbit_r251_c48 bl_48 br_48 wl_251 vdd gnd cell_6t
Xbit_r252_c48 bl_48 br_48 wl_252 vdd gnd cell_6t
Xbit_r253_c48 bl_48 br_48 wl_253 vdd gnd cell_6t
Xbit_r254_c48 bl_48 br_48 wl_254 vdd gnd cell_6t
Xbit_r255_c48 bl_48 br_48 wl_255 vdd gnd cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd cell_6t
Xbit_r1_c49 bl_49 br_49 wl_1 vdd gnd cell_6t
Xbit_r2_c49 bl_49 br_49 wl_2 vdd gnd cell_6t
Xbit_r3_c49 bl_49 br_49 wl_3 vdd gnd cell_6t
Xbit_r4_c49 bl_49 br_49 wl_4 vdd gnd cell_6t
Xbit_r5_c49 bl_49 br_49 wl_5 vdd gnd cell_6t
Xbit_r6_c49 bl_49 br_49 wl_6 vdd gnd cell_6t
Xbit_r7_c49 bl_49 br_49 wl_7 vdd gnd cell_6t
Xbit_r8_c49 bl_49 br_49 wl_8 vdd gnd cell_6t
Xbit_r9_c49 bl_49 br_49 wl_9 vdd gnd cell_6t
Xbit_r10_c49 bl_49 br_49 wl_10 vdd gnd cell_6t
Xbit_r11_c49 bl_49 br_49 wl_11 vdd gnd cell_6t
Xbit_r12_c49 bl_49 br_49 wl_12 vdd gnd cell_6t
Xbit_r13_c49 bl_49 br_49 wl_13 vdd gnd cell_6t
Xbit_r14_c49 bl_49 br_49 wl_14 vdd gnd cell_6t
Xbit_r15_c49 bl_49 br_49 wl_15 vdd gnd cell_6t
Xbit_r16_c49 bl_49 br_49 wl_16 vdd gnd cell_6t
Xbit_r17_c49 bl_49 br_49 wl_17 vdd gnd cell_6t
Xbit_r18_c49 bl_49 br_49 wl_18 vdd gnd cell_6t
Xbit_r19_c49 bl_49 br_49 wl_19 vdd gnd cell_6t
Xbit_r20_c49 bl_49 br_49 wl_20 vdd gnd cell_6t
Xbit_r21_c49 bl_49 br_49 wl_21 vdd gnd cell_6t
Xbit_r22_c49 bl_49 br_49 wl_22 vdd gnd cell_6t
Xbit_r23_c49 bl_49 br_49 wl_23 vdd gnd cell_6t
Xbit_r24_c49 bl_49 br_49 wl_24 vdd gnd cell_6t
Xbit_r25_c49 bl_49 br_49 wl_25 vdd gnd cell_6t
Xbit_r26_c49 bl_49 br_49 wl_26 vdd gnd cell_6t
Xbit_r27_c49 bl_49 br_49 wl_27 vdd gnd cell_6t
Xbit_r28_c49 bl_49 br_49 wl_28 vdd gnd cell_6t
Xbit_r29_c49 bl_49 br_49 wl_29 vdd gnd cell_6t
Xbit_r30_c49 bl_49 br_49 wl_30 vdd gnd cell_6t
Xbit_r31_c49 bl_49 br_49 wl_31 vdd gnd cell_6t
Xbit_r32_c49 bl_49 br_49 wl_32 vdd gnd cell_6t
Xbit_r33_c49 bl_49 br_49 wl_33 vdd gnd cell_6t
Xbit_r34_c49 bl_49 br_49 wl_34 vdd gnd cell_6t
Xbit_r35_c49 bl_49 br_49 wl_35 vdd gnd cell_6t
Xbit_r36_c49 bl_49 br_49 wl_36 vdd gnd cell_6t
Xbit_r37_c49 bl_49 br_49 wl_37 vdd gnd cell_6t
Xbit_r38_c49 bl_49 br_49 wl_38 vdd gnd cell_6t
Xbit_r39_c49 bl_49 br_49 wl_39 vdd gnd cell_6t
Xbit_r40_c49 bl_49 br_49 wl_40 vdd gnd cell_6t
Xbit_r41_c49 bl_49 br_49 wl_41 vdd gnd cell_6t
Xbit_r42_c49 bl_49 br_49 wl_42 vdd gnd cell_6t
Xbit_r43_c49 bl_49 br_49 wl_43 vdd gnd cell_6t
Xbit_r44_c49 bl_49 br_49 wl_44 vdd gnd cell_6t
Xbit_r45_c49 bl_49 br_49 wl_45 vdd gnd cell_6t
Xbit_r46_c49 bl_49 br_49 wl_46 vdd gnd cell_6t
Xbit_r47_c49 bl_49 br_49 wl_47 vdd gnd cell_6t
Xbit_r48_c49 bl_49 br_49 wl_48 vdd gnd cell_6t
Xbit_r49_c49 bl_49 br_49 wl_49 vdd gnd cell_6t
Xbit_r50_c49 bl_49 br_49 wl_50 vdd gnd cell_6t
Xbit_r51_c49 bl_49 br_49 wl_51 vdd gnd cell_6t
Xbit_r52_c49 bl_49 br_49 wl_52 vdd gnd cell_6t
Xbit_r53_c49 bl_49 br_49 wl_53 vdd gnd cell_6t
Xbit_r54_c49 bl_49 br_49 wl_54 vdd gnd cell_6t
Xbit_r55_c49 bl_49 br_49 wl_55 vdd gnd cell_6t
Xbit_r56_c49 bl_49 br_49 wl_56 vdd gnd cell_6t
Xbit_r57_c49 bl_49 br_49 wl_57 vdd gnd cell_6t
Xbit_r58_c49 bl_49 br_49 wl_58 vdd gnd cell_6t
Xbit_r59_c49 bl_49 br_49 wl_59 vdd gnd cell_6t
Xbit_r60_c49 bl_49 br_49 wl_60 vdd gnd cell_6t
Xbit_r61_c49 bl_49 br_49 wl_61 vdd gnd cell_6t
Xbit_r62_c49 bl_49 br_49 wl_62 vdd gnd cell_6t
Xbit_r63_c49 bl_49 br_49 wl_63 vdd gnd cell_6t
Xbit_r64_c49 bl_49 br_49 wl_64 vdd gnd cell_6t
Xbit_r65_c49 bl_49 br_49 wl_65 vdd gnd cell_6t
Xbit_r66_c49 bl_49 br_49 wl_66 vdd gnd cell_6t
Xbit_r67_c49 bl_49 br_49 wl_67 vdd gnd cell_6t
Xbit_r68_c49 bl_49 br_49 wl_68 vdd gnd cell_6t
Xbit_r69_c49 bl_49 br_49 wl_69 vdd gnd cell_6t
Xbit_r70_c49 bl_49 br_49 wl_70 vdd gnd cell_6t
Xbit_r71_c49 bl_49 br_49 wl_71 vdd gnd cell_6t
Xbit_r72_c49 bl_49 br_49 wl_72 vdd gnd cell_6t
Xbit_r73_c49 bl_49 br_49 wl_73 vdd gnd cell_6t
Xbit_r74_c49 bl_49 br_49 wl_74 vdd gnd cell_6t
Xbit_r75_c49 bl_49 br_49 wl_75 vdd gnd cell_6t
Xbit_r76_c49 bl_49 br_49 wl_76 vdd gnd cell_6t
Xbit_r77_c49 bl_49 br_49 wl_77 vdd gnd cell_6t
Xbit_r78_c49 bl_49 br_49 wl_78 vdd gnd cell_6t
Xbit_r79_c49 bl_49 br_49 wl_79 vdd gnd cell_6t
Xbit_r80_c49 bl_49 br_49 wl_80 vdd gnd cell_6t
Xbit_r81_c49 bl_49 br_49 wl_81 vdd gnd cell_6t
Xbit_r82_c49 bl_49 br_49 wl_82 vdd gnd cell_6t
Xbit_r83_c49 bl_49 br_49 wl_83 vdd gnd cell_6t
Xbit_r84_c49 bl_49 br_49 wl_84 vdd gnd cell_6t
Xbit_r85_c49 bl_49 br_49 wl_85 vdd gnd cell_6t
Xbit_r86_c49 bl_49 br_49 wl_86 vdd gnd cell_6t
Xbit_r87_c49 bl_49 br_49 wl_87 vdd gnd cell_6t
Xbit_r88_c49 bl_49 br_49 wl_88 vdd gnd cell_6t
Xbit_r89_c49 bl_49 br_49 wl_89 vdd gnd cell_6t
Xbit_r90_c49 bl_49 br_49 wl_90 vdd gnd cell_6t
Xbit_r91_c49 bl_49 br_49 wl_91 vdd gnd cell_6t
Xbit_r92_c49 bl_49 br_49 wl_92 vdd gnd cell_6t
Xbit_r93_c49 bl_49 br_49 wl_93 vdd gnd cell_6t
Xbit_r94_c49 bl_49 br_49 wl_94 vdd gnd cell_6t
Xbit_r95_c49 bl_49 br_49 wl_95 vdd gnd cell_6t
Xbit_r96_c49 bl_49 br_49 wl_96 vdd gnd cell_6t
Xbit_r97_c49 bl_49 br_49 wl_97 vdd gnd cell_6t
Xbit_r98_c49 bl_49 br_49 wl_98 vdd gnd cell_6t
Xbit_r99_c49 bl_49 br_49 wl_99 vdd gnd cell_6t
Xbit_r100_c49 bl_49 br_49 wl_100 vdd gnd cell_6t
Xbit_r101_c49 bl_49 br_49 wl_101 vdd gnd cell_6t
Xbit_r102_c49 bl_49 br_49 wl_102 vdd gnd cell_6t
Xbit_r103_c49 bl_49 br_49 wl_103 vdd gnd cell_6t
Xbit_r104_c49 bl_49 br_49 wl_104 vdd gnd cell_6t
Xbit_r105_c49 bl_49 br_49 wl_105 vdd gnd cell_6t
Xbit_r106_c49 bl_49 br_49 wl_106 vdd gnd cell_6t
Xbit_r107_c49 bl_49 br_49 wl_107 vdd gnd cell_6t
Xbit_r108_c49 bl_49 br_49 wl_108 vdd gnd cell_6t
Xbit_r109_c49 bl_49 br_49 wl_109 vdd gnd cell_6t
Xbit_r110_c49 bl_49 br_49 wl_110 vdd gnd cell_6t
Xbit_r111_c49 bl_49 br_49 wl_111 vdd gnd cell_6t
Xbit_r112_c49 bl_49 br_49 wl_112 vdd gnd cell_6t
Xbit_r113_c49 bl_49 br_49 wl_113 vdd gnd cell_6t
Xbit_r114_c49 bl_49 br_49 wl_114 vdd gnd cell_6t
Xbit_r115_c49 bl_49 br_49 wl_115 vdd gnd cell_6t
Xbit_r116_c49 bl_49 br_49 wl_116 vdd gnd cell_6t
Xbit_r117_c49 bl_49 br_49 wl_117 vdd gnd cell_6t
Xbit_r118_c49 bl_49 br_49 wl_118 vdd gnd cell_6t
Xbit_r119_c49 bl_49 br_49 wl_119 vdd gnd cell_6t
Xbit_r120_c49 bl_49 br_49 wl_120 vdd gnd cell_6t
Xbit_r121_c49 bl_49 br_49 wl_121 vdd gnd cell_6t
Xbit_r122_c49 bl_49 br_49 wl_122 vdd gnd cell_6t
Xbit_r123_c49 bl_49 br_49 wl_123 vdd gnd cell_6t
Xbit_r124_c49 bl_49 br_49 wl_124 vdd gnd cell_6t
Xbit_r125_c49 bl_49 br_49 wl_125 vdd gnd cell_6t
Xbit_r126_c49 bl_49 br_49 wl_126 vdd gnd cell_6t
Xbit_r127_c49 bl_49 br_49 wl_127 vdd gnd cell_6t
Xbit_r128_c49 bl_49 br_49 wl_128 vdd gnd cell_6t
Xbit_r129_c49 bl_49 br_49 wl_129 vdd gnd cell_6t
Xbit_r130_c49 bl_49 br_49 wl_130 vdd gnd cell_6t
Xbit_r131_c49 bl_49 br_49 wl_131 vdd gnd cell_6t
Xbit_r132_c49 bl_49 br_49 wl_132 vdd gnd cell_6t
Xbit_r133_c49 bl_49 br_49 wl_133 vdd gnd cell_6t
Xbit_r134_c49 bl_49 br_49 wl_134 vdd gnd cell_6t
Xbit_r135_c49 bl_49 br_49 wl_135 vdd gnd cell_6t
Xbit_r136_c49 bl_49 br_49 wl_136 vdd gnd cell_6t
Xbit_r137_c49 bl_49 br_49 wl_137 vdd gnd cell_6t
Xbit_r138_c49 bl_49 br_49 wl_138 vdd gnd cell_6t
Xbit_r139_c49 bl_49 br_49 wl_139 vdd gnd cell_6t
Xbit_r140_c49 bl_49 br_49 wl_140 vdd gnd cell_6t
Xbit_r141_c49 bl_49 br_49 wl_141 vdd gnd cell_6t
Xbit_r142_c49 bl_49 br_49 wl_142 vdd gnd cell_6t
Xbit_r143_c49 bl_49 br_49 wl_143 vdd gnd cell_6t
Xbit_r144_c49 bl_49 br_49 wl_144 vdd gnd cell_6t
Xbit_r145_c49 bl_49 br_49 wl_145 vdd gnd cell_6t
Xbit_r146_c49 bl_49 br_49 wl_146 vdd gnd cell_6t
Xbit_r147_c49 bl_49 br_49 wl_147 vdd gnd cell_6t
Xbit_r148_c49 bl_49 br_49 wl_148 vdd gnd cell_6t
Xbit_r149_c49 bl_49 br_49 wl_149 vdd gnd cell_6t
Xbit_r150_c49 bl_49 br_49 wl_150 vdd gnd cell_6t
Xbit_r151_c49 bl_49 br_49 wl_151 vdd gnd cell_6t
Xbit_r152_c49 bl_49 br_49 wl_152 vdd gnd cell_6t
Xbit_r153_c49 bl_49 br_49 wl_153 vdd gnd cell_6t
Xbit_r154_c49 bl_49 br_49 wl_154 vdd gnd cell_6t
Xbit_r155_c49 bl_49 br_49 wl_155 vdd gnd cell_6t
Xbit_r156_c49 bl_49 br_49 wl_156 vdd gnd cell_6t
Xbit_r157_c49 bl_49 br_49 wl_157 vdd gnd cell_6t
Xbit_r158_c49 bl_49 br_49 wl_158 vdd gnd cell_6t
Xbit_r159_c49 bl_49 br_49 wl_159 vdd gnd cell_6t
Xbit_r160_c49 bl_49 br_49 wl_160 vdd gnd cell_6t
Xbit_r161_c49 bl_49 br_49 wl_161 vdd gnd cell_6t
Xbit_r162_c49 bl_49 br_49 wl_162 vdd gnd cell_6t
Xbit_r163_c49 bl_49 br_49 wl_163 vdd gnd cell_6t
Xbit_r164_c49 bl_49 br_49 wl_164 vdd gnd cell_6t
Xbit_r165_c49 bl_49 br_49 wl_165 vdd gnd cell_6t
Xbit_r166_c49 bl_49 br_49 wl_166 vdd gnd cell_6t
Xbit_r167_c49 bl_49 br_49 wl_167 vdd gnd cell_6t
Xbit_r168_c49 bl_49 br_49 wl_168 vdd gnd cell_6t
Xbit_r169_c49 bl_49 br_49 wl_169 vdd gnd cell_6t
Xbit_r170_c49 bl_49 br_49 wl_170 vdd gnd cell_6t
Xbit_r171_c49 bl_49 br_49 wl_171 vdd gnd cell_6t
Xbit_r172_c49 bl_49 br_49 wl_172 vdd gnd cell_6t
Xbit_r173_c49 bl_49 br_49 wl_173 vdd gnd cell_6t
Xbit_r174_c49 bl_49 br_49 wl_174 vdd gnd cell_6t
Xbit_r175_c49 bl_49 br_49 wl_175 vdd gnd cell_6t
Xbit_r176_c49 bl_49 br_49 wl_176 vdd gnd cell_6t
Xbit_r177_c49 bl_49 br_49 wl_177 vdd gnd cell_6t
Xbit_r178_c49 bl_49 br_49 wl_178 vdd gnd cell_6t
Xbit_r179_c49 bl_49 br_49 wl_179 vdd gnd cell_6t
Xbit_r180_c49 bl_49 br_49 wl_180 vdd gnd cell_6t
Xbit_r181_c49 bl_49 br_49 wl_181 vdd gnd cell_6t
Xbit_r182_c49 bl_49 br_49 wl_182 vdd gnd cell_6t
Xbit_r183_c49 bl_49 br_49 wl_183 vdd gnd cell_6t
Xbit_r184_c49 bl_49 br_49 wl_184 vdd gnd cell_6t
Xbit_r185_c49 bl_49 br_49 wl_185 vdd gnd cell_6t
Xbit_r186_c49 bl_49 br_49 wl_186 vdd gnd cell_6t
Xbit_r187_c49 bl_49 br_49 wl_187 vdd gnd cell_6t
Xbit_r188_c49 bl_49 br_49 wl_188 vdd gnd cell_6t
Xbit_r189_c49 bl_49 br_49 wl_189 vdd gnd cell_6t
Xbit_r190_c49 bl_49 br_49 wl_190 vdd gnd cell_6t
Xbit_r191_c49 bl_49 br_49 wl_191 vdd gnd cell_6t
Xbit_r192_c49 bl_49 br_49 wl_192 vdd gnd cell_6t
Xbit_r193_c49 bl_49 br_49 wl_193 vdd gnd cell_6t
Xbit_r194_c49 bl_49 br_49 wl_194 vdd gnd cell_6t
Xbit_r195_c49 bl_49 br_49 wl_195 vdd gnd cell_6t
Xbit_r196_c49 bl_49 br_49 wl_196 vdd gnd cell_6t
Xbit_r197_c49 bl_49 br_49 wl_197 vdd gnd cell_6t
Xbit_r198_c49 bl_49 br_49 wl_198 vdd gnd cell_6t
Xbit_r199_c49 bl_49 br_49 wl_199 vdd gnd cell_6t
Xbit_r200_c49 bl_49 br_49 wl_200 vdd gnd cell_6t
Xbit_r201_c49 bl_49 br_49 wl_201 vdd gnd cell_6t
Xbit_r202_c49 bl_49 br_49 wl_202 vdd gnd cell_6t
Xbit_r203_c49 bl_49 br_49 wl_203 vdd gnd cell_6t
Xbit_r204_c49 bl_49 br_49 wl_204 vdd gnd cell_6t
Xbit_r205_c49 bl_49 br_49 wl_205 vdd gnd cell_6t
Xbit_r206_c49 bl_49 br_49 wl_206 vdd gnd cell_6t
Xbit_r207_c49 bl_49 br_49 wl_207 vdd gnd cell_6t
Xbit_r208_c49 bl_49 br_49 wl_208 vdd gnd cell_6t
Xbit_r209_c49 bl_49 br_49 wl_209 vdd gnd cell_6t
Xbit_r210_c49 bl_49 br_49 wl_210 vdd gnd cell_6t
Xbit_r211_c49 bl_49 br_49 wl_211 vdd gnd cell_6t
Xbit_r212_c49 bl_49 br_49 wl_212 vdd gnd cell_6t
Xbit_r213_c49 bl_49 br_49 wl_213 vdd gnd cell_6t
Xbit_r214_c49 bl_49 br_49 wl_214 vdd gnd cell_6t
Xbit_r215_c49 bl_49 br_49 wl_215 vdd gnd cell_6t
Xbit_r216_c49 bl_49 br_49 wl_216 vdd gnd cell_6t
Xbit_r217_c49 bl_49 br_49 wl_217 vdd gnd cell_6t
Xbit_r218_c49 bl_49 br_49 wl_218 vdd gnd cell_6t
Xbit_r219_c49 bl_49 br_49 wl_219 vdd gnd cell_6t
Xbit_r220_c49 bl_49 br_49 wl_220 vdd gnd cell_6t
Xbit_r221_c49 bl_49 br_49 wl_221 vdd gnd cell_6t
Xbit_r222_c49 bl_49 br_49 wl_222 vdd gnd cell_6t
Xbit_r223_c49 bl_49 br_49 wl_223 vdd gnd cell_6t
Xbit_r224_c49 bl_49 br_49 wl_224 vdd gnd cell_6t
Xbit_r225_c49 bl_49 br_49 wl_225 vdd gnd cell_6t
Xbit_r226_c49 bl_49 br_49 wl_226 vdd gnd cell_6t
Xbit_r227_c49 bl_49 br_49 wl_227 vdd gnd cell_6t
Xbit_r228_c49 bl_49 br_49 wl_228 vdd gnd cell_6t
Xbit_r229_c49 bl_49 br_49 wl_229 vdd gnd cell_6t
Xbit_r230_c49 bl_49 br_49 wl_230 vdd gnd cell_6t
Xbit_r231_c49 bl_49 br_49 wl_231 vdd gnd cell_6t
Xbit_r232_c49 bl_49 br_49 wl_232 vdd gnd cell_6t
Xbit_r233_c49 bl_49 br_49 wl_233 vdd gnd cell_6t
Xbit_r234_c49 bl_49 br_49 wl_234 vdd gnd cell_6t
Xbit_r235_c49 bl_49 br_49 wl_235 vdd gnd cell_6t
Xbit_r236_c49 bl_49 br_49 wl_236 vdd gnd cell_6t
Xbit_r237_c49 bl_49 br_49 wl_237 vdd gnd cell_6t
Xbit_r238_c49 bl_49 br_49 wl_238 vdd gnd cell_6t
Xbit_r239_c49 bl_49 br_49 wl_239 vdd gnd cell_6t
Xbit_r240_c49 bl_49 br_49 wl_240 vdd gnd cell_6t
Xbit_r241_c49 bl_49 br_49 wl_241 vdd gnd cell_6t
Xbit_r242_c49 bl_49 br_49 wl_242 vdd gnd cell_6t
Xbit_r243_c49 bl_49 br_49 wl_243 vdd gnd cell_6t
Xbit_r244_c49 bl_49 br_49 wl_244 vdd gnd cell_6t
Xbit_r245_c49 bl_49 br_49 wl_245 vdd gnd cell_6t
Xbit_r246_c49 bl_49 br_49 wl_246 vdd gnd cell_6t
Xbit_r247_c49 bl_49 br_49 wl_247 vdd gnd cell_6t
Xbit_r248_c49 bl_49 br_49 wl_248 vdd gnd cell_6t
Xbit_r249_c49 bl_49 br_49 wl_249 vdd gnd cell_6t
Xbit_r250_c49 bl_49 br_49 wl_250 vdd gnd cell_6t
Xbit_r251_c49 bl_49 br_49 wl_251 vdd gnd cell_6t
Xbit_r252_c49 bl_49 br_49 wl_252 vdd gnd cell_6t
Xbit_r253_c49 bl_49 br_49 wl_253 vdd gnd cell_6t
Xbit_r254_c49 bl_49 br_49 wl_254 vdd gnd cell_6t
Xbit_r255_c49 bl_49 br_49 wl_255 vdd gnd cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd cell_6t
Xbit_r1_c50 bl_50 br_50 wl_1 vdd gnd cell_6t
Xbit_r2_c50 bl_50 br_50 wl_2 vdd gnd cell_6t
Xbit_r3_c50 bl_50 br_50 wl_3 vdd gnd cell_6t
Xbit_r4_c50 bl_50 br_50 wl_4 vdd gnd cell_6t
Xbit_r5_c50 bl_50 br_50 wl_5 vdd gnd cell_6t
Xbit_r6_c50 bl_50 br_50 wl_6 vdd gnd cell_6t
Xbit_r7_c50 bl_50 br_50 wl_7 vdd gnd cell_6t
Xbit_r8_c50 bl_50 br_50 wl_8 vdd gnd cell_6t
Xbit_r9_c50 bl_50 br_50 wl_9 vdd gnd cell_6t
Xbit_r10_c50 bl_50 br_50 wl_10 vdd gnd cell_6t
Xbit_r11_c50 bl_50 br_50 wl_11 vdd gnd cell_6t
Xbit_r12_c50 bl_50 br_50 wl_12 vdd gnd cell_6t
Xbit_r13_c50 bl_50 br_50 wl_13 vdd gnd cell_6t
Xbit_r14_c50 bl_50 br_50 wl_14 vdd gnd cell_6t
Xbit_r15_c50 bl_50 br_50 wl_15 vdd gnd cell_6t
Xbit_r16_c50 bl_50 br_50 wl_16 vdd gnd cell_6t
Xbit_r17_c50 bl_50 br_50 wl_17 vdd gnd cell_6t
Xbit_r18_c50 bl_50 br_50 wl_18 vdd gnd cell_6t
Xbit_r19_c50 bl_50 br_50 wl_19 vdd gnd cell_6t
Xbit_r20_c50 bl_50 br_50 wl_20 vdd gnd cell_6t
Xbit_r21_c50 bl_50 br_50 wl_21 vdd gnd cell_6t
Xbit_r22_c50 bl_50 br_50 wl_22 vdd gnd cell_6t
Xbit_r23_c50 bl_50 br_50 wl_23 vdd gnd cell_6t
Xbit_r24_c50 bl_50 br_50 wl_24 vdd gnd cell_6t
Xbit_r25_c50 bl_50 br_50 wl_25 vdd gnd cell_6t
Xbit_r26_c50 bl_50 br_50 wl_26 vdd gnd cell_6t
Xbit_r27_c50 bl_50 br_50 wl_27 vdd gnd cell_6t
Xbit_r28_c50 bl_50 br_50 wl_28 vdd gnd cell_6t
Xbit_r29_c50 bl_50 br_50 wl_29 vdd gnd cell_6t
Xbit_r30_c50 bl_50 br_50 wl_30 vdd gnd cell_6t
Xbit_r31_c50 bl_50 br_50 wl_31 vdd gnd cell_6t
Xbit_r32_c50 bl_50 br_50 wl_32 vdd gnd cell_6t
Xbit_r33_c50 bl_50 br_50 wl_33 vdd gnd cell_6t
Xbit_r34_c50 bl_50 br_50 wl_34 vdd gnd cell_6t
Xbit_r35_c50 bl_50 br_50 wl_35 vdd gnd cell_6t
Xbit_r36_c50 bl_50 br_50 wl_36 vdd gnd cell_6t
Xbit_r37_c50 bl_50 br_50 wl_37 vdd gnd cell_6t
Xbit_r38_c50 bl_50 br_50 wl_38 vdd gnd cell_6t
Xbit_r39_c50 bl_50 br_50 wl_39 vdd gnd cell_6t
Xbit_r40_c50 bl_50 br_50 wl_40 vdd gnd cell_6t
Xbit_r41_c50 bl_50 br_50 wl_41 vdd gnd cell_6t
Xbit_r42_c50 bl_50 br_50 wl_42 vdd gnd cell_6t
Xbit_r43_c50 bl_50 br_50 wl_43 vdd gnd cell_6t
Xbit_r44_c50 bl_50 br_50 wl_44 vdd gnd cell_6t
Xbit_r45_c50 bl_50 br_50 wl_45 vdd gnd cell_6t
Xbit_r46_c50 bl_50 br_50 wl_46 vdd gnd cell_6t
Xbit_r47_c50 bl_50 br_50 wl_47 vdd gnd cell_6t
Xbit_r48_c50 bl_50 br_50 wl_48 vdd gnd cell_6t
Xbit_r49_c50 bl_50 br_50 wl_49 vdd gnd cell_6t
Xbit_r50_c50 bl_50 br_50 wl_50 vdd gnd cell_6t
Xbit_r51_c50 bl_50 br_50 wl_51 vdd gnd cell_6t
Xbit_r52_c50 bl_50 br_50 wl_52 vdd gnd cell_6t
Xbit_r53_c50 bl_50 br_50 wl_53 vdd gnd cell_6t
Xbit_r54_c50 bl_50 br_50 wl_54 vdd gnd cell_6t
Xbit_r55_c50 bl_50 br_50 wl_55 vdd gnd cell_6t
Xbit_r56_c50 bl_50 br_50 wl_56 vdd gnd cell_6t
Xbit_r57_c50 bl_50 br_50 wl_57 vdd gnd cell_6t
Xbit_r58_c50 bl_50 br_50 wl_58 vdd gnd cell_6t
Xbit_r59_c50 bl_50 br_50 wl_59 vdd gnd cell_6t
Xbit_r60_c50 bl_50 br_50 wl_60 vdd gnd cell_6t
Xbit_r61_c50 bl_50 br_50 wl_61 vdd gnd cell_6t
Xbit_r62_c50 bl_50 br_50 wl_62 vdd gnd cell_6t
Xbit_r63_c50 bl_50 br_50 wl_63 vdd gnd cell_6t
Xbit_r64_c50 bl_50 br_50 wl_64 vdd gnd cell_6t
Xbit_r65_c50 bl_50 br_50 wl_65 vdd gnd cell_6t
Xbit_r66_c50 bl_50 br_50 wl_66 vdd gnd cell_6t
Xbit_r67_c50 bl_50 br_50 wl_67 vdd gnd cell_6t
Xbit_r68_c50 bl_50 br_50 wl_68 vdd gnd cell_6t
Xbit_r69_c50 bl_50 br_50 wl_69 vdd gnd cell_6t
Xbit_r70_c50 bl_50 br_50 wl_70 vdd gnd cell_6t
Xbit_r71_c50 bl_50 br_50 wl_71 vdd gnd cell_6t
Xbit_r72_c50 bl_50 br_50 wl_72 vdd gnd cell_6t
Xbit_r73_c50 bl_50 br_50 wl_73 vdd gnd cell_6t
Xbit_r74_c50 bl_50 br_50 wl_74 vdd gnd cell_6t
Xbit_r75_c50 bl_50 br_50 wl_75 vdd gnd cell_6t
Xbit_r76_c50 bl_50 br_50 wl_76 vdd gnd cell_6t
Xbit_r77_c50 bl_50 br_50 wl_77 vdd gnd cell_6t
Xbit_r78_c50 bl_50 br_50 wl_78 vdd gnd cell_6t
Xbit_r79_c50 bl_50 br_50 wl_79 vdd gnd cell_6t
Xbit_r80_c50 bl_50 br_50 wl_80 vdd gnd cell_6t
Xbit_r81_c50 bl_50 br_50 wl_81 vdd gnd cell_6t
Xbit_r82_c50 bl_50 br_50 wl_82 vdd gnd cell_6t
Xbit_r83_c50 bl_50 br_50 wl_83 vdd gnd cell_6t
Xbit_r84_c50 bl_50 br_50 wl_84 vdd gnd cell_6t
Xbit_r85_c50 bl_50 br_50 wl_85 vdd gnd cell_6t
Xbit_r86_c50 bl_50 br_50 wl_86 vdd gnd cell_6t
Xbit_r87_c50 bl_50 br_50 wl_87 vdd gnd cell_6t
Xbit_r88_c50 bl_50 br_50 wl_88 vdd gnd cell_6t
Xbit_r89_c50 bl_50 br_50 wl_89 vdd gnd cell_6t
Xbit_r90_c50 bl_50 br_50 wl_90 vdd gnd cell_6t
Xbit_r91_c50 bl_50 br_50 wl_91 vdd gnd cell_6t
Xbit_r92_c50 bl_50 br_50 wl_92 vdd gnd cell_6t
Xbit_r93_c50 bl_50 br_50 wl_93 vdd gnd cell_6t
Xbit_r94_c50 bl_50 br_50 wl_94 vdd gnd cell_6t
Xbit_r95_c50 bl_50 br_50 wl_95 vdd gnd cell_6t
Xbit_r96_c50 bl_50 br_50 wl_96 vdd gnd cell_6t
Xbit_r97_c50 bl_50 br_50 wl_97 vdd gnd cell_6t
Xbit_r98_c50 bl_50 br_50 wl_98 vdd gnd cell_6t
Xbit_r99_c50 bl_50 br_50 wl_99 vdd gnd cell_6t
Xbit_r100_c50 bl_50 br_50 wl_100 vdd gnd cell_6t
Xbit_r101_c50 bl_50 br_50 wl_101 vdd gnd cell_6t
Xbit_r102_c50 bl_50 br_50 wl_102 vdd gnd cell_6t
Xbit_r103_c50 bl_50 br_50 wl_103 vdd gnd cell_6t
Xbit_r104_c50 bl_50 br_50 wl_104 vdd gnd cell_6t
Xbit_r105_c50 bl_50 br_50 wl_105 vdd gnd cell_6t
Xbit_r106_c50 bl_50 br_50 wl_106 vdd gnd cell_6t
Xbit_r107_c50 bl_50 br_50 wl_107 vdd gnd cell_6t
Xbit_r108_c50 bl_50 br_50 wl_108 vdd gnd cell_6t
Xbit_r109_c50 bl_50 br_50 wl_109 vdd gnd cell_6t
Xbit_r110_c50 bl_50 br_50 wl_110 vdd gnd cell_6t
Xbit_r111_c50 bl_50 br_50 wl_111 vdd gnd cell_6t
Xbit_r112_c50 bl_50 br_50 wl_112 vdd gnd cell_6t
Xbit_r113_c50 bl_50 br_50 wl_113 vdd gnd cell_6t
Xbit_r114_c50 bl_50 br_50 wl_114 vdd gnd cell_6t
Xbit_r115_c50 bl_50 br_50 wl_115 vdd gnd cell_6t
Xbit_r116_c50 bl_50 br_50 wl_116 vdd gnd cell_6t
Xbit_r117_c50 bl_50 br_50 wl_117 vdd gnd cell_6t
Xbit_r118_c50 bl_50 br_50 wl_118 vdd gnd cell_6t
Xbit_r119_c50 bl_50 br_50 wl_119 vdd gnd cell_6t
Xbit_r120_c50 bl_50 br_50 wl_120 vdd gnd cell_6t
Xbit_r121_c50 bl_50 br_50 wl_121 vdd gnd cell_6t
Xbit_r122_c50 bl_50 br_50 wl_122 vdd gnd cell_6t
Xbit_r123_c50 bl_50 br_50 wl_123 vdd gnd cell_6t
Xbit_r124_c50 bl_50 br_50 wl_124 vdd gnd cell_6t
Xbit_r125_c50 bl_50 br_50 wl_125 vdd gnd cell_6t
Xbit_r126_c50 bl_50 br_50 wl_126 vdd gnd cell_6t
Xbit_r127_c50 bl_50 br_50 wl_127 vdd gnd cell_6t
Xbit_r128_c50 bl_50 br_50 wl_128 vdd gnd cell_6t
Xbit_r129_c50 bl_50 br_50 wl_129 vdd gnd cell_6t
Xbit_r130_c50 bl_50 br_50 wl_130 vdd gnd cell_6t
Xbit_r131_c50 bl_50 br_50 wl_131 vdd gnd cell_6t
Xbit_r132_c50 bl_50 br_50 wl_132 vdd gnd cell_6t
Xbit_r133_c50 bl_50 br_50 wl_133 vdd gnd cell_6t
Xbit_r134_c50 bl_50 br_50 wl_134 vdd gnd cell_6t
Xbit_r135_c50 bl_50 br_50 wl_135 vdd gnd cell_6t
Xbit_r136_c50 bl_50 br_50 wl_136 vdd gnd cell_6t
Xbit_r137_c50 bl_50 br_50 wl_137 vdd gnd cell_6t
Xbit_r138_c50 bl_50 br_50 wl_138 vdd gnd cell_6t
Xbit_r139_c50 bl_50 br_50 wl_139 vdd gnd cell_6t
Xbit_r140_c50 bl_50 br_50 wl_140 vdd gnd cell_6t
Xbit_r141_c50 bl_50 br_50 wl_141 vdd gnd cell_6t
Xbit_r142_c50 bl_50 br_50 wl_142 vdd gnd cell_6t
Xbit_r143_c50 bl_50 br_50 wl_143 vdd gnd cell_6t
Xbit_r144_c50 bl_50 br_50 wl_144 vdd gnd cell_6t
Xbit_r145_c50 bl_50 br_50 wl_145 vdd gnd cell_6t
Xbit_r146_c50 bl_50 br_50 wl_146 vdd gnd cell_6t
Xbit_r147_c50 bl_50 br_50 wl_147 vdd gnd cell_6t
Xbit_r148_c50 bl_50 br_50 wl_148 vdd gnd cell_6t
Xbit_r149_c50 bl_50 br_50 wl_149 vdd gnd cell_6t
Xbit_r150_c50 bl_50 br_50 wl_150 vdd gnd cell_6t
Xbit_r151_c50 bl_50 br_50 wl_151 vdd gnd cell_6t
Xbit_r152_c50 bl_50 br_50 wl_152 vdd gnd cell_6t
Xbit_r153_c50 bl_50 br_50 wl_153 vdd gnd cell_6t
Xbit_r154_c50 bl_50 br_50 wl_154 vdd gnd cell_6t
Xbit_r155_c50 bl_50 br_50 wl_155 vdd gnd cell_6t
Xbit_r156_c50 bl_50 br_50 wl_156 vdd gnd cell_6t
Xbit_r157_c50 bl_50 br_50 wl_157 vdd gnd cell_6t
Xbit_r158_c50 bl_50 br_50 wl_158 vdd gnd cell_6t
Xbit_r159_c50 bl_50 br_50 wl_159 vdd gnd cell_6t
Xbit_r160_c50 bl_50 br_50 wl_160 vdd gnd cell_6t
Xbit_r161_c50 bl_50 br_50 wl_161 vdd gnd cell_6t
Xbit_r162_c50 bl_50 br_50 wl_162 vdd gnd cell_6t
Xbit_r163_c50 bl_50 br_50 wl_163 vdd gnd cell_6t
Xbit_r164_c50 bl_50 br_50 wl_164 vdd gnd cell_6t
Xbit_r165_c50 bl_50 br_50 wl_165 vdd gnd cell_6t
Xbit_r166_c50 bl_50 br_50 wl_166 vdd gnd cell_6t
Xbit_r167_c50 bl_50 br_50 wl_167 vdd gnd cell_6t
Xbit_r168_c50 bl_50 br_50 wl_168 vdd gnd cell_6t
Xbit_r169_c50 bl_50 br_50 wl_169 vdd gnd cell_6t
Xbit_r170_c50 bl_50 br_50 wl_170 vdd gnd cell_6t
Xbit_r171_c50 bl_50 br_50 wl_171 vdd gnd cell_6t
Xbit_r172_c50 bl_50 br_50 wl_172 vdd gnd cell_6t
Xbit_r173_c50 bl_50 br_50 wl_173 vdd gnd cell_6t
Xbit_r174_c50 bl_50 br_50 wl_174 vdd gnd cell_6t
Xbit_r175_c50 bl_50 br_50 wl_175 vdd gnd cell_6t
Xbit_r176_c50 bl_50 br_50 wl_176 vdd gnd cell_6t
Xbit_r177_c50 bl_50 br_50 wl_177 vdd gnd cell_6t
Xbit_r178_c50 bl_50 br_50 wl_178 vdd gnd cell_6t
Xbit_r179_c50 bl_50 br_50 wl_179 vdd gnd cell_6t
Xbit_r180_c50 bl_50 br_50 wl_180 vdd gnd cell_6t
Xbit_r181_c50 bl_50 br_50 wl_181 vdd gnd cell_6t
Xbit_r182_c50 bl_50 br_50 wl_182 vdd gnd cell_6t
Xbit_r183_c50 bl_50 br_50 wl_183 vdd gnd cell_6t
Xbit_r184_c50 bl_50 br_50 wl_184 vdd gnd cell_6t
Xbit_r185_c50 bl_50 br_50 wl_185 vdd gnd cell_6t
Xbit_r186_c50 bl_50 br_50 wl_186 vdd gnd cell_6t
Xbit_r187_c50 bl_50 br_50 wl_187 vdd gnd cell_6t
Xbit_r188_c50 bl_50 br_50 wl_188 vdd gnd cell_6t
Xbit_r189_c50 bl_50 br_50 wl_189 vdd gnd cell_6t
Xbit_r190_c50 bl_50 br_50 wl_190 vdd gnd cell_6t
Xbit_r191_c50 bl_50 br_50 wl_191 vdd gnd cell_6t
Xbit_r192_c50 bl_50 br_50 wl_192 vdd gnd cell_6t
Xbit_r193_c50 bl_50 br_50 wl_193 vdd gnd cell_6t
Xbit_r194_c50 bl_50 br_50 wl_194 vdd gnd cell_6t
Xbit_r195_c50 bl_50 br_50 wl_195 vdd gnd cell_6t
Xbit_r196_c50 bl_50 br_50 wl_196 vdd gnd cell_6t
Xbit_r197_c50 bl_50 br_50 wl_197 vdd gnd cell_6t
Xbit_r198_c50 bl_50 br_50 wl_198 vdd gnd cell_6t
Xbit_r199_c50 bl_50 br_50 wl_199 vdd gnd cell_6t
Xbit_r200_c50 bl_50 br_50 wl_200 vdd gnd cell_6t
Xbit_r201_c50 bl_50 br_50 wl_201 vdd gnd cell_6t
Xbit_r202_c50 bl_50 br_50 wl_202 vdd gnd cell_6t
Xbit_r203_c50 bl_50 br_50 wl_203 vdd gnd cell_6t
Xbit_r204_c50 bl_50 br_50 wl_204 vdd gnd cell_6t
Xbit_r205_c50 bl_50 br_50 wl_205 vdd gnd cell_6t
Xbit_r206_c50 bl_50 br_50 wl_206 vdd gnd cell_6t
Xbit_r207_c50 bl_50 br_50 wl_207 vdd gnd cell_6t
Xbit_r208_c50 bl_50 br_50 wl_208 vdd gnd cell_6t
Xbit_r209_c50 bl_50 br_50 wl_209 vdd gnd cell_6t
Xbit_r210_c50 bl_50 br_50 wl_210 vdd gnd cell_6t
Xbit_r211_c50 bl_50 br_50 wl_211 vdd gnd cell_6t
Xbit_r212_c50 bl_50 br_50 wl_212 vdd gnd cell_6t
Xbit_r213_c50 bl_50 br_50 wl_213 vdd gnd cell_6t
Xbit_r214_c50 bl_50 br_50 wl_214 vdd gnd cell_6t
Xbit_r215_c50 bl_50 br_50 wl_215 vdd gnd cell_6t
Xbit_r216_c50 bl_50 br_50 wl_216 vdd gnd cell_6t
Xbit_r217_c50 bl_50 br_50 wl_217 vdd gnd cell_6t
Xbit_r218_c50 bl_50 br_50 wl_218 vdd gnd cell_6t
Xbit_r219_c50 bl_50 br_50 wl_219 vdd gnd cell_6t
Xbit_r220_c50 bl_50 br_50 wl_220 vdd gnd cell_6t
Xbit_r221_c50 bl_50 br_50 wl_221 vdd gnd cell_6t
Xbit_r222_c50 bl_50 br_50 wl_222 vdd gnd cell_6t
Xbit_r223_c50 bl_50 br_50 wl_223 vdd gnd cell_6t
Xbit_r224_c50 bl_50 br_50 wl_224 vdd gnd cell_6t
Xbit_r225_c50 bl_50 br_50 wl_225 vdd gnd cell_6t
Xbit_r226_c50 bl_50 br_50 wl_226 vdd gnd cell_6t
Xbit_r227_c50 bl_50 br_50 wl_227 vdd gnd cell_6t
Xbit_r228_c50 bl_50 br_50 wl_228 vdd gnd cell_6t
Xbit_r229_c50 bl_50 br_50 wl_229 vdd gnd cell_6t
Xbit_r230_c50 bl_50 br_50 wl_230 vdd gnd cell_6t
Xbit_r231_c50 bl_50 br_50 wl_231 vdd gnd cell_6t
Xbit_r232_c50 bl_50 br_50 wl_232 vdd gnd cell_6t
Xbit_r233_c50 bl_50 br_50 wl_233 vdd gnd cell_6t
Xbit_r234_c50 bl_50 br_50 wl_234 vdd gnd cell_6t
Xbit_r235_c50 bl_50 br_50 wl_235 vdd gnd cell_6t
Xbit_r236_c50 bl_50 br_50 wl_236 vdd gnd cell_6t
Xbit_r237_c50 bl_50 br_50 wl_237 vdd gnd cell_6t
Xbit_r238_c50 bl_50 br_50 wl_238 vdd gnd cell_6t
Xbit_r239_c50 bl_50 br_50 wl_239 vdd gnd cell_6t
Xbit_r240_c50 bl_50 br_50 wl_240 vdd gnd cell_6t
Xbit_r241_c50 bl_50 br_50 wl_241 vdd gnd cell_6t
Xbit_r242_c50 bl_50 br_50 wl_242 vdd gnd cell_6t
Xbit_r243_c50 bl_50 br_50 wl_243 vdd gnd cell_6t
Xbit_r244_c50 bl_50 br_50 wl_244 vdd gnd cell_6t
Xbit_r245_c50 bl_50 br_50 wl_245 vdd gnd cell_6t
Xbit_r246_c50 bl_50 br_50 wl_246 vdd gnd cell_6t
Xbit_r247_c50 bl_50 br_50 wl_247 vdd gnd cell_6t
Xbit_r248_c50 bl_50 br_50 wl_248 vdd gnd cell_6t
Xbit_r249_c50 bl_50 br_50 wl_249 vdd gnd cell_6t
Xbit_r250_c50 bl_50 br_50 wl_250 vdd gnd cell_6t
Xbit_r251_c50 bl_50 br_50 wl_251 vdd gnd cell_6t
Xbit_r252_c50 bl_50 br_50 wl_252 vdd gnd cell_6t
Xbit_r253_c50 bl_50 br_50 wl_253 vdd gnd cell_6t
Xbit_r254_c50 bl_50 br_50 wl_254 vdd gnd cell_6t
Xbit_r255_c50 bl_50 br_50 wl_255 vdd gnd cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd cell_6t
Xbit_r1_c51 bl_51 br_51 wl_1 vdd gnd cell_6t
Xbit_r2_c51 bl_51 br_51 wl_2 vdd gnd cell_6t
Xbit_r3_c51 bl_51 br_51 wl_3 vdd gnd cell_6t
Xbit_r4_c51 bl_51 br_51 wl_4 vdd gnd cell_6t
Xbit_r5_c51 bl_51 br_51 wl_5 vdd gnd cell_6t
Xbit_r6_c51 bl_51 br_51 wl_6 vdd gnd cell_6t
Xbit_r7_c51 bl_51 br_51 wl_7 vdd gnd cell_6t
Xbit_r8_c51 bl_51 br_51 wl_8 vdd gnd cell_6t
Xbit_r9_c51 bl_51 br_51 wl_9 vdd gnd cell_6t
Xbit_r10_c51 bl_51 br_51 wl_10 vdd gnd cell_6t
Xbit_r11_c51 bl_51 br_51 wl_11 vdd gnd cell_6t
Xbit_r12_c51 bl_51 br_51 wl_12 vdd gnd cell_6t
Xbit_r13_c51 bl_51 br_51 wl_13 vdd gnd cell_6t
Xbit_r14_c51 bl_51 br_51 wl_14 vdd gnd cell_6t
Xbit_r15_c51 bl_51 br_51 wl_15 vdd gnd cell_6t
Xbit_r16_c51 bl_51 br_51 wl_16 vdd gnd cell_6t
Xbit_r17_c51 bl_51 br_51 wl_17 vdd gnd cell_6t
Xbit_r18_c51 bl_51 br_51 wl_18 vdd gnd cell_6t
Xbit_r19_c51 bl_51 br_51 wl_19 vdd gnd cell_6t
Xbit_r20_c51 bl_51 br_51 wl_20 vdd gnd cell_6t
Xbit_r21_c51 bl_51 br_51 wl_21 vdd gnd cell_6t
Xbit_r22_c51 bl_51 br_51 wl_22 vdd gnd cell_6t
Xbit_r23_c51 bl_51 br_51 wl_23 vdd gnd cell_6t
Xbit_r24_c51 bl_51 br_51 wl_24 vdd gnd cell_6t
Xbit_r25_c51 bl_51 br_51 wl_25 vdd gnd cell_6t
Xbit_r26_c51 bl_51 br_51 wl_26 vdd gnd cell_6t
Xbit_r27_c51 bl_51 br_51 wl_27 vdd gnd cell_6t
Xbit_r28_c51 bl_51 br_51 wl_28 vdd gnd cell_6t
Xbit_r29_c51 bl_51 br_51 wl_29 vdd gnd cell_6t
Xbit_r30_c51 bl_51 br_51 wl_30 vdd gnd cell_6t
Xbit_r31_c51 bl_51 br_51 wl_31 vdd gnd cell_6t
Xbit_r32_c51 bl_51 br_51 wl_32 vdd gnd cell_6t
Xbit_r33_c51 bl_51 br_51 wl_33 vdd gnd cell_6t
Xbit_r34_c51 bl_51 br_51 wl_34 vdd gnd cell_6t
Xbit_r35_c51 bl_51 br_51 wl_35 vdd gnd cell_6t
Xbit_r36_c51 bl_51 br_51 wl_36 vdd gnd cell_6t
Xbit_r37_c51 bl_51 br_51 wl_37 vdd gnd cell_6t
Xbit_r38_c51 bl_51 br_51 wl_38 vdd gnd cell_6t
Xbit_r39_c51 bl_51 br_51 wl_39 vdd gnd cell_6t
Xbit_r40_c51 bl_51 br_51 wl_40 vdd gnd cell_6t
Xbit_r41_c51 bl_51 br_51 wl_41 vdd gnd cell_6t
Xbit_r42_c51 bl_51 br_51 wl_42 vdd gnd cell_6t
Xbit_r43_c51 bl_51 br_51 wl_43 vdd gnd cell_6t
Xbit_r44_c51 bl_51 br_51 wl_44 vdd gnd cell_6t
Xbit_r45_c51 bl_51 br_51 wl_45 vdd gnd cell_6t
Xbit_r46_c51 bl_51 br_51 wl_46 vdd gnd cell_6t
Xbit_r47_c51 bl_51 br_51 wl_47 vdd gnd cell_6t
Xbit_r48_c51 bl_51 br_51 wl_48 vdd gnd cell_6t
Xbit_r49_c51 bl_51 br_51 wl_49 vdd gnd cell_6t
Xbit_r50_c51 bl_51 br_51 wl_50 vdd gnd cell_6t
Xbit_r51_c51 bl_51 br_51 wl_51 vdd gnd cell_6t
Xbit_r52_c51 bl_51 br_51 wl_52 vdd gnd cell_6t
Xbit_r53_c51 bl_51 br_51 wl_53 vdd gnd cell_6t
Xbit_r54_c51 bl_51 br_51 wl_54 vdd gnd cell_6t
Xbit_r55_c51 bl_51 br_51 wl_55 vdd gnd cell_6t
Xbit_r56_c51 bl_51 br_51 wl_56 vdd gnd cell_6t
Xbit_r57_c51 bl_51 br_51 wl_57 vdd gnd cell_6t
Xbit_r58_c51 bl_51 br_51 wl_58 vdd gnd cell_6t
Xbit_r59_c51 bl_51 br_51 wl_59 vdd gnd cell_6t
Xbit_r60_c51 bl_51 br_51 wl_60 vdd gnd cell_6t
Xbit_r61_c51 bl_51 br_51 wl_61 vdd gnd cell_6t
Xbit_r62_c51 bl_51 br_51 wl_62 vdd gnd cell_6t
Xbit_r63_c51 bl_51 br_51 wl_63 vdd gnd cell_6t
Xbit_r64_c51 bl_51 br_51 wl_64 vdd gnd cell_6t
Xbit_r65_c51 bl_51 br_51 wl_65 vdd gnd cell_6t
Xbit_r66_c51 bl_51 br_51 wl_66 vdd gnd cell_6t
Xbit_r67_c51 bl_51 br_51 wl_67 vdd gnd cell_6t
Xbit_r68_c51 bl_51 br_51 wl_68 vdd gnd cell_6t
Xbit_r69_c51 bl_51 br_51 wl_69 vdd gnd cell_6t
Xbit_r70_c51 bl_51 br_51 wl_70 vdd gnd cell_6t
Xbit_r71_c51 bl_51 br_51 wl_71 vdd gnd cell_6t
Xbit_r72_c51 bl_51 br_51 wl_72 vdd gnd cell_6t
Xbit_r73_c51 bl_51 br_51 wl_73 vdd gnd cell_6t
Xbit_r74_c51 bl_51 br_51 wl_74 vdd gnd cell_6t
Xbit_r75_c51 bl_51 br_51 wl_75 vdd gnd cell_6t
Xbit_r76_c51 bl_51 br_51 wl_76 vdd gnd cell_6t
Xbit_r77_c51 bl_51 br_51 wl_77 vdd gnd cell_6t
Xbit_r78_c51 bl_51 br_51 wl_78 vdd gnd cell_6t
Xbit_r79_c51 bl_51 br_51 wl_79 vdd gnd cell_6t
Xbit_r80_c51 bl_51 br_51 wl_80 vdd gnd cell_6t
Xbit_r81_c51 bl_51 br_51 wl_81 vdd gnd cell_6t
Xbit_r82_c51 bl_51 br_51 wl_82 vdd gnd cell_6t
Xbit_r83_c51 bl_51 br_51 wl_83 vdd gnd cell_6t
Xbit_r84_c51 bl_51 br_51 wl_84 vdd gnd cell_6t
Xbit_r85_c51 bl_51 br_51 wl_85 vdd gnd cell_6t
Xbit_r86_c51 bl_51 br_51 wl_86 vdd gnd cell_6t
Xbit_r87_c51 bl_51 br_51 wl_87 vdd gnd cell_6t
Xbit_r88_c51 bl_51 br_51 wl_88 vdd gnd cell_6t
Xbit_r89_c51 bl_51 br_51 wl_89 vdd gnd cell_6t
Xbit_r90_c51 bl_51 br_51 wl_90 vdd gnd cell_6t
Xbit_r91_c51 bl_51 br_51 wl_91 vdd gnd cell_6t
Xbit_r92_c51 bl_51 br_51 wl_92 vdd gnd cell_6t
Xbit_r93_c51 bl_51 br_51 wl_93 vdd gnd cell_6t
Xbit_r94_c51 bl_51 br_51 wl_94 vdd gnd cell_6t
Xbit_r95_c51 bl_51 br_51 wl_95 vdd gnd cell_6t
Xbit_r96_c51 bl_51 br_51 wl_96 vdd gnd cell_6t
Xbit_r97_c51 bl_51 br_51 wl_97 vdd gnd cell_6t
Xbit_r98_c51 bl_51 br_51 wl_98 vdd gnd cell_6t
Xbit_r99_c51 bl_51 br_51 wl_99 vdd gnd cell_6t
Xbit_r100_c51 bl_51 br_51 wl_100 vdd gnd cell_6t
Xbit_r101_c51 bl_51 br_51 wl_101 vdd gnd cell_6t
Xbit_r102_c51 bl_51 br_51 wl_102 vdd gnd cell_6t
Xbit_r103_c51 bl_51 br_51 wl_103 vdd gnd cell_6t
Xbit_r104_c51 bl_51 br_51 wl_104 vdd gnd cell_6t
Xbit_r105_c51 bl_51 br_51 wl_105 vdd gnd cell_6t
Xbit_r106_c51 bl_51 br_51 wl_106 vdd gnd cell_6t
Xbit_r107_c51 bl_51 br_51 wl_107 vdd gnd cell_6t
Xbit_r108_c51 bl_51 br_51 wl_108 vdd gnd cell_6t
Xbit_r109_c51 bl_51 br_51 wl_109 vdd gnd cell_6t
Xbit_r110_c51 bl_51 br_51 wl_110 vdd gnd cell_6t
Xbit_r111_c51 bl_51 br_51 wl_111 vdd gnd cell_6t
Xbit_r112_c51 bl_51 br_51 wl_112 vdd gnd cell_6t
Xbit_r113_c51 bl_51 br_51 wl_113 vdd gnd cell_6t
Xbit_r114_c51 bl_51 br_51 wl_114 vdd gnd cell_6t
Xbit_r115_c51 bl_51 br_51 wl_115 vdd gnd cell_6t
Xbit_r116_c51 bl_51 br_51 wl_116 vdd gnd cell_6t
Xbit_r117_c51 bl_51 br_51 wl_117 vdd gnd cell_6t
Xbit_r118_c51 bl_51 br_51 wl_118 vdd gnd cell_6t
Xbit_r119_c51 bl_51 br_51 wl_119 vdd gnd cell_6t
Xbit_r120_c51 bl_51 br_51 wl_120 vdd gnd cell_6t
Xbit_r121_c51 bl_51 br_51 wl_121 vdd gnd cell_6t
Xbit_r122_c51 bl_51 br_51 wl_122 vdd gnd cell_6t
Xbit_r123_c51 bl_51 br_51 wl_123 vdd gnd cell_6t
Xbit_r124_c51 bl_51 br_51 wl_124 vdd gnd cell_6t
Xbit_r125_c51 bl_51 br_51 wl_125 vdd gnd cell_6t
Xbit_r126_c51 bl_51 br_51 wl_126 vdd gnd cell_6t
Xbit_r127_c51 bl_51 br_51 wl_127 vdd gnd cell_6t
Xbit_r128_c51 bl_51 br_51 wl_128 vdd gnd cell_6t
Xbit_r129_c51 bl_51 br_51 wl_129 vdd gnd cell_6t
Xbit_r130_c51 bl_51 br_51 wl_130 vdd gnd cell_6t
Xbit_r131_c51 bl_51 br_51 wl_131 vdd gnd cell_6t
Xbit_r132_c51 bl_51 br_51 wl_132 vdd gnd cell_6t
Xbit_r133_c51 bl_51 br_51 wl_133 vdd gnd cell_6t
Xbit_r134_c51 bl_51 br_51 wl_134 vdd gnd cell_6t
Xbit_r135_c51 bl_51 br_51 wl_135 vdd gnd cell_6t
Xbit_r136_c51 bl_51 br_51 wl_136 vdd gnd cell_6t
Xbit_r137_c51 bl_51 br_51 wl_137 vdd gnd cell_6t
Xbit_r138_c51 bl_51 br_51 wl_138 vdd gnd cell_6t
Xbit_r139_c51 bl_51 br_51 wl_139 vdd gnd cell_6t
Xbit_r140_c51 bl_51 br_51 wl_140 vdd gnd cell_6t
Xbit_r141_c51 bl_51 br_51 wl_141 vdd gnd cell_6t
Xbit_r142_c51 bl_51 br_51 wl_142 vdd gnd cell_6t
Xbit_r143_c51 bl_51 br_51 wl_143 vdd gnd cell_6t
Xbit_r144_c51 bl_51 br_51 wl_144 vdd gnd cell_6t
Xbit_r145_c51 bl_51 br_51 wl_145 vdd gnd cell_6t
Xbit_r146_c51 bl_51 br_51 wl_146 vdd gnd cell_6t
Xbit_r147_c51 bl_51 br_51 wl_147 vdd gnd cell_6t
Xbit_r148_c51 bl_51 br_51 wl_148 vdd gnd cell_6t
Xbit_r149_c51 bl_51 br_51 wl_149 vdd gnd cell_6t
Xbit_r150_c51 bl_51 br_51 wl_150 vdd gnd cell_6t
Xbit_r151_c51 bl_51 br_51 wl_151 vdd gnd cell_6t
Xbit_r152_c51 bl_51 br_51 wl_152 vdd gnd cell_6t
Xbit_r153_c51 bl_51 br_51 wl_153 vdd gnd cell_6t
Xbit_r154_c51 bl_51 br_51 wl_154 vdd gnd cell_6t
Xbit_r155_c51 bl_51 br_51 wl_155 vdd gnd cell_6t
Xbit_r156_c51 bl_51 br_51 wl_156 vdd gnd cell_6t
Xbit_r157_c51 bl_51 br_51 wl_157 vdd gnd cell_6t
Xbit_r158_c51 bl_51 br_51 wl_158 vdd gnd cell_6t
Xbit_r159_c51 bl_51 br_51 wl_159 vdd gnd cell_6t
Xbit_r160_c51 bl_51 br_51 wl_160 vdd gnd cell_6t
Xbit_r161_c51 bl_51 br_51 wl_161 vdd gnd cell_6t
Xbit_r162_c51 bl_51 br_51 wl_162 vdd gnd cell_6t
Xbit_r163_c51 bl_51 br_51 wl_163 vdd gnd cell_6t
Xbit_r164_c51 bl_51 br_51 wl_164 vdd gnd cell_6t
Xbit_r165_c51 bl_51 br_51 wl_165 vdd gnd cell_6t
Xbit_r166_c51 bl_51 br_51 wl_166 vdd gnd cell_6t
Xbit_r167_c51 bl_51 br_51 wl_167 vdd gnd cell_6t
Xbit_r168_c51 bl_51 br_51 wl_168 vdd gnd cell_6t
Xbit_r169_c51 bl_51 br_51 wl_169 vdd gnd cell_6t
Xbit_r170_c51 bl_51 br_51 wl_170 vdd gnd cell_6t
Xbit_r171_c51 bl_51 br_51 wl_171 vdd gnd cell_6t
Xbit_r172_c51 bl_51 br_51 wl_172 vdd gnd cell_6t
Xbit_r173_c51 bl_51 br_51 wl_173 vdd gnd cell_6t
Xbit_r174_c51 bl_51 br_51 wl_174 vdd gnd cell_6t
Xbit_r175_c51 bl_51 br_51 wl_175 vdd gnd cell_6t
Xbit_r176_c51 bl_51 br_51 wl_176 vdd gnd cell_6t
Xbit_r177_c51 bl_51 br_51 wl_177 vdd gnd cell_6t
Xbit_r178_c51 bl_51 br_51 wl_178 vdd gnd cell_6t
Xbit_r179_c51 bl_51 br_51 wl_179 vdd gnd cell_6t
Xbit_r180_c51 bl_51 br_51 wl_180 vdd gnd cell_6t
Xbit_r181_c51 bl_51 br_51 wl_181 vdd gnd cell_6t
Xbit_r182_c51 bl_51 br_51 wl_182 vdd gnd cell_6t
Xbit_r183_c51 bl_51 br_51 wl_183 vdd gnd cell_6t
Xbit_r184_c51 bl_51 br_51 wl_184 vdd gnd cell_6t
Xbit_r185_c51 bl_51 br_51 wl_185 vdd gnd cell_6t
Xbit_r186_c51 bl_51 br_51 wl_186 vdd gnd cell_6t
Xbit_r187_c51 bl_51 br_51 wl_187 vdd gnd cell_6t
Xbit_r188_c51 bl_51 br_51 wl_188 vdd gnd cell_6t
Xbit_r189_c51 bl_51 br_51 wl_189 vdd gnd cell_6t
Xbit_r190_c51 bl_51 br_51 wl_190 vdd gnd cell_6t
Xbit_r191_c51 bl_51 br_51 wl_191 vdd gnd cell_6t
Xbit_r192_c51 bl_51 br_51 wl_192 vdd gnd cell_6t
Xbit_r193_c51 bl_51 br_51 wl_193 vdd gnd cell_6t
Xbit_r194_c51 bl_51 br_51 wl_194 vdd gnd cell_6t
Xbit_r195_c51 bl_51 br_51 wl_195 vdd gnd cell_6t
Xbit_r196_c51 bl_51 br_51 wl_196 vdd gnd cell_6t
Xbit_r197_c51 bl_51 br_51 wl_197 vdd gnd cell_6t
Xbit_r198_c51 bl_51 br_51 wl_198 vdd gnd cell_6t
Xbit_r199_c51 bl_51 br_51 wl_199 vdd gnd cell_6t
Xbit_r200_c51 bl_51 br_51 wl_200 vdd gnd cell_6t
Xbit_r201_c51 bl_51 br_51 wl_201 vdd gnd cell_6t
Xbit_r202_c51 bl_51 br_51 wl_202 vdd gnd cell_6t
Xbit_r203_c51 bl_51 br_51 wl_203 vdd gnd cell_6t
Xbit_r204_c51 bl_51 br_51 wl_204 vdd gnd cell_6t
Xbit_r205_c51 bl_51 br_51 wl_205 vdd gnd cell_6t
Xbit_r206_c51 bl_51 br_51 wl_206 vdd gnd cell_6t
Xbit_r207_c51 bl_51 br_51 wl_207 vdd gnd cell_6t
Xbit_r208_c51 bl_51 br_51 wl_208 vdd gnd cell_6t
Xbit_r209_c51 bl_51 br_51 wl_209 vdd gnd cell_6t
Xbit_r210_c51 bl_51 br_51 wl_210 vdd gnd cell_6t
Xbit_r211_c51 bl_51 br_51 wl_211 vdd gnd cell_6t
Xbit_r212_c51 bl_51 br_51 wl_212 vdd gnd cell_6t
Xbit_r213_c51 bl_51 br_51 wl_213 vdd gnd cell_6t
Xbit_r214_c51 bl_51 br_51 wl_214 vdd gnd cell_6t
Xbit_r215_c51 bl_51 br_51 wl_215 vdd gnd cell_6t
Xbit_r216_c51 bl_51 br_51 wl_216 vdd gnd cell_6t
Xbit_r217_c51 bl_51 br_51 wl_217 vdd gnd cell_6t
Xbit_r218_c51 bl_51 br_51 wl_218 vdd gnd cell_6t
Xbit_r219_c51 bl_51 br_51 wl_219 vdd gnd cell_6t
Xbit_r220_c51 bl_51 br_51 wl_220 vdd gnd cell_6t
Xbit_r221_c51 bl_51 br_51 wl_221 vdd gnd cell_6t
Xbit_r222_c51 bl_51 br_51 wl_222 vdd gnd cell_6t
Xbit_r223_c51 bl_51 br_51 wl_223 vdd gnd cell_6t
Xbit_r224_c51 bl_51 br_51 wl_224 vdd gnd cell_6t
Xbit_r225_c51 bl_51 br_51 wl_225 vdd gnd cell_6t
Xbit_r226_c51 bl_51 br_51 wl_226 vdd gnd cell_6t
Xbit_r227_c51 bl_51 br_51 wl_227 vdd gnd cell_6t
Xbit_r228_c51 bl_51 br_51 wl_228 vdd gnd cell_6t
Xbit_r229_c51 bl_51 br_51 wl_229 vdd gnd cell_6t
Xbit_r230_c51 bl_51 br_51 wl_230 vdd gnd cell_6t
Xbit_r231_c51 bl_51 br_51 wl_231 vdd gnd cell_6t
Xbit_r232_c51 bl_51 br_51 wl_232 vdd gnd cell_6t
Xbit_r233_c51 bl_51 br_51 wl_233 vdd gnd cell_6t
Xbit_r234_c51 bl_51 br_51 wl_234 vdd gnd cell_6t
Xbit_r235_c51 bl_51 br_51 wl_235 vdd gnd cell_6t
Xbit_r236_c51 bl_51 br_51 wl_236 vdd gnd cell_6t
Xbit_r237_c51 bl_51 br_51 wl_237 vdd gnd cell_6t
Xbit_r238_c51 bl_51 br_51 wl_238 vdd gnd cell_6t
Xbit_r239_c51 bl_51 br_51 wl_239 vdd gnd cell_6t
Xbit_r240_c51 bl_51 br_51 wl_240 vdd gnd cell_6t
Xbit_r241_c51 bl_51 br_51 wl_241 vdd gnd cell_6t
Xbit_r242_c51 bl_51 br_51 wl_242 vdd gnd cell_6t
Xbit_r243_c51 bl_51 br_51 wl_243 vdd gnd cell_6t
Xbit_r244_c51 bl_51 br_51 wl_244 vdd gnd cell_6t
Xbit_r245_c51 bl_51 br_51 wl_245 vdd gnd cell_6t
Xbit_r246_c51 bl_51 br_51 wl_246 vdd gnd cell_6t
Xbit_r247_c51 bl_51 br_51 wl_247 vdd gnd cell_6t
Xbit_r248_c51 bl_51 br_51 wl_248 vdd gnd cell_6t
Xbit_r249_c51 bl_51 br_51 wl_249 vdd gnd cell_6t
Xbit_r250_c51 bl_51 br_51 wl_250 vdd gnd cell_6t
Xbit_r251_c51 bl_51 br_51 wl_251 vdd gnd cell_6t
Xbit_r252_c51 bl_51 br_51 wl_252 vdd gnd cell_6t
Xbit_r253_c51 bl_51 br_51 wl_253 vdd gnd cell_6t
Xbit_r254_c51 bl_51 br_51 wl_254 vdd gnd cell_6t
Xbit_r255_c51 bl_51 br_51 wl_255 vdd gnd cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd cell_6t
Xbit_r1_c52 bl_52 br_52 wl_1 vdd gnd cell_6t
Xbit_r2_c52 bl_52 br_52 wl_2 vdd gnd cell_6t
Xbit_r3_c52 bl_52 br_52 wl_3 vdd gnd cell_6t
Xbit_r4_c52 bl_52 br_52 wl_4 vdd gnd cell_6t
Xbit_r5_c52 bl_52 br_52 wl_5 vdd gnd cell_6t
Xbit_r6_c52 bl_52 br_52 wl_6 vdd gnd cell_6t
Xbit_r7_c52 bl_52 br_52 wl_7 vdd gnd cell_6t
Xbit_r8_c52 bl_52 br_52 wl_8 vdd gnd cell_6t
Xbit_r9_c52 bl_52 br_52 wl_9 vdd gnd cell_6t
Xbit_r10_c52 bl_52 br_52 wl_10 vdd gnd cell_6t
Xbit_r11_c52 bl_52 br_52 wl_11 vdd gnd cell_6t
Xbit_r12_c52 bl_52 br_52 wl_12 vdd gnd cell_6t
Xbit_r13_c52 bl_52 br_52 wl_13 vdd gnd cell_6t
Xbit_r14_c52 bl_52 br_52 wl_14 vdd gnd cell_6t
Xbit_r15_c52 bl_52 br_52 wl_15 vdd gnd cell_6t
Xbit_r16_c52 bl_52 br_52 wl_16 vdd gnd cell_6t
Xbit_r17_c52 bl_52 br_52 wl_17 vdd gnd cell_6t
Xbit_r18_c52 bl_52 br_52 wl_18 vdd gnd cell_6t
Xbit_r19_c52 bl_52 br_52 wl_19 vdd gnd cell_6t
Xbit_r20_c52 bl_52 br_52 wl_20 vdd gnd cell_6t
Xbit_r21_c52 bl_52 br_52 wl_21 vdd gnd cell_6t
Xbit_r22_c52 bl_52 br_52 wl_22 vdd gnd cell_6t
Xbit_r23_c52 bl_52 br_52 wl_23 vdd gnd cell_6t
Xbit_r24_c52 bl_52 br_52 wl_24 vdd gnd cell_6t
Xbit_r25_c52 bl_52 br_52 wl_25 vdd gnd cell_6t
Xbit_r26_c52 bl_52 br_52 wl_26 vdd gnd cell_6t
Xbit_r27_c52 bl_52 br_52 wl_27 vdd gnd cell_6t
Xbit_r28_c52 bl_52 br_52 wl_28 vdd gnd cell_6t
Xbit_r29_c52 bl_52 br_52 wl_29 vdd gnd cell_6t
Xbit_r30_c52 bl_52 br_52 wl_30 vdd gnd cell_6t
Xbit_r31_c52 bl_52 br_52 wl_31 vdd gnd cell_6t
Xbit_r32_c52 bl_52 br_52 wl_32 vdd gnd cell_6t
Xbit_r33_c52 bl_52 br_52 wl_33 vdd gnd cell_6t
Xbit_r34_c52 bl_52 br_52 wl_34 vdd gnd cell_6t
Xbit_r35_c52 bl_52 br_52 wl_35 vdd gnd cell_6t
Xbit_r36_c52 bl_52 br_52 wl_36 vdd gnd cell_6t
Xbit_r37_c52 bl_52 br_52 wl_37 vdd gnd cell_6t
Xbit_r38_c52 bl_52 br_52 wl_38 vdd gnd cell_6t
Xbit_r39_c52 bl_52 br_52 wl_39 vdd gnd cell_6t
Xbit_r40_c52 bl_52 br_52 wl_40 vdd gnd cell_6t
Xbit_r41_c52 bl_52 br_52 wl_41 vdd gnd cell_6t
Xbit_r42_c52 bl_52 br_52 wl_42 vdd gnd cell_6t
Xbit_r43_c52 bl_52 br_52 wl_43 vdd gnd cell_6t
Xbit_r44_c52 bl_52 br_52 wl_44 vdd gnd cell_6t
Xbit_r45_c52 bl_52 br_52 wl_45 vdd gnd cell_6t
Xbit_r46_c52 bl_52 br_52 wl_46 vdd gnd cell_6t
Xbit_r47_c52 bl_52 br_52 wl_47 vdd gnd cell_6t
Xbit_r48_c52 bl_52 br_52 wl_48 vdd gnd cell_6t
Xbit_r49_c52 bl_52 br_52 wl_49 vdd gnd cell_6t
Xbit_r50_c52 bl_52 br_52 wl_50 vdd gnd cell_6t
Xbit_r51_c52 bl_52 br_52 wl_51 vdd gnd cell_6t
Xbit_r52_c52 bl_52 br_52 wl_52 vdd gnd cell_6t
Xbit_r53_c52 bl_52 br_52 wl_53 vdd gnd cell_6t
Xbit_r54_c52 bl_52 br_52 wl_54 vdd gnd cell_6t
Xbit_r55_c52 bl_52 br_52 wl_55 vdd gnd cell_6t
Xbit_r56_c52 bl_52 br_52 wl_56 vdd gnd cell_6t
Xbit_r57_c52 bl_52 br_52 wl_57 vdd gnd cell_6t
Xbit_r58_c52 bl_52 br_52 wl_58 vdd gnd cell_6t
Xbit_r59_c52 bl_52 br_52 wl_59 vdd gnd cell_6t
Xbit_r60_c52 bl_52 br_52 wl_60 vdd gnd cell_6t
Xbit_r61_c52 bl_52 br_52 wl_61 vdd gnd cell_6t
Xbit_r62_c52 bl_52 br_52 wl_62 vdd gnd cell_6t
Xbit_r63_c52 bl_52 br_52 wl_63 vdd gnd cell_6t
Xbit_r64_c52 bl_52 br_52 wl_64 vdd gnd cell_6t
Xbit_r65_c52 bl_52 br_52 wl_65 vdd gnd cell_6t
Xbit_r66_c52 bl_52 br_52 wl_66 vdd gnd cell_6t
Xbit_r67_c52 bl_52 br_52 wl_67 vdd gnd cell_6t
Xbit_r68_c52 bl_52 br_52 wl_68 vdd gnd cell_6t
Xbit_r69_c52 bl_52 br_52 wl_69 vdd gnd cell_6t
Xbit_r70_c52 bl_52 br_52 wl_70 vdd gnd cell_6t
Xbit_r71_c52 bl_52 br_52 wl_71 vdd gnd cell_6t
Xbit_r72_c52 bl_52 br_52 wl_72 vdd gnd cell_6t
Xbit_r73_c52 bl_52 br_52 wl_73 vdd gnd cell_6t
Xbit_r74_c52 bl_52 br_52 wl_74 vdd gnd cell_6t
Xbit_r75_c52 bl_52 br_52 wl_75 vdd gnd cell_6t
Xbit_r76_c52 bl_52 br_52 wl_76 vdd gnd cell_6t
Xbit_r77_c52 bl_52 br_52 wl_77 vdd gnd cell_6t
Xbit_r78_c52 bl_52 br_52 wl_78 vdd gnd cell_6t
Xbit_r79_c52 bl_52 br_52 wl_79 vdd gnd cell_6t
Xbit_r80_c52 bl_52 br_52 wl_80 vdd gnd cell_6t
Xbit_r81_c52 bl_52 br_52 wl_81 vdd gnd cell_6t
Xbit_r82_c52 bl_52 br_52 wl_82 vdd gnd cell_6t
Xbit_r83_c52 bl_52 br_52 wl_83 vdd gnd cell_6t
Xbit_r84_c52 bl_52 br_52 wl_84 vdd gnd cell_6t
Xbit_r85_c52 bl_52 br_52 wl_85 vdd gnd cell_6t
Xbit_r86_c52 bl_52 br_52 wl_86 vdd gnd cell_6t
Xbit_r87_c52 bl_52 br_52 wl_87 vdd gnd cell_6t
Xbit_r88_c52 bl_52 br_52 wl_88 vdd gnd cell_6t
Xbit_r89_c52 bl_52 br_52 wl_89 vdd gnd cell_6t
Xbit_r90_c52 bl_52 br_52 wl_90 vdd gnd cell_6t
Xbit_r91_c52 bl_52 br_52 wl_91 vdd gnd cell_6t
Xbit_r92_c52 bl_52 br_52 wl_92 vdd gnd cell_6t
Xbit_r93_c52 bl_52 br_52 wl_93 vdd gnd cell_6t
Xbit_r94_c52 bl_52 br_52 wl_94 vdd gnd cell_6t
Xbit_r95_c52 bl_52 br_52 wl_95 vdd gnd cell_6t
Xbit_r96_c52 bl_52 br_52 wl_96 vdd gnd cell_6t
Xbit_r97_c52 bl_52 br_52 wl_97 vdd gnd cell_6t
Xbit_r98_c52 bl_52 br_52 wl_98 vdd gnd cell_6t
Xbit_r99_c52 bl_52 br_52 wl_99 vdd gnd cell_6t
Xbit_r100_c52 bl_52 br_52 wl_100 vdd gnd cell_6t
Xbit_r101_c52 bl_52 br_52 wl_101 vdd gnd cell_6t
Xbit_r102_c52 bl_52 br_52 wl_102 vdd gnd cell_6t
Xbit_r103_c52 bl_52 br_52 wl_103 vdd gnd cell_6t
Xbit_r104_c52 bl_52 br_52 wl_104 vdd gnd cell_6t
Xbit_r105_c52 bl_52 br_52 wl_105 vdd gnd cell_6t
Xbit_r106_c52 bl_52 br_52 wl_106 vdd gnd cell_6t
Xbit_r107_c52 bl_52 br_52 wl_107 vdd gnd cell_6t
Xbit_r108_c52 bl_52 br_52 wl_108 vdd gnd cell_6t
Xbit_r109_c52 bl_52 br_52 wl_109 vdd gnd cell_6t
Xbit_r110_c52 bl_52 br_52 wl_110 vdd gnd cell_6t
Xbit_r111_c52 bl_52 br_52 wl_111 vdd gnd cell_6t
Xbit_r112_c52 bl_52 br_52 wl_112 vdd gnd cell_6t
Xbit_r113_c52 bl_52 br_52 wl_113 vdd gnd cell_6t
Xbit_r114_c52 bl_52 br_52 wl_114 vdd gnd cell_6t
Xbit_r115_c52 bl_52 br_52 wl_115 vdd gnd cell_6t
Xbit_r116_c52 bl_52 br_52 wl_116 vdd gnd cell_6t
Xbit_r117_c52 bl_52 br_52 wl_117 vdd gnd cell_6t
Xbit_r118_c52 bl_52 br_52 wl_118 vdd gnd cell_6t
Xbit_r119_c52 bl_52 br_52 wl_119 vdd gnd cell_6t
Xbit_r120_c52 bl_52 br_52 wl_120 vdd gnd cell_6t
Xbit_r121_c52 bl_52 br_52 wl_121 vdd gnd cell_6t
Xbit_r122_c52 bl_52 br_52 wl_122 vdd gnd cell_6t
Xbit_r123_c52 bl_52 br_52 wl_123 vdd gnd cell_6t
Xbit_r124_c52 bl_52 br_52 wl_124 vdd gnd cell_6t
Xbit_r125_c52 bl_52 br_52 wl_125 vdd gnd cell_6t
Xbit_r126_c52 bl_52 br_52 wl_126 vdd gnd cell_6t
Xbit_r127_c52 bl_52 br_52 wl_127 vdd gnd cell_6t
Xbit_r128_c52 bl_52 br_52 wl_128 vdd gnd cell_6t
Xbit_r129_c52 bl_52 br_52 wl_129 vdd gnd cell_6t
Xbit_r130_c52 bl_52 br_52 wl_130 vdd gnd cell_6t
Xbit_r131_c52 bl_52 br_52 wl_131 vdd gnd cell_6t
Xbit_r132_c52 bl_52 br_52 wl_132 vdd gnd cell_6t
Xbit_r133_c52 bl_52 br_52 wl_133 vdd gnd cell_6t
Xbit_r134_c52 bl_52 br_52 wl_134 vdd gnd cell_6t
Xbit_r135_c52 bl_52 br_52 wl_135 vdd gnd cell_6t
Xbit_r136_c52 bl_52 br_52 wl_136 vdd gnd cell_6t
Xbit_r137_c52 bl_52 br_52 wl_137 vdd gnd cell_6t
Xbit_r138_c52 bl_52 br_52 wl_138 vdd gnd cell_6t
Xbit_r139_c52 bl_52 br_52 wl_139 vdd gnd cell_6t
Xbit_r140_c52 bl_52 br_52 wl_140 vdd gnd cell_6t
Xbit_r141_c52 bl_52 br_52 wl_141 vdd gnd cell_6t
Xbit_r142_c52 bl_52 br_52 wl_142 vdd gnd cell_6t
Xbit_r143_c52 bl_52 br_52 wl_143 vdd gnd cell_6t
Xbit_r144_c52 bl_52 br_52 wl_144 vdd gnd cell_6t
Xbit_r145_c52 bl_52 br_52 wl_145 vdd gnd cell_6t
Xbit_r146_c52 bl_52 br_52 wl_146 vdd gnd cell_6t
Xbit_r147_c52 bl_52 br_52 wl_147 vdd gnd cell_6t
Xbit_r148_c52 bl_52 br_52 wl_148 vdd gnd cell_6t
Xbit_r149_c52 bl_52 br_52 wl_149 vdd gnd cell_6t
Xbit_r150_c52 bl_52 br_52 wl_150 vdd gnd cell_6t
Xbit_r151_c52 bl_52 br_52 wl_151 vdd gnd cell_6t
Xbit_r152_c52 bl_52 br_52 wl_152 vdd gnd cell_6t
Xbit_r153_c52 bl_52 br_52 wl_153 vdd gnd cell_6t
Xbit_r154_c52 bl_52 br_52 wl_154 vdd gnd cell_6t
Xbit_r155_c52 bl_52 br_52 wl_155 vdd gnd cell_6t
Xbit_r156_c52 bl_52 br_52 wl_156 vdd gnd cell_6t
Xbit_r157_c52 bl_52 br_52 wl_157 vdd gnd cell_6t
Xbit_r158_c52 bl_52 br_52 wl_158 vdd gnd cell_6t
Xbit_r159_c52 bl_52 br_52 wl_159 vdd gnd cell_6t
Xbit_r160_c52 bl_52 br_52 wl_160 vdd gnd cell_6t
Xbit_r161_c52 bl_52 br_52 wl_161 vdd gnd cell_6t
Xbit_r162_c52 bl_52 br_52 wl_162 vdd gnd cell_6t
Xbit_r163_c52 bl_52 br_52 wl_163 vdd gnd cell_6t
Xbit_r164_c52 bl_52 br_52 wl_164 vdd gnd cell_6t
Xbit_r165_c52 bl_52 br_52 wl_165 vdd gnd cell_6t
Xbit_r166_c52 bl_52 br_52 wl_166 vdd gnd cell_6t
Xbit_r167_c52 bl_52 br_52 wl_167 vdd gnd cell_6t
Xbit_r168_c52 bl_52 br_52 wl_168 vdd gnd cell_6t
Xbit_r169_c52 bl_52 br_52 wl_169 vdd gnd cell_6t
Xbit_r170_c52 bl_52 br_52 wl_170 vdd gnd cell_6t
Xbit_r171_c52 bl_52 br_52 wl_171 vdd gnd cell_6t
Xbit_r172_c52 bl_52 br_52 wl_172 vdd gnd cell_6t
Xbit_r173_c52 bl_52 br_52 wl_173 vdd gnd cell_6t
Xbit_r174_c52 bl_52 br_52 wl_174 vdd gnd cell_6t
Xbit_r175_c52 bl_52 br_52 wl_175 vdd gnd cell_6t
Xbit_r176_c52 bl_52 br_52 wl_176 vdd gnd cell_6t
Xbit_r177_c52 bl_52 br_52 wl_177 vdd gnd cell_6t
Xbit_r178_c52 bl_52 br_52 wl_178 vdd gnd cell_6t
Xbit_r179_c52 bl_52 br_52 wl_179 vdd gnd cell_6t
Xbit_r180_c52 bl_52 br_52 wl_180 vdd gnd cell_6t
Xbit_r181_c52 bl_52 br_52 wl_181 vdd gnd cell_6t
Xbit_r182_c52 bl_52 br_52 wl_182 vdd gnd cell_6t
Xbit_r183_c52 bl_52 br_52 wl_183 vdd gnd cell_6t
Xbit_r184_c52 bl_52 br_52 wl_184 vdd gnd cell_6t
Xbit_r185_c52 bl_52 br_52 wl_185 vdd gnd cell_6t
Xbit_r186_c52 bl_52 br_52 wl_186 vdd gnd cell_6t
Xbit_r187_c52 bl_52 br_52 wl_187 vdd gnd cell_6t
Xbit_r188_c52 bl_52 br_52 wl_188 vdd gnd cell_6t
Xbit_r189_c52 bl_52 br_52 wl_189 vdd gnd cell_6t
Xbit_r190_c52 bl_52 br_52 wl_190 vdd gnd cell_6t
Xbit_r191_c52 bl_52 br_52 wl_191 vdd gnd cell_6t
Xbit_r192_c52 bl_52 br_52 wl_192 vdd gnd cell_6t
Xbit_r193_c52 bl_52 br_52 wl_193 vdd gnd cell_6t
Xbit_r194_c52 bl_52 br_52 wl_194 vdd gnd cell_6t
Xbit_r195_c52 bl_52 br_52 wl_195 vdd gnd cell_6t
Xbit_r196_c52 bl_52 br_52 wl_196 vdd gnd cell_6t
Xbit_r197_c52 bl_52 br_52 wl_197 vdd gnd cell_6t
Xbit_r198_c52 bl_52 br_52 wl_198 vdd gnd cell_6t
Xbit_r199_c52 bl_52 br_52 wl_199 vdd gnd cell_6t
Xbit_r200_c52 bl_52 br_52 wl_200 vdd gnd cell_6t
Xbit_r201_c52 bl_52 br_52 wl_201 vdd gnd cell_6t
Xbit_r202_c52 bl_52 br_52 wl_202 vdd gnd cell_6t
Xbit_r203_c52 bl_52 br_52 wl_203 vdd gnd cell_6t
Xbit_r204_c52 bl_52 br_52 wl_204 vdd gnd cell_6t
Xbit_r205_c52 bl_52 br_52 wl_205 vdd gnd cell_6t
Xbit_r206_c52 bl_52 br_52 wl_206 vdd gnd cell_6t
Xbit_r207_c52 bl_52 br_52 wl_207 vdd gnd cell_6t
Xbit_r208_c52 bl_52 br_52 wl_208 vdd gnd cell_6t
Xbit_r209_c52 bl_52 br_52 wl_209 vdd gnd cell_6t
Xbit_r210_c52 bl_52 br_52 wl_210 vdd gnd cell_6t
Xbit_r211_c52 bl_52 br_52 wl_211 vdd gnd cell_6t
Xbit_r212_c52 bl_52 br_52 wl_212 vdd gnd cell_6t
Xbit_r213_c52 bl_52 br_52 wl_213 vdd gnd cell_6t
Xbit_r214_c52 bl_52 br_52 wl_214 vdd gnd cell_6t
Xbit_r215_c52 bl_52 br_52 wl_215 vdd gnd cell_6t
Xbit_r216_c52 bl_52 br_52 wl_216 vdd gnd cell_6t
Xbit_r217_c52 bl_52 br_52 wl_217 vdd gnd cell_6t
Xbit_r218_c52 bl_52 br_52 wl_218 vdd gnd cell_6t
Xbit_r219_c52 bl_52 br_52 wl_219 vdd gnd cell_6t
Xbit_r220_c52 bl_52 br_52 wl_220 vdd gnd cell_6t
Xbit_r221_c52 bl_52 br_52 wl_221 vdd gnd cell_6t
Xbit_r222_c52 bl_52 br_52 wl_222 vdd gnd cell_6t
Xbit_r223_c52 bl_52 br_52 wl_223 vdd gnd cell_6t
Xbit_r224_c52 bl_52 br_52 wl_224 vdd gnd cell_6t
Xbit_r225_c52 bl_52 br_52 wl_225 vdd gnd cell_6t
Xbit_r226_c52 bl_52 br_52 wl_226 vdd gnd cell_6t
Xbit_r227_c52 bl_52 br_52 wl_227 vdd gnd cell_6t
Xbit_r228_c52 bl_52 br_52 wl_228 vdd gnd cell_6t
Xbit_r229_c52 bl_52 br_52 wl_229 vdd gnd cell_6t
Xbit_r230_c52 bl_52 br_52 wl_230 vdd gnd cell_6t
Xbit_r231_c52 bl_52 br_52 wl_231 vdd gnd cell_6t
Xbit_r232_c52 bl_52 br_52 wl_232 vdd gnd cell_6t
Xbit_r233_c52 bl_52 br_52 wl_233 vdd gnd cell_6t
Xbit_r234_c52 bl_52 br_52 wl_234 vdd gnd cell_6t
Xbit_r235_c52 bl_52 br_52 wl_235 vdd gnd cell_6t
Xbit_r236_c52 bl_52 br_52 wl_236 vdd gnd cell_6t
Xbit_r237_c52 bl_52 br_52 wl_237 vdd gnd cell_6t
Xbit_r238_c52 bl_52 br_52 wl_238 vdd gnd cell_6t
Xbit_r239_c52 bl_52 br_52 wl_239 vdd gnd cell_6t
Xbit_r240_c52 bl_52 br_52 wl_240 vdd gnd cell_6t
Xbit_r241_c52 bl_52 br_52 wl_241 vdd gnd cell_6t
Xbit_r242_c52 bl_52 br_52 wl_242 vdd gnd cell_6t
Xbit_r243_c52 bl_52 br_52 wl_243 vdd gnd cell_6t
Xbit_r244_c52 bl_52 br_52 wl_244 vdd gnd cell_6t
Xbit_r245_c52 bl_52 br_52 wl_245 vdd gnd cell_6t
Xbit_r246_c52 bl_52 br_52 wl_246 vdd gnd cell_6t
Xbit_r247_c52 bl_52 br_52 wl_247 vdd gnd cell_6t
Xbit_r248_c52 bl_52 br_52 wl_248 vdd gnd cell_6t
Xbit_r249_c52 bl_52 br_52 wl_249 vdd gnd cell_6t
Xbit_r250_c52 bl_52 br_52 wl_250 vdd gnd cell_6t
Xbit_r251_c52 bl_52 br_52 wl_251 vdd gnd cell_6t
Xbit_r252_c52 bl_52 br_52 wl_252 vdd gnd cell_6t
Xbit_r253_c52 bl_52 br_52 wl_253 vdd gnd cell_6t
Xbit_r254_c52 bl_52 br_52 wl_254 vdd gnd cell_6t
Xbit_r255_c52 bl_52 br_52 wl_255 vdd gnd cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd cell_6t
Xbit_r1_c53 bl_53 br_53 wl_1 vdd gnd cell_6t
Xbit_r2_c53 bl_53 br_53 wl_2 vdd gnd cell_6t
Xbit_r3_c53 bl_53 br_53 wl_3 vdd gnd cell_6t
Xbit_r4_c53 bl_53 br_53 wl_4 vdd gnd cell_6t
Xbit_r5_c53 bl_53 br_53 wl_5 vdd gnd cell_6t
Xbit_r6_c53 bl_53 br_53 wl_6 vdd gnd cell_6t
Xbit_r7_c53 bl_53 br_53 wl_7 vdd gnd cell_6t
Xbit_r8_c53 bl_53 br_53 wl_8 vdd gnd cell_6t
Xbit_r9_c53 bl_53 br_53 wl_9 vdd gnd cell_6t
Xbit_r10_c53 bl_53 br_53 wl_10 vdd gnd cell_6t
Xbit_r11_c53 bl_53 br_53 wl_11 vdd gnd cell_6t
Xbit_r12_c53 bl_53 br_53 wl_12 vdd gnd cell_6t
Xbit_r13_c53 bl_53 br_53 wl_13 vdd gnd cell_6t
Xbit_r14_c53 bl_53 br_53 wl_14 vdd gnd cell_6t
Xbit_r15_c53 bl_53 br_53 wl_15 vdd gnd cell_6t
Xbit_r16_c53 bl_53 br_53 wl_16 vdd gnd cell_6t
Xbit_r17_c53 bl_53 br_53 wl_17 vdd gnd cell_6t
Xbit_r18_c53 bl_53 br_53 wl_18 vdd gnd cell_6t
Xbit_r19_c53 bl_53 br_53 wl_19 vdd gnd cell_6t
Xbit_r20_c53 bl_53 br_53 wl_20 vdd gnd cell_6t
Xbit_r21_c53 bl_53 br_53 wl_21 vdd gnd cell_6t
Xbit_r22_c53 bl_53 br_53 wl_22 vdd gnd cell_6t
Xbit_r23_c53 bl_53 br_53 wl_23 vdd gnd cell_6t
Xbit_r24_c53 bl_53 br_53 wl_24 vdd gnd cell_6t
Xbit_r25_c53 bl_53 br_53 wl_25 vdd gnd cell_6t
Xbit_r26_c53 bl_53 br_53 wl_26 vdd gnd cell_6t
Xbit_r27_c53 bl_53 br_53 wl_27 vdd gnd cell_6t
Xbit_r28_c53 bl_53 br_53 wl_28 vdd gnd cell_6t
Xbit_r29_c53 bl_53 br_53 wl_29 vdd gnd cell_6t
Xbit_r30_c53 bl_53 br_53 wl_30 vdd gnd cell_6t
Xbit_r31_c53 bl_53 br_53 wl_31 vdd gnd cell_6t
Xbit_r32_c53 bl_53 br_53 wl_32 vdd gnd cell_6t
Xbit_r33_c53 bl_53 br_53 wl_33 vdd gnd cell_6t
Xbit_r34_c53 bl_53 br_53 wl_34 vdd gnd cell_6t
Xbit_r35_c53 bl_53 br_53 wl_35 vdd gnd cell_6t
Xbit_r36_c53 bl_53 br_53 wl_36 vdd gnd cell_6t
Xbit_r37_c53 bl_53 br_53 wl_37 vdd gnd cell_6t
Xbit_r38_c53 bl_53 br_53 wl_38 vdd gnd cell_6t
Xbit_r39_c53 bl_53 br_53 wl_39 vdd gnd cell_6t
Xbit_r40_c53 bl_53 br_53 wl_40 vdd gnd cell_6t
Xbit_r41_c53 bl_53 br_53 wl_41 vdd gnd cell_6t
Xbit_r42_c53 bl_53 br_53 wl_42 vdd gnd cell_6t
Xbit_r43_c53 bl_53 br_53 wl_43 vdd gnd cell_6t
Xbit_r44_c53 bl_53 br_53 wl_44 vdd gnd cell_6t
Xbit_r45_c53 bl_53 br_53 wl_45 vdd gnd cell_6t
Xbit_r46_c53 bl_53 br_53 wl_46 vdd gnd cell_6t
Xbit_r47_c53 bl_53 br_53 wl_47 vdd gnd cell_6t
Xbit_r48_c53 bl_53 br_53 wl_48 vdd gnd cell_6t
Xbit_r49_c53 bl_53 br_53 wl_49 vdd gnd cell_6t
Xbit_r50_c53 bl_53 br_53 wl_50 vdd gnd cell_6t
Xbit_r51_c53 bl_53 br_53 wl_51 vdd gnd cell_6t
Xbit_r52_c53 bl_53 br_53 wl_52 vdd gnd cell_6t
Xbit_r53_c53 bl_53 br_53 wl_53 vdd gnd cell_6t
Xbit_r54_c53 bl_53 br_53 wl_54 vdd gnd cell_6t
Xbit_r55_c53 bl_53 br_53 wl_55 vdd gnd cell_6t
Xbit_r56_c53 bl_53 br_53 wl_56 vdd gnd cell_6t
Xbit_r57_c53 bl_53 br_53 wl_57 vdd gnd cell_6t
Xbit_r58_c53 bl_53 br_53 wl_58 vdd gnd cell_6t
Xbit_r59_c53 bl_53 br_53 wl_59 vdd gnd cell_6t
Xbit_r60_c53 bl_53 br_53 wl_60 vdd gnd cell_6t
Xbit_r61_c53 bl_53 br_53 wl_61 vdd gnd cell_6t
Xbit_r62_c53 bl_53 br_53 wl_62 vdd gnd cell_6t
Xbit_r63_c53 bl_53 br_53 wl_63 vdd gnd cell_6t
Xbit_r64_c53 bl_53 br_53 wl_64 vdd gnd cell_6t
Xbit_r65_c53 bl_53 br_53 wl_65 vdd gnd cell_6t
Xbit_r66_c53 bl_53 br_53 wl_66 vdd gnd cell_6t
Xbit_r67_c53 bl_53 br_53 wl_67 vdd gnd cell_6t
Xbit_r68_c53 bl_53 br_53 wl_68 vdd gnd cell_6t
Xbit_r69_c53 bl_53 br_53 wl_69 vdd gnd cell_6t
Xbit_r70_c53 bl_53 br_53 wl_70 vdd gnd cell_6t
Xbit_r71_c53 bl_53 br_53 wl_71 vdd gnd cell_6t
Xbit_r72_c53 bl_53 br_53 wl_72 vdd gnd cell_6t
Xbit_r73_c53 bl_53 br_53 wl_73 vdd gnd cell_6t
Xbit_r74_c53 bl_53 br_53 wl_74 vdd gnd cell_6t
Xbit_r75_c53 bl_53 br_53 wl_75 vdd gnd cell_6t
Xbit_r76_c53 bl_53 br_53 wl_76 vdd gnd cell_6t
Xbit_r77_c53 bl_53 br_53 wl_77 vdd gnd cell_6t
Xbit_r78_c53 bl_53 br_53 wl_78 vdd gnd cell_6t
Xbit_r79_c53 bl_53 br_53 wl_79 vdd gnd cell_6t
Xbit_r80_c53 bl_53 br_53 wl_80 vdd gnd cell_6t
Xbit_r81_c53 bl_53 br_53 wl_81 vdd gnd cell_6t
Xbit_r82_c53 bl_53 br_53 wl_82 vdd gnd cell_6t
Xbit_r83_c53 bl_53 br_53 wl_83 vdd gnd cell_6t
Xbit_r84_c53 bl_53 br_53 wl_84 vdd gnd cell_6t
Xbit_r85_c53 bl_53 br_53 wl_85 vdd gnd cell_6t
Xbit_r86_c53 bl_53 br_53 wl_86 vdd gnd cell_6t
Xbit_r87_c53 bl_53 br_53 wl_87 vdd gnd cell_6t
Xbit_r88_c53 bl_53 br_53 wl_88 vdd gnd cell_6t
Xbit_r89_c53 bl_53 br_53 wl_89 vdd gnd cell_6t
Xbit_r90_c53 bl_53 br_53 wl_90 vdd gnd cell_6t
Xbit_r91_c53 bl_53 br_53 wl_91 vdd gnd cell_6t
Xbit_r92_c53 bl_53 br_53 wl_92 vdd gnd cell_6t
Xbit_r93_c53 bl_53 br_53 wl_93 vdd gnd cell_6t
Xbit_r94_c53 bl_53 br_53 wl_94 vdd gnd cell_6t
Xbit_r95_c53 bl_53 br_53 wl_95 vdd gnd cell_6t
Xbit_r96_c53 bl_53 br_53 wl_96 vdd gnd cell_6t
Xbit_r97_c53 bl_53 br_53 wl_97 vdd gnd cell_6t
Xbit_r98_c53 bl_53 br_53 wl_98 vdd gnd cell_6t
Xbit_r99_c53 bl_53 br_53 wl_99 vdd gnd cell_6t
Xbit_r100_c53 bl_53 br_53 wl_100 vdd gnd cell_6t
Xbit_r101_c53 bl_53 br_53 wl_101 vdd gnd cell_6t
Xbit_r102_c53 bl_53 br_53 wl_102 vdd gnd cell_6t
Xbit_r103_c53 bl_53 br_53 wl_103 vdd gnd cell_6t
Xbit_r104_c53 bl_53 br_53 wl_104 vdd gnd cell_6t
Xbit_r105_c53 bl_53 br_53 wl_105 vdd gnd cell_6t
Xbit_r106_c53 bl_53 br_53 wl_106 vdd gnd cell_6t
Xbit_r107_c53 bl_53 br_53 wl_107 vdd gnd cell_6t
Xbit_r108_c53 bl_53 br_53 wl_108 vdd gnd cell_6t
Xbit_r109_c53 bl_53 br_53 wl_109 vdd gnd cell_6t
Xbit_r110_c53 bl_53 br_53 wl_110 vdd gnd cell_6t
Xbit_r111_c53 bl_53 br_53 wl_111 vdd gnd cell_6t
Xbit_r112_c53 bl_53 br_53 wl_112 vdd gnd cell_6t
Xbit_r113_c53 bl_53 br_53 wl_113 vdd gnd cell_6t
Xbit_r114_c53 bl_53 br_53 wl_114 vdd gnd cell_6t
Xbit_r115_c53 bl_53 br_53 wl_115 vdd gnd cell_6t
Xbit_r116_c53 bl_53 br_53 wl_116 vdd gnd cell_6t
Xbit_r117_c53 bl_53 br_53 wl_117 vdd gnd cell_6t
Xbit_r118_c53 bl_53 br_53 wl_118 vdd gnd cell_6t
Xbit_r119_c53 bl_53 br_53 wl_119 vdd gnd cell_6t
Xbit_r120_c53 bl_53 br_53 wl_120 vdd gnd cell_6t
Xbit_r121_c53 bl_53 br_53 wl_121 vdd gnd cell_6t
Xbit_r122_c53 bl_53 br_53 wl_122 vdd gnd cell_6t
Xbit_r123_c53 bl_53 br_53 wl_123 vdd gnd cell_6t
Xbit_r124_c53 bl_53 br_53 wl_124 vdd gnd cell_6t
Xbit_r125_c53 bl_53 br_53 wl_125 vdd gnd cell_6t
Xbit_r126_c53 bl_53 br_53 wl_126 vdd gnd cell_6t
Xbit_r127_c53 bl_53 br_53 wl_127 vdd gnd cell_6t
Xbit_r128_c53 bl_53 br_53 wl_128 vdd gnd cell_6t
Xbit_r129_c53 bl_53 br_53 wl_129 vdd gnd cell_6t
Xbit_r130_c53 bl_53 br_53 wl_130 vdd gnd cell_6t
Xbit_r131_c53 bl_53 br_53 wl_131 vdd gnd cell_6t
Xbit_r132_c53 bl_53 br_53 wl_132 vdd gnd cell_6t
Xbit_r133_c53 bl_53 br_53 wl_133 vdd gnd cell_6t
Xbit_r134_c53 bl_53 br_53 wl_134 vdd gnd cell_6t
Xbit_r135_c53 bl_53 br_53 wl_135 vdd gnd cell_6t
Xbit_r136_c53 bl_53 br_53 wl_136 vdd gnd cell_6t
Xbit_r137_c53 bl_53 br_53 wl_137 vdd gnd cell_6t
Xbit_r138_c53 bl_53 br_53 wl_138 vdd gnd cell_6t
Xbit_r139_c53 bl_53 br_53 wl_139 vdd gnd cell_6t
Xbit_r140_c53 bl_53 br_53 wl_140 vdd gnd cell_6t
Xbit_r141_c53 bl_53 br_53 wl_141 vdd gnd cell_6t
Xbit_r142_c53 bl_53 br_53 wl_142 vdd gnd cell_6t
Xbit_r143_c53 bl_53 br_53 wl_143 vdd gnd cell_6t
Xbit_r144_c53 bl_53 br_53 wl_144 vdd gnd cell_6t
Xbit_r145_c53 bl_53 br_53 wl_145 vdd gnd cell_6t
Xbit_r146_c53 bl_53 br_53 wl_146 vdd gnd cell_6t
Xbit_r147_c53 bl_53 br_53 wl_147 vdd gnd cell_6t
Xbit_r148_c53 bl_53 br_53 wl_148 vdd gnd cell_6t
Xbit_r149_c53 bl_53 br_53 wl_149 vdd gnd cell_6t
Xbit_r150_c53 bl_53 br_53 wl_150 vdd gnd cell_6t
Xbit_r151_c53 bl_53 br_53 wl_151 vdd gnd cell_6t
Xbit_r152_c53 bl_53 br_53 wl_152 vdd gnd cell_6t
Xbit_r153_c53 bl_53 br_53 wl_153 vdd gnd cell_6t
Xbit_r154_c53 bl_53 br_53 wl_154 vdd gnd cell_6t
Xbit_r155_c53 bl_53 br_53 wl_155 vdd gnd cell_6t
Xbit_r156_c53 bl_53 br_53 wl_156 vdd gnd cell_6t
Xbit_r157_c53 bl_53 br_53 wl_157 vdd gnd cell_6t
Xbit_r158_c53 bl_53 br_53 wl_158 vdd gnd cell_6t
Xbit_r159_c53 bl_53 br_53 wl_159 vdd gnd cell_6t
Xbit_r160_c53 bl_53 br_53 wl_160 vdd gnd cell_6t
Xbit_r161_c53 bl_53 br_53 wl_161 vdd gnd cell_6t
Xbit_r162_c53 bl_53 br_53 wl_162 vdd gnd cell_6t
Xbit_r163_c53 bl_53 br_53 wl_163 vdd gnd cell_6t
Xbit_r164_c53 bl_53 br_53 wl_164 vdd gnd cell_6t
Xbit_r165_c53 bl_53 br_53 wl_165 vdd gnd cell_6t
Xbit_r166_c53 bl_53 br_53 wl_166 vdd gnd cell_6t
Xbit_r167_c53 bl_53 br_53 wl_167 vdd gnd cell_6t
Xbit_r168_c53 bl_53 br_53 wl_168 vdd gnd cell_6t
Xbit_r169_c53 bl_53 br_53 wl_169 vdd gnd cell_6t
Xbit_r170_c53 bl_53 br_53 wl_170 vdd gnd cell_6t
Xbit_r171_c53 bl_53 br_53 wl_171 vdd gnd cell_6t
Xbit_r172_c53 bl_53 br_53 wl_172 vdd gnd cell_6t
Xbit_r173_c53 bl_53 br_53 wl_173 vdd gnd cell_6t
Xbit_r174_c53 bl_53 br_53 wl_174 vdd gnd cell_6t
Xbit_r175_c53 bl_53 br_53 wl_175 vdd gnd cell_6t
Xbit_r176_c53 bl_53 br_53 wl_176 vdd gnd cell_6t
Xbit_r177_c53 bl_53 br_53 wl_177 vdd gnd cell_6t
Xbit_r178_c53 bl_53 br_53 wl_178 vdd gnd cell_6t
Xbit_r179_c53 bl_53 br_53 wl_179 vdd gnd cell_6t
Xbit_r180_c53 bl_53 br_53 wl_180 vdd gnd cell_6t
Xbit_r181_c53 bl_53 br_53 wl_181 vdd gnd cell_6t
Xbit_r182_c53 bl_53 br_53 wl_182 vdd gnd cell_6t
Xbit_r183_c53 bl_53 br_53 wl_183 vdd gnd cell_6t
Xbit_r184_c53 bl_53 br_53 wl_184 vdd gnd cell_6t
Xbit_r185_c53 bl_53 br_53 wl_185 vdd gnd cell_6t
Xbit_r186_c53 bl_53 br_53 wl_186 vdd gnd cell_6t
Xbit_r187_c53 bl_53 br_53 wl_187 vdd gnd cell_6t
Xbit_r188_c53 bl_53 br_53 wl_188 vdd gnd cell_6t
Xbit_r189_c53 bl_53 br_53 wl_189 vdd gnd cell_6t
Xbit_r190_c53 bl_53 br_53 wl_190 vdd gnd cell_6t
Xbit_r191_c53 bl_53 br_53 wl_191 vdd gnd cell_6t
Xbit_r192_c53 bl_53 br_53 wl_192 vdd gnd cell_6t
Xbit_r193_c53 bl_53 br_53 wl_193 vdd gnd cell_6t
Xbit_r194_c53 bl_53 br_53 wl_194 vdd gnd cell_6t
Xbit_r195_c53 bl_53 br_53 wl_195 vdd gnd cell_6t
Xbit_r196_c53 bl_53 br_53 wl_196 vdd gnd cell_6t
Xbit_r197_c53 bl_53 br_53 wl_197 vdd gnd cell_6t
Xbit_r198_c53 bl_53 br_53 wl_198 vdd gnd cell_6t
Xbit_r199_c53 bl_53 br_53 wl_199 vdd gnd cell_6t
Xbit_r200_c53 bl_53 br_53 wl_200 vdd gnd cell_6t
Xbit_r201_c53 bl_53 br_53 wl_201 vdd gnd cell_6t
Xbit_r202_c53 bl_53 br_53 wl_202 vdd gnd cell_6t
Xbit_r203_c53 bl_53 br_53 wl_203 vdd gnd cell_6t
Xbit_r204_c53 bl_53 br_53 wl_204 vdd gnd cell_6t
Xbit_r205_c53 bl_53 br_53 wl_205 vdd gnd cell_6t
Xbit_r206_c53 bl_53 br_53 wl_206 vdd gnd cell_6t
Xbit_r207_c53 bl_53 br_53 wl_207 vdd gnd cell_6t
Xbit_r208_c53 bl_53 br_53 wl_208 vdd gnd cell_6t
Xbit_r209_c53 bl_53 br_53 wl_209 vdd gnd cell_6t
Xbit_r210_c53 bl_53 br_53 wl_210 vdd gnd cell_6t
Xbit_r211_c53 bl_53 br_53 wl_211 vdd gnd cell_6t
Xbit_r212_c53 bl_53 br_53 wl_212 vdd gnd cell_6t
Xbit_r213_c53 bl_53 br_53 wl_213 vdd gnd cell_6t
Xbit_r214_c53 bl_53 br_53 wl_214 vdd gnd cell_6t
Xbit_r215_c53 bl_53 br_53 wl_215 vdd gnd cell_6t
Xbit_r216_c53 bl_53 br_53 wl_216 vdd gnd cell_6t
Xbit_r217_c53 bl_53 br_53 wl_217 vdd gnd cell_6t
Xbit_r218_c53 bl_53 br_53 wl_218 vdd gnd cell_6t
Xbit_r219_c53 bl_53 br_53 wl_219 vdd gnd cell_6t
Xbit_r220_c53 bl_53 br_53 wl_220 vdd gnd cell_6t
Xbit_r221_c53 bl_53 br_53 wl_221 vdd gnd cell_6t
Xbit_r222_c53 bl_53 br_53 wl_222 vdd gnd cell_6t
Xbit_r223_c53 bl_53 br_53 wl_223 vdd gnd cell_6t
Xbit_r224_c53 bl_53 br_53 wl_224 vdd gnd cell_6t
Xbit_r225_c53 bl_53 br_53 wl_225 vdd gnd cell_6t
Xbit_r226_c53 bl_53 br_53 wl_226 vdd gnd cell_6t
Xbit_r227_c53 bl_53 br_53 wl_227 vdd gnd cell_6t
Xbit_r228_c53 bl_53 br_53 wl_228 vdd gnd cell_6t
Xbit_r229_c53 bl_53 br_53 wl_229 vdd gnd cell_6t
Xbit_r230_c53 bl_53 br_53 wl_230 vdd gnd cell_6t
Xbit_r231_c53 bl_53 br_53 wl_231 vdd gnd cell_6t
Xbit_r232_c53 bl_53 br_53 wl_232 vdd gnd cell_6t
Xbit_r233_c53 bl_53 br_53 wl_233 vdd gnd cell_6t
Xbit_r234_c53 bl_53 br_53 wl_234 vdd gnd cell_6t
Xbit_r235_c53 bl_53 br_53 wl_235 vdd gnd cell_6t
Xbit_r236_c53 bl_53 br_53 wl_236 vdd gnd cell_6t
Xbit_r237_c53 bl_53 br_53 wl_237 vdd gnd cell_6t
Xbit_r238_c53 bl_53 br_53 wl_238 vdd gnd cell_6t
Xbit_r239_c53 bl_53 br_53 wl_239 vdd gnd cell_6t
Xbit_r240_c53 bl_53 br_53 wl_240 vdd gnd cell_6t
Xbit_r241_c53 bl_53 br_53 wl_241 vdd gnd cell_6t
Xbit_r242_c53 bl_53 br_53 wl_242 vdd gnd cell_6t
Xbit_r243_c53 bl_53 br_53 wl_243 vdd gnd cell_6t
Xbit_r244_c53 bl_53 br_53 wl_244 vdd gnd cell_6t
Xbit_r245_c53 bl_53 br_53 wl_245 vdd gnd cell_6t
Xbit_r246_c53 bl_53 br_53 wl_246 vdd gnd cell_6t
Xbit_r247_c53 bl_53 br_53 wl_247 vdd gnd cell_6t
Xbit_r248_c53 bl_53 br_53 wl_248 vdd gnd cell_6t
Xbit_r249_c53 bl_53 br_53 wl_249 vdd gnd cell_6t
Xbit_r250_c53 bl_53 br_53 wl_250 vdd gnd cell_6t
Xbit_r251_c53 bl_53 br_53 wl_251 vdd gnd cell_6t
Xbit_r252_c53 bl_53 br_53 wl_252 vdd gnd cell_6t
Xbit_r253_c53 bl_53 br_53 wl_253 vdd gnd cell_6t
Xbit_r254_c53 bl_53 br_53 wl_254 vdd gnd cell_6t
Xbit_r255_c53 bl_53 br_53 wl_255 vdd gnd cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd cell_6t
Xbit_r1_c54 bl_54 br_54 wl_1 vdd gnd cell_6t
Xbit_r2_c54 bl_54 br_54 wl_2 vdd gnd cell_6t
Xbit_r3_c54 bl_54 br_54 wl_3 vdd gnd cell_6t
Xbit_r4_c54 bl_54 br_54 wl_4 vdd gnd cell_6t
Xbit_r5_c54 bl_54 br_54 wl_5 vdd gnd cell_6t
Xbit_r6_c54 bl_54 br_54 wl_6 vdd gnd cell_6t
Xbit_r7_c54 bl_54 br_54 wl_7 vdd gnd cell_6t
Xbit_r8_c54 bl_54 br_54 wl_8 vdd gnd cell_6t
Xbit_r9_c54 bl_54 br_54 wl_9 vdd gnd cell_6t
Xbit_r10_c54 bl_54 br_54 wl_10 vdd gnd cell_6t
Xbit_r11_c54 bl_54 br_54 wl_11 vdd gnd cell_6t
Xbit_r12_c54 bl_54 br_54 wl_12 vdd gnd cell_6t
Xbit_r13_c54 bl_54 br_54 wl_13 vdd gnd cell_6t
Xbit_r14_c54 bl_54 br_54 wl_14 vdd gnd cell_6t
Xbit_r15_c54 bl_54 br_54 wl_15 vdd gnd cell_6t
Xbit_r16_c54 bl_54 br_54 wl_16 vdd gnd cell_6t
Xbit_r17_c54 bl_54 br_54 wl_17 vdd gnd cell_6t
Xbit_r18_c54 bl_54 br_54 wl_18 vdd gnd cell_6t
Xbit_r19_c54 bl_54 br_54 wl_19 vdd gnd cell_6t
Xbit_r20_c54 bl_54 br_54 wl_20 vdd gnd cell_6t
Xbit_r21_c54 bl_54 br_54 wl_21 vdd gnd cell_6t
Xbit_r22_c54 bl_54 br_54 wl_22 vdd gnd cell_6t
Xbit_r23_c54 bl_54 br_54 wl_23 vdd gnd cell_6t
Xbit_r24_c54 bl_54 br_54 wl_24 vdd gnd cell_6t
Xbit_r25_c54 bl_54 br_54 wl_25 vdd gnd cell_6t
Xbit_r26_c54 bl_54 br_54 wl_26 vdd gnd cell_6t
Xbit_r27_c54 bl_54 br_54 wl_27 vdd gnd cell_6t
Xbit_r28_c54 bl_54 br_54 wl_28 vdd gnd cell_6t
Xbit_r29_c54 bl_54 br_54 wl_29 vdd gnd cell_6t
Xbit_r30_c54 bl_54 br_54 wl_30 vdd gnd cell_6t
Xbit_r31_c54 bl_54 br_54 wl_31 vdd gnd cell_6t
Xbit_r32_c54 bl_54 br_54 wl_32 vdd gnd cell_6t
Xbit_r33_c54 bl_54 br_54 wl_33 vdd gnd cell_6t
Xbit_r34_c54 bl_54 br_54 wl_34 vdd gnd cell_6t
Xbit_r35_c54 bl_54 br_54 wl_35 vdd gnd cell_6t
Xbit_r36_c54 bl_54 br_54 wl_36 vdd gnd cell_6t
Xbit_r37_c54 bl_54 br_54 wl_37 vdd gnd cell_6t
Xbit_r38_c54 bl_54 br_54 wl_38 vdd gnd cell_6t
Xbit_r39_c54 bl_54 br_54 wl_39 vdd gnd cell_6t
Xbit_r40_c54 bl_54 br_54 wl_40 vdd gnd cell_6t
Xbit_r41_c54 bl_54 br_54 wl_41 vdd gnd cell_6t
Xbit_r42_c54 bl_54 br_54 wl_42 vdd gnd cell_6t
Xbit_r43_c54 bl_54 br_54 wl_43 vdd gnd cell_6t
Xbit_r44_c54 bl_54 br_54 wl_44 vdd gnd cell_6t
Xbit_r45_c54 bl_54 br_54 wl_45 vdd gnd cell_6t
Xbit_r46_c54 bl_54 br_54 wl_46 vdd gnd cell_6t
Xbit_r47_c54 bl_54 br_54 wl_47 vdd gnd cell_6t
Xbit_r48_c54 bl_54 br_54 wl_48 vdd gnd cell_6t
Xbit_r49_c54 bl_54 br_54 wl_49 vdd gnd cell_6t
Xbit_r50_c54 bl_54 br_54 wl_50 vdd gnd cell_6t
Xbit_r51_c54 bl_54 br_54 wl_51 vdd gnd cell_6t
Xbit_r52_c54 bl_54 br_54 wl_52 vdd gnd cell_6t
Xbit_r53_c54 bl_54 br_54 wl_53 vdd gnd cell_6t
Xbit_r54_c54 bl_54 br_54 wl_54 vdd gnd cell_6t
Xbit_r55_c54 bl_54 br_54 wl_55 vdd gnd cell_6t
Xbit_r56_c54 bl_54 br_54 wl_56 vdd gnd cell_6t
Xbit_r57_c54 bl_54 br_54 wl_57 vdd gnd cell_6t
Xbit_r58_c54 bl_54 br_54 wl_58 vdd gnd cell_6t
Xbit_r59_c54 bl_54 br_54 wl_59 vdd gnd cell_6t
Xbit_r60_c54 bl_54 br_54 wl_60 vdd gnd cell_6t
Xbit_r61_c54 bl_54 br_54 wl_61 vdd gnd cell_6t
Xbit_r62_c54 bl_54 br_54 wl_62 vdd gnd cell_6t
Xbit_r63_c54 bl_54 br_54 wl_63 vdd gnd cell_6t
Xbit_r64_c54 bl_54 br_54 wl_64 vdd gnd cell_6t
Xbit_r65_c54 bl_54 br_54 wl_65 vdd gnd cell_6t
Xbit_r66_c54 bl_54 br_54 wl_66 vdd gnd cell_6t
Xbit_r67_c54 bl_54 br_54 wl_67 vdd gnd cell_6t
Xbit_r68_c54 bl_54 br_54 wl_68 vdd gnd cell_6t
Xbit_r69_c54 bl_54 br_54 wl_69 vdd gnd cell_6t
Xbit_r70_c54 bl_54 br_54 wl_70 vdd gnd cell_6t
Xbit_r71_c54 bl_54 br_54 wl_71 vdd gnd cell_6t
Xbit_r72_c54 bl_54 br_54 wl_72 vdd gnd cell_6t
Xbit_r73_c54 bl_54 br_54 wl_73 vdd gnd cell_6t
Xbit_r74_c54 bl_54 br_54 wl_74 vdd gnd cell_6t
Xbit_r75_c54 bl_54 br_54 wl_75 vdd gnd cell_6t
Xbit_r76_c54 bl_54 br_54 wl_76 vdd gnd cell_6t
Xbit_r77_c54 bl_54 br_54 wl_77 vdd gnd cell_6t
Xbit_r78_c54 bl_54 br_54 wl_78 vdd gnd cell_6t
Xbit_r79_c54 bl_54 br_54 wl_79 vdd gnd cell_6t
Xbit_r80_c54 bl_54 br_54 wl_80 vdd gnd cell_6t
Xbit_r81_c54 bl_54 br_54 wl_81 vdd gnd cell_6t
Xbit_r82_c54 bl_54 br_54 wl_82 vdd gnd cell_6t
Xbit_r83_c54 bl_54 br_54 wl_83 vdd gnd cell_6t
Xbit_r84_c54 bl_54 br_54 wl_84 vdd gnd cell_6t
Xbit_r85_c54 bl_54 br_54 wl_85 vdd gnd cell_6t
Xbit_r86_c54 bl_54 br_54 wl_86 vdd gnd cell_6t
Xbit_r87_c54 bl_54 br_54 wl_87 vdd gnd cell_6t
Xbit_r88_c54 bl_54 br_54 wl_88 vdd gnd cell_6t
Xbit_r89_c54 bl_54 br_54 wl_89 vdd gnd cell_6t
Xbit_r90_c54 bl_54 br_54 wl_90 vdd gnd cell_6t
Xbit_r91_c54 bl_54 br_54 wl_91 vdd gnd cell_6t
Xbit_r92_c54 bl_54 br_54 wl_92 vdd gnd cell_6t
Xbit_r93_c54 bl_54 br_54 wl_93 vdd gnd cell_6t
Xbit_r94_c54 bl_54 br_54 wl_94 vdd gnd cell_6t
Xbit_r95_c54 bl_54 br_54 wl_95 vdd gnd cell_6t
Xbit_r96_c54 bl_54 br_54 wl_96 vdd gnd cell_6t
Xbit_r97_c54 bl_54 br_54 wl_97 vdd gnd cell_6t
Xbit_r98_c54 bl_54 br_54 wl_98 vdd gnd cell_6t
Xbit_r99_c54 bl_54 br_54 wl_99 vdd gnd cell_6t
Xbit_r100_c54 bl_54 br_54 wl_100 vdd gnd cell_6t
Xbit_r101_c54 bl_54 br_54 wl_101 vdd gnd cell_6t
Xbit_r102_c54 bl_54 br_54 wl_102 vdd gnd cell_6t
Xbit_r103_c54 bl_54 br_54 wl_103 vdd gnd cell_6t
Xbit_r104_c54 bl_54 br_54 wl_104 vdd gnd cell_6t
Xbit_r105_c54 bl_54 br_54 wl_105 vdd gnd cell_6t
Xbit_r106_c54 bl_54 br_54 wl_106 vdd gnd cell_6t
Xbit_r107_c54 bl_54 br_54 wl_107 vdd gnd cell_6t
Xbit_r108_c54 bl_54 br_54 wl_108 vdd gnd cell_6t
Xbit_r109_c54 bl_54 br_54 wl_109 vdd gnd cell_6t
Xbit_r110_c54 bl_54 br_54 wl_110 vdd gnd cell_6t
Xbit_r111_c54 bl_54 br_54 wl_111 vdd gnd cell_6t
Xbit_r112_c54 bl_54 br_54 wl_112 vdd gnd cell_6t
Xbit_r113_c54 bl_54 br_54 wl_113 vdd gnd cell_6t
Xbit_r114_c54 bl_54 br_54 wl_114 vdd gnd cell_6t
Xbit_r115_c54 bl_54 br_54 wl_115 vdd gnd cell_6t
Xbit_r116_c54 bl_54 br_54 wl_116 vdd gnd cell_6t
Xbit_r117_c54 bl_54 br_54 wl_117 vdd gnd cell_6t
Xbit_r118_c54 bl_54 br_54 wl_118 vdd gnd cell_6t
Xbit_r119_c54 bl_54 br_54 wl_119 vdd gnd cell_6t
Xbit_r120_c54 bl_54 br_54 wl_120 vdd gnd cell_6t
Xbit_r121_c54 bl_54 br_54 wl_121 vdd gnd cell_6t
Xbit_r122_c54 bl_54 br_54 wl_122 vdd gnd cell_6t
Xbit_r123_c54 bl_54 br_54 wl_123 vdd gnd cell_6t
Xbit_r124_c54 bl_54 br_54 wl_124 vdd gnd cell_6t
Xbit_r125_c54 bl_54 br_54 wl_125 vdd gnd cell_6t
Xbit_r126_c54 bl_54 br_54 wl_126 vdd gnd cell_6t
Xbit_r127_c54 bl_54 br_54 wl_127 vdd gnd cell_6t
Xbit_r128_c54 bl_54 br_54 wl_128 vdd gnd cell_6t
Xbit_r129_c54 bl_54 br_54 wl_129 vdd gnd cell_6t
Xbit_r130_c54 bl_54 br_54 wl_130 vdd gnd cell_6t
Xbit_r131_c54 bl_54 br_54 wl_131 vdd gnd cell_6t
Xbit_r132_c54 bl_54 br_54 wl_132 vdd gnd cell_6t
Xbit_r133_c54 bl_54 br_54 wl_133 vdd gnd cell_6t
Xbit_r134_c54 bl_54 br_54 wl_134 vdd gnd cell_6t
Xbit_r135_c54 bl_54 br_54 wl_135 vdd gnd cell_6t
Xbit_r136_c54 bl_54 br_54 wl_136 vdd gnd cell_6t
Xbit_r137_c54 bl_54 br_54 wl_137 vdd gnd cell_6t
Xbit_r138_c54 bl_54 br_54 wl_138 vdd gnd cell_6t
Xbit_r139_c54 bl_54 br_54 wl_139 vdd gnd cell_6t
Xbit_r140_c54 bl_54 br_54 wl_140 vdd gnd cell_6t
Xbit_r141_c54 bl_54 br_54 wl_141 vdd gnd cell_6t
Xbit_r142_c54 bl_54 br_54 wl_142 vdd gnd cell_6t
Xbit_r143_c54 bl_54 br_54 wl_143 vdd gnd cell_6t
Xbit_r144_c54 bl_54 br_54 wl_144 vdd gnd cell_6t
Xbit_r145_c54 bl_54 br_54 wl_145 vdd gnd cell_6t
Xbit_r146_c54 bl_54 br_54 wl_146 vdd gnd cell_6t
Xbit_r147_c54 bl_54 br_54 wl_147 vdd gnd cell_6t
Xbit_r148_c54 bl_54 br_54 wl_148 vdd gnd cell_6t
Xbit_r149_c54 bl_54 br_54 wl_149 vdd gnd cell_6t
Xbit_r150_c54 bl_54 br_54 wl_150 vdd gnd cell_6t
Xbit_r151_c54 bl_54 br_54 wl_151 vdd gnd cell_6t
Xbit_r152_c54 bl_54 br_54 wl_152 vdd gnd cell_6t
Xbit_r153_c54 bl_54 br_54 wl_153 vdd gnd cell_6t
Xbit_r154_c54 bl_54 br_54 wl_154 vdd gnd cell_6t
Xbit_r155_c54 bl_54 br_54 wl_155 vdd gnd cell_6t
Xbit_r156_c54 bl_54 br_54 wl_156 vdd gnd cell_6t
Xbit_r157_c54 bl_54 br_54 wl_157 vdd gnd cell_6t
Xbit_r158_c54 bl_54 br_54 wl_158 vdd gnd cell_6t
Xbit_r159_c54 bl_54 br_54 wl_159 vdd gnd cell_6t
Xbit_r160_c54 bl_54 br_54 wl_160 vdd gnd cell_6t
Xbit_r161_c54 bl_54 br_54 wl_161 vdd gnd cell_6t
Xbit_r162_c54 bl_54 br_54 wl_162 vdd gnd cell_6t
Xbit_r163_c54 bl_54 br_54 wl_163 vdd gnd cell_6t
Xbit_r164_c54 bl_54 br_54 wl_164 vdd gnd cell_6t
Xbit_r165_c54 bl_54 br_54 wl_165 vdd gnd cell_6t
Xbit_r166_c54 bl_54 br_54 wl_166 vdd gnd cell_6t
Xbit_r167_c54 bl_54 br_54 wl_167 vdd gnd cell_6t
Xbit_r168_c54 bl_54 br_54 wl_168 vdd gnd cell_6t
Xbit_r169_c54 bl_54 br_54 wl_169 vdd gnd cell_6t
Xbit_r170_c54 bl_54 br_54 wl_170 vdd gnd cell_6t
Xbit_r171_c54 bl_54 br_54 wl_171 vdd gnd cell_6t
Xbit_r172_c54 bl_54 br_54 wl_172 vdd gnd cell_6t
Xbit_r173_c54 bl_54 br_54 wl_173 vdd gnd cell_6t
Xbit_r174_c54 bl_54 br_54 wl_174 vdd gnd cell_6t
Xbit_r175_c54 bl_54 br_54 wl_175 vdd gnd cell_6t
Xbit_r176_c54 bl_54 br_54 wl_176 vdd gnd cell_6t
Xbit_r177_c54 bl_54 br_54 wl_177 vdd gnd cell_6t
Xbit_r178_c54 bl_54 br_54 wl_178 vdd gnd cell_6t
Xbit_r179_c54 bl_54 br_54 wl_179 vdd gnd cell_6t
Xbit_r180_c54 bl_54 br_54 wl_180 vdd gnd cell_6t
Xbit_r181_c54 bl_54 br_54 wl_181 vdd gnd cell_6t
Xbit_r182_c54 bl_54 br_54 wl_182 vdd gnd cell_6t
Xbit_r183_c54 bl_54 br_54 wl_183 vdd gnd cell_6t
Xbit_r184_c54 bl_54 br_54 wl_184 vdd gnd cell_6t
Xbit_r185_c54 bl_54 br_54 wl_185 vdd gnd cell_6t
Xbit_r186_c54 bl_54 br_54 wl_186 vdd gnd cell_6t
Xbit_r187_c54 bl_54 br_54 wl_187 vdd gnd cell_6t
Xbit_r188_c54 bl_54 br_54 wl_188 vdd gnd cell_6t
Xbit_r189_c54 bl_54 br_54 wl_189 vdd gnd cell_6t
Xbit_r190_c54 bl_54 br_54 wl_190 vdd gnd cell_6t
Xbit_r191_c54 bl_54 br_54 wl_191 vdd gnd cell_6t
Xbit_r192_c54 bl_54 br_54 wl_192 vdd gnd cell_6t
Xbit_r193_c54 bl_54 br_54 wl_193 vdd gnd cell_6t
Xbit_r194_c54 bl_54 br_54 wl_194 vdd gnd cell_6t
Xbit_r195_c54 bl_54 br_54 wl_195 vdd gnd cell_6t
Xbit_r196_c54 bl_54 br_54 wl_196 vdd gnd cell_6t
Xbit_r197_c54 bl_54 br_54 wl_197 vdd gnd cell_6t
Xbit_r198_c54 bl_54 br_54 wl_198 vdd gnd cell_6t
Xbit_r199_c54 bl_54 br_54 wl_199 vdd gnd cell_6t
Xbit_r200_c54 bl_54 br_54 wl_200 vdd gnd cell_6t
Xbit_r201_c54 bl_54 br_54 wl_201 vdd gnd cell_6t
Xbit_r202_c54 bl_54 br_54 wl_202 vdd gnd cell_6t
Xbit_r203_c54 bl_54 br_54 wl_203 vdd gnd cell_6t
Xbit_r204_c54 bl_54 br_54 wl_204 vdd gnd cell_6t
Xbit_r205_c54 bl_54 br_54 wl_205 vdd gnd cell_6t
Xbit_r206_c54 bl_54 br_54 wl_206 vdd gnd cell_6t
Xbit_r207_c54 bl_54 br_54 wl_207 vdd gnd cell_6t
Xbit_r208_c54 bl_54 br_54 wl_208 vdd gnd cell_6t
Xbit_r209_c54 bl_54 br_54 wl_209 vdd gnd cell_6t
Xbit_r210_c54 bl_54 br_54 wl_210 vdd gnd cell_6t
Xbit_r211_c54 bl_54 br_54 wl_211 vdd gnd cell_6t
Xbit_r212_c54 bl_54 br_54 wl_212 vdd gnd cell_6t
Xbit_r213_c54 bl_54 br_54 wl_213 vdd gnd cell_6t
Xbit_r214_c54 bl_54 br_54 wl_214 vdd gnd cell_6t
Xbit_r215_c54 bl_54 br_54 wl_215 vdd gnd cell_6t
Xbit_r216_c54 bl_54 br_54 wl_216 vdd gnd cell_6t
Xbit_r217_c54 bl_54 br_54 wl_217 vdd gnd cell_6t
Xbit_r218_c54 bl_54 br_54 wl_218 vdd gnd cell_6t
Xbit_r219_c54 bl_54 br_54 wl_219 vdd gnd cell_6t
Xbit_r220_c54 bl_54 br_54 wl_220 vdd gnd cell_6t
Xbit_r221_c54 bl_54 br_54 wl_221 vdd gnd cell_6t
Xbit_r222_c54 bl_54 br_54 wl_222 vdd gnd cell_6t
Xbit_r223_c54 bl_54 br_54 wl_223 vdd gnd cell_6t
Xbit_r224_c54 bl_54 br_54 wl_224 vdd gnd cell_6t
Xbit_r225_c54 bl_54 br_54 wl_225 vdd gnd cell_6t
Xbit_r226_c54 bl_54 br_54 wl_226 vdd gnd cell_6t
Xbit_r227_c54 bl_54 br_54 wl_227 vdd gnd cell_6t
Xbit_r228_c54 bl_54 br_54 wl_228 vdd gnd cell_6t
Xbit_r229_c54 bl_54 br_54 wl_229 vdd gnd cell_6t
Xbit_r230_c54 bl_54 br_54 wl_230 vdd gnd cell_6t
Xbit_r231_c54 bl_54 br_54 wl_231 vdd gnd cell_6t
Xbit_r232_c54 bl_54 br_54 wl_232 vdd gnd cell_6t
Xbit_r233_c54 bl_54 br_54 wl_233 vdd gnd cell_6t
Xbit_r234_c54 bl_54 br_54 wl_234 vdd gnd cell_6t
Xbit_r235_c54 bl_54 br_54 wl_235 vdd gnd cell_6t
Xbit_r236_c54 bl_54 br_54 wl_236 vdd gnd cell_6t
Xbit_r237_c54 bl_54 br_54 wl_237 vdd gnd cell_6t
Xbit_r238_c54 bl_54 br_54 wl_238 vdd gnd cell_6t
Xbit_r239_c54 bl_54 br_54 wl_239 vdd gnd cell_6t
Xbit_r240_c54 bl_54 br_54 wl_240 vdd gnd cell_6t
Xbit_r241_c54 bl_54 br_54 wl_241 vdd gnd cell_6t
Xbit_r242_c54 bl_54 br_54 wl_242 vdd gnd cell_6t
Xbit_r243_c54 bl_54 br_54 wl_243 vdd gnd cell_6t
Xbit_r244_c54 bl_54 br_54 wl_244 vdd gnd cell_6t
Xbit_r245_c54 bl_54 br_54 wl_245 vdd gnd cell_6t
Xbit_r246_c54 bl_54 br_54 wl_246 vdd gnd cell_6t
Xbit_r247_c54 bl_54 br_54 wl_247 vdd gnd cell_6t
Xbit_r248_c54 bl_54 br_54 wl_248 vdd gnd cell_6t
Xbit_r249_c54 bl_54 br_54 wl_249 vdd gnd cell_6t
Xbit_r250_c54 bl_54 br_54 wl_250 vdd gnd cell_6t
Xbit_r251_c54 bl_54 br_54 wl_251 vdd gnd cell_6t
Xbit_r252_c54 bl_54 br_54 wl_252 vdd gnd cell_6t
Xbit_r253_c54 bl_54 br_54 wl_253 vdd gnd cell_6t
Xbit_r254_c54 bl_54 br_54 wl_254 vdd gnd cell_6t
Xbit_r255_c54 bl_54 br_54 wl_255 vdd gnd cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd cell_6t
Xbit_r1_c55 bl_55 br_55 wl_1 vdd gnd cell_6t
Xbit_r2_c55 bl_55 br_55 wl_2 vdd gnd cell_6t
Xbit_r3_c55 bl_55 br_55 wl_3 vdd gnd cell_6t
Xbit_r4_c55 bl_55 br_55 wl_4 vdd gnd cell_6t
Xbit_r5_c55 bl_55 br_55 wl_5 vdd gnd cell_6t
Xbit_r6_c55 bl_55 br_55 wl_6 vdd gnd cell_6t
Xbit_r7_c55 bl_55 br_55 wl_7 vdd gnd cell_6t
Xbit_r8_c55 bl_55 br_55 wl_8 vdd gnd cell_6t
Xbit_r9_c55 bl_55 br_55 wl_9 vdd gnd cell_6t
Xbit_r10_c55 bl_55 br_55 wl_10 vdd gnd cell_6t
Xbit_r11_c55 bl_55 br_55 wl_11 vdd gnd cell_6t
Xbit_r12_c55 bl_55 br_55 wl_12 vdd gnd cell_6t
Xbit_r13_c55 bl_55 br_55 wl_13 vdd gnd cell_6t
Xbit_r14_c55 bl_55 br_55 wl_14 vdd gnd cell_6t
Xbit_r15_c55 bl_55 br_55 wl_15 vdd gnd cell_6t
Xbit_r16_c55 bl_55 br_55 wl_16 vdd gnd cell_6t
Xbit_r17_c55 bl_55 br_55 wl_17 vdd gnd cell_6t
Xbit_r18_c55 bl_55 br_55 wl_18 vdd gnd cell_6t
Xbit_r19_c55 bl_55 br_55 wl_19 vdd gnd cell_6t
Xbit_r20_c55 bl_55 br_55 wl_20 vdd gnd cell_6t
Xbit_r21_c55 bl_55 br_55 wl_21 vdd gnd cell_6t
Xbit_r22_c55 bl_55 br_55 wl_22 vdd gnd cell_6t
Xbit_r23_c55 bl_55 br_55 wl_23 vdd gnd cell_6t
Xbit_r24_c55 bl_55 br_55 wl_24 vdd gnd cell_6t
Xbit_r25_c55 bl_55 br_55 wl_25 vdd gnd cell_6t
Xbit_r26_c55 bl_55 br_55 wl_26 vdd gnd cell_6t
Xbit_r27_c55 bl_55 br_55 wl_27 vdd gnd cell_6t
Xbit_r28_c55 bl_55 br_55 wl_28 vdd gnd cell_6t
Xbit_r29_c55 bl_55 br_55 wl_29 vdd gnd cell_6t
Xbit_r30_c55 bl_55 br_55 wl_30 vdd gnd cell_6t
Xbit_r31_c55 bl_55 br_55 wl_31 vdd gnd cell_6t
Xbit_r32_c55 bl_55 br_55 wl_32 vdd gnd cell_6t
Xbit_r33_c55 bl_55 br_55 wl_33 vdd gnd cell_6t
Xbit_r34_c55 bl_55 br_55 wl_34 vdd gnd cell_6t
Xbit_r35_c55 bl_55 br_55 wl_35 vdd gnd cell_6t
Xbit_r36_c55 bl_55 br_55 wl_36 vdd gnd cell_6t
Xbit_r37_c55 bl_55 br_55 wl_37 vdd gnd cell_6t
Xbit_r38_c55 bl_55 br_55 wl_38 vdd gnd cell_6t
Xbit_r39_c55 bl_55 br_55 wl_39 vdd gnd cell_6t
Xbit_r40_c55 bl_55 br_55 wl_40 vdd gnd cell_6t
Xbit_r41_c55 bl_55 br_55 wl_41 vdd gnd cell_6t
Xbit_r42_c55 bl_55 br_55 wl_42 vdd gnd cell_6t
Xbit_r43_c55 bl_55 br_55 wl_43 vdd gnd cell_6t
Xbit_r44_c55 bl_55 br_55 wl_44 vdd gnd cell_6t
Xbit_r45_c55 bl_55 br_55 wl_45 vdd gnd cell_6t
Xbit_r46_c55 bl_55 br_55 wl_46 vdd gnd cell_6t
Xbit_r47_c55 bl_55 br_55 wl_47 vdd gnd cell_6t
Xbit_r48_c55 bl_55 br_55 wl_48 vdd gnd cell_6t
Xbit_r49_c55 bl_55 br_55 wl_49 vdd gnd cell_6t
Xbit_r50_c55 bl_55 br_55 wl_50 vdd gnd cell_6t
Xbit_r51_c55 bl_55 br_55 wl_51 vdd gnd cell_6t
Xbit_r52_c55 bl_55 br_55 wl_52 vdd gnd cell_6t
Xbit_r53_c55 bl_55 br_55 wl_53 vdd gnd cell_6t
Xbit_r54_c55 bl_55 br_55 wl_54 vdd gnd cell_6t
Xbit_r55_c55 bl_55 br_55 wl_55 vdd gnd cell_6t
Xbit_r56_c55 bl_55 br_55 wl_56 vdd gnd cell_6t
Xbit_r57_c55 bl_55 br_55 wl_57 vdd gnd cell_6t
Xbit_r58_c55 bl_55 br_55 wl_58 vdd gnd cell_6t
Xbit_r59_c55 bl_55 br_55 wl_59 vdd gnd cell_6t
Xbit_r60_c55 bl_55 br_55 wl_60 vdd gnd cell_6t
Xbit_r61_c55 bl_55 br_55 wl_61 vdd gnd cell_6t
Xbit_r62_c55 bl_55 br_55 wl_62 vdd gnd cell_6t
Xbit_r63_c55 bl_55 br_55 wl_63 vdd gnd cell_6t
Xbit_r64_c55 bl_55 br_55 wl_64 vdd gnd cell_6t
Xbit_r65_c55 bl_55 br_55 wl_65 vdd gnd cell_6t
Xbit_r66_c55 bl_55 br_55 wl_66 vdd gnd cell_6t
Xbit_r67_c55 bl_55 br_55 wl_67 vdd gnd cell_6t
Xbit_r68_c55 bl_55 br_55 wl_68 vdd gnd cell_6t
Xbit_r69_c55 bl_55 br_55 wl_69 vdd gnd cell_6t
Xbit_r70_c55 bl_55 br_55 wl_70 vdd gnd cell_6t
Xbit_r71_c55 bl_55 br_55 wl_71 vdd gnd cell_6t
Xbit_r72_c55 bl_55 br_55 wl_72 vdd gnd cell_6t
Xbit_r73_c55 bl_55 br_55 wl_73 vdd gnd cell_6t
Xbit_r74_c55 bl_55 br_55 wl_74 vdd gnd cell_6t
Xbit_r75_c55 bl_55 br_55 wl_75 vdd gnd cell_6t
Xbit_r76_c55 bl_55 br_55 wl_76 vdd gnd cell_6t
Xbit_r77_c55 bl_55 br_55 wl_77 vdd gnd cell_6t
Xbit_r78_c55 bl_55 br_55 wl_78 vdd gnd cell_6t
Xbit_r79_c55 bl_55 br_55 wl_79 vdd gnd cell_6t
Xbit_r80_c55 bl_55 br_55 wl_80 vdd gnd cell_6t
Xbit_r81_c55 bl_55 br_55 wl_81 vdd gnd cell_6t
Xbit_r82_c55 bl_55 br_55 wl_82 vdd gnd cell_6t
Xbit_r83_c55 bl_55 br_55 wl_83 vdd gnd cell_6t
Xbit_r84_c55 bl_55 br_55 wl_84 vdd gnd cell_6t
Xbit_r85_c55 bl_55 br_55 wl_85 vdd gnd cell_6t
Xbit_r86_c55 bl_55 br_55 wl_86 vdd gnd cell_6t
Xbit_r87_c55 bl_55 br_55 wl_87 vdd gnd cell_6t
Xbit_r88_c55 bl_55 br_55 wl_88 vdd gnd cell_6t
Xbit_r89_c55 bl_55 br_55 wl_89 vdd gnd cell_6t
Xbit_r90_c55 bl_55 br_55 wl_90 vdd gnd cell_6t
Xbit_r91_c55 bl_55 br_55 wl_91 vdd gnd cell_6t
Xbit_r92_c55 bl_55 br_55 wl_92 vdd gnd cell_6t
Xbit_r93_c55 bl_55 br_55 wl_93 vdd gnd cell_6t
Xbit_r94_c55 bl_55 br_55 wl_94 vdd gnd cell_6t
Xbit_r95_c55 bl_55 br_55 wl_95 vdd gnd cell_6t
Xbit_r96_c55 bl_55 br_55 wl_96 vdd gnd cell_6t
Xbit_r97_c55 bl_55 br_55 wl_97 vdd gnd cell_6t
Xbit_r98_c55 bl_55 br_55 wl_98 vdd gnd cell_6t
Xbit_r99_c55 bl_55 br_55 wl_99 vdd gnd cell_6t
Xbit_r100_c55 bl_55 br_55 wl_100 vdd gnd cell_6t
Xbit_r101_c55 bl_55 br_55 wl_101 vdd gnd cell_6t
Xbit_r102_c55 bl_55 br_55 wl_102 vdd gnd cell_6t
Xbit_r103_c55 bl_55 br_55 wl_103 vdd gnd cell_6t
Xbit_r104_c55 bl_55 br_55 wl_104 vdd gnd cell_6t
Xbit_r105_c55 bl_55 br_55 wl_105 vdd gnd cell_6t
Xbit_r106_c55 bl_55 br_55 wl_106 vdd gnd cell_6t
Xbit_r107_c55 bl_55 br_55 wl_107 vdd gnd cell_6t
Xbit_r108_c55 bl_55 br_55 wl_108 vdd gnd cell_6t
Xbit_r109_c55 bl_55 br_55 wl_109 vdd gnd cell_6t
Xbit_r110_c55 bl_55 br_55 wl_110 vdd gnd cell_6t
Xbit_r111_c55 bl_55 br_55 wl_111 vdd gnd cell_6t
Xbit_r112_c55 bl_55 br_55 wl_112 vdd gnd cell_6t
Xbit_r113_c55 bl_55 br_55 wl_113 vdd gnd cell_6t
Xbit_r114_c55 bl_55 br_55 wl_114 vdd gnd cell_6t
Xbit_r115_c55 bl_55 br_55 wl_115 vdd gnd cell_6t
Xbit_r116_c55 bl_55 br_55 wl_116 vdd gnd cell_6t
Xbit_r117_c55 bl_55 br_55 wl_117 vdd gnd cell_6t
Xbit_r118_c55 bl_55 br_55 wl_118 vdd gnd cell_6t
Xbit_r119_c55 bl_55 br_55 wl_119 vdd gnd cell_6t
Xbit_r120_c55 bl_55 br_55 wl_120 vdd gnd cell_6t
Xbit_r121_c55 bl_55 br_55 wl_121 vdd gnd cell_6t
Xbit_r122_c55 bl_55 br_55 wl_122 vdd gnd cell_6t
Xbit_r123_c55 bl_55 br_55 wl_123 vdd gnd cell_6t
Xbit_r124_c55 bl_55 br_55 wl_124 vdd gnd cell_6t
Xbit_r125_c55 bl_55 br_55 wl_125 vdd gnd cell_6t
Xbit_r126_c55 bl_55 br_55 wl_126 vdd gnd cell_6t
Xbit_r127_c55 bl_55 br_55 wl_127 vdd gnd cell_6t
Xbit_r128_c55 bl_55 br_55 wl_128 vdd gnd cell_6t
Xbit_r129_c55 bl_55 br_55 wl_129 vdd gnd cell_6t
Xbit_r130_c55 bl_55 br_55 wl_130 vdd gnd cell_6t
Xbit_r131_c55 bl_55 br_55 wl_131 vdd gnd cell_6t
Xbit_r132_c55 bl_55 br_55 wl_132 vdd gnd cell_6t
Xbit_r133_c55 bl_55 br_55 wl_133 vdd gnd cell_6t
Xbit_r134_c55 bl_55 br_55 wl_134 vdd gnd cell_6t
Xbit_r135_c55 bl_55 br_55 wl_135 vdd gnd cell_6t
Xbit_r136_c55 bl_55 br_55 wl_136 vdd gnd cell_6t
Xbit_r137_c55 bl_55 br_55 wl_137 vdd gnd cell_6t
Xbit_r138_c55 bl_55 br_55 wl_138 vdd gnd cell_6t
Xbit_r139_c55 bl_55 br_55 wl_139 vdd gnd cell_6t
Xbit_r140_c55 bl_55 br_55 wl_140 vdd gnd cell_6t
Xbit_r141_c55 bl_55 br_55 wl_141 vdd gnd cell_6t
Xbit_r142_c55 bl_55 br_55 wl_142 vdd gnd cell_6t
Xbit_r143_c55 bl_55 br_55 wl_143 vdd gnd cell_6t
Xbit_r144_c55 bl_55 br_55 wl_144 vdd gnd cell_6t
Xbit_r145_c55 bl_55 br_55 wl_145 vdd gnd cell_6t
Xbit_r146_c55 bl_55 br_55 wl_146 vdd gnd cell_6t
Xbit_r147_c55 bl_55 br_55 wl_147 vdd gnd cell_6t
Xbit_r148_c55 bl_55 br_55 wl_148 vdd gnd cell_6t
Xbit_r149_c55 bl_55 br_55 wl_149 vdd gnd cell_6t
Xbit_r150_c55 bl_55 br_55 wl_150 vdd gnd cell_6t
Xbit_r151_c55 bl_55 br_55 wl_151 vdd gnd cell_6t
Xbit_r152_c55 bl_55 br_55 wl_152 vdd gnd cell_6t
Xbit_r153_c55 bl_55 br_55 wl_153 vdd gnd cell_6t
Xbit_r154_c55 bl_55 br_55 wl_154 vdd gnd cell_6t
Xbit_r155_c55 bl_55 br_55 wl_155 vdd gnd cell_6t
Xbit_r156_c55 bl_55 br_55 wl_156 vdd gnd cell_6t
Xbit_r157_c55 bl_55 br_55 wl_157 vdd gnd cell_6t
Xbit_r158_c55 bl_55 br_55 wl_158 vdd gnd cell_6t
Xbit_r159_c55 bl_55 br_55 wl_159 vdd gnd cell_6t
Xbit_r160_c55 bl_55 br_55 wl_160 vdd gnd cell_6t
Xbit_r161_c55 bl_55 br_55 wl_161 vdd gnd cell_6t
Xbit_r162_c55 bl_55 br_55 wl_162 vdd gnd cell_6t
Xbit_r163_c55 bl_55 br_55 wl_163 vdd gnd cell_6t
Xbit_r164_c55 bl_55 br_55 wl_164 vdd gnd cell_6t
Xbit_r165_c55 bl_55 br_55 wl_165 vdd gnd cell_6t
Xbit_r166_c55 bl_55 br_55 wl_166 vdd gnd cell_6t
Xbit_r167_c55 bl_55 br_55 wl_167 vdd gnd cell_6t
Xbit_r168_c55 bl_55 br_55 wl_168 vdd gnd cell_6t
Xbit_r169_c55 bl_55 br_55 wl_169 vdd gnd cell_6t
Xbit_r170_c55 bl_55 br_55 wl_170 vdd gnd cell_6t
Xbit_r171_c55 bl_55 br_55 wl_171 vdd gnd cell_6t
Xbit_r172_c55 bl_55 br_55 wl_172 vdd gnd cell_6t
Xbit_r173_c55 bl_55 br_55 wl_173 vdd gnd cell_6t
Xbit_r174_c55 bl_55 br_55 wl_174 vdd gnd cell_6t
Xbit_r175_c55 bl_55 br_55 wl_175 vdd gnd cell_6t
Xbit_r176_c55 bl_55 br_55 wl_176 vdd gnd cell_6t
Xbit_r177_c55 bl_55 br_55 wl_177 vdd gnd cell_6t
Xbit_r178_c55 bl_55 br_55 wl_178 vdd gnd cell_6t
Xbit_r179_c55 bl_55 br_55 wl_179 vdd gnd cell_6t
Xbit_r180_c55 bl_55 br_55 wl_180 vdd gnd cell_6t
Xbit_r181_c55 bl_55 br_55 wl_181 vdd gnd cell_6t
Xbit_r182_c55 bl_55 br_55 wl_182 vdd gnd cell_6t
Xbit_r183_c55 bl_55 br_55 wl_183 vdd gnd cell_6t
Xbit_r184_c55 bl_55 br_55 wl_184 vdd gnd cell_6t
Xbit_r185_c55 bl_55 br_55 wl_185 vdd gnd cell_6t
Xbit_r186_c55 bl_55 br_55 wl_186 vdd gnd cell_6t
Xbit_r187_c55 bl_55 br_55 wl_187 vdd gnd cell_6t
Xbit_r188_c55 bl_55 br_55 wl_188 vdd gnd cell_6t
Xbit_r189_c55 bl_55 br_55 wl_189 vdd gnd cell_6t
Xbit_r190_c55 bl_55 br_55 wl_190 vdd gnd cell_6t
Xbit_r191_c55 bl_55 br_55 wl_191 vdd gnd cell_6t
Xbit_r192_c55 bl_55 br_55 wl_192 vdd gnd cell_6t
Xbit_r193_c55 bl_55 br_55 wl_193 vdd gnd cell_6t
Xbit_r194_c55 bl_55 br_55 wl_194 vdd gnd cell_6t
Xbit_r195_c55 bl_55 br_55 wl_195 vdd gnd cell_6t
Xbit_r196_c55 bl_55 br_55 wl_196 vdd gnd cell_6t
Xbit_r197_c55 bl_55 br_55 wl_197 vdd gnd cell_6t
Xbit_r198_c55 bl_55 br_55 wl_198 vdd gnd cell_6t
Xbit_r199_c55 bl_55 br_55 wl_199 vdd gnd cell_6t
Xbit_r200_c55 bl_55 br_55 wl_200 vdd gnd cell_6t
Xbit_r201_c55 bl_55 br_55 wl_201 vdd gnd cell_6t
Xbit_r202_c55 bl_55 br_55 wl_202 vdd gnd cell_6t
Xbit_r203_c55 bl_55 br_55 wl_203 vdd gnd cell_6t
Xbit_r204_c55 bl_55 br_55 wl_204 vdd gnd cell_6t
Xbit_r205_c55 bl_55 br_55 wl_205 vdd gnd cell_6t
Xbit_r206_c55 bl_55 br_55 wl_206 vdd gnd cell_6t
Xbit_r207_c55 bl_55 br_55 wl_207 vdd gnd cell_6t
Xbit_r208_c55 bl_55 br_55 wl_208 vdd gnd cell_6t
Xbit_r209_c55 bl_55 br_55 wl_209 vdd gnd cell_6t
Xbit_r210_c55 bl_55 br_55 wl_210 vdd gnd cell_6t
Xbit_r211_c55 bl_55 br_55 wl_211 vdd gnd cell_6t
Xbit_r212_c55 bl_55 br_55 wl_212 vdd gnd cell_6t
Xbit_r213_c55 bl_55 br_55 wl_213 vdd gnd cell_6t
Xbit_r214_c55 bl_55 br_55 wl_214 vdd gnd cell_6t
Xbit_r215_c55 bl_55 br_55 wl_215 vdd gnd cell_6t
Xbit_r216_c55 bl_55 br_55 wl_216 vdd gnd cell_6t
Xbit_r217_c55 bl_55 br_55 wl_217 vdd gnd cell_6t
Xbit_r218_c55 bl_55 br_55 wl_218 vdd gnd cell_6t
Xbit_r219_c55 bl_55 br_55 wl_219 vdd gnd cell_6t
Xbit_r220_c55 bl_55 br_55 wl_220 vdd gnd cell_6t
Xbit_r221_c55 bl_55 br_55 wl_221 vdd gnd cell_6t
Xbit_r222_c55 bl_55 br_55 wl_222 vdd gnd cell_6t
Xbit_r223_c55 bl_55 br_55 wl_223 vdd gnd cell_6t
Xbit_r224_c55 bl_55 br_55 wl_224 vdd gnd cell_6t
Xbit_r225_c55 bl_55 br_55 wl_225 vdd gnd cell_6t
Xbit_r226_c55 bl_55 br_55 wl_226 vdd gnd cell_6t
Xbit_r227_c55 bl_55 br_55 wl_227 vdd gnd cell_6t
Xbit_r228_c55 bl_55 br_55 wl_228 vdd gnd cell_6t
Xbit_r229_c55 bl_55 br_55 wl_229 vdd gnd cell_6t
Xbit_r230_c55 bl_55 br_55 wl_230 vdd gnd cell_6t
Xbit_r231_c55 bl_55 br_55 wl_231 vdd gnd cell_6t
Xbit_r232_c55 bl_55 br_55 wl_232 vdd gnd cell_6t
Xbit_r233_c55 bl_55 br_55 wl_233 vdd gnd cell_6t
Xbit_r234_c55 bl_55 br_55 wl_234 vdd gnd cell_6t
Xbit_r235_c55 bl_55 br_55 wl_235 vdd gnd cell_6t
Xbit_r236_c55 bl_55 br_55 wl_236 vdd gnd cell_6t
Xbit_r237_c55 bl_55 br_55 wl_237 vdd gnd cell_6t
Xbit_r238_c55 bl_55 br_55 wl_238 vdd gnd cell_6t
Xbit_r239_c55 bl_55 br_55 wl_239 vdd gnd cell_6t
Xbit_r240_c55 bl_55 br_55 wl_240 vdd gnd cell_6t
Xbit_r241_c55 bl_55 br_55 wl_241 vdd gnd cell_6t
Xbit_r242_c55 bl_55 br_55 wl_242 vdd gnd cell_6t
Xbit_r243_c55 bl_55 br_55 wl_243 vdd gnd cell_6t
Xbit_r244_c55 bl_55 br_55 wl_244 vdd gnd cell_6t
Xbit_r245_c55 bl_55 br_55 wl_245 vdd gnd cell_6t
Xbit_r246_c55 bl_55 br_55 wl_246 vdd gnd cell_6t
Xbit_r247_c55 bl_55 br_55 wl_247 vdd gnd cell_6t
Xbit_r248_c55 bl_55 br_55 wl_248 vdd gnd cell_6t
Xbit_r249_c55 bl_55 br_55 wl_249 vdd gnd cell_6t
Xbit_r250_c55 bl_55 br_55 wl_250 vdd gnd cell_6t
Xbit_r251_c55 bl_55 br_55 wl_251 vdd gnd cell_6t
Xbit_r252_c55 bl_55 br_55 wl_252 vdd gnd cell_6t
Xbit_r253_c55 bl_55 br_55 wl_253 vdd gnd cell_6t
Xbit_r254_c55 bl_55 br_55 wl_254 vdd gnd cell_6t
Xbit_r255_c55 bl_55 br_55 wl_255 vdd gnd cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd cell_6t
Xbit_r1_c56 bl_56 br_56 wl_1 vdd gnd cell_6t
Xbit_r2_c56 bl_56 br_56 wl_2 vdd gnd cell_6t
Xbit_r3_c56 bl_56 br_56 wl_3 vdd gnd cell_6t
Xbit_r4_c56 bl_56 br_56 wl_4 vdd gnd cell_6t
Xbit_r5_c56 bl_56 br_56 wl_5 vdd gnd cell_6t
Xbit_r6_c56 bl_56 br_56 wl_6 vdd gnd cell_6t
Xbit_r7_c56 bl_56 br_56 wl_7 vdd gnd cell_6t
Xbit_r8_c56 bl_56 br_56 wl_8 vdd gnd cell_6t
Xbit_r9_c56 bl_56 br_56 wl_9 vdd gnd cell_6t
Xbit_r10_c56 bl_56 br_56 wl_10 vdd gnd cell_6t
Xbit_r11_c56 bl_56 br_56 wl_11 vdd gnd cell_6t
Xbit_r12_c56 bl_56 br_56 wl_12 vdd gnd cell_6t
Xbit_r13_c56 bl_56 br_56 wl_13 vdd gnd cell_6t
Xbit_r14_c56 bl_56 br_56 wl_14 vdd gnd cell_6t
Xbit_r15_c56 bl_56 br_56 wl_15 vdd gnd cell_6t
Xbit_r16_c56 bl_56 br_56 wl_16 vdd gnd cell_6t
Xbit_r17_c56 bl_56 br_56 wl_17 vdd gnd cell_6t
Xbit_r18_c56 bl_56 br_56 wl_18 vdd gnd cell_6t
Xbit_r19_c56 bl_56 br_56 wl_19 vdd gnd cell_6t
Xbit_r20_c56 bl_56 br_56 wl_20 vdd gnd cell_6t
Xbit_r21_c56 bl_56 br_56 wl_21 vdd gnd cell_6t
Xbit_r22_c56 bl_56 br_56 wl_22 vdd gnd cell_6t
Xbit_r23_c56 bl_56 br_56 wl_23 vdd gnd cell_6t
Xbit_r24_c56 bl_56 br_56 wl_24 vdd gnd cell_6t
Xbit_r25_c56 bl_56 br_56 wl_25 vdd gnd cell_6t
Xbit_r26_c56 bl_56 br_56 wl_26 vdd gnd cell_6t
Xbit_r27_c56 bl_56 br_56 wl_27 vdd gnd cell_6t
Xbit_r28_c56 bl_56 br_56 wl_28 vdd gnd cell_6t
Xbit_r29_c56 bl_56 br_56 wl_29 vdd gnd cell_6t
Xbit_r30_c56 bl_56 br_56 wl_30 vdd gnd cell_6t
Xbit_r31_c56 bl_56 br_56 wl_31 vdd gnd cell_6t
Xbit_r32_c56 bl_56 br_56 wl_32 vdd gnd cell_6t
Xbit_r33_c56 bl_56 br_56 wl_33 vdd gnd cell_6t
Xbit_r34_c56 bl_56 br_56 wl_34 vdd gnd cell_6t
Xbit_r35_c56 bl_56 br_56 wl_35 vdd gnd cell_6t
Xbit_r36_c56 bl_56 br_56 wl_36 vdd gnd cell_6t
Xbit_r37_c56 bl_56 br_56 wl_37 vdd gnd cell_6t
Xbit_r38_c56 bl_56 br_56 wl_38 vdd gnd cell_6t
Xbit_r39_c56 bl_56 br_56 wl_39 vdd gnd cell_6t
Xbit_r40_c56 bl_56 br_56 wl_40 vdd gnd cell_6t
Xbit_r41_c56 bl_56 br_56 wl_41 vdd gnd cell_6t
Xbit_r42_c56 bl_56 br_56 wl_42 vdd gnd cell_6t
Xbit_r43_c56 bl_56 br_56 wl_43 vdd gnd cell_6t
Xbit_r44_c56 bl_56 br_56 wl_44 vdd gnd cell_6t
Xbit_r45_c56 bl_56 br_56 wl_45 vdd gnd cell_6t
Xbit_r46_c56 bl_56 br_56 wl_46 vdd gnd cell_6t
Xbit_r47_c56 bl_56 br_56 wl_47 vdd gnd cell_6t
Xbit_r48_c56 bl_56 br_56 wl_48 vdd gnd cell_6t
Xbit_r49_c56 bl_56 br_56 wl_49 vdd gnd cell_6t
Xbit_r50_c56 bl_56 br_56 wl_50 vdd gnd cell_6t
Xbit_r51_c56 bl_56 br_56 wl_51 vdd gnd cell_6t
Xbit_r52_c56 bl_56 br_56 wl_52 vdd gnd cell_6t
Xbit_r53_c56 bl_56 br_56 wl_53 vdd gnd cell_6t
Xbit_r54_c56 bl_56 br_56 wl_54 vdd gnd cell_6t
Xbit_r55_c56 bl_56 br_56 wl_55 vdd gnd cell_6t
Xbit_r56_c56 bl_56 br_56 wl_56 vdd gnd cell_6t
Xbit_r57_c56 bl_56 br_56 wl_57 vdd gnd cell_6t
Xbit_r58_c56 bl_56 br_56 wl_58 vdd gnd cell_6t
Xbit_r59_c56 bl_56 br_56 wl_59 vdd gnd cell_6t
Xbit_r60_c56 bl_56 br_56 wl_60 vdd gnd cell_6t
Xbit_r61_c56 bl_56 br_56 wl_61 vdd gnd cell_6t
Xbit_r62_c56 bl_56 br_56 wl_62 vdd gnd cell_6t
Xbit_r63_c56 bl_56 br_56 wl_63 vdd gnd cell_6t
Xbit_r64_c56 bl_56 br_56 wl_64 vdd gnd cell_6t
Xbit_r65_c56 bl_56 br_56 wl_65 vdd gnd cell_6t
Xbit_r66_c56 bl_56 br_56 wl_66 vdd gnd cell_6t
Xbit_r67_c56 bl_56 br_56 wl_67 vdd gnd cell_6t
Xbit_r68_c56 bl_56 br_56 wl_68 vdd gnd cell_6t
Xbit_r69_c56 bl_56 br_56 wl_69 vdd gnd cell_6t
Xbit_r70_c56 bl_56 br_56 wl_70 vdd gnd cell_6t
Xbit_r71_c56 bl_56 br_56 wl_71 vdd gnd cell_6t
Xbit_r72_c56 bl_56 br_56 wl_72 vdd gnd cell_6t
Xbit_r73_c56 bl_56 br_56 wl_73 vdd gnd cell_6t
Xbit_r74_c56 bl_56 br_56 wl_74 vdd gnd cell_6t
Xbit_r75_c56 bl_56 br_56 wl_75 vdd gnd cell_6t
Xbit_r76_c56 bl_56 br_56 wl_76 vdd gnd cell_6t
Xbit_r77_c56 bl_56 br_56 wl_77 vdd gnd cell_6t
Xbit_r78_c56 bl_56 br_56 wl_78 vdd gnd cell_6t
Xbit_r79_c56 bl_56 br_56 wl_79 vdd gnd cell_6t
Xbit_r80_c56 bl_56 br_56 wl_80 vdd gnd cell_6t
Xbit_r81_c56 bl_56 br_56 wl_81 vdd gnd cell_6t
Xbit_r82_c56 bl_56 br_56 wl_82 vdd gnd cell_6t
Xbit_r83_c56 bl_56 br_56 wl_83 vdd gnd cell_6t
Xbit_r84_c56 bl_56 br_56 wl_84 vdd gnd cell_6t
Xbit_r85_c56 bl_56 br_56 wl_85 vdd gnd cell_6t
Xbit_r86_c56 bl_56 br_56 wl_86 vdd gnd cell_6t
Xbit_r87_c56 bl_56 br_56 wl_87 vdd gnd cell_6t
Xbit_r88_c56 bl_56 br_56 wl_88 vdd gnd cell_6t
Xbit_r89_c56 bl_56 br_56 wl_89 vdd gnd cell_6t
Xbit_r90_c56 bl_56 br_56 wl_90 vdd gnd cell_6t
Xbit_r91_c56 bl_56 br_56 wl_91 vdd gnd cell_6t
Xbit_r92_c56 bl_56 br_56 wl_92 vdd gnd cell_6t
Xbit_r93_c56 bl_56 br_56 wl_93 vdd gnd cell_6t
Xbit_r94_c56 bl_56 br_56 wl_94 vdd gnd cell_6t
Xbit_r95_c56 bl_56 br_56 wl_95 vdd gnd cell_6t
Xbit_r96_c56 bl_56 br_56 wl_96 vdd gnd cell_6t
Xbit_r97_c56 bl_56 br_56 wl_97 vdd gnd cell_6t
Xbit_r98_c56 bl_56 br_56 wl_98 vdd gnd cell_6t
Xbit_r99_c56 bl_56 br_56 wl_99 vdd gnd cell_6t
Xbit_r100_c56 bl_56 br_56 wl_100 vdd gnd cell_6t
Xbit_r101_c56 bl_56 br_56 wl_101 vdd gnd cell_6t
Xbit_r102_c56 bl_56 br_56 wl_102 vdd gnd cell_6t
Xbit_r103_c56 bl_56 br_56 wl_103 vdd gnd cell_6t
Xbit_r104_c56 bl_56 br_56 wl_104 vdd gnd cell_6t
Xbit_r105_c56 bl_56 br_56 wl_105 vdd gnd cell_6t
Xbit_r106_c56 bl_56 br_56 wl_106 vdd gnd cell_6t
Xbit_r107_c56 bl_56 br_56 wl_107 vdd gnd cell_6t
Xbit_r108_c56 bl_56 br_56 wl_108 vdd gnd cell_6t
Xbit_r109_c56 bl_56 br_56 wl_109 vdd gnd cell_6t
Xbit_r110_c56 bl_56 br_56 wl_110 vdd gnd cell_6t
Xbit_r111_c56 bl_56 br_56 wl_111 vdd gnd cell_6t
Xbit_r112_c56 bl_56 br_56 wl_112 vdd gnd cell_6t
Xbit_r113_c56 bl_56 br_56 wl_113 vdd gnd cell_6t
Xbit_r114_c56 bl_56 br_56 wl_114 vdd gnd cell_6t
Xbit_r115_c56 bl_56 br_56 wl_115 vdd gnd cell_6t
Xbit_r116_c56 bl_56 br_56 wl_116 vdd gnd cell_6t
Xbit_r117_c56 bl_56 br_56 wl_117 vdd gnd cell_6t
Xbit_r118_c56 bl_56 br_56 wl_118 vdd gnd cell_6t
Xbit_r119_c56 bl_56 br_56 wl_119 vdd gnd cell_6t
Xbit_r120_c56 bl_56 br_56 wl_120 vdd gnd cell_6t
Xbit_r121_c56 bl_56 br_56 wl_121 vdd gnd cell_6t
Xbit_r122_c56 bl_56 br_56 wl_122 vdd gnd cell_6t
Xbit_r123_c56 bl_56 br_56 wl_123 vdd gnd cell_6t
Xbit_r124_c56 bl_56 br_56 wl_124 vdd gnd cell_6t
Xbit_r125_c56 bl_56 br_56 wl_125 vdd gnd cell_6t
Xbit_r126_c56 bl_56 br_56 wl_126 vdd gnd cell_6t
Xbit_r127_c56 bl_56 br_56 wl_127 vdd gnd cell_6t
Xbit_r128_c56 bl_56 br_56 wl_128 vdd gnd cell_6t
Xbit_r129_c56 bl_56 br_56 wl_129 vdd gnd cell_6t
Xbit_r130_c56 bl_56 br_56 wl_130 vdd gnd cell_6t
Xbit_r131_c56 bl_56 br_56 wl_131 vdd gnd cell_6t
Xbit_r132_c56 bl_56 br_56 wl_132 vdd gnd cell_6t
Xbit_r133_c56 bl_56 br_56 wl_133 vdd gnd cell_6t
Xbit_r134_c56 bl_56 br_56 wl_134 vdd gnd cell_6t
Xbit_r135_c56 bl_56 br_56 wl_135 vdd gnd cell_6t
Xbit_r136_c56 bl_56 br_56 wl_136 vdd gnd cell_6t
Xbit_r137_c56 bl_56 br_56 wl_137 vdd gnd cell_6t
Xbit_r138_c56 bl_56 br_56 wl_138 vdd gnd cell_6t
Xbit_r139_c56 bl_56 br_56 wl_139 vdd gnd cell_6t
Xbit_r140_c56 bl_56 br_56 wl_140 vdd gnd cell_6t
Xbit_r141_c56 bl_56 br_56 wl_141 vdd gnd cell_6t
Xbit_r142_c56 bl_56 br_56 wl_142 vdd gnd cell_6t
Xbit_r143_c56 bl_56 br_56 wl_143 vdd gnd cell_6t
Xbit_r144_c56 bl_56 br_56 wl_144 vdd gnd cell_6t
Xbit_r145_c56 bl_56 br_56 wl_145 vdd gnd cell_6t
Xbit_r146_c56 bl_56 br_56 wl_146 vdd gnd cell_6t
Xbit_r147_c56 bl_56 br_56 wl_147 vdd gnd cell_6t
Xbit_r148_c56 bl_56 br_56 wl_148 vdd gnd cell_6t
Xbit_r149_c56 bl_56 br_56 wl_149 vdd gnd cell_6t
Xbit_r150_c56 bl_56 br_56 wl_150 vdd gnd cell_6t
Xbit_r151_c56 bl_56 br_56 wl_151 vdd gnd cell_6t
Xbit_r152_c56 bl_56 br_56 wl_152 vdd gnd cell_6t
Xbit_r153_c56 bl_56 br_56 wl_153 vdd gnd cell_6t
Xbit_r154_c56 bl_56 br_56 wl_154 vdd gnd cell_6t
Xbit_r155_c56 bl_56 br_56 wl_155 vdd gnd cell_6t
Xbit_r156_c56 bl_56 br_56 wl_156 vdd gnd cell_6t
Xbit_r157_c56 bl_56 br_56 wl_157 vdd gnd cell_6t
Xbit_r158_c56 bl_56 br_56 wl_158 vdd gnd cell_6t
Xbit_r159_c56 bl_56 br_56 wl_159 vdd gnd cell_6t
Xbit_r160_c56 bl_56 br_56 wl_160 vdd gnd cell_6t
Xbit_r161_c56 bl_56 br_56 wl_161 vdd gnd cell_6t
Xbit_r162_c56 bl_56 br_56 wl_162 vdd gnd cell_6t
Xbit_r163_c56 bl_56 br_56 wl_163 vdd gnd cell_6t
Xbit_r164_c56 bl_56 br_56 wl_164 vdd gnd cell_6t
Xbit_r165_c56 bl_56 br_56 wl_165 vdd gnd cell_6t
Xbit_r166_c56 bl_56 br_56 wl_166 vdd gnd cell_6t
Xbit_r167_c56 bl_56 br_56 wl_167 vdd gnd cell_6t
Xbit_r168_c56 bl_56 br_56 wl_168 vdd gnd cell_6t
Xbit_r169_c56 bl_56 br_56 wl_169 vdd gnd cell_6t
Xbit_r170_c56 bl_56 br_56 wl_170 vdd gnd cell_6t
Xbit_r171_c56 bl_56 br_56 wl_171 vdd gnd cell_6t
Xbit_r172_c56 bl_56 br_56 wl_172 vdd gnd cell_6t
Xbit_r173_c56 bl_56 br_56 wl_173 vdd gnd cell_6t
Xbit_r174_c56 bl_56 br_56 wl_174 vdd gnd cell_6t
Xbit_r175_c56 bl_56 br_56 wl_175 vdd gnd cell_6t
Xbit_r176_c56 bl_56 br_56 wl_176 vdd gnd cell_6t
Xbit_r177_c56 bl_56 br_56 wl_177 vdd gnd cell_6t
Xbit_r178_c56 bl_56 br_56 wl_178 vdd gnd cell_6t
Xbit_r179_c56 bl_56 br_56 wl_179 vdd gnd cell_6t
Xbit_r180_c56 bl_56 br_56 wl_180 vdd gnd cell_6t
Xbit_r181_c56 bl_56 br_56 wl_181 vdd gnd cell_6t
Xbit_r182_c56 bl_56 br_56 wl_182 vdd gnd cell_6t
Xbit_r183_c56 bl_56 br_56 wl_183 vdd gnd cell_6t
Xbit_r184_c56 bl_56 br_56 wl_184 vdd gnd cell_6t
Xbit_r185_c56 bl_56 br_56 wl_185 vdd gnd cell_6t
Xbit_r186_c56 bl_56 br_56 wl_186 vdd gnd cell_6t
Xbit_r187_c56 bl_56 br_56 wl_187 vdd gnd cell_6t
Xbit_r188_c56 bl_56 br_56 wl_188 vdd gnd cell_6t
Xbit_r189_c56 bl_56 br_56 wl_189 vdd gnd cell_6t
Xbit_r190_c56 bl_56 br_56 wl_190 vdd gnd cell_6t
Xbit_r191_c56 bl_56 br_56 wl_191 vdd gnd cell_6t
Xbit_r192_c56 bl_56 br_56 wl_192 vdd gnd cell_6t
Xbit_r193_c56 bl_56 br_56 wl_193 vdd gnd cell_6t
Xbit_r194_c56 bl_56 br_56 wl_194 vdd gnd cell_6t
Xbit_r195_c56 bl_56 br_56 wl_195 vdd gnd cell_6t
Xbit_r196_c56 bl_56 br_56 wl_196 vdd gnd cell_6t
Xbit_r197_c56 bl_56 br_56 wl_197 vdd gnd cell_6t
Xbit_r198_c56 bl_56 br_56 wl_198 vdd gnd cell_6t
Xbit_r199_c56 bl_56 br_56 wl_199 vdd gnd cell_6t
Xbit_r200_c56 bl_56 br_56 wl_200 vdd gnd cell_6t
Xbit_r201_c56 bl_56 br_56 wl_201 vdd gnd cell_6t
Xbit_r202_c56 bl_56 br_56 wl_202 vdd gnd cell_6t
Xbit_r203_c56 bl_56 br_56 wl_203 vdd gnd cell_6t
Xbit_r204_c56 bl_56 br_56 wl_204 vdd gnd cell_6t
Xbit_r205_c56 bl_56 br_56 wl_205 vdd gnd cell_6t
Xbit_r206_c56 bl_56 br_56 wl_206 vdd gnd cell_6t
Xbit_r207_c56 bl_56 br_56 wl_207 vdd gnd cell_6t
Xbit_r208_c56 bl_56 br_56 wl_208 vdd gnd cell_6t
Xbit_r209_c56 bl_56 br_56 wl_209 vdd gnd cell_6t
Xbit_r210_c56 bl_56 br_56 wl_210 vdd gnd cell_6t
Xbit_r211_c56 bl_56 br_56 wl_211 vdd gnd cell_6t
Xbit_r212_c56 bl_56 br_56 wl_212 vdd gnd cell_6t
Xbit_r213_c56 bl_56 br_56 wl_213 vdd gnd cell_6t
Xbit_r214_c56 bl_56 br_56 wl_214 vdd gnd cell_6t
Xbit_r215_c56 bl_56 br_56 wl_215 vdd gnd cell_6t
Xbit_r216_c56 bl_56 br_56 wl_216 vdd gnd cell_6t
Xbit_r217_c56 bl_56 br_56 wl_217 vdd gnd cell_6t
Xbit_r218_c56 bl_56 br_56 wl_218 vdd gnd cell_6t
Xbit_r219_c56 bl_56 br_56 wl_219 vdd gnd cell_6t
Xbit_r220_c56 bl_56 br_56 wl_220 vdd gnd cell_6t
Xbit_r221_c56 bl_56 br_56 wl_221 vdd gnd cell_6t
Xbit_r222_c56 bl_56 br_56 wl_222 vdd gnd cell_6t
Xbit_r223_c56 bl_56 br_56 wl_223 vdd gnd cell_6t
Xbit_r224_c56 bl_56 br_56 wl_224 vdd gnd cell_6t
Xbit_r225_c56 bl_56 br_56 wl_225 vdd gnd cell_6t
Xbit_r226_c56 bl_56 br_56 wl_226 vdd gnd cell_6t
Xbit_r227_c56 bl_56 br_56 wl_227 vdd gnd cell_6t
Xbit_r228_c56 bl_56 br_56 wl_228 vdd gnd cell_6t
Xbit_r229_c56 bl_56 br_56 wl_229 vdd gnd cell_6t
Xbit_r230_c56 bl_56 br_56 wl_230 vdd gnd cell_6t
Xbit_r231_c56 bl_56 br_56 wl_231 vdd gnd cell_6t
Xbit_r232_c56 bl_56 br_56 wl_232 vdd gnd cell_6t
Xbit_r233_c56 bl_56 br_56 wl_233 vdd gnd cell_6t
Xbit_r234_c56 bl_56 br_56 wl_234 vdd gnd cell_6t
Xbit_r235_c56 bl_56 br_56 wl_235 vdd gnd cell_6t
Xbit_r236_c56 bl_56 br_56 wl_236 vdd gnd cell_6t
Xbit_r237_c56 bl_56 br_56 wl_237 vdd gnd cell_6t
Xbit_r238_c56 bl_56 br_56 wl_238 vdd gnd cell_6t
Xbit_r239_c56 bl_56 br_56 wl_239 vdd gnd cell_6t
Xbit_r240_c56 bl_56 br_56 wl_240 vdd gnd cell_6t
Xbit_r241_c56 bl_56 br_56 wl_241 vdd gnd cell_6t
Xbit_r242_c56 bl_56 br_56 wl_242 vdd gnd cell_6t
Xbit_r243_c56 bl_56 br_56 wl_243 vdd gnd cell_6t
Xbit_r244_c56 bl_56 br_56 wl_244 vdd gnd cell_6t
Xbit_r245_c56 bl_56 br_56 wl_245 vdd gnd cell_6t
Xbit_r246_c56 bl_56 br_56 wl_246 vdd gnd cell_6t
Xbit_r247_c56 bl_56 br_56 wl_247 vdd gnd cell_6t
Xbit_r248_c56 bl_56 br_56 wl_248 vdd gnd cell_6t
Xbit_r249_c56 bl_56 br_56 wl_249 vdd gnd cell_6t
Xbit_r250_c56 bl_56 br_56 wl_250 vdd gnd cell_6t
Xbit_r251_c56 bl_56 br_56 wl_251 vdd gnd cell_6t
Xbit_r252_c56 bl_56 br_56 wl_252 vdd gnd cell_6t
Xbit_r253_c56 bl_56 br_56 wl_253 vdd gnd cell_6t
Xbit_r254_c56 bl_56 br_56 wl_254 vdd gnd cell_6t
Xbit_r255_c56 bl_56 br_56 wl_255 vdd gnd cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd cell_6t
Xbit_r1_c57 bl_57 br_57 wl_1 vdd gnd cell_6t
Xbit_r2_c57 bl_57 br_57 wl_2 vdd gnd cell_6t
Xbit_r3_c57 bl_57 br_57 wl_3 vdd gnd cell_6t
Xbit_r4_c57 bl_57 br_57 wl_4 vdd gnd cell_6t
Xbit_r5_c57 bl_57 br_57 wl_5 vdd gnd cell_6t
Xbit_r6_c57 bl_57 br_57 wl_6 vdd gnd cell_6t
Xbit_r7_c57 bl_57 br_57 wl_7 vdd gnd cell_6t
Xbit_r8_c57 bl_57 br_57 wl_8 vdd gnd cell_6t
Xbit_r9_c57 bl_57 br_57 wl_9 vdd gnd cell_6t
Xbit_r10_c57 bl_57 br_57 wl_10 vdd gnd cell_6t
Xbit_r11_c57 bl_57 br_57 wl_11 vdd gnd cell_6t
Xbit_r12_c57 bl_57 br_57 wl_12 vdd gnd cell_6t
Xbit_r13_c57 bl_57 br_57 wl_13 vdd gnd cell_6t
Xbit_r14_c57 bl_57 br_57 wl_14 vdd gnd cell_6t
Xbit_r15_c57 bl_57 br_57 wl_15 vdd gnd cell_6t
Xbit_r16_c57 bl_57 br_57 wl_16 vdd gnd cell_6t
Xbit_r17_c57 bl_57 br_57 wl_17 vdd gnd cell_6t
Xbit_r18_c57 bl_57 br_57 wl_18 vdd gnd cell_6t
Xbit_r19_c57 bl_57 br_57 wl_19 vdd gnd cell_6t
Xbit_r20_c57 bl_57 br_57 wl_20 vdd gnd cell_6t
Xbit_r21_c57 bl_57 br_57 wl_21 vdd gnd cell_6t
Xbit_r22_c57 bl_57 br_57 wl_22 vdd gnd cell_6t
Xbit_r23_c57 bl_57 br_57 wl_23 vdd gnd cell_6t
Xbit_r24_c57 bl_57 br_57 wl_24 vdd gnd cell_6t
Xbit_r25_c57 bl_57 br_57 wl_25 vdd gnd cell_6t
Xbit_r26_c57 bl_57 br_57 wl_26 vdd gnd cell_6t
Xbit_r27_c57 bl_57 br_57 wl_27 vdd gnd cell_6t
Xbit_r28_c57 bl_57 br_57 wl_28 vdd gnd cell_6t
Xbit_r29_c57 bl_57 br_57 wl_29 vdd gnd cell_6t
Xbit_r30_c57 bl_57 br_57 wl_30 vdd gnd cell_6t
Xbit_r31_c57 bl_57 br_57 wl_31 vdd gnd cell_6t
Xbit_r32_c57 bl_57 br_57 wl_32 vdd gnd cell_6t
Xbit_r33_c57 bl_57 br_57 wl_33 vdd gnd cell_6t
Xbit_r34_c57 bl_57 br_57 wl_34 vdd gnd cell_6t
Xbit_r35_c57 bl_57 br_57 wl_35 vdd gnd cell_6t
Xbit_r36_c57 bl_57 br_57 wl_36 vdd gnd cell_6t
Xbit_r37_c57 bl_57 br_57 wl_37 vdd gnd cell_6t
Xbit_r38_c57 bl_57 br_57 wl_38 vdd gnd cell_6t
Xbit_r39_c57 bl_57 br_57 wl_39 vdd gnd cell_6t
Xbit_r40_c57 bl_57 br_57 wl_40 vdd gnd cell_6t
Xbit_r41_c57 bl_57 br_57 wl_41 vdd gnd cell_6t
Xbit_r42_c57 bl_57 br_57 wl_42 vdd gnd cell_6t
Xbit_r43_c57 bl_57 br_57 wl_43 vdd gnd cell_6t
Xbit_r44_c57 bl_57 br_57 wl_44 vdd gnd cell_6t
Xbit_r45_c57 bl_57 br_57 wl_45 vdd gnd cell_6t
Xbit_r46_c57 bl_57 br_57 wl_46 vdd gnd cell_6t
Xbit_r47_c57 bl_57 br_57 wl_47 vdd gnd cell_6t
Xbit_r48_c57 bl_57 br_57 wl_48 vdd gnd cell_6t
Xbit_r49_c57 bl_57 br_57 wl_49 vdd gnd cell_6t
Xbit_r50_c57 bl_57 br_57 wl_50 vdd gnd cell_6t
Xbit_r51_c57 bl_57 br_57 wl_51 vdd gnd cell_6t
Xbit_r52_c57 bl_57 br_57 wl_52 vdd gnd cell_6t
Xbit_r53_c57 bl_57 br_57 wl_53 vdd gnd cell_6t
Xbit_r54_c57 bl_57 br_57 wl_54 vdd gnd cell_6t
Xbit_r55_c57 bl_57 br_57 wl_55 vdd gnd cell_6t
Xbit_r56_c57 bl_57 br_57 wl_56 vdd gnd cell_6t
Xbit_r57_c57 bl_57 br_57 wl_57 vdd gnd cell_6t
Xbit_r58_c57 bl_57 br_57 wl_58 vdd gnd cell_6t
Xbit_r59_c57 bl_57 br_57 wl_59 vdd gnd cell_6t
Xbit_r60_c57 bl_57 br_57 wl_60 vdd gnd cell_6t
Xbit_r61_c57 bl_57 br_57 wl_61 vdd gnd cell_6t
Xbit_r62_c57 bl_57 br_57 wl_62 vdd gnd cell_6t
Xbit_r63_c57 bl_57 br_57 wl_63 vdd gnd cell_6t
Xbit_r64_c57 bl_57 br_57 wl_64 vdd gnd cell_6t
Xbit_r65_c57 bl_57 br_57 wl_65 vdd gnd cell_6t
Xbit_r66_c57 bl_57 br_57 wl_66 vdd gnd cell_6t
Xbit_r67_c57 bl_57 br_57 wl_67 vdd gnd cell_6t
Xbit_r68_c57 bl_57 br_57 wl_68 vdd gnd cell_6t
Xbit_r69_c57 bl_57 br_57 wl_69 vdd gnd cell_6t
Xbit_r70_c57 bl_57 br_57 wl_70 vdd gnd cell_6t
Xbit_r71_c57 bl_57 br_57 wl_71 vdd gnd cell_6t
Xbit_r72_c57 bl_57 br_57 wl_72 vdd gnd cell_6t
Xbit_r73_c57 bl_57 br_57 wl_73 vdd gnd cell_6t
Xbit_r74_c57 bl_57 br_57 wl_74 vdd gnd cell_6t
Xbit_r75_c57 bl_57 br_57 wl_75 vdd gnd cell_6t
Xbit_r76_c57 bl_57 br_57 wl_76 vdd gnd cell_6t
Xbit_r77_c57 bl_57 br_57 wl_77 vdd gnd cell_6t
Xbit_r78_c57 bl_57 br_57 wl_78 vdd gnd cell_6t
Xbit_r79_c57 bl_57 br_57 wl_79 vdd gnd cell_6t
Xbit_r80_c57 bl_57 br_57 wl_80 vdd gnd cell_6t
Xbit_r81_c57 bl_57 br_57 wl_81 vdd gnd cell_6t
Xbit_r82_c57 bl_57 br_57 wl_82 vdd gnd cell_6t
Xbit_r83_c57 bl_57 br_57 wl_83 vdd gnd cell_6t
Xbit_r84_c57 bl_57 br_57 wl_84 vdd gnd cell_6t
Xbit_r85_c57 bl_57 br_57 wl_85 vdd gnd cell_6t
Xbit_r86_c57 bl_57 br_57 wl_86 vdd gnd cell_6t
Xbit_r87_c57 bl_57 br_57 wl_87 vdd gnd cell_6t
Xbit_r88_c57 bl_57 br_57 wl_88 vdd gnd cell_6t
Xbit_r89_c57 bl_57 br_57 wl_89 vdd gnd cell_6t
Xbit_r90_c57 bl_57 br_57 wl_90 vdd gnd cell_6t
Xbit_r91_c57 bl_57 br_57 wl_91 vdd gnd cell_6t
Xbit_r92_c57 bl_57 br_57 wl_92 vdd gnd cell_6t
Xbit_r93_c57 bl_57 br_57 wl_93 vdd gnd cell_6t
Xbit_r94_c57 bl_57 br_57 wl_94 vdd gnd cell_6t
Xbit_r95_c57 bl_57 br_57 wl_95 vdd gnd cell_6t
Xbit_r96_c57 bl_57 br_57 wl_96 vdd gnd cell_6t
Xbit_r97_c57 bl_57 br_57 wl_97 vdd gnd cell_6t
Xbit_r98_c57 bl_57 br_57 wl_98 vdd gnd cell_6t
Xbit_r99_c57 bl_57 br_57 wl_99 vdd gnd cell_6t
Xbit_r100_c57 bl_57 br_57 wl_100 vdd gnd cell_6t
Xbit_r101_c57 bl_57 br_57 wl_101 vdd gnd cell_6t
Xbit_r102_c57 bl_57 br_57 wl_102 vdd gnd cell_6t
Xbit_r103_c57 bl_57 br_57 wl_103 vdd gnd cell_6t
Xbit_r104_c57 bl_57 br_57 wl_104 vdd gnd cell_6t
Xbit_r105_c57 bl_57 br_57 wl_105 vdd gnd cell_6t
Xbit_r106_c57 bl_57 br_57 wl_106 vdd gnd cell_6t
Xbit_r107_c57 bl_57 br_57 wl_107 vdd gnd cell_6t
Xbit_r108_c57 bl_57 br_57 wl_108 vdd gnd cell_6t
Xbit_r109_c57 bl_57 br_57 wl_109 vdd gnd cell_6t
Xbit_r110_c57 bl_57 br_57 wl_110 vdd gnd cell_6t
Xbit_r111_c57 bl_57 br_57 wl_111 vdd gnd cell_6t
Xbit_r112_c57 bl_57 br_57 wl_112 vdd gnd cell_6t
Xbit_r113_c57 bl_57 br_57 wl_113 vdd gnd cell_6t
Xbit_r114_c57 bl_57 br_57 wl_114 vdd gnd cell_6t
Xbit_r115_c57 bl_57 br_57 wl_115 vdd gnd cell_6t
Xbit_r116_c57 bl_57 br_57 wl_116 vdd gnd cell_6t
Xbit_r117_c57 bl_57 br_57 wl_117 vdd gnd cell_6t
Xbit_r118_c57 bl_57 br_57 wl_118 vdd gnd cell_6t
Xbit_r119_c57 bl_57 br_57 wl_119 vdd gnd cell_6t
Xbit_r120_c57 bl_57 br_57 wl_120 vdd gnd cell_6t
Xbit_r121_c57 bl_57 br_57 wl_121 vdd gnd cell_6t
Xbit_r122_c57 bl_57 br_57 wl_122 vdd gnd cell_6t
Xbit_r123_c57 bl_57 br_57 wl_123 vdd gnd cell_6t
Xbit_r124_c57 bl_57 br_57 wl_124 vdd gnd cell_6t
Xbit_r125_c57 bl_57 br_57 wl_125 vdd gnd cell_6t
Xbit_r126_c57 bl_57 br_57 wl_126 vdd gnd cell_6t
Xbit_r127_c57 bl_57 br_57 wl_127 vdd gnd cell_6t
Xbit_r128_c57 bl_57 br_57 wl_128 vdd gnd cell_6t
Xbit_r129_c57 bl_57 br_57 wl_129 vdd gnd cell_6t
Xbit_r130_c57 bl_57 br_57 wl_130 vdd gnd cell_6t
Xbit_r131_c57 bl_57 br_57 wl_131 vdd gnd cell_6t
Xbit_r132_c57 bl_57 br_57 wl_132 vdd gnd cell_6t
Xbit_r133_c57 bl_57 br_57 wl_133 vdd gnd cell_6t
Xbit_r134_c57 bl_57 br_57 wl_134 vdd gnd cell_6t
Xbit_r135_c57 bl_57 br_57 wl_135 vdd gnd cell_6t
Xbit_r136_c57 bl_57 br_57 wl_136 vdd gnd cell_6t
Xbit_r137_c57 bl_57 br_57 wl_137 vdd gnd cell_6t
Xbit_r138_c57 bl_57 br_57 wl_138 vdd gnd cell_6t
Xbit_r139_c57 bl_57 br_57 wl_139 vdd gnd cell_6t
Xbit_r140_c57 bl_57 br_57 wl_140 vdd gnd cell_6t
Xbit_r141_c57 bl_57 br_57 wl_141 vdd gnd cell_6t
Xbit_r142_c57 bl_57 br_57 wl_142 vdd gnd cell_6t
Xbit_r143_c57 bl_57 br_57 wl_143 vdd gnd cell_6t
Xbit_r144_c57 bl_57 br_57 wl_144 vdd gnd cell_6t
Xbit_r145_c57 bl_57 br_57 wl_145 vdd gnd cell_6t
Xbit_r146_c57 bl_57 br_57 wl_146 vdd gnd cell_6t
Xbit_r147_c57 bl_57 br_57 wl_147 vdd gnd cell_6t
Xbit_r148_c57 bl_57 br_57 wl_148 vdd gnd cell_6t
Xbit_r149_c57 bl_57 br_57 wl_149 vdd gnd cell_6t
Xbit_r150_c57 bl_57 br_57 wl_150 vdd gnd cell_6t
Xbit_r151_c57 bl_57 br_57 wl_151 vdd gnd cell_6t
Xbit_r152_c57 bl_57 br_57 wl_152 vdd gnd cell_6t
Xbit_r153_c57 bl_57 br_57 wl_153 vdd gnd cell_6t
Xbit_r154_c57 bl_57 br_57 wl_154 vdd gnd cell_6t
Xbit_r155_c57 bl_57 br_57 wl_155 vdd gnd cell_6t
Xbit_r156_c57 bl_57 br_57 wl_156 vdd gnd cell_6t
Xbit_r157_c57 bl_57 br_57 wl_157 vdd gnd cell_6t
Xbit_r158_c57 bl_57 br_57 wl_158 vdd gnd cell_6t
Xbit_r159_c57 bl_57 br_57 wl_159 vdd gnd cell_6t
Xbit_r160_c57 bl_57 br_57 wl_160 vdd gnd cell_6t
Xbit_r161_c57 bl_57 br_57 wl_161 vdd gnd cell_6t
Xbit_r162_c57 bl_57 br_57 wl_162 vdd gnd cell_6t
Xbit_r163_c57 bl_57 br_57 wl_163 vdd gnd cell_6t
Xbit_r164_c57 bl_57 br_57 wl_164 vdd gnd cell_6t
Xbit_r165_c57 bl_57 br_57 wl_165 vdd gnd cell_6t
Xbit_r166_c57 bl_57 br_57 wl_166 vdd gnd cell_6t
Xbit_r167_c57 bl_57 br_57 wl_167 vdd gnd cell_6t
Xbit_r168_c57 bl_57 br_57 wl_168 vdd gnd cell_6t
Xbit_r169_c57 bl_57 br_57 wl_169 vdd gnd cell_6t
Xbit_r170_c57 bl_57 br_57 wl_170 vdd gnd cell_6t
Xbit_r171_c57 bl_57 br_57 wl_171 vdd gnd cell_6t
Xbit_r172_c57 bl_57 br_57 wl_172 vdd gnd cell_6t
Xbit_r173_c57 bl_57 br_57 wl_173 vdd gnd cell_6t
Xbit_r174_c57 bl_57 br_57 wl_174 vdd gnd cell_6t
Xbit_r175_c57 bl_57 br_57 wl_175 vdd gnd cell_6t
Xbit_r176_c57 bl_57 br_57 wl_176 vdd gnd cell_6t
Xbit_r177_c57 bl_57 br_57 wl_177 vdd gnd cell_6t
Xbit_r178_c57 bl_57 br_57 wl_178 vdd gnd cell_6t
Xbit_r179_c57 bl_57 br_57 wl_179 vdd gnd cell_6t
Xbit_r180_c57 bl_57 br_57 wl_180 vdd gnd cell_6t
Xbit_r181_c57 bl_57 br_57 wl_181 vdd gnd cell_6t
Xbit_r182_c57 bl_57 br_57 wl_182 vdd gnd cell_6t
Xbit_r183_c57 bl_57 br_57 wl_183 vdd gnd cell_6t
Xbit_r184_c57 bl_57 br_57 wl_184 vdd gnd cell_6t
Xbit_r185_c57 bl_57 br_57 wl_185 vdd gnd cell_6t
Xbit_r186_c57 bl_57 br_57 wl_186 vdd gnd cell_6t
Xbit_r187_c57 bl_57 br_57 wl_187 vdd gnd cell_6t
Xbit_r188_c57 bl_57 br_57 wl_188 vdd gnd cell_6t
Xbit_r189_c57 bl_57 br_57 wl_189 vdd gnd cell_6t
Xbit_r190_c57 bl_57 br_57 wl_190 vdd gnd cell_6t
Xbit_r191_c57 bl_57 br_57 wl_191 vdd gnd cell_6t
Xbit_r192_c57 bl_57 br_57 wl_192 vdd gnd cell_6t
Xbit_r193_c57 bl_57 br_57 wl_193 vdd gnd cell_6t
Xbit_r194_c57 bl_57 br_57 wl_194 vdd gnd cell_6t
Xbit_r195_c57 bl_57 br_57 wl_195 vdd gnd cell_6t
Xbit_r196_c57 bl_57 br_57 wl_196 vdd gnd cell_6t
Xbit_r197_c57 bl_57 br_57 wl_197 vdd gnd cell_6t
Xbit_r198_c57 bl_57 br_57 wl_198 vdd gnd cell_6t
Xbit_r199_c57 bl_57 br_57 wl_199 vdd gnd cell_6t
Xbit_r200_c57 bl_57 br_57 wl_200 vdd gnd cell_6t
Xbit_r201_c57 bl_57 br_57 wl_201 vdd gnd cell_6t
Xbit_r202_c57 bl_57 br_57 wl_202 vdd gnd cell_6t
Xbit_r203_c57 bl_57 br_57 wl_203 vdd gnd cell_6t
Xbit_r204_c57 bl_57 br_57 wl_204 vdd gnd cell_6t
Xbit_r205_c57 bl_57 br_57 wl_205 vdd gnd cell_6t
Xbit_r206_c57 bl_57 br_57 wl_206 vdd gnd cell_6t
Xbit_r207_c57 bl_57 br_57 wl_207 vdd gnd cell_6t
Xbit_r208_c57 bl_57 br_57 wl_208 vdd gnd cell_6t
Xbit_r209_c57 bl_57 br_57 wl_209 vdd gnd cell_6t
Xbit_r210_c57 bl_57 br_57 wl_210 vdd gnd cell_6t
Xbit_r211_c57 bl_57 br_57 wl_211 vdd gnd cell_6t
Xbit_r212_c57 bl_57 br_57 wl_212 vdd gnd cell_6t
Xbit_r213_c57 bl_57 br_57 wl_213 vdd gnd cell_6t
Xbit_r214_c57 bl_57 br_57 wl_214 vdd gnd cell_6t
Xbit_r215_c57 bl_57 br_57 wl_215 vdd gnd cell_6t
Xbit_r216_c57 bl_57 br_57 wl_216 vdd gnd cell_6t
Xbit_r217_c57 bl_57 br_57 wl_217 vdd gnd cell_6t
Xbit_r218_c57 bl_57 br_57 wl_218 vdd gnd cell_6t
Xbit_r219_c57 bl_57 br_57 wl_219 vdd gnd cell_6t
Xbit_r220_c57 bl_57 br_57 wl_220 vdd gnd cell_6t
Xbit_r221_c57 bl_57 br_57 wl_221 vdd gnd cell_6t
Xbit_r222_c57 bl_57 br_57 wl_222 vdd gnd cell_6t
Xbit_r223_c57 bl_57 br_57 wl_223 vdd gnd cell_6t
Xbit_r224_c57 bl_57 br_57 wl_224 vdd gnd cell_6t
Xbit_r225_c57 bl_57 br_57 wl_225 vdd gnd cell_6t
Xbit_r226_c57 bl_57 br_57 wl_226 vdd gnd cell_6t
Xbit_r227_c57 bl_57 br_57 wl_227 vdd gnd cell_6t
Xbit_r228_c57 bl_57 br_57 wl_228 vdd gnd cell_6t
Xbit_r229_c57 bl_57 br_57 wl_229 vdd gnd cell_6t
Xbit_r230_c57 bl_57 br_57 wl_230 vdd gnd cell_6t
Xbit_r231_c57 bl_57 br_57 wl_231 vdd gnd cell_6t
Xbit_r232_c57 bl_57 br_57 wl_232 vdd gnd cell_6t
Xbit_r233_c57 bl_57 br_57 wl_233 vdd gnd cell_6t
Xbit_r234_c57 bl_57 br_57 wl_234 vdd gnd cell_6t
Xbit_r235_c57 bl_57 br_57 wl_235 vdd gnd cell_6t
Xbit_r236_c57 bl_57 br_57 wl_236 vdd gnd cell_6t
Xbit_r237_c57 bl_57 br_57 wl_237 vdd gnd cell_6t
Xbit_r238_c57 bl_57 br_57 wl_238 vdd gnd cell_6t
Xbit_r239_c57 bl_57 br_57 wl_239 vdd gnd cell_6t
Xbit_r240_c57 bl_57 br_57 wl_240 vdd gnd cell_6t
Xbit_r241_c57 bl_57 br_57 wl_241 vdd gnd cell_6t
Xbit_r242_c57 bl_57 br_57 wl_242 vdd gnd cell_6t
Xbit_r243_c57 bl_57 br_57 wl_243 vdd gnd cell_6t
Xbit_r244_c57 bl_57 br_57 wl_244 vdd gnd cell_6t
Xbit_r245_c57 bl_57 br_57 wl_245 vdd gnd cell_6t
Xbit_r246_c57 bl_57 br_57 wl_246 vdd gnd cell_6t
Xbit_r247_c57 bl_57 br_57 wl_247 vdd gnd cell_6t
Xbit_r248_c57 bl_57 br_57 wl_248 vdd gnd cell_6t
Xbit_r249_c57 bl_57 br_57 wl_249 vdd gnd cell_6t
Xbit_r250_c57 bl_57 br_57 wl_250 vdd gnd cell_6t
Xbit_r251_c57 bl_57 br_57 wl_251 vdd gnd cell_6t
Xbit_r252_c57 bl_57 br_57 wl_252 vdd gnd cell_6t
Xbit_r253_c57 bl_57 br_57 wl_253 vdd gnd cell_6t
Xbit_r254_c57 bl_57 br_57 wl_254 vdd gnd cell_6t
Xbit_r255_c57 bl_57 br_57 wl_255 vdd gnd cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd cell_6t
Xbit_r1_c58 bl_58 br_58 wl_1 vdd gnd cell_6t
Xbit_r2_c58 bl_58 br_58 wl_2 vdd gnd cell_6t
Xbit_r3_c58 bl_58 br_58 wl_3 vdd gnd cell_6t
Xbit_r4_c58 bl_58 br_58 wl_4 vdd gnd cell_6t
Xbit_r5_c58 bl_58 br_58 wl_5 vdd gnd cell_6t
Xbit_r6_c58 bl_58 br_58 wl_6 vdd gnd cell_6t
Xbit_r7_c58 bl_58 br_58 wl_7 vdd gnd cell_6t
Xbit_r8_c58 bl_58 br_58 wl_8 vdd gnd cell_6t
Xbit_r9_c58 bl_58 br_58 wl_9 vdd gnd cell_6t
Xbit_r10_c58 bl_58 br_58 wl_10 vdd gnd cell_6t
Xbit_r11_c58 bl_58 br_58 wl_11 vdd gnd cell_6t
Xbit_r12_c58 bl_58 br_58 wl_12 vdd gnd cell_6t
Xbit_r13_c58 bl_58 br_58 wl_13 vdd gnd cell_6t
Xbit_r14_c58 bl_58 br_58 wl_14 vdd gnd cell_6t
Xbit_r15_c58 bl_58 br_58 wl_15 vdd gnd cell_6t
Xbit_r16_c58 bl_58 br_58 wl_16 vdd gnd cell_6t
Xbit_r17_c58 bl_58 br_58 wl_17 vdd gnd cell_6t
Xbit_r18_c58 bl_58 br_58 wl_18 vdd gnd cell_6t
Xbit_r19_c58 bl_58 br_58 wl_19 vdd gnd cell_6t
Xbit_r20_c58 bl_58 br_58 wl_20 vdd gnd cell_6t
Xbit_r21_c58 bl_58 br_58 wl_21 vdd gnd cell_6t
Xbit_r22_c58 bl_58 br_58 wl_22 vdd gnd cell_6t
Xbit_r23_c58 bl_58 br_58 wl_23 vdd gnd cell_6t
Xbit_r24_c58 bl_58 br_58 wl_24 vdd gnd cell_6t
Xbit_r25_c58 bl_58 br_58 wl_25 vdd gnd cell_6t
Xbit_r26_c58 bl_58 br_58 wl_26 vdd gnd cell_6t
Xbit_r27_c58 bl_58 br_58 wl_27 vdd gnd cell_6t
Xbit_r28_c58 bl_58 br_58 wl_28 vdd gnd cell_6t
Xbit_r29_c58 bl_58 br_58 wl_29 vdd gnd cell_6t
Xbit_r30_c58 bl_58 br_58 wl_30 vdd gnd cell_6t
Xbit_r31_c58 bl_58 br_58 wl_31 vdd gnd cell_6t
Xbit_r32_c58 bl_58 br_58 wl_32 vdd gnd cell_6t
Xbit_r33_c58 bl_58 br_58 wl_33 vdd gnd cell_6t
Xbit_r34_c58 bl_58 br_58 wl_34 vdd gnd cell_6t
Xbit_r35_c58 bl_58 br_58 wl_35 vdd gnd cell_6t
Xbit_r36_c58 bl_58 br_58 wl_36 vdd gnd cell_6t
Xbit_r37_c58 bl_58 br_58 wl_37 vdd gnd cell_6t
Xbit_r38_c58 bl_58 br_58 wl_38 vdd gnd cell_6t
Xbit_r39_c58 bl_58 br_58 wl_39 vdd gnd cell_6t
Xbit_r40_c58 bl_58 br_58 wl_40 vdd gnd cell_6t
Xbit_r41_c58 bl_58 br_58 wl_41 vdd gnd cell_6t
Xbit_r42_c58 bl_58 br_58 wl_42 vdd gnd cell_6t
Xbit_r43_c58 bl_58 br_58 wl_43 vdd gnd cell_6t
Xbit_r44_c58 bl_58 br_58 wl_44 vdd gnd cell_6t
Xbit_r45_c58 bl_58 br_58 wl_45 vdd gnd cell_6t
Xbit_r46_c58 bl_58 br_58 wl_46 vdd gnd cell_6t
Xbit_r47_c58 bl_58 br_58 wl_47 vdd gnd cell_6t
Xbit_r48_c58 bl_58 br_58 wl_48 vdd gnd cell_6t
Xbit_r49_c58 bl_58 br_58 wl_49 vdd gnd cell_6t
Xbit_r50_c58 bl_58 br_58 wl_50 vdd gnd cell_6t
Xbit_r51_c58 bl_58 br_58 wl_51 vdd gnd cell_6t
Xbit_r52_c58 bl_58 br_58 wl_52 vdd gnd cell_6t
Xbit_r53_c58 bl_58 br_58 wl_53 vdd gnd cell_6t
Xbit_r54_c58 bl_58 br_58 wl_54 vdd gnd cell_6t
Xbit_r55_c58 bl_58 br_58 wl_55 vdd gnd cell_6t
Xbit_r56_c58 bl_58 br_58 wl_56 vdd gnd cell_6t
Xbit_r57_c58 bl_58 br_58 wl_57 vdd gnd cell_6t
Xbit_r58_c58 bl_58 br_58 wl_58 vdd gnd cell_6t
Xbit_r59_c58 bl_58 br_58 wl_59 vdd gnd cell_6t
Xbit_r60_c58 bl_58 br_58 wl_60 vdd gnd cell_6t
Xbit_r61_c58 bl_58 br_58 wl_61 vdd gnd cell_6t
Xbit_r62_c58 bl_58 br_58 wl_62 vdd gnd cell_6t
Xbit_r63_c58 bl_58 br_58 wl_63 vdd gnd cell_6t
Xbit_r64_c58 bl_58 br_58 wl_64 vdd gnd cell_6t
Xbit_r65_c58 bl_58 br_58 wl_65 vdd gnd cell_6t
Xbit_r66_c58 bl_58 br_58 wl_66 vdd gnd cell_6t
Xbit_r67_c58 bl_58 br_58 wl_67 vdd gnd cell_6t
Xbit_r68_c58 bl_58 br_58 wl_68 vdd gnd cell_6t
Xbit_r69_c58 bl_58 br_58 wl_69 vdd gnd cell_6t
Xbit_r70_c58 bl_58 br_58 wl_70 vdd gnd cell_6t
Xbit_r71_c58 bl_58 br_58 wl_71 vdd gnd cell_6t
Xbit_r72_c58 bl_58 br_58 wl_72 vdd gnd cell_6t
Xbit_r73_c58 bl_58 br_58 wl_73 vdd gnd cell_6t
Xbit_r74_c58 bl_58 br_58 wl_74 vdd gnd cell_6t
Xbit_r75_c58 bl_58 br_58 wl_75 vdd gnd cell_6t
Xbit_r76_c58 bl_58 br_58 wl_76 vdd gnd cell_6t
Xbit_r77_c58 bl_58 br_58 wl_77 vdd gnd cell_6t
Xbit_r78_c58 bl_58 br_58 wl_78 vdd gnd cell_6t
Xbit_r79_c58 bl_58 br_58 wl_79 vdd gnd cell_6t
Xbit_r80_c58 bl_58 br_58 wl_80 vdd gnd cell_6t
Xbit_r81_c58 bl_58 br_58 wl_81 vdd gnd cell_6t
Xbit_r82_c58 bl_58 br_58 wl_82 vdd gnd cell_6t
Xbit_r83_c58 bl_58 br_58 wl_83 vdd gnd cell_6t
Xbit_r84_c58 bl_58 br_58 wl_84 vdd gnd cell_6t
Xbit_r85_c58 bl_58 br_58 wl_85 vdd gnd cell_6t
Xbit_r86_c58 bl_58 br_58 wl_86 vdd gnd cell_6t
Xbit_r87_c58 bl_58 br_58 wl_87 vdd gnd cell_6t
Xbit_r88_c58 bl_58 br_58 wl_88 vdd gnd cell_6t
Xbit_r89_c58 bl_58 br_58 wl_89 vdd gnd cell_6t
Xbit_r90_c58 bl_58 br_58 wl_90 vdd gnd cell_6t
Xbit_r91_c58 bl_58 br_58 wl_91 vdd gnd cell_6t
Xbit_r92_c58 bl_58 br_58 wl_92 vdd gnd cell_6t
Xbit_r93_c58 bl_58 br_58 wl_93 vdd gnd cell_6t
Xbit_r94_c58 bl_58 br_58 wl_94 vdd gnd cell_6t
Xbit_r95_c58 bl_58 br_58 wl_95 vdd gnd cell_6t
Xbit_r96_c58 bl_58 br_58 wl_96 vdd gnd cell_6t
Xbit_r97_c58 bl_58 br_58 wl_97 vdd gnd cell_6t
Xbit_r98_c58 bl_58 br_58 wl_98 vdd gnd cell_6t
Xbit_r99_c58 bl_58 br_58 wl_99 vdd gnd cell_6t
Xbit_r100_c58 bl_58 br_58 wl_100 vdd gnd cell_6t
Xbit_r101_c58 bl_58 br_58 wl_101 vdd gnd cell_6t
Xbit_r102_c58 bl_58 br_58 wl_102 vdd gnd cell_6t
Xbit_r103_c58 bl_58 br_58 wl_103 vdd gnd cell_6t
Xbit_r104_c58 bl_58 br_58 wl_104 vdd gnd cell_6t
Xbit_r105_c58 bl_58 br_58 wl_105 vdd gnd cell_6t
Xbit_r106_c58 bl_58 br_58 wl_106 vdd gnd cell_6t
Xbit_r107_c58 bl_58 br_58 wl_107 vdd gnd cell_6t
Xbit_r108_c58 bl_58 br_58 wl_108 vdd gnd cell_6t
Xbit_r109_c58 bl_58 br_58 wl_109 vdd gnd cell_6t
Xbit_r110_c58 bl_58 br_58 wl_110 vdd gnd cell_6t
Xbit_r111_c58 bl_58 br_58 wl_111 vdd gnd cell_6t
Xbit_r112_c58 bl_58 br_58 wl_112 vdd gnd cell_6t
Xbit_r113_c58 bl_58 br_58 wl_113 vdd gnd cell_6t
Xbit_r114_c58 bl_58 br_58 wl_114 vdd gnd cell_6t
Xbit_r115_c58 bl_58 br_58 wl_115 vdd gnd cell_6t
Xbit_r116_c58 bl_58 br_58 wl_116 vdd gnd cell_6t
Xbit_r117_c58 bl_58 br_58 wl_117 vdd gnd cell_6t
Xbit_r118_c58 bl_58 br_58 wl_118 vdd gnd cell_6t
Xbit_r119_c58 bl_58 br_58 wl_119 vdd gnd cell_6t
Xbit_r120_c58 bl_58 br_58 wl_120 vdd gnd cell_6t
Xbit_r121_c58 bl_58 br_58 wl_121 vdd gnd cell_6t
Xbit_r122_c58 bl_58 br_58 wl_122 vdd gnd cell_6t
Xbit_r123_c58 bl_58 br_58 wl_123 vdd gnd cell_6t
Xbit_r124_c58 bl_58 br_58 wl_124 vdd gnd cell_6t
Xbit_r125_c58 bl_58 br_58 wl_125 vdd gnd cell_6t
Xbit_r126_c58 bl_58 br_58 wl_126 vdd gnd cell_6t
Xbit_r127_c58 bl_58 br_58 wl_127 vdd gnd cell_6t
Xbit_r128_c58 bl_58 br_58 wl_128 vdd gnd cell_6t
Xbit_r129_c58 bl_58 br_58 wl_129 vdd gnd cell_6t
Xbit_r130_c58 bl_58 br_58 wl_130 vdd gnd cell_6t
Xbit_r131_c58 bl_58 br_58 wl_131 vdd gnd cell_6t
Xbit_r132_c58 bl_58 br_58 wl_132 vdd gnd cell_6t
Xbit_r133_c58 bl_58 br_58 wl_133 vdd gnd cell_6t
Xbit_r134_c58 bl_58 br_58 wl_134 vdd gnd cell_6t
Xbit_r135_c58 bl_58 br_58 wl_135 vdd gnd cell_6t
Xbit_r136_c58 bl_58 br_58 wl_136 vdd gnd cell_6t
Xbit_r137_c58 bl_58 br_58 wl_137 vdd gnd cell_6t
Xbit_r138_c58 bl_58 br_58 wl_138 vdd gnd cell_6t
Xbit_r139_c58 bl_58 br_58 wl_139 vdd gnd cell_6t
Xbit_r140_c58 bl_58 br_58 wl_140 vdd gnd cell_6t
Xbit_r141_c58 bl_58 br_58 wl_141 vdd gnd cell_6t
Xbit_r142_c58 bl_58 br_58 wl_142 vdd gnd cell_6t
Xbit_r143_c58 bl_58 br_58 wl_143 vdd gnd cell_6t
Xbit_r144_c58 bl_58 br_58 wl_144 vdd gnd cell_6t
Xbit_r145_c58 bl_58 br_58 wl_145 vdd gnd cell_6t
Xbit_r146_c58 bl_58 br_58 wl_146 vdd gnd cell_6t
Xbit_r147_c58 bl_58 br_58 wl_147 vdd gnd cell_6t
Xbit_r148_c58 bl_58 br_58 wl_148 vdd gnd cell_6t
Xbit_r149_c58 bl_58 br_58 wl_149 vdd gnd cell_6t
Xbit_r150_c58 bl_58 br_58 wl_150 vdd gnd cell_6t
Xbit_r151_c58 bl_58 br_58 wl_151 vdd gnd cell_6t
Xbit_r152_c58 bl_58 br_58 wl_152 vdd gnd cell_6t
Xbit_r153_c58 bl_58 br_58 wl_153 vdd gnd cell_6t
Xbit_r154_c58 bl_58 br_58 wl_154 vdd gnd cell_6t
Xbit_r155_c58 bl_58 br_58 wl_155 vdd gnd cell_6t
Xbit_r156_c58 bl_58 br_58 wl_156 vdd gnd cell_6t
Xbit_r157_c58 bl_58 br_58 wl_157 vdd gnd cell_6t
Xbit_r158_c58 bl_58 br_58 wl_158 vdd gnd cell_6t
Xbit_r159_c58 bl_58 br_58 wl_159 vdd gnd cell_6t
Xbit_r160_c58 bl_58 br_58 wl_160 vdd gnd cell_6t
Xbit_r161_c58 bl_58 br_58 wl_161 vdd gnd cell_6t
Xbit_r162_c58 bl_58 br_58 wl_162 vdd gnd cell_6t
Xbit_r163_c58 bl_58 br_58 wl_163 vdd gnd cell_6t
Xbit_r164_c58 bl_58 br_58 wl_164 vdd gnd cell_6t
Xbit_r165_c58 bl_58 br_58 wl_165 vdd gnd cell_6t
Xbit_r166_c58 bl_58 br_58 wl_166 vdd gnd cell_6t
Xbit_r167_c58 bl_58 br_58 wl_167 vdd gnd cell_6t
Xbit_r168_c58 bl_58 br_58 wl_168 vdd gnd cell_6t
Xbit_r169_c58 bl_58 br_58 wl_169 vdd gnd cell_6t
Xbit_r170_c58 bl_58 br_58 wl_170 vdd gnd cell_6t
Xbit_r171_c58 bl_58 br_58 wl_171 vdd gnd cell_6t
Xbit_r172_c58 bl_58 br_58 wl_172 vdd gnd cell_6t
Xbit_r173_c58 bl_58 br_58 wl_173 vdd gnd cell_6t
Xbit_r174_c58 bl_58 br_58 wl_174 vdd gnd cell_6t
Xbit_r175_c58 bl_58 br_58 wl_175 vdd gnd cell_6t
Xbit_r176_c58 bl_58 br_58 wl_176 vdd gnd cell_6t
Xbit_r177_c58 bl_58 br_58 wl_177 vdd gnd cell_6t
Xbit_r178_c58 bl_58 br_58 wl_178 vdd gnd cell_6t
Xbit_r179_c58 bl_58 br_58 wl_179 vdd gnd cell_6t
Xbit_r180_c58 bl_58 br_58 wl_180 vdd gnd cell_6t
Xbit_r181_c58 bl_58 br_58 wl_181 vdd gnd cell_6t
Xbit_r182_c58 bl_58 br_58 wl_182 vdd gnd cell_6t
Xbit_r183_c58 bl_58 br_58 wl_183 vdd gnd cell_6t
Xbit_r184_c58 bl_58 br_58 wl_184 vdd gnd cell_6t
Xbit_r185_c58 bl_58 br_58 wl_185 vdd gnd cell_6t
Xbit_r186_c58 bl_58 br_58 wl_186 vdd gnd cell_6t
Xbit_r187_c58 bl_58 br_58 wl_187 vdd gnd cell_6t
Xbit_r188_c58 bl_58 br_58 wl_188 vdd gnd cell_6t
Xbit_r189_c58 bl_58 br_58 wl_189 vdd gnd cell_6t
Xbit_r190_c58 bl_58 br_58 wl_190 vdd gnd cell_6t
Xbit_r191_c58 bl_58 br_58 wl_191 vdd gnd cell_6t
Xbit_r192_c58 bl_58 br_58 wl_192 vdd gnd cell_6t
Xbit_r193_c58 bl_58 br_58 wl_193 vdd gnd cell_6t
Xbit_r194_c58 bl_58 br_58 wl_194 vdd gnd cell_6t
Xbit_r195_c58 bl_58 br_58 wl_195 vdd gnd cell_6t
Xbit_r196_c58 bl_58 br_58 wl_196 vdd gnd cell_6t
Xbit_r197_c58 bl_58 br_58 wl_197 vdd gnd cell_6t
Xbit_r198_c58 bl_58 br_58 wl_198 vdd gnd cell_6t
Xbit_r199_c58 bl_58 br_58 wl_199 vdd gnd cell_6t
Xbit_r200_c58 bl_58 br_58 wl_200 vdd gnd cell_6t
Xbit_r201_c58 bl_58 br_58 wl_201 vdd gnd cell_6t
Xbit_r202_c58 bl_58 br_58 wl_202 vdd gnd cell_6t
Xbit_r203_c58 bl_58 br_58 wl_203 vdd gnd cell_6t
Xbit_r204_c58 bl_58 br_58 wl_204 vdd gnd cell_6t
Xbit_r205_c58 bl_58 br_58 wl_205 vdd gnd cell_6t
Xbit_r206_c58 bl_58 br_58 wl_206 vdd gnd cell_6t
Xbit_r207_c58 bl_58 br_58 wl_207 vdd gnd cell_6t
Xbit_r208_c58 bl_58 br_58 wl_208 vdd gnd cell_6t
Xbit_r209_c58 bl_58 br_58 wl_209 vdd gnd cell_6t
Xbit_r210_c58 bl_58 br_58 wl_210 vdd gnd cell_6t
Xbit_r211_c58 bl_58 br_58 wl_211 vdd gnd cell_6t
Xbit_r212_c58 bl_58 br_58 wl_212 vdd gnd cell_6t
Xbit_r213_c58 bl_58 br_58 wl_213 vdd gnd cell_6t
Xbit_r214_c58 bl_58 br_58 wl_214 vdd gnd cell_6t
Xbit_r215_c58 bl_58 br_58 wl_215 vdd gnd cell_6t
Xbit_r216_c58 bl_58 br_58 wl_216 vdd gnd cell_6t
Xbit_r217_c58 bl_58 br_58 wl_217 vdd gnd cell_6t
Xbit_r218_c58 bl_58 br_58 wl_218 vdd gnd cell_6t
Xbit_r219_c58 bl_58 br_58 wl_219 vdd gnd cell_6t
Xbit_r220_c58 bl_58 br_58 wl_220 vdd gnd cell_6t
Xbit_r221_c58 bl_58 br_58 wl_221 vdd gnd cell_6t
Xbit_r222_c58 bl_58 br_58 wl_222 vdd gnd cell_6t
Xbit_r223_c58 bl_58 br_58 wl_223 vdd gnd cell_6t
Xbit_r224_c58 bl_58 br_58 wl_224 vdd gnd cell_6t
Xbit_r225_c58 bl_58 br_58 wl_225 vdd gnd cell_6t
Xbit_r226_c58 bl_58 br_58 wl_226 vdd gnd cell_6t
Xbit_r227_c58 bl_58 br_58 wl_227 vdd gnd cell_6t
Xbit_r228_c58 bl_58 br_58 wl_228 vdd gnd cell_6t
Xbit_r229_c58 bl_58 br_58 wl_229 vdd gnd cell_6t
Xbit_r230_c58 bl_58 br_58 wl_230 vdd gnd cell_6t
Xbit_r231_c58 bl_58 br_58 wl_231 vdd gnd cell_6t
Xbit_r232_c58 bl_58 br_58 wl_232 vdd gnd cell_6t
Xbit_r233_c58 bl_58 br_58 wl_233 vdd gnd cell_6t
Xbit_r234_c58 bl_58 br_58 wl_234 vdd gnd cell_6t
Xbit_r235_c58 bl_58 br_58 wl_235 vdd gnd cell_6t
Xbit_r236_c58 bl_58 br_58 wl_236 vdd gnd cell_6t
Xbit_r237_c58 bl_58 br_58 wl_237 vdd gnd cell_6t
Xbit_r238_c58 bl_58 br_58 wl_238 vdd gnd cell_6t
Xbit_r239_c58 bl_58 br_58 wl_239 vdd gnd cell_6t
Xbit_r240_c58 bl_58 br_58 wl_240 vdd gnd cell_6t
Xbit_r241_c58 bl_58 br_58 wl_241 vdd gnd cell_6t
Xbit_r242_c58 bl_58 br_58 wl_242 vdd gnd cell_6t
Xbit_r243_c58 bl_58 br_58 wl_243 vdd gnd cell_6t
Xbit_r244_c58 bl_58 br_58 wl_244 vdd gnd cell_6t
Xbit_r245_c58 bl_58 br_58 wl_245 vdd gnd cell_6t
Xbit_r246_c58 bl_58 br_58 wl_246 vdd gnd cell_6t
Xbit_r247_c58 bl_58 br_58 wl_247 vdd gnd cell_6t
Xbit_r248_c58 bl_58 br_58 wl_248 vdd gnd cell_6t
Xbit_r249_c58 bl_58 br_58 wl_249 vdd gnd cell_6t
Xbit_r250_c58 bl_58 br_58 wl_250 vdd gnd cell_6t
Xbit_r251_c58 bl_58 br_58 wl_251 vdd gnd cell_6t
Xbit_r252_c58 bl_58 br_58 wl_252 vdd gnd cell_6t
Xbit_r253_c58 bl_58 br_58 wl_253 vdd gnd cell_6t
Xbit_r254_c58 bl_58 br_58 wl_254 vdd gnd cell_6t
Xbit_r255_c58 bl_58 br_58 wl_255 vdd gnd cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd cell_6t
Xbit_r1_c59 bl_59 br_59 wl_1 vdd gnd cell_6t
Xbit_r2_c59 bl_59 br_59 wl_2 vdd gnd cell_6t
Xbit_r3_c59 bl_59 br_59 wl_3 vdd gnd cell_6t
Xbit_r4_c59 bl_59 br_59 wl_4 vdd gnd cell_6t
Xbit_r5_c59 bl_59 br_59 wl_5 vdd gnd cell_6t
Xbit_r6_c59 bl_59 br_59 wl_6 vdd gnd cell_6t
Xbit_r7_c59 bl_59 br_59 wl_7 vdd gnd cell_6t
Xbit_r8_c59 bl_59 br_59 wl_8 vdd gnd cell_6t
Xbit_r9_c59 bl_59 br_59 wl_9 vdd gnd cell_6t
Xbit_r10_c59 bl_59 br_59 wl_10 vdd gnd cell_6t
Xbit_r11_c59 bl_59 br_59 wl_11 vdd gnd cell_6t
Xbit_r12_c59 bl_59 br_59 wl_12 vdd gnd cell_6t
Xbit_r13_c59 bl_59 br_59 wl_13 vdd gnd cell_6t
Xbit_r14_c59 bl_59 br_59 wl_14 vdd gnd cell_6t
Xbit_r15_c59 bl_59 br_59 wl_15 vdd gnd cell_6t
Xbit_r16_c59 bl_59 br_59 wl_16 vdd gnd cell_6t
Xbit_r17_c59 bl_59 br_59 wl_17 vdd gnd cell_6t
Xbit_r18_c59 bl_59 br_59 wl_18 vdd gnd cell_6t
Xbit_r19_c59 bl_59 br_59 wl_19 vdd gnd cell_6t
Xbit_r20_c59 bl_59 br_59 wl_20 vdd gnd cell_6t
Xbit_r21_c59 bl_59 br_59 wl_21 vdd gnd cell_6t
Xbit_r22_c59 bl_59 br_59 wl_22 vdd gnd cell_6t
Xbit_r23_c59 bl_59 br_59 wl_23 vdd gnd cell_6t
Xbit_r24_c59 bl_59 br_59 wl_24 vdd gnd cell_6t
Xbit_r25_c59 bl_59 br_59 wl_25 vdd gnd cell_6t
Xbit_r26_c59 bl_59 br_59 wl_26 vdd gnd cell_6t
Xbit_r27_c59 bl_59 br_59 wl_27 vdd gnd cell_6t
Xbit_r28_c59 bl_59 br_59 wl_28 vdd gnd cell_6t
Xbit_r29_c59 bl_59 br_59 wl_29 vdd gnd cell_6t
Xbit_r30_c59 bl_59 br_59 wl_30 vdd gnd cell_6t
Xbit_r31_c59 bl_59 br_59 wl_31 vdd gnd cell_6t
Xbit_r32_c59 bl_59 br_59 wl_32 vdd gnd cell_6t
Xbit_r33_c59 bl_59 br_59 wl_33 vdd gnd cell_6t
Xbit_r34_c59 bl_59 br_59 wl_34 vdd gnd cell_6t
Xbit_r35_c59 bl_59 br_59 wl_35 vdd gnd cell_6t
Xbit_r36_c59 bl_59 br_59 wl_36 vdd gnd cell_6t
Xbit_r37_c59 bl_59 br_59 wl_37 vdd gnd cell_6t
Xbit_r38_c59 bl_59 br_59 wl_38 vdd gnd cell_6t
Xbit_r39_c59 bl_59 br_59 wl_39 vdd gnd cell_6t
Xbit_r40_c59 bl_59 br_59 wl_40 vdd gnd cell_6t
Xbit_r41_c59 bl_59 br_59 wl_41 vdd gnd cell_6t
Xbit_r42_c59 bl_59 br_59 wl_42 vdd gnd cell_6t
Xbit_r43_c59 bl_59 br_59 wl_43 vdd gnd cell_6t
Xbit_r44_c59 bl_59 br_59 wl_44 vdd gnd cell_6t
Xbit_r45_c59 bl_59 br_59 wl_45 vdd gnd cell_6t
Xbit_r46_c59 bl_59 br_59 wl_46 vdd gnd cell_6t
Xbit_r47_c59 bl_59 br_59 wl_47 vdd gnd cell_6t
Xbit_r48_c59 bl_59 br_59 wl_48 vdd gnd cell_6t
Xbit_r49_c59 bl_59 br_59 wl_49 vdd gnd cell_6t
Xbit_r50_c59 bl_59 br_59 wl_50 vdd gnd cell_6t
Xbit_r51_c59 bl_59 br_59 wl_51 vdd gnd cell_6t
Xbit_r52_c59 bl_59 br_59 wl_52 vdd gnd cell_6t
Xbit_r53_c59 bl_59 br_59 wl_53 vdd gnd cell_6t
Xbit_r54_c59 bl_59 br_59 wl_54 vdd gnd cell_6t
Xbit_r55_c59 bl_59 br_59 wl_55 vdd gnd cell_6t
Xbit_r56_c59 bl_59 br_59 wl_56 vdd gnd cell_6t
Xbit_r57_c59 bl_59 br_59 wl_57 vdd gnd cell_6t
Xbit_r58_c59 bl_59 br_59 wl_58 vdd gnd cell_6t
Xbit_r59_c59 bl_59 br_59 wl_59 vdd gnd cell_6t
Xbit_r60_c59 bl_59 br_59 wl_60 vdd gnd cell_6t
Xbit_r61_c59 bl_59 br_59 wl_61 vdd gnd cell_6t
Xbit_r62_c59 bl_59 br_59 wl_62 vdd gnd cell_6t
Xbit_r63_c59 bl_59 br_59 wl_63 vdd gnd cell_6t
Xbit_r64_c59 bl_59 br_59 wl_64 vdd gnd cell_6t
Xbit_r65_c59 bl_59 br_59 wl_65 vdd gnd cell_6t
Xbit_r66_c59 bl_59 br_59 wl_66 vdd gnd cell_6t
Xbit_r67_c59 bl_59 br_59 wl_67 vdd gnd cell_6t
Xbit_r68_c59 bl_59 br_59 wl_68 vdd gnd cell_6t
Xbit_r69_c59 bl_59 br_59 wl_69 vdd gnd cell_6t
Xbit_r70_c59 bl_59 br_59 wl_70 vdd gnd cell_6t
Xbit_r71_c59 bl_59 br_59 wl_71 vdd gnd cell_6t
Xbit_r72_c59 bl_59 br_59 wl_72 vdd gnd cell_6t
Xbit_r73_c59 bl_59 br_59 wl_73 vdd gnd cell_6t
Xbit_r74_c59 bl_59 br_59 wl_74 vdd gnd cell_6t
Xbit_r75_c59 bl_59 br_59 wl_75 vdd gnd cell_6t
Xbit_r76_c59 bl_59 br_59 wl_76 vdd gnd cell_6t
Xbit_r77_c59 bl_59 br_59 wl_77 vdd gnd cell_6t
Xbit_r78_c59 bl_59 br_59 wl_78 vdd gnd cell_6t
Xbit_r79_c59 bl_59 br_59 wl_79 vdd gnd cell_6t
Xbit_r80_c59 bl_59 br_59 wl_80 vdd gnd cell_6t
Xbit_r81_c59 bl_59 br_59 wl_81 vdd gnd cell_6t
Xbit_r82_c59 bl_59 br_59 wl_82 vdd gnd cell_6t
Xbit_r83_c59 bl_59 br_59 wl_83 vdd gnd cell_6t
Xbit_r84_c59 bl_59 br_59 wl_84 vdd gnd cell_6t
Xbit_r85_c59 bl_59 br_59 wl_85 vdd gnd cell_6t
Xbit_r86_c59 bl_59 br_59 wl_86 vdd gnd cell_6t
Xbit_r87_c59 bl_59 br_59 wl_87 vdd gnd cell_6t
Xbit_r88_c59 bl_59 br_59 wl_88 vdd gnd cell_6t
Xbit_r89_c59 bl_59 br_59 wl_89 vdd gnd cell_6t
Xbit_r90_c59 bl_59 br_59 wl_90 vdd gnd cell_6t
Xbit_r91_c59 bl_59 br_59 wl_91 vdd gnd cell_6t
Xbit_r92_c59 bl_59 br_59 wl_92 vdd gnd cell_6t
Xbit_r93_c59 bl_59 br_59 wl_93 vdd gnd cell_6t
Xbit_r94_c59 bl_59 br_59 wl_94 vdd gnd cell_6t
Xbit_r95_c59 bl_59 br_59 wl_95 vdd gnd cell_6t
Xbit_r96_c59 bl_59 br_59 wl_96 vdd gnd cell_6t
Xbit_r97_c59 bl_59 br_59 wl_97 vdd gnd cell_6t
Xbit_r98_c59 bl_59 br_59 wl_98 vdd gnd cell_6t
Xbit_r99_c59 bl_59 br_59 wl_99 vdd gnd cell_6t
Xbit_r100_c59 bl_59 br_59 wl_100 vdd gnd cell_6t
Xbit_r101_c59 bl_59 br_59 wl_101 vdd gnd cell_6t
Xbit_r102_c59 bl_59 br_59 wl_102 vdd gnd cell_6t
Xbit_r103_c59 bl_59 br_59 wl_103 vdd gnd cell_6t
Xbit_r104_c59 bl_59 br_59 wl_104 vdd gnd cell_6t
Xbit_r105_c59 bl_59 br_59 wl_105 vdd gnd cell_6t
Xbit_r106_c59 bl_59 br_59 wl_106 vdd gnd cell_6t
Xbit_r107_c59 bl_59 br_59 wl_107 vdd gnd cell_6t
Xbit_r108_c59 bl_59 br_59 wl_108 vdd gnd cell_6t
Xbit_r109_c59 bl_59 br_59 wl_109 vdd gnd cell_6t
Xbit_r110_c59 bl_59 br_59 wl_110 vdd gnd cell_6t
Xbit_r111_c59 bl_59 br_59 wl_111 vdd gnd cell_6t
Xbit_r112_c59 bl_59 br_59 wl_112 vdd gnd cell_6t
Xbit_r113_c59 bl_59 br_59 wl_113 vdd gnd cell_6t
Xbit_r114_c59 bl_59 br_59 wl_114 vdd gnd cell_6t
Xbit_r115_c59 bl_59 br_59 wl_115 vdd gnd cell_6t
Xbit_r116_c59 bl_59 br_59 wl_116 vdd gnd cell_6t
Xbit_r117_c59 bl_59 br_59 wl_117 vdd gnd cell_6t
Xbit_r118_c59 bl_59 br_59 wl_118 vdd gnd cell_6t
Xbit_r119_c59 bl_59 br_59 wl_119 vdd gnd cell_6t
Xbit_r120_c59 bl_59 br_59 wl_120 vdd gnd cell_6t
Xbit_r121_c59 bl_59 br_59 wl_121 vdd gnd cell_6t
Xbit_r122_c59 bl_59 br_59 wl_122 vdd gnd cell_6t
Xbit_r123_c59 bl_59 br_59 wl_123 vdd gnd cell_6t
Xbit_r124_c59 bl_59 br_59 wl_124 vdd gnd cell_6t
Xbit_r125_c59 bl_59 br_59 wl_125 vdd gnd cell_6t
Xbit_r126_c59 bl_59 br_59 wl_126 vdd gnd cell_6t
Xbit_r127_c59 bl_59 br_59 wl_127 vdd gnd cell_6t
Xbit_r128_c59 bl_59 br_59 wl_128 vdd gnd cell_6t
Xbit_r129_c59 bl_59 br_59 wl_129 vdd gnd cell_6t
Xbit_r130_c59 bl_59 br_59 wl_130 vdd gnd cell_6t
Xbit_r131_c59 bl_59 br_59 wl_131 vdd gnd cell_6t
Xbit_r132_c59 bl_59 br_59 wl_132 vdd gnd cell_6t
Xbit_r133_c59 bl_59 br_59 wl_133 vdd gnd cell_6t
Xbit_r134_c59 bl_59 br_59 wl_134 vdd gnd cell_6t
Xbit_r135_c59 bl_59 br_59 wl_135 vdd gnd cell_6t
Xbit_r136_c59 bl_59 br_59 wl_136 vdd gnd cell_6t
Xbit_r137_c59 bl_59 br_59 wl_137 vdd gnd cell_6t
Xbit_r138_c59 bl_59 br_59 wl_138 vdd gnd cell_6t
Xbit_r139_c59 bl_59 br_59 wl_139 vdd gnd cell_6t
Xbit_r140_c59 bl_59 br_59 wl_140 vdd gnd cell_6t
Xbit_r141_c59 bl_59 br_59 wl_141 vdd gnd cell_6t
Xbit_r142_c59 bl_59 br_59 wl_142 vdd gnd cell_6t
Xbit_r143_c59 bl_59 br_59 wl_143 vdd gnd cell_6t
Xbit_r144_c59 bl_59 br_59 wl_144 vdd gnd cell_6t
Xbit_r145_c59 bl_59 br_59 wl_145 vdd gnd cell_6t
Xbit_r146_c59 bl_59 br_59 wl_146 vdd gnd cell_6t
Xbit_r147_c59 bl_59 br_59 wl_147 vdd gnd cell_6t
Xbit_r148_c59 bl_59 br_59 wl_148 vdd gnd cell_6t
Xbit_r149_c59 bl_59 br_59 wl_149 vdd gnd cell_6t
Xbit_r150_c59 bl_59 br_59 wl_150 vdd gnd cell_6t
Xbit_r151_c59 bl_59 br_59 wl_151 vdd gnd cell_6t
Xbit_r152_c59 bl_59 br_59 wl_152 vdd gnd cell_6t
Xbit_r153_c59 bl_59 br_59 wl_153 vdd gnd cell_6t
Xbit_r154_c59 bl_59 br_59 wl_154 vdd gnd cell_6t
Xbit_r155_c59 bl_59 br_59 wl_155 vdd gnd cell_6t
Xbit_r156_c59 bl_59 br_59 wl_156 vdd gnd cell_6t
Xbit_r157_c59 bl_59 br_59 wl_157 vdd gnd cell_6t
Xbit_r158_c59 bl_59 br_59 wl_158 vdd gnd cell_6t
Xbit_r159_c59 bl_59 br_59 wl_159 vdd gnd cell_6t
Xbit_r160_c59 bl_59 br_59 wl_160 vdd gnd cell_6t
Xbit_r161_c59 bl_59 br_59 wl_161 vdd gnd cell_6t
Xbit_r162_c59 bl_59 br_59 wl_162 vdd gnd cell_6t
Xbit_r163_c59 bl_59 br_59 wl_163 vdd gnd cell_6t
Xbit_r164_c59 bl_59 br_59 wl_164 vdd gnd cell_6t
Xbit_r165_c59 bl_59 br_59 wl_165 vdd gnd cell_6t
Xbit_r166_c59 bl_59 br_59 wl_166 vdd gnd cell_6t
Xbit_r167_c59 bl_59 br_59 wl_167 vdd gnd cell_6t
Xbit_r168_c59 bl_59 br_59 wl_168 vdd gnd cell_6t
Xbit_r169_c59 bl_59 br_59 wl_169 vdd gnd cell_6t
Xbit_r170_c59 bl_59 br_59 wl_170 vdd gnd cell_6t
Xbit_r171_c59 bl_59 br_59 wl_171 vdd gnd cell_6t
Xbit_r172_c59 bl_59 br_59 wl_172 vdd gnd cell_6t
Xbit_r173_c59 bl_59 br_59 wl_173 vdd gnd cell_6t
Xbit_r174_c59 bl_59 br_59 wl_174 vdd gnd cell_6t
Xbit_r175_c59 bl_59 br_59 wl_175 vdd gnd cell_6t
Xbit_r176_c59 bl_59 br_59 wl_176 vdd gnd cell_6t
Xbit_r177_c59 bl_59 br_59 wl_177 vdd gnd cell_6t
Xbit_r178_c59 bl_59 br_59 wl_178 vdd gnd cell_6t
Xbit_r179_c59 bl_59 br_59 wl_179 vdd gnd cell_6t
Xbit_r180_c59 bl_59 br_59 wl_180 vdd gnd cell_6t
Xbit_r181_c59 bl_59 br_59 wl_181 vdd gnd cell_6t
Xbit_r182_c59 bl_59 br_59 wl_182 vdd gnd cell_6t
Xbit_r183_c59 bl_59 br_59 wl_183 vdd gnd cell_6t
Xbit_r184_c59 bl_59 br_59 wl_184 vdd gnd cell_6t
Xbit_r185_c59 bl_59 br_59 wl_185 vdd gnd cell_6t
Xbit_r186_c59 bl_59 br_59 wl_186 vdd gnd cell_6t
Xbit_r187_c59 bl_59 br_59 wl_187 vdd gnd cell_6t
Xbit_r188_c59 bl_59 br_59 wl_188 vdd gnd cell_6t
Xbit_r189_c59 bl_59 br_59 wl_189 vdd gnd cell_6t
Xbit_r190_c59 bl_59 br_59 wl_190 vdd gnd cell_6t
Xbit_r191_c59 bl_59 br_59 wl_191 vdd gnd cell_6t
Xbit_r192_c59 bl_59 br_59 wl_192 vdd gnd cell_6t
Xbit_r193_c59 bl_59 br_59 wl_193 vdd gnd cell_6t
Xbit_r194_c59 bl_59 br_59 wl_194 vdd gnd cell_6t
Xbit_r195_c59 bl_59 br_59 wl_195 vdd gnd cell_6t
Xbit_r196_c59 bl_59 br_59 wl_196 vdd gnd cell_6t
Xbit_r197_c59 bl_59 br_59 wl_197 vdd gnd cell_6t
Xbit_r198_c59 bl_59 br_59 wl_198 vdd gnd cell_6t
Xbit_r199_c59 bl_59 br_59 wl_199 vdd gnd cell_6t
Xbit_r200_c59 bl_59 br_59 wl_200 vdd gnd cell_6t
Xbit_r201_c59 bl_59 br_59 wl_201 vdd gnd cell_6t
Xbit_r202_c59 bl_59 br_59 wl_202 vdd gnd cell_6t
Xbit_r203_c59 bl_59 br_59 wl_203 vdd gnd cell_6t
Xbit_r204_c59 bl_59 br_59 wl_204 vdd gnd cell_6t
Xbit_r205_c59 bl_59 br_59 wl_205 vdd gnd cell_6t
Xbit_r206_c59 bl_59 br_59 wl_206 vdd gnd cell_6t
Xbit_r207_c59 bl_59 br_59 wl_207 vdd gnd cell_6t
Xbit_r208_c59 bl_59 br_59 wl_208 vdd gnd cell_6t
Xbit_r209_c59 bl_59 br_59 wl_209 vdd gnd cell_6t
Xbit_r210_c59 bl_59 br_59 wl_210 vdd gnd cell_6t
Xbit_r211_c59 bl_59 br_59 wl_211 vdd gnd cell_6t
Xbit_r212_c59 bl_59 br_59 wl_212 vdd gnd cell_6t
Xbit_r213_c59 bl_59 br_59 wl_213 vdd gnd cell_6t
Xbit_r214_c59 bl_59 br_59 wl_214 vdd gnd cell_6t
Xbit_r215_c59 bl_59 br_59 wl_215 vdd gnd cell_6t
Xbit_r216_c59 bl_59 br_59 wl_216 vdd gnd cell_6t
Xbit_r217_c59 bl_59 br_59 wl_217 vdd gnd cell_6t
Xbit_r218_c59 bl_59 br_59 wl_218 vdd gnd cell_6t
Xbit_r219_c59 bl_59 br_59 wl_219 vdd gnd cell_6t
Xbit_r220_c59 bl_59 br_59 wl_220 vdd gnd cell_6t
Xbit_r221_c59 bl_59 br_59 wl_221 vdd gnd cell_6t
Xbit_r222_c59 bl_59 br_59 wl_222 vdd gnd cell_6t
Xbit_r223_c59 bl_59 br_59 wl_223 vdd gnd cell_6t
Xbit_r224_c59 bl_59 br_59 wl_224 vdd gnd cell_6t
Xbit_r225_c59 bl_59 br_59 wl_225 vdd gnd cell_6t
Xbit_r226_c59 bl_59 br_59 wl_226 vdd gnd cell_6t
Xbit_r227_c59 bl_59 br_59 wl_227 vdd gnd cell_6t
Xbit_r228_c59 bl_59 br_59 wl_228 vdd gnd cell_6t
Xbit_r229_c59 bl_59 br_59 wl_229 vdd gnd cell_6t
Xbit_r230_c59 bl_59 br_59 wl_230 vdd gnd cell_6t
Xbit_r231_c59 bl_59 br_59 wl_231 vdd gnd cell_6t
Xbit_r232_c59 bl_59 br_59 wl_232 vdd gnd cell_6t
Xbit_r233_c59 bl_59 br_59 wl_233 vdd gnd cell_6t
Xbit_r234_c59 bl_59 br_59 wl_234 vdd gnd cell_6t
Xbit_r235_c59 bl_59 br_59 wl_235 vdd gnd cell_6t
Xbit_r236_c59 bl_59 br_59 wl_236 vdd gnd cell_6t
Xbit_r237_c59 bl_59 br_59 wl_237 vdd gnd cell_6t
Xbit_r238_c59 bl_59 br_59 wl_238 vdd gnd cell_6t
Xbit_r239_c59 bl_59 br_59 wl_239 vdd gnd cell_6t
Xbit_r240_c59 bl_59 br_59 wl_240 vdd gnd cell_6t
Xbit_r241_c59 bl_59 br_59 wl_241 vdd gnd cell_6t
Xbit_r242_c59 bl_59 br_59 wl_242 vdd gnd cell_6t
Xbit_r243_c59 bl_59 br_59 wl_243 vdd gnd cell_6t
Xbit_r244_c59 bl_59 br_59 wl_244 vdd gnd cell_6t
Xbit_r245_c59 bl_59 br_59 wl_245 vdd gnd cell_6t
Xbit_r246_c59 bl_59 br_59 wl_246 vdd gnd cell_6t
Xbit_r247_c59 bl_59 br_59 wl_247 vdd gnd cell_6t
Xbit_r248_c59 bl_59 br_59 wl_248 vdd gnd cell_6t
Xbit_r249_c59 bl_59 br_59 wl_249 vdd gnd cell_6t
Xbit_r250_c59 bl_59 br_59 wl_250 vdd gnd cell_6t
Xbit_r251_c59 bl_59 br_59 wl_251 vdd gnd cell_6t
Xbit_r252_c59 bl_59 br_59 wl_252 vdd gnd cell_6t
Xbit_r253_c59 bl_59 br_59 wl_253 vdd gnd cell_6t
Xbit_r254_c59 bl_59 br_59 wl_254 vdd gnd cell_6t
Xbit_r255_c59 bl_59 br_59 wl_255 vdd gnd cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd cell_6t
Xbit_r1_c60 bl_60 br_60 wl_1 vdd gnd cell_6t
Xbit_r2_c60 bl_60 br_60 wl_2 vdd gnd cell_6t
Xbit_r3_c60 bl_60 br_60 wl_3 vdd gnd cell_6t
Xbit_r4_c60 bl_60 br_60 wl_4 vdd gnd cell_6t
Xbit_r5_c60 bl_60 br_60 wl_5 vdd gnd cell_6t
Xbit_r6_c60 bl_60 br_60 wl_6 vdd gnd cell_6t
Xbit_r7_c60 bl_60 br_60 wl_7 vdd gnd cell_6t
Xbit_r8_c60 bl_60 br_60 wl_8 vdd gnd cell_6t
Xbit_r9_c60 bl_60 br_60 wl_9 vdd gnd cell_6t
Xbit_r10_c60 bl_60 br_60 wl_10 vdd gnd cell_6t
Xbit_r11_c60 bl_60 br_60 wl_11 vdd gnd cell_6t
Xbit_r12_c60 bl_60 br_60 wl_12 vdd gnd cell_6t
Xbit_r13_c60 bl_60 br_60 wl_13 vdd gnd cell_6t
Xbit_r14_c60 bl_60 br_60 wl_14 vdd gnd cell_6t
Xbit_r15_c60 bl_60 br_60 wl_15 vdd gnd cell_6t
Xbit_r16_c60 bl_60 br_60 wl_16 vdd gnd cell_6t
Xbit_r17_c60 bl_60 br_60 wl_17 vdd gnd cell_6t
Xbit_r18_c60 bl_60 br_60 wl_18 vdd gnd cell_6t
Xbit_r19_c60 bl_60 br_60 wl_19 vdd gnd cell_6t
Xbit_r20_c60 bl_60 br_60 wl_20 vdd gnd cell_6t
Xbit_r21_c60 bl_60 br_60 wl_21 vdd gnd cell_6t
Xbit_r22_c60 bl_60 br_60 wl_22 vdd gnd cell_6t
Xbit_r23_c60 bl_60 br_60 wl_23 vdd gnd cell_6t
Xbit_r24_c60 bl_60 br_60 wl_24 vdd gnd cell_6t
Xbit_r25_c60 bl_60 br_60 wl_25 vdd gnd cell_6t
Xbit_r26_c60 bl_60 br_60 wl_26 vdd gnd cell_6t
Xbit_r27_c60 bl_60 br_60 wl_27 vdd gnd cell_6t
Xbit_r28_c60 bl_60 br_60 wl_28 vdd gnd cell_6t
Xbit_r29_c60 bl_60 br_60 wl_29 vdd gnd cell_6t
Xbit_r30_c60 bl_60 br_60 wl_30 vdd gnd cell_6t
Xbit_r31_c60 bl_60 br_60 wl_31 vdd gnd cell_6t
Xbit_r32_c60 bl_60 br_60 wl_32 vdd gnd cell_6t
Xbit_r33_c60 bl_60 br_60 wl_33 vdd gnd cell_6t
Xbit_r34_c60 bl_60 br_60 wl_34 vdd gnd cell_6t
Xbit_r35_c60 bl_60 br_60 wl_35 vdd gnd cell_6t
Xbit_r36_c60 bl_60 br_60 wl_36 vdd gnd cell_6t
Xbit_r37_c60 bl_60 br_60 wl_37 vdd gnd cell_6t
Xbit_r38_c60 bl_60 br_60 wl_38 vdd gnd cell_6t
Xbit_r39_c60 bl_60 br_60 wl_39 vdd gnd cell_6t
Xbit_r40_c60 bl_60 br_60 wl_40 vdd gnd cell_6t
Xbit_r41_c60 bl_60 br_60 wl_41 vdd gnd cell_6t
Xbit_r42_c60 bl_60 br_60 wl_42 vdd gnd cell_6t
Xbit_r43_c60 bl_60 br_60 wl_43 vdd gnd cell_6t
Xbit_r44_c60 bl_60 br_60 wl_44 vdd gnd cell_6t
Xbit_r45_c60 bl_60 br_60 wl_45 vdd gnd cell_6t
Xbit_r46_c60 bl_60 br_60 wl_46 vdd gnd cell_6t
Xbit_r47_c60 bl_60 br_60 wl_47 vdd gnd cell_6t
Xbit_r48_c60 bl_60 br_60 wl_48 vdd gnd cell_6t
Xbit_r49_c60 bl_60 br_60 wl_49 vdd gnd cell_6t
Xbit_r50_c60 bl_60 br_60 wl_50 vdd gnd cell_6t
Xbit_r51_c60 bl_60 br_60 wl_51 vdd gnd cell_6t
Xbit_r52_c60 bl_60 br_60 wl_52 vdd gnd cell_6t
Xbit_r53_c60 bl_60 br_60 wl_53 vdd gnd cell_6t
Xbit_r54_c60 bl_60 br_60 wl_54 vdd gnd cell_6t
Xbit_r55_c60 bl_60 br_60 wl_55 vdd gnd cell_6t
Xbit_r56_c60 bl_60 br_60 wl_56 vdd gnd cell_6t
Xbit_r57_c60 bl_60 br_60 wl_57 vdd gnd cell_6t
Xbit_r58_c60 bl_60 br_60 wl_58 vdd gnd cell_6t
Xbit_r59_c60 bl_60 br_60 wl_59 vdd gnd cell_6t
Xbit_r60_c60 bl_60 br_60 wl_60 vdd gnd cell_6t
Xbit_r61_c60 bl_60 br_60 wl_61 vdd gnd cell_6t
Xbit_r62_c60 bl_60 br_60 wl_62 vdd gnd cell_6t
Xbit_r63_c60 bl_60 br_60 wl_63 vdd gnd cell_6t
Xbit_r64_c60 bl_60 br_60 wl_64 vdd gnd cell_6t
Xbit_r65_c60 bl_60 br_60 wl_65 vdd gnd cell_6t
Xbit_r66_c60 bl_60 br_60 wl_66 vdd gnd cell_6t
Xbit_r67_c60 bl_60 br_60 wl_67 vdd gnd cell_6t
Xbit_r68_c60 bl_60 br_60 wl_68 vdd gnd cell_6t
Xbit_r69_c60 bl_60 br_60 wl_69 vdd gnd cell_6t
Xbit_r70_c60 bl_60 br_60 wl_70 vdd gnd cell_6t
Xbit_r71_c60 bl_60 br_60 wl_71 vdd gnd cell_6t
Xbit_r72_c60 bl_60 br_60 wl_72 vdd gnd cell_6t
Xbit_r73_c60 bl_60 br_60 wl_73 vdd gnd cell_6t
Xbit_r74_c60 bl_60 br_60 wl_74 vdd gnd cell_6t
Xbit_r75_c60 bl_60 br_60 wl_75 vdd gnd cell_6t
Xbit_r76_c60 bl_60 br_60 wl_76 vdd gnd cell_6t
Xbit_r77_c60 bl_60 br_60 wl_77 vdd gnd cell_6t
Xbit_r78_c60 bl_60 br_60 wl_78 vdd gnd cell_6t
Xbit_r79_c60 bl_60 br_60 wl_79 vdd gnd cell_6t
Xbit_r80_c60 bl_60 br_60 wl_80 vdd gnd cell_6t
Xbit_r81_c60 bl_60 br_60 wl_81 vdd gnd cell_6t
Xbit_r82_c60 bl_60 br_60 wl_82 vdd gnd cell_6t
Xbit_r83_c60 bl_60 br_60 wl_83 vdd gnd cell_6t
Xbit_r84_c60 bl_60 br_60 wl_84 vdd gnd cell_6t
Xbit_r85_c60 bl_60 br_60 wl_85 vdd gnd cell_6t
Xbit_r86_c60 bl_60 br_60 wl_86 vdd gnd cell_6t
Xbit_r87_c60 bl_60 br_60 wl_87 vdd gnd cell_6t
Xbit_r88_c60 bl_60 br_60 wl_88 vdd gnd cell_6t
Xbit_r89_c60 bl_60 br_60 wl_89 vdd gnd cell_6t
Xbit_r90_c60 bl_60 br_60 wl_90 vdd gnd cell_6t
Xbit_r91_c60 bl_60 br_60 wl_91 vdd gnd cell_6t
Xbit_r92_c60 bl_60 br_60 wl_92 vdd gnd cell_6t
Xbit_r93_c60 bl_60 br_60 wl_93 vdd gnd cell_6t
Xbit_r94_c60 bl_60 br_60 wl_94 vdd gnd cell_6t
Xbit_r95_c60 bl_60 br_60 wl_95 vdd gnd cell_6t
Xbit_r96_c60 bl_60 br_60 wl_96 vdd gnd cell_6t
Xbit_r97_c60 bl_60 br_60 wl_97 vdd gnd cell_6t
Xbit_r98_c60 bl_60 br_60 wl_98 vdd gnd cell_6t
Xbit_r99_c60 bl_60 br_60 wl_99 vdd gnd cell_6t
Xbit_r100_c60 bl_60 br_60 wl_100 vdd gnd cell_6t
Xbit_r101_c60 bl_60 br_60 wl_101 vdd gnd cell_6t
Xbit_r102_c60 bl_60 br_60 wl_102 vdd gnd cell_6t
Xbit_r103_c60 bl_60 br_60 wl_103 vdd gnd cell_6t
Xbit_r104_c60 bl_60 br_60 wl_104 vdd gnd cell_6t
Xbit_r105_c60 bl_60 br_60 wl_105 vdd gnd cell_6t
Xbit_r106_c60 bl_60 br_60 wl_106 vdd gnd cell_6t
Xbit_r107_c60 bl_60 br_60 wl_107 vdd gnd cell_6t
Xbit_r108_c60 bl_60 br_60 wl_108 vdd gnd cell_6t
Xbit_r109_c60 bl_60 br_60 wl_109 vdd gnd cell_6t
Xbit_r110_c60 bl_60 br_60 wl_110 vdd gnd cell_6t
Xbit_r111_c60 bl_60 br_60 wl_111 vdd gnd cell_6t
Xbit_r112_c60 bl_60 br_60 wl_112 vdd gnd cell_6t
Xbit_r113_c60 bl_60 br_60 wl_113 vdd gnd cell_6t
Xbit_r114_c60 bl_60 br_60 wl_114 vdd gnd cell_6t
Xbit_r115_c60 bl_60 br_60 wl_115 vdd gnd cell_6t
Xbit_r116_c60 bl_60 br_60 wl_116 vdd gnd cell_6t
Xbit_r117_c60 bl_60 br_60 wl_117 vdd gnd cell_6t
Xbit_r118_c60 bl_60 br_60 wl_118 vdd gnd cell_6t
Xbit_r119_c60 bl_60 br_60 wl_119 vdd gnd cell_6t
Xbit_r120_c60 bl_60 br_60 wl_120 vdd gnd cell_6t
Xbit_r121_c60 bl_60 br_60 wl_121 vdd gnd cell_6t
Xbit_r122_c60 bl_60 br_60 wl_122 vdd gnd cell_6t
Xbit_r123_c60 bl_60 br_60 wl_123 vdd gnd cell_6t
Xbit_r124_c60 bl_60 br_60 wl_124 vdd gnd cell_6t
Xbit_r125_c60 bl_60 br_60 wl_125 vdd gnd cell_6t
Xbit_r126_c60 bl_60 br_60 wl_126 vdd gnd cell_6t
Xbit_r127_c60 bl_60 br_60 wl_127 vdd gnd cell_6t
Xbit_r128_c60 bl_60 br_60 wl_128 vdd gnd cell_6t
Xbit_r129_c60 bl_60 br_60 wl_129 vdd gnd cell_6t
Xbit_r130_c60 bl_60 br_60 wl_130 vdd gnd cell_6t
Xbit_r131_c60 bl_60 br_60 wl_131 vdd gnd cell_6t
Xbit_r132_c60 bl_60 br_60 wl_132 vdd gnd cell_6t
Xbit_r133_c60 bl_60 br_60 wl_133 vdd gnd cell_6t
Xbit_r134_c60 bl_60 br_60 wl_134 vdd gnd cell_6t
Xbit_r135_c60 bl_60 br_60 wl_135 vdd gnd cell_6t
Xbit_r136_c60 bl_60 br_60 wl_136 vdd gnd cell_6t
Xbit_r137_c60 bl_60 br_60 wl_137 vdd gnd cell_6t
Xbit_r138_c60 bl_60 br_60 wl_138 vdd gnd cell_6t
Xbit_r139_c60 bl_60 br_60 wl_139 vdd gnd cell_6t
Xbit_r140_c60 bl_60 br_60 wl_140 vdd gnd cell_6t
Xbit_r141_c60 bl_60 br_60 wl_141 vdd gnd cell_6t
Xbit_r142_c60 bl_60 br_60 wl_142 vdd gnd cell_6t
Xbit_r143_c60 bl_60 br_60 wl_143 vdd gnd cell_6t
Xbit_r144_c60 bl_60 br_60 wl_144 vdd gnd cell_6t
Xbit_r145_c60 bl_60 br_60 wl_145 vdd gnd cell_6t
Xbit_r146_c60 bl_60 br_60 wl_146 vdd gnd cell_6t
Xbit_r147_c60 bl_60 br_60 wl_147 vdd gnd cell_6t
Xbit_r148_c60 bl_60 br_60 wl_148 vdd gnd cell_6t
Xbit_r149_c60 bl_60 br_60 wl_149 vdd gnd cell_6t
Xbit_r150_c60 bl_60 br_60 wl_150 vdd gnd cell_6t
Xbit_r151_c60 bl_60 br_60 wl_151 vdd gnd cell_6t
Xbit_r152_c60 bl_60 br_60 wl_152 vdd gnd cell_6t
Xbit_r153_c60 bl_60 br_60 wl_153 vdd gnd cell_6t
Xbit_r154_c60 bl_60 br_60 wl_154 vdd gnd cell_6t
Xbit_r155_c60 bl_60 br_60 wl_155 vdd gnd cell_6t
Xbit_r156_c60 bl_60 br_60 wl_156 vdd gnd cell_6t
Xbit_r157_c60 bl_60 br_60 wl_157 vdd gnd cell_6t
Xbit_r158_c60 bl_60 br_60 wl_158 vdd gnd cell_6t
Xbit_r159_c60 bl_60 br_60 wl_159 vdd gnd cell_6t
Xbit_r160_c60 bl_60 br_60 wl_160 vdd gnd cell_6t
Xbit_r161_c60 bl_60 br_60 wl_161 vdd gnd cell_6t
Xbit_r162_c60 bl_60 br_60 wl_162 vdd gnd cell_6t
Xbit_r163_c60 bl_60 br_60 wl_163 vdd gnd cell_6t
Xbit_r164_c60 bl_60 br_60 wl_164 vdd gnd cell_6t
Xbit_r165_c60 bl_60 br_60 wl_165 vdd gnd cell_6t
Xbit_r166_c60 bl_60 br_60 wl_166 vdd gnd cell_6t
Xbit_r167_c60 bl_60 br_60 wl_167 vdd gnd cell_6t
Xbit_r168_c60 bl_60 br_60 wl_168 vdd gnd cell_6t
Xbit_r169_c60 bl_60 br_60 wl_169 vdd gnd cell_6t
Xbit_r170_c60 bl_60 br_60 wl_170 vdd gnd cell_6t
Xbit_r171_c60 bl_60 br_60 wl_171 vdd gnd cell_6t
Xbit_r172_c60 bl_60 br_60 wl_172 vdd gnd cell_6t
Xbit_r173_c60 bl_60 br_60 wl_173 vdd gnd cell_6t
Xbit_r174_c60 bl_60 br_60 wl_174 vdd gnd cell_6t
Xbit_r175_c60 bl_60 br_60 wl_175 vdd gnd cell_6t
Xbit_r176_c60 bl_60 br_60 wl_176 vdd gnd cell_6t
Xbit_r177_c60 bl_60 br_60 wl_177 vdd gnd cell_6t
Xbit_r178_c60 bl_60 br_60 wl_178 vdd gnd cell_6t
Xbit_r179_c60 bl_60 br_60 wl_179 vdd gnd cell_6t
Xbit_r180_c60 bl_60 br_60 wl_180 vdd gnd cell_6t
Xbit_r181_c60 bl_60 br_60 wl_181 vdd gnd cell_6t
Xbit_r182_c60 bl_60 br_60 wl_182 vdd gnd cell_6t
Xbit_r183_c60 bl_60 br_60 wl_183 vdd gnd cell_6t
Xbit_r184_c60 bl_60 br_60 wl_184 vdd gnd cell_6t
Xbit_r185_c60 bl_60 br_60 wl_185 vdd gnd cell_6t
Xbit_r186_c60 bl_60 br_60 wl_186 vdd gnd cell_6t
Xbit_r187_c60 bl_60 br_60 wl_187 vdd gnd cell_6t
Xbit_r188_c60 bl_60 br_60 wl_188 vdd gnd cell_6t
Xbit_r189_c60 bl_60 br_60 wl_189 vdd gnd cell_6t
Xbit_r190_c60 bl_60 br_60 wl_190 vdd gnd cell_6t
Xbit_r191_c60 bl_60 br_60 wl_191 vdd gnd cell_6t
Xbit_r192_c60 bl_60 br_60 wl_192 vdd gnd cell_6t
Xbit_r193_c60 bl_60 br_60 wl_193 vdd gnd cell_6t
Xbit_r194_c60 bl_60 br_60 wl_194 vdd gnd cell_6t
Xbit_r195_c60 bl_60 br_60 wl_195 vdd gnd cell_6t
Xbit_r196_c60 bl_60 br_60 wl_196 vdd gnd cell_6t
Xbit_r197_c60 bl_60 br_60 wl_197 vdd gnd cell_6t
Xbit_r198_c60 bl_60 br_60 wl_198 vdd gnd cell_6t
Xbit_r199_c60 bl_60 br_60 wl_199 vdd gnd cell_6t
Xbit_r200_c60 bl_60 br_60 wl_200 vdd gnd cell_6t
Xbit_r201_c60 bl_60 br_60 wl_201 vdd gnd cell_6t
Xbit_r202_c60 bl_60 br_60 wl_202 vdd gnd cell_6t
Xbit_r203_c60 bl_60 br_60 wl_203 vdd gnd cell_6t
Xbit_r204_c60 bl_60 br_60 wl_204 vdd gnd cell_6t
Xbit_r205_c60 bl_60 br_60 wl_205 vdd gnd cell_6t
Xbit_r206_c60 bl_60 br_60 wl_206 vdd gnd cell_6t
Xbit_r207_c60 bl_60 br_60 wl_207 vdd gnd cell_6t
Xbit_r208_c60 bl_60 br_60 wl_208 vdd gnd cell_6t
Xbit_r209_c60 bl_60 br_60 wl_209 vdd gnd cell_6t
Xbit_r210_c60 bl_60 br_60 wl_210 vdd gnd cell_6t
Xbit_r211_c60 bl_60 br_60 wl_211 vdd gnd cell_6t
Xbit_r212_c60 bl_60 br_60 wl_212 vdd gnd cell_6t
Xbit_r213_c60 bl_60 br_60 wl_213 vdd gnd cell_6t
Xbit_r214_c60 bl_60 br_60 wl_214 vdd gnd cell_6t
Xbit_r215_c60 bl_60 br_60 wl_215 vdd gnd cell_6t
Xbit_r216_c60 bl_60 br_60 wl_216 vdd gnd cell_6t
Xbit_r217_c60 bl_60 br_60 wl_217 vdd gnd cell_6t
Xbit_r218_c60 bl_60 br_60 wl_218 vdd gnd cell_6t
Xbit_r219_c60 bl_60 br_60 wl_219 vdd gnd cell_6t
Xbit_r220_c60 bl_60 br_60 wl_220 vdd gnd cell_6t
Xbit_r221_c60 bl_60 br_60 wl_221 vdd gnd cell_6t
Xbit_r222_c60 bl_60 br_60 wl_222 vdd gnd cell_6t
Xbit_r223_c60 bl_60 br_60 wl_223 vdd gnd cell_6t
Xbit_r224_c60 bl_60 br_60 wl_224 vdd gnd cell_6t
Xbit_r225_c60 bl_60 br_60 wl_225 vdd gnd cell_6t
Xbit_r226_c60 bl_60 br_60 wl_226 vdd gnd cell_6t
Xbit_r227_c60 bl_60 br_60 wl_227 vdd gnd cell_6t
Xbit_r228_c60 bl_60 br_60 wl_228 vdd gnd cell_6t
Xbit_r229_c60 bl_60 br_60 wl_229 vdd gnd cell_6t
Xbit_r230_c60 bl_60 br_60 wl_230 vdd gnd cell_6t
Xbit_r231_c60 bl_60 br_60 wl_231 vdd gnd cell_6t
Xbit_r232_c60 bl_60 br_60 wl_232 vdd gnd cell_6t
Xbit_r233_c60 bl_60 br_60 wl_233 vdd gnd cell_6t
Xbit_r234_c60 bl_60 br_60 wl_234 vdd gnd cell_6t
Xbit_r235_c60 bl_60 br_60 wl_235 vdd gnd cell_6t
Xbit_r236_c60 bl_60 br_60 wl_236 vdd gnd cell_6t
Xbit_r237_c60 bl_60 br_60 wl_237 vdd gnd cell_6t
Xbit_r238_c60 bl_60 br_60 wl_238 vdd gnd cell_6t
Xbit_r239_c60 bl_60 br_60 wl_239 vdd gnd cell_6t
Xbit_r240_c60 bl_60 br_60 wl_240 vdd gnd cell_6t
Xbit_r241_c60 bl_60 br_60 wl_241 vdd gnd cell_6t
Xbit_r242_c60 bl_60 br_60 wl_242 vdd gnd cell_6t
Xbit_r243_c60 bl_60 br_60 wl_243 vdd gnd cell_6t
Xbit_r244_c60 bl_60 br_60 wl_244 vdd gnd cell_6t
Xbit_r245_c60 bl_60 br_60 wl_245 vdd gnd cell_6t
Xbit_r246_c60 bl_60 br_60 wl_246 vdd gnd cell_6t
Xbit_r247_c60 bl_60 br_60 wl_247 vdd gnd cell_6t
Xbit_r248_c60 bl_60 br_60 wl_248 vdd gnd cell_6t
Xbit_r249_c60 bl_60 br_60 wl_249 vdd gnd cell_6t
Xbit_r250_c60 bl_60 br_60 wl_250 vdd gnd cell_6t
Xbit_r251_c60 bl_60 br_60 wl_251 vdd gnd cell_6t
Xbit_r252_c60 bl_60 br_60 wl_252 vdd gnd cell_6t
Xbit_r253_c60 bl_60 br_60 wl_253 vdd gnd cell_6t
Xbit_r254_c60 bl_60 br_60 wl_254 vdd gnd cell_6t
Xbit_r255_c60 bl_60 br_60 wl_255 vdd gnd cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd cell_6t
Xbit_r1_c61 bl_61 br_61 wl_1 vdd gnd cell_6t
Xbit_r2_c61 bl_61 br_61 wl_2 vdd gnd cell_6t
Xbit_r3_c61 bl_61 br_61 wl_3 vdd gnd cell_6t
Xbit_r4_c61 bl_61 br_61 wl_4 vdd gnd cell_6t
Xbit_r5_c61 bl_61 br_61 wl_5 vdd gnd cell_6t
Xbit_r6_c61 bl_61 br_61 wl_6 vdd gnd cell_6t
Xbit_r7_c61 bl_61 br_61 wl_7 vdd gnd cell_6t
Xbit_r8_c61 bl_61 br_61 wl_8 vdd gnd cell_6t
Xbit_r9_c61 bl_61 br_61 wl_9 vdd gnd cell_6t
Xbit_r10_c61 bl_61 br_61 wl_10 vdd gnd cell_6t
Xbit_r11_c61 bl_61 br_61 wl_11 vdd gnd cell_6t
Xbit_r12_c61 bl_61 br_61 wl_12 vdd gnd cell_6t
Xbit_r13_c61 bl_61 br_61 wl_13 vdd gnd cell_6t
Xbit_r14_c61 bl_61 br_61 wl_14 vdd gnd cell_6t
Xbit_r15_c61 bl_61 br_61 wl_15 vdd gnd cell_6t
Xbit_r16_c61 bl_61 br_61 wl_16 vdd gnd cell_6t
Xbit_r17_c61 bl_61 br_61 wl_17 vdd gnd cell_6t
Xbit_r18_c61 bl_61 br_61 wl_18 vdd gnd cell_6t
Xbit_r19_c61 bl_61 br_61 wl_19 vdd gnd cell_6t
Xbit_r20_c61 bl_61 br_61 wl_20 vdd gnd cell_6t
Xbit_r21_c61 bl_61 br_61 wl_21 vdd gnd cell_6t
Xbit_r22_c61 bl_61 br_61 wl_22 vdd gnd cell_6t
Xbit_r23_c61 bl_61 br_61 wl_23 vdd gnd cell_6t
Xbit_r24_c61 bl_61 br_61 wl_24 vdd gnd cell_6t
Xbit_r25_c61 bl_61 br_61 wl_25 vdd gnd cell_6t
Xbit_r26_c61 bl_61 br_61 wl_26 vdd gnd cell_6t
Xbit_r27_c61 bl_61 br_61 wl_27 vdd gnd cell_6t
Xbit_r28_c61 bl_61 br_61 wl_28 vdd gnd cell_6t
Xbit_r29_c61 bl_61 br_61 wl_29 vdd gnd cell_6t
Xbit_r30_c61 bl_61 br_61 wl_30 vdd gnd cell_6t
Xbit_r31_c61 bl_61 br_61 wl_31 vdd gnd cell_6t
Xbit_r32_c61 bl_61 br_61 wl_32 vdd gnd cell_6t
Xbit_r33_c61 bl_61 br_61 wl_33 vdd gnd cell_6t
Xbit_r34_c61 bl_61 br_61 wl_34 vdd gnd cell_6t
Xbit_r35_c61 bl_61 br_61 wl_35 vdd gnd cell_6t
Xbit_r36_c61 bl_61 br_61 wl_36 vdd gnd cell_6t
Xbit_r37_c61 bl_61 br_61 wl_37 vdd gnd cell_6t
Xbit_r38_c61 bl_61 br_61 wl_38 vdd gnd cell_6t
Xbit_r39_c61 bl_61 br_61 wl_39 vdd gnd cell_6t
Xbit_r40_c61 bl_61 br_61 wl_40 vdd gnd cell_6t
Xbit_r41_c61 bl_61 br_61 wl_41 vdd gnd cell_6t
Xbit_r42_c61 bl_61 br_61 wl_42 vdd gnd cell_6t
Xbit_r43_c61 bl_61 br_61 wl_43 vdd gnd cell_6t
Xbit_r44_c61 bl_61 br_61 wl_44 vdd gnd cell_6t
Xbit_r45_c61 bl_61 br_61 wl_45 vdd gnd cell_6t
Xbit_r46_c61 bl_61 br_61 wl_46 vdd gnd cell_6t
Xbit_r47_c61 bl_61 br_61 wl_47 vdd gnd cell_6t
Xbit_r48_c61 bl_61 br_61 wl_48 vdd gnd cell_6t
Xbit_r49_c61 bl_61 br_61 wl_49 vdd gnd cell_6t
Xbit_r50_c61 bl_61 br_61 wl_50 vdd gnd cell_6t
Xbit_r51_c61 bl_61 br_61 wl_51 vdd gnd cell_6t
Xbit_r52_c61 bl_61 br_61 wl_52 vdd gnd cell_6t
Xbit_r53_c61 bl_61 br_61 wl_53 vdd gnd cell_6t
Xbit_r54_c61 bl_61 br_61 wl_54 vdd gnd cell_6t
Xbit_r55_c61 bl_61 br_61 wl_55 vdd gnd cell_6t
Xbit_r56_c61 bl_61 br_61 wl_56 vdd gnd cell_6t
Xbit_r57_c61 bl_61 br_61 wl_57 vdd gnd cell_6t
Xbit_r58_c61 bl_61 br_61 wl_58 vdd gnd cell_6t
Xbit_r59_c61 bl_61 br_61 wl_59 vdd gnd cell_6t
Xbit_r60_c61 bl_61 br_61 wl_60 vdd gnd cell_6t
Xbit_r61_c61 bl_61 br_61 wl_61 vdd gnd cell_6t
Xbit_r62_c61 bl_61 br_61 wl_62 vdd gnd cell_6t
Xbit_r63_c61 bl_61 br_61 wl_63 vdd gnd cell_6t
Xbit_r64_c61 bl_61 br_61 wl_64 vdd gnd cell_6t
Xbit_r65_c61 bl_61 br_61 wl_65 vdd gnd cell_6t
Xbit_r66_c61 bl_61 br_61 wl_66 vdd gnd cell_6t
Xbit_r67_c61 bl_61 br_61 wl_67 vdd gnd cell_6t
Xbit_r68_c61 bl_61 br_61 wl_68 vdd gnd cell_6t
Xbit_r69_c61 bl_61 br_61 wl_69 vdd gnd cell_6t
Xbit_r70_c61 bl_61 br_61 wl_70 vdd gnd cell_6t
Xbit_r71_c61 bl_61 br_61 wl_71 vdd gnd cell_6t
Xbit_r72_c61 bl_61 br_61 wl_72 vdd gnd cell_6t
Xbit_r73_c61 bl_61 br_61 wl_73 vdd gnd cell_6t
Xbit_r74_c61 bl_61 br_61 wl_74 vdd gnd cell_6t
Xbit_r75_c61 bl_61 br_61 wl_75 vdd gnd cell_6t
Xbit_r76_c61 bl_61 br_61 wl_76 vdd gnd cell_6t
Xbit_r77_c61 bl_61 br_61 wl_77 vdd gnd cell_6t
Xbit_r78_c61 bl_61 br_61 wl_78 vdd gnd cell_6t
Xbit_r79_c61 bl_61 br_61 wl_79 vdd gnd cell_6t
Xbit_r80_c61 bl_61 br_61 wl_80 vdd gnd cell_6t
Xbit_r81_c61 bl_61 br_61 wl_81 vdd gnd cell_6t
Xbit_r82_c61 bl_61 br_61 wl_82 vdd gnd cell_6t
Xbit_r83_c61 bl_61 br_61 wl_83 vdd gnd cell_6t
Xbit_r84_c61 bl_61 br_61 wl_84 vdd gnd cell_6t
Xbit_r85_c61 bl_61 br_61 wl_85 vdd gnd cell_6t
Xbit_r86_c61 bl_61 br_61 wl_86 vdd gnd cell_6t
Xbit_r87_c61 bl_61 br_61 wl_87 vdd gnd cell_6t
Xbit_r88_c61 bl_61 br_61 wl_88 vdd gnd cell_6t
Xbit_r89_c61 bl_61 br_61 wl_89 vdd gnd cell_6t
Xbit_r90_c61 bl_61 br_61 wl_90 vdd gnd cell_6t
Xbit_r91_c61 bl_61 br_61 wl_91 vdd gnd cell_6t
Xbit_r92_c61 bl_61 br_61 wl_92 vdd gnd cell_6t
Xbit_r93_c61 bl_61 br_61 wl_93 vdd gnd cell_6t
Xbit_r94_c61 bl_61 br_61 wl_94 vdd gnd cell_6t
Xbit_r95_c61 bl_61 br_61 wl_95 vdd gnd cell_6t
Xbit_r96_c61 bl_61 br_61 wl_96 vdd gnd cell_6t
Xbit_r97_c61 bl_61 br_61 wl_97 vdd gnd cell_6t
Xbit_r98_c61 bl_61 br_61 wl_98 vdd gnd cell_6t
Xbit_r99_c61 bl_61 br_61 wl_99 vdd gnd cell_6t
Xbit_r100_c61 bl_61 br_61 wl_100 vdd gnd cell_6t
Xbit_r101_c61 bl_61 br_61 wl_101 vdd gnd cell_6t
Xbit_r102_c61 bl_61 br_61 wl_102 vdd gnd cell_6t
Xbit_r103_c61 bl_61 br_61 wl_103 vdd gnd cell_6t
Xbit_r104_c61 bl_61 br_61 wl_104 vdd gnd cell_6t
Xbit_r105_c61 bl_61 br_61 wl_105 vdd gnd cell_6t
Xbit_r106_c61 bl_61 br_61 wl_106 vdd gnd cell_6t
Xbit_r107_c61 bl_61 br_61 wl_107 vdd gnd cell_6t
Xbit_r108_c61 bl_61 br_61 wl_108 vdd gnd cell_6t
Xbit_r109_c61 bl_61 br_61 wl_109 vdd gnd cell_6t
Xbit_r110_c61 bl_61 br_61 wl_110 vdd gnd cell_6t
Xbit_r111_c61 bl_61 br_61 wl_111 vdd gnd cell_6t
Xbit_r112_c61 bl_61 br_61 wl_112 vdd gnd cell_6t
Xbit_r113_c61 bl_61 br_61 wl_113 vdd gnd cell_6t
Xbit_r114_c61 bl_61 br_61 wl_114 vdd gnd cell_6t
Xbit_r115_c61 bl_61 br_61 wl_115 vdd gnd cell_6t
Xbit_r116_c61 bl_61 br_61 wl_116 vdd gnd cell_6t
Xbit_r117_c61 bl_61 br_61 wl_117 vdd gnd cell_6t
Xbit_r118_c61 bl_61 br_61 wl_118 vdd gnd cell_6t
Xbit_r119_c61 bl_61 br_61 wl_119 vdd gnd cell_6t
Xbit_r120_c61 bl_61 br_61 wl_120 vdd gnd cell_6t
Xbit_r121_c61 bl_61 br_61 wl_121 vdd gnd cell_6t
Xbit_r122_c61 bl_61 br_61 wl_122 vdd gnd cell_6t
Xbit_r123_c61 bl_61 br_61 wl_123 vdd gnd cell_6t
Xbit_r124_c61 bl_61 br_61 wl_124 vdd gnd cell_6t
Xbit_r125_c61 bl_61 br_61 wl_125 vdd gnd cell_6t
Xbit_r126_c61 bl_61 br_61 wl_126 vdd gnd cell_6t
Xbit_r127_c61 bl_61 br_61 wl_127 vdd gnd cell_6t
Xbit_r128_c61 bl_61 br_61 wl_128 vdd gnd cell_6t
Xbit_r129_c61 bl_61 br_61 wl_129 vdd gnd cell_6t
Xbit_r130_c61 bl_61 br_61 wl_130 vdd gnd cell_6t
Xbit_r131_c61 bl_61 br_61 wl_131 vdd gnd cell_6t
Xbit_r132_c61 bl_61 br_61 wl_132 vdd gnd cell_6t
Xbit_r133_c61 bl_61 br_61 wl_133 vdd gnd cell_6t
Xbit_r134_c61 bl_61 br_61 wl_134 vdd gnd cell_6t
Xbit_r135_c61 bl_61 br_61 wl_135 vdd gnd cell_6t
Xbit_r136_c61 bl_61 br_61 wl_136 vdd gnd cell_6t
Xbit_r137_c61 bl_61 br_61 wl_137 vdd gnd cell_6t
Xbit_r138_c61 bl_61 br_61 wl_138 vdd gnd cell_6t
Xbit_r139_c61 bl_61 br_61 wl_139 vdd gnd cell_6t
Xbit_r140_c61 bl_61 br_61 wl_140 vdd gnd cell_6t
Xbit_r141_c61 bl_61 br_61 wl_141 vdd gnd cell_6t
Xbit_r142_c61 bl_61 br_61 wl_142 vdd gnd cell_6t
Xbit_r143_c61 bl_61 br_61 wl_143 vdd gnd cell_6t
Xbit_r144_c61 bl_61 br_61 wl_144 vdd gnd cell_6t
Xbit_r145_c61 bl_61 br_61 wl_145 vdd gnd cell_6t
Xbit_r146_c61 bl_61 br_61 wl_146 vdd gnd cell_6t
Xbit_r147_c61 bl_61 br_61 wl_147 vdd gnd cell_6t
Xbit_r148_c61 bl_61 br_61 wl_148 vdd gnd cell_6t
Xbit_r149_c61 bl_61 br_61 wl_149 vdd gnd cell_6t
Xbit_r150_c61 bl_61 br_61 wl_150 vdd gnd cell_6t
Xbit_r151_c61 bl_61 br_61 wl_151 vdd gnd cell_6t
Xbit_r152_c61 bl_61 br_61 wl_152 vdd gnd cell_6t
Xbit_r153_c61 bl_61 br_61 wl_153 vdd gnd cell_6t
Xbit_r154_c61 bl_61 br_61 wl_154 vdd gnd cell_6t
Xbit_r155_c61 bl_61 br_61 wl_155 vdd gnd cell_6t
Xbit_r156_c61 bl_61 br_61 wl_156 vdd gnd cell_6t
Xbit_r157_c61 bl_61 br_61 wl_157 vdd gnd cell_6t
Xbit_r158_c61 bl_61 br_61 wl_158 vdd gnd cell_6t
Xbit_r159_c61 bl_61 br_61 wl_159 vdd gnd cell_6t
Xbit_r160_c61 bl_61 br_61 wl_160 vdd gnd cell_6t
Xbit_r161_c61 bl_61 br_61 wl_161 vdd gnd cell_6t
Xbit_r162_c61 bl_61 br_61 wl_162 vdd gnd cell_6t
Xbit_r163_c61 bl_61 br_61 wl_163 vdd gnd cell_6t
Xbit_r164_c61 bl_61 br_61 wl_164 vdd gnd cell_6t
Xbit_r165_c61 bl_61 br_61 wl_165 vdd gnd cell_6t
Xbit_r166_c61 bl_61 br_61 wl_166 vdd gnd cell_6t
Xbit_r167_c61 bl_61 br_61 wl_167 vdd gnd cell_6t
Xbit_r168_c61 bl_61 br_61 wl_168 vdd gnd cell_6t
Xbit_r169_c61 bl_61 br_61 wl_169 vdd gnd cell_6t
Xbit_r170_c61 bl_61 br_61 wl_170 vdd gnd cell_6t
Xbit_r171_c61 bl_61 br_61 wl_171 vdd gnd cell_6t
Xbit_r172_c61 bl_61 br_61 wl_172 vdd gnd cell_6t
Xbit_r173_c61 bl_61 br_61 wl_173 vdd gnd cell_6t
Xbit_r174_c61 bl_61 br_61 wl_174 vdd gnd cell_6t
Xbit_r175_c61 bl_61 br_61 wl_175 vdd gnd cell_6t
Xbit_r176_c61 bl_61 br_61 wl_176 vdd gnd cell_6t
Xbit_r177_c61 bl_61 br_61 wl_177 vdd gnd cell_6t
Xbit_r178_c61 bl_61 br_61 wl_178 vdd gnd cell_6t
Xbit_r179_c61 bl_61 br_61 wl_179 vdd gnd cell_6t
Xbit_r180_c61 bl_61 br_61 wl_180 vdd gnd cell_6t
Xbit_r181_c61 bl_61 br_61 wl_181 vdd gnd cell_6t
Xbit_r182_c61 bl_61 br_61 wl_182 vdd gnd cell_6t
Xbit_r183_c61 bl_61 br_61 wl_183 vdd gnd cell_6t
Xbit_r184_c61 bl_61 br_61 wl_184 vdd gnd cell_6t
Xbit_r185_c61 bl_61 br_61 wl_185 vdd gnd cell_6t
Xbit_r186_c61 bl_61 br_61 wl_186 vdd gnd cell_6t
Xbit_r187_c61 bl_61 br_61 wl_187 vdd gnd cell_6t
Xbit_r188_c61 bl_61 br_61 wl_188 vdd gnd cell_6t
Xbit_r189_c61 bl_61 br_61 wl_189 vdd gnd cell_6t
Xbit_r190_c61 bl_61 br_61 wl_190 vdd gnd cell_6t
Xbit_r191_c61 bl_61 br_61 wl_191 vdd gnd cell_6t
Xbit_r192_c61 bl_61 br_61 wl_192 vdd gnd cell_6t
Xbit_r193_c61 bl_61 br_61 wl_193 vdd gnd cell_6t
Xbit_r194_c61 bl_61 br_61 wl_194 vdd gnd cell_6t
Xbit_r195_c61 bl_61 br_61 wl_195 vdd gnd cell_6t
Xbit_r196_c61 bl_61 br_61 wl_196 vdd gnd cell_6t
Xbit_r197_c61 bl_61 br_61 wl_197 vdd gnd cell_6t
Xbit_r198_c61 bl_61 br_61 wl_198 vdd gnd cell_6t
Xbit_r199_c61 bl_61 br_61 wl_199 vdd gnd cell_6t
Xbit_r200_c61 bl_61 br_61 wl_200 vdd gnd cell_6t
Xbit_r201_c61 bl_61 br_61 wl_201 vdd gnd cell_6t
Xbit_r202_c61 bl_61 br_61 wl_202 vdd gnd cell_6t
Xbit_r203_c61 bl_61 br_61 wl_203 vdd gnd cell_6t
Xbit_r204_c61 bl_61 br_61 wl_204 vdd gnd cell_6t
Xbit_r205_c61 bl_61 br_61 wl_205 vdd gnd cell_6t
Xbit_r206_c61 bl_61 br_61 wl_206 vdd gnd cell_6t
Xbit_r207_c61 bl_61 br_61 wl_207 vdd gnd cell_6t
Xbit_r208_c61 bl_61 br_61 wl_208 vdd gnd cell_6t
Xbit_r209_c61 bl_61 br_61 wl_209 vdd gnd cell_6t
Xbit_r210_c61 bl_61 br_61 wl_210 vdd gnd cell_6t
Xbit_r211_c61 bl_61 br_61 wl_211 vdd gnd cell_6t
Xbit_r212_c61 bl_61 br_61 wl_212 vdd gnd cell_6t
Xbit_r213_c61 bl_61 br_61 wl_213 vdd gnd cell_6t
Xbit_r214_c61 bl_61 br_61 wl_214 vdd gnd cell_6t
Xbit_r215_c61 bl_61 br_61 wl_215 vdd gnd cell_6t
Xbit_r216_c61 bl_61 br_61 wl_216 vdd gnd cell_6t
Xbit_r217_c61 bl_61 br_61 wl_217 vdd gnd cell_6t
Xbit_r218_c61 bl_61 br_61 wl_218 vdd gnd cell_6t
Xbit_r219_c61 bl_61 br_61 wl_219 vdd gnd cell_6t
Xbit_r220_c61 bl_61 br_61 wl_220 vdd gnd cell_6t
Xbit_r221_c61 bl_61 br_61 wl_221 vdd gnd cell_6t
Xbit_r222_c61 bl_61 br_61 wl_222 vdd gnd cell_6t
Xbit_r223_c61 bl_61 br_61 wl_223 vdd gnd cell_6t
Xbit_r224_c61 bl_61 br_61 wl_224 vdd gnd cell_6t
Xbit_r225_c61 bl_61 br_61 wl_225 vdd gnd cell_6t
Xbit_r226_c61 bl_61 br_61 wl_226 vdd gnd cell_6t
Xbit_r227_c61 bl_61 br_61 wl_227 vdd gnd cell_6t
Xbit_r228_c61 bl_61 br_61 wl_228 vdd gnd cell_6t
Xbit_r229_c61 bl_61 br_61 wl_229 vdd gnd cell_6t
Xbit_r230_c61 bl_61 br_61 wl_230 vdd gnd cell_6t
Xbit_r231_c61 bl_61 br_61 wl_231 vdd gnd cell_6t
Xbit_r232_c61 bl_61 br_61 wl_232 vdd gnd cell_6t
Xbit_r233_c61 bl_61 br_61 wl_233 vdd gnd cell_6t
Xbit_r234_c61 bl_61 br_61 wl_234 vdd gnd cell_6t
Xbit_r235_c61 bl_61 br_61 wl_235 vdd gnd cell_6t
Xbit_r236_c61 bl_61 br_61 wl_236 vdd gnd cell_6t
Xbit_r237_c61 bl_61 br_61 wl_237 vdd gnd cell_6t
Xbit_r238_c61 bl_61 br_61 wl_238 vdd gnd cell_6t
Xbit_r239_c61 bl_61 br_61 wl_239 vdd gnd cell_6t
Xbit_r240_c61 bl_61 br_61 wl_240 vdd gnd cell_6t
Xbit_r241_c61 bl_61 br_61 wl_241 vdd gnd cell_6t
Xbit_r242_c61 bl_61 br_61 wl_242 vdd gnd cell_6t
Xbit_r243_c61 bl_61 br_61 wl_243 vdd gnd cell_6t
Xbit_r244_c61 bl_61 br_61 wl_244 vdd gnd cell_6t
Xbit_r245_c61 bl_61 br_61 wl_245 vdd gnd cell_6t
Xbit_r246_c61 bl_61 br_61 wl_246 vdd gnd cell_6t
Xbit_r247_c61 bl_61 br_61 wl_247 vdd gnd cell_6t
Xbit_r248_c61 bl_61 br_61 wl_248 vdd gnd cell_6t
Xbit_r249_c61 bl_61 br_61 wl_249 vdd gnd cell_6t
Xbit_r250_c61 bl_61 br_61 wl_250 vdd gnd cell_6t
Xbit_r251_c61 bl_61 br_61 wl_251 vdd gnd cell_6t
Xbit_r252_c61 bl_61 br_61 wl_252 vdd gnd cell_6t
Xbit_r253_c61 bl_61 br_61 wl_253 vdd gnd cell_6t
Xbit_r254_c61 bl_61 br_61 wl_254 vdd gnd cell_6t
Xbit_r255_c61 bl_61 br_61 wl_255 vdd gnd cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd cell_6t
Xbit_r1_c62 bl_62 br_62 wl_1 vdd gnd cell_6t
Xbit_r2_c62 bl_62 br_62 wl_2 vdd gnd cell_6t
Xbit_r3_c62 bl_62 br_62 wl_3 vdd gnd cell_6t
Xbit_r4_c62 bl_62 br_62 wl_4 vdd gnd cell_6t
Xbit_r5_c62 bl_62 br_62 wl_5 vdd gnd cell_6t
Xbit_r6_c62 bl_62 br_62 wl_6 vdd gnd cell_6t
Xbit_r7_c62 bl_62 br_62 wl_7 vdd gnd cell_6t
Xbit_r8_c62 bl_62 br_62 wl_8 vdd gnd cell_6t
Xbit_r9_c62 bl_62 br_62 wl_9 vdd gnd cell_6t
Xbit_r10_c62 bl_62 br_62 wl_10 vdd gnd cell_6t
Xbit_r11_c62 bl_62 br_62 wl_11 vdd gnd cell_6t
Xbit_r12_c62 bl_62 br_62 wl_12 vdd gnd cell_6t
Xbit_r13_c62 bl_62 br_62 wl_13 vdd gnd cell_6t
Xbit_r14_c62 bl_62 br_62 wl_14 vdd gnd cell_6t
Xbit_r15_c62 bl_62 br_62 wl_15 vdd gnd cell_6t
Xbit_r16_c62 bl_62 br_62 wl_16 vdd gnd cell_6t
Xbit_r17_c62 bl_62 br_62 wl_17 vdd gnd cell_6t
Xbit_r18_c62 bl_62 br_62 wl_18 vdd gnd cell_6t
Xbit_r19_c62 bl_62 br_62 wl_19 vdd gnd cell_6t
Xbit_r20_c62 bl_62 br_62 wl_20 vdd gnd cell_6t
Xbit_r21_c62 bl_62 br_62 wl_21 vdd gnd cell_6t
Xbit_r22_c62 bl_62 br_62 wl_22 vdd gnd cell_6t
Xbit_r23_c62 bl_62 br_62 wl_23 vdd gnd cell_6t
Xbit_r24_c62 bl_62 br_62 wl_24 vdd gnd cell_6t
Xbit_r25_c62 bl_62 br_62 wl_25 vdd gnd cell_6t
Xbit_r26_c62 bl_62 br_62 wl_26 vdd gnd cell_6t
Xbit_r27_c62 bl_62 br_62 wl_27 vdd gnd cell_6t
Xbit_r28_c62 bl_62 br_62 wl_28 vdd gnd cell_6t
Xbit_r29_c62 bl_62 br_62 wl_29 vdd gnd cell_6t
Xbit_r30_c62 bl_62 br_62 wl_30 vdd gnd cell_6t
Xbit_r31_c62 bl_62 br_62 wl_31 vdd gnd cell_6t
Xbit_r32_c62 bl_62 br_62 wl_32 vdd gnd cell_6t
Xbit_r33_c62 bl_62 br_62 wl_33 vdd gnd cell_6t
Xbit_r34_c62 bl_62 br_62 wl_34 vdd gnd cell_6t
Xbit_r35_c62 bl_62 br_62 wl_35 vdd gnd cell_6t
Xbit_r36_c62 bl_62 br_62 wl_36 vdd gnd cell_6t
Xbit_r37_c62 bl_62 br_62 wl_37 vdd gnd cell_6t
Xbit_r38_c62 bl_62 br_62 wl_38 vdd gnd cell_6t
Xbit_r39_c62 bl_62 br_62 wl_39 vdd gnd cell_6t
Xbit_r40_c62 bl_62 br_62 wl_40 vdd gnd cell_6t
Xbit_r41_c62 bl_62 br_62 wl_41 vdd gnd cell_6t
Xbit_r42_c62 bl_62 br_62 wl_42 vdd gnd cell_6t
Xbit_r43_c62 bl_62 br_62 wl_43 vdd gnd cell_6t
Xbit_r44_c62 bl_62 br_62 wl_44 vdd gnd cell_6t
Xbit_r45_c62 bl_62 br_62 wl_45 vdd gnd cell_6t
Xbit_r46_c62 bl_62 br_62 wl_46 vdd gnd cell_6t
Xbit_r47_c62 bl_62 br_62 wl_47 vdd gnd cell_6t
Xbit_r48_c62 bl_62 br_62 wl_48 vdd gnd cell_6t
Xbit_r49_c62 bl_62 br_62 wl_49 vdd gnd cell_6t
Xbit_r50_c62 bl_62 br_62 wl_50 vdd gnd cell_6t
Xbit_r51_c62 bl_62 br_62 wl_51 vdd gnd cell_6t
Xbit_r52_c62 bl_62 br_62 wl_52 vdd gnd cell_6t
Xbit_r53_c62 bl_62 br_62 wl_53 vdd gnd cell_6t
Xbit_r54_c62 bl_62 br_62 wl_54 vdd gnd cell_6t
Xbit_r55_c62 bl_62 br_62 wl_55 vdd gnd cell_6t
Xbit_r56_c62 bl_62 br_62 wl_56 vdd gnd cell_6t
Xbit_r57_c62 bl_62 br_62 wl_57 vdd gnd cell_6t
Xbit_r58_c62 bl_62 br_62 wl_58 vdd gnd cell_6t
Xbit_r59_c62 bl_62 br_62 wl_59 vdd gnd cell_6t
Xbit_r60_c62 bl_62 br_62 wl_60 vdd gnd cell_6t
Xbit_r61_c62 bl_62 br_62 wl_61 vdd gnd cell_6t
Xbit_r62_c62 bl_62 br_62 wl_62 vdd gnd cell_6t
Xbit_r63_c62 bl_62 br_62 wl_63 vdd gnd cell_6t
Xbit_r64_c62 bl_62 br_62 wl_64 vdd gnd cell_6t
Xbit_r65_c62 bl_62 br_62 wl_65 vdd gnd cell_6t
Xbit_r66_c62 bl_62 br_62 wl_66 vdd gnd cell_6t
Xbit_r67_c62 bl_62 br_62 wl_67 vdd gnd cell_6t
Xbit_r68_c62 bl_62 br_62 wl_68 vdd gnd cell_6t
Xbit_r69_c62 bl_62 br_62 wl_69 vdd gnd cell_6t
Xbit_r70_c62 bl_62 br_62 wl_70 vdd gnd cell_6t
Xbit_r71_c62 bl_62 br_62 wl_71 vdd gnd cell_6t
Xbit_r72_c62 bl_62 br_62 wl_72 vdd gnd cell_6t
Xbit_r73_c62 bl_62 br_62 wl_73 vdd gnd cell_6t
Xbit_r74_c62 bl_62 br_62 wl_74 vdd gnd cell_6t
Xbit_r75_c62 bl_62 br_62 wl_75 vdd gnd cell_6t
Xbit_r76_c62 bl_62 br_62 wl_76 vdd gnd cell_6t
Xbit_r77_c62 bl_62 br_62 wl_77 vdd gnd cell_6t
Xbit_r78_c62 bl_62 br_62 wl_78 vdd gnd cell_6t
Xbit_r79_c62 bl_62 br_62 wl_79 vdd gnd cell_6t
Xbit_r80_c62 bl_62 br_62 wl_80 vdd gnd cell_6t
Xbit_r81_c62 bl_62 br_62 wl_81 vdd gnd cell_6t
Xbit_r82_c62 bl_62 br_62 wl_82 vdd gnd cell_6t
Xbit_r83_c62 bl_62 br_62 wl_83 vdd gnd cell_6t
Xbit_r84_c62 bl_62 br_62 wl_84 vdd gnd cell_6t
Xbit_r85_c62 bl_62 br_62 wl_85 vdd gnd cell_6t
Xbit_r86_c62 bl_62 br_62 wl_86 vdd gnd cell_6t
Xbit_r87_c62 bl_62 br_62 wl_87 vdd gnd cell_6t
Xbit_r88_c62 bl_62 br_62 wl_88 vdd gnd cell_6t
Xbit_r89_c62 bl_62 br_62 wl_89 vdd gnd cell_6t
Xbit_r90_c62 bl_62 br_62 wl_90 vdd gnd cell_6t
Xbit_r91_c62 bl_62 br_62 wl_91 vdd gnd cell_6t
Xbit_r92_c62 bl_62 br_62 wl_92 vdd gnd cell_6t
Xbit_r93_c62 bl_62 br_62 wl_93 vdd gnd cell_6t
Xbit_r94_c62 bl_62 br_62 wl_94 vdd gnd cell_6t
Xbit_r95_c62 bl_62 br_62 wl_95 vdd gnd cell_6t
Xbit_r96_c62 bl_62 br_62 wl_96 vdd gnd cell_6t
Xbit_r97_c62 bl_62 br_62 wl_97 vdd gnd cell_6t
Xbit_r98_c62 bl_62 br_62 wl_98 vdd gnd cell_6t
Xbit_r99_c62 bl_62 br_62 wl_99 vdd gnd cell_6t
Xbit_r100_c62 bl_62 br_62 wl_100 vdd gnd cell_6t
Xbit_r101_c62 bl_62 br_62 wl_101 vdd gnd cell_6t
Xbit_r102_c62 bl_62 br_62 wl_102 vdd gnd cell_6t
Xbit_r103_c62 bl_62 br_62 wl_103 vdd gnd cell_6t
Xbit_r104_c62 bl_62 br_62 wl_104 vdd gnd cell_6t
Xbit_r105_c62 bl_62 br_62 wl_105 vdd gnd cell_6t
Xbit_r106_c62 bl_62 br_62 wl_106 vdd gnd cell_6t
Xbit_r107_c62 bl_62 br_62 wl_107 vdd gnd cell_6t
Xbit_r108_c62 bl_62 br_62 wl_108 vdd gnd cell_6t
Xbit_r109_c62 bl_62 br_62 wl_109 vdd gnd cell_6t
Xbit_r110_c62 bl_62 br_62 wl_110 vdd gnd cell_6t
Xbit_r111_c62 bl_62 br_62 wl_111 vdd gnd cell_6t
Xbit_r112_c62 bl_62 br_62 wl_112 vdd gnd cell_6t
Xbit_r113_c62 bl_62 br_62 wl_113 vdd gnd cell_6t
Xbit_r114_c62 bl_62 br_62 wl_114 vdd gnd cell_6t
Xbit_r115_c62 bl_62 br_62 wl_115 vdd gnd cell_6t
Xbit_r116_c62 bl_62 br_62 wl_116 vdd gnd cell_6t
Xbit_r117_c62 bl_62 br_62 wl_117 vdd gnd cell_6t
Xbit_r118_c62 bl_62 br_62 wl_118 vdd gnd cell_6t
Xbit_r119_c62 bl_62 br_62 wl_119 vdd gnd cell_6t
Xbit_r120_c62 bl_62 br_62 wl_120 vdd gnd cell_6t
Xbit_r121_c62 bl_62 br_62 wl_121 vdd gnd cell_6t
Xbit_r122_c62 bl_62 br_62 wl_122 vdd gnd cell_6t
Xbit_r123_c62 bl_62 br_62 wl_123 vdd gnd cell_6t
Xbit_r124_c62 bl_62 br_62 wl_124 vdd gnd cell_6t
Xbit_r125_c62 bl_62 br_62 wl_125 vdd gnd cell_6t
Xbit_r126_c62 bl_62 br_62 wl_126 vdd gnd cell_6t
Xbit_r127_c62 bl_62 br_62 wl_127 vdd gnd cell_6t
Xbit_r128_c62 bl_62 br_62 wl_128 vdd gnd cell_6t
Xbit_r129_c62 bl_62 br_62 wl_129 vdd gnd cell_6t
Xbit_r130_c62 bl_62 br_62 wl_130 vdd gnd cell_6t
Xbit_r131_c62 bl_62 br_62 wl_131 vdd gnd cell_6t
Xbit_r132_c62 bl_62 br_62 wl_132 vdd gnd cell_6t
Xbit_r133_c62 bl_62 br_62 wl_133 vdd gnd cell_6t
Xbit_r134_c62 bl_62 br_62 wl_134 vdd gnd cell_6t
Xbit_r135_c62 bl_62 br_62 wl_135 vdd gnd cell_6t
Xbit_r136_c62 bl_62 br_62 wl_136 vdd gnd cell_6t
Xbit_r137_c62 bl_62 br_62 wl_137 vdd gnd cell_6t
Xbit_r138_c62 bl_62 br_62 wl_138 vdd gnd cell_6t
Xbit_r139_c62 bl_62 br_62 wl_139 vdd gnd cell_6t
Xbit_r140_c62 bl_62 br_62 wl_140 vdd gnd cell_6t
Xbit_r141_c62 bl_62 br_62 wl_141 vdd gnd cell_6t
Xbit_r142_c62 bl_62 br_62 wl_142 vdd gnd cell_6t
Xbit_r143_c62 bl_62 br_62 wl_143 vdd gnd cell_6t
Xbit_r144_c62 bl_62 br_62 wl_144 vdd gnd cell_6t
Xbit_r145_c62 bl_62 br_62 wl_145 vdd gnd cell_6t
Xbit_r146_c62 bl_62 br_62 wl_146 vdd gnd cell_6t
Xbit_r147_c62 bl_62 br_62 wl_147 vdd gnd cell_6t
Xbit_r148_c62 bl_62 br_62 wl_148 vdd gnd cell_6t
Xbit_r149_c62 bl_62 br_62 wl_149 vdd gnd cell_6t
Xbit_r150_c62 bl_62 br_62 wl_150 vdd gnd cell_6t
Xbit_r151_c62 bl_62 br_62 wl_151 vdd gnd cell_6t
Xbit_r152_c62 bl_62 br_62 wl_152 vdd gnd cell_6t
Xbit_r153_c62 bl_62 br_62 wl_153 vdd gnd cell_6t
Xbit_r154_c62 bl_62 br_62 wl_154 vdd gnd cell_6t
Xbit_r155_c62 bl_62 br_62 wl_155 vdd gnd cell_6t
Xbit_r156_c62 bl_62 br_62 wl_156 vdd gnd cell_6t
Xbit_r157_c62 bl_62 br_62 wl_157 vdd gnd cell_6t
Xbit_r158_c62 bl_62 br_62 wl_158 vdd gnd cell_6t
Xbit_r159_c62 bl_62 br_62 wl_159 vdd gnd cell_6t
Xbit_r160_c62 bl_62 br_62 wl_160 vdd gnd cell_6t
Xbit_r161_c62 bl_62 br_62 wl_161 vdd gnd cell_6t
Xbit_r162_c62 bl_62 br_62 wl_162 vdd gnd cell_6t
Xbit_r163_c62 bl_62 br_62 wl_163 vdd gnd cell_6t
Xbit_r164_c62 bl_62 br_62 wl_164 vdd gnd cell_6t
Xbit_r165_c62 bl_62 br_62 wl_165 vdd gnd cell_6t
Xbit_r166_c62 bl_62 br_62 wl_166 vdd gnd cell_6t
Xbit_r167_c62 bl_62 br_62 wl_167 vdd gnd cell_6t
Xbit_r168_c62 bl_62 br_62 wl_168 vdd gnd cell_6t
Xbit_r169_c62 bl_62 br_62 wl_169 vdd gnd cell_6t
Xbit_r170_c62 bl_62 br_62 wl_170 vdd gnd cell_6t
Xbit_r171_c62 bl_62 br_62 wl_171 vdd gnd cell_6t
Xbit_r172_c62 bl_62 br_62 wl_172 vdd gnd cell_6t
Xbit_r173_c62 bl_62 br_62 wl_173 vdd gnd cell_6t
Xbit_r174_c62 bl_62 br_62 wl_174 vdd gnd cell_6t
Xbit_r175_c62 bl_62 br_62 wl_175 vdd gnd cell_6t
Xbit_r176_c62 bl_62 br_62 wl_176 vdd gnd cell_6t
Xbit_r177_c62 bl_62 br_62 wl_177 vdd gnd cell_6t
Xbit_r178_c62 bl_62 br_62 wl_178 vdd gnd cell_6t
Xbit_r179_c62 bl_62 br_62 wl_179 vdd gnd cell_6t
Xbit_r180_c62 bl_62 br_62 wl_180 vdd gnd cell_6t
Xbit_r181_c62 bl_62 br_62 wl_181 vdd gnd cell_6t
Xbit_r182_c62 bl_62 br_62 wl_182 vdd gnd cell_6t
Xbit_r183_c62 bl_62 br_62 wl_183 vdd gnd cell_6t
Xbit_r184_c62 bl_62 br_62 wl_184 vdd gnd cell_6t
Xbit_r185_c62 bl_62 br_62 wl_185 vdd gnd cell_6t
Xbit_r186_c62 bl_62 br_62 wl_186 vdd gnd cell_6t
Xbit_r187_c62 bl_62 br_62 wl_187 vdd gnd cell_6t
Xbit_r188_c62 bl_62 br_62 wl_188 vdd gnd cell_6t
Xbit_r189_c62 bl_62 br_62 wl_189 vdd gnd cell_6t
Xbit_r190_c62 bl_62 br_62 wl_190 vdd gnd cell_6t
Xbit_r191_c62 bl_62 br_62 wl_191 vdd gnd cell_6t
Xbit_r192_c62 bl_62 br_62 wl_192 vdd gnd cell_6t
Xbit_r193_c62 bl_62 br_62 wl_193 vdd gnd cell_6t
Xbit_r194_c62 bl_62 br_62 wl_194 vdd gnd cell_6t
Xbit_r195_c62 bl_62 br_62 wl_195 vdd gnd cell_6t
Xbit_r196_c62 bl_62 br_62 wl_196 vdd gnd cell_6t
Xbit_r197_c62 bl_62 br_62 wl_197 vdd gnd cell_6t
Xbit_r198_c62 bl_62 br_62 wl_198 vdd gnd cell_6t
Xbit_r199_c62 bl_62 br_62 wl_199 vdd gnd cell_6t
Xbit_r200_c62 bl_62 br_62 wl_200 vdd gnd cell_6t
Xbit_r201_c62 bl_62 br_62 wl_201 vdd gnd cell_6t
Xbit_r202_c62 bl_62 br_62 wl_202 vdd gnd cell_6t
Xbit_r203_c62 bl_62 br_62 wl_203 vdd gnd cell_6t
Xbit_r204_c62 bl_62 br_62 wl_204 vdd gnd cell_6t
Xbit_r205_c62 bl_62 br_62 wl_205 vdd gnd cell_6t
Xbit_r206_c62 bl_62 br_62 wl_206 vdd gnd cell_6t
Xbit_r207_c62 bl_62 br_62 wl_207 vdd gnd cell_6t
Xbit_r208_c62 bl_62 br_62 wl_208 vdd gnd cell_6t
Xbit_r209_c62 bl_62 br_62 wl_209 vdd gnd cell_6t
Xbit_r210_c62 bl_62 br_62 wl_210 vdd gnd cell_6t
Xbit_r211_c62 bl_62 br_62 wl_211 vdd gnd cell_6t
Xbit_r212_c62 bl_62 br_62 wl_212 vdd gnd cell_6t
Xbit_r213_c62 bl_62 br_62 wl_213 vdd gnd cell_6t
Xbit_r214_c62 bl_62 br_62 wl_214 vdd gnd cell_6t
Xbit_r215_c62 bl_62 br_62 wl_215 vdd gnd cell_6t
Xbit_r216_c62 bl_62 br_62 wl_216 vdd gnd cell_6t
Xbit_r217_c62 bl_62 br_62 wl_217 vdd gnd cell_6t
Xbit_r218_c62 bl_62 br_62 wl_218 vdd gnd cell_6t
Xbit_r219_c62 bl_62 br_62 wl_219 vdd gnd cell_6t
Xbit_r220_c62 bl_62 br_62 wl_220 vdd gnd cell_6t
Xbit_r221_c62 bl_62 br_62 wl_221 vdd gnd cell_6t
Xbit_r222_c62 bl_62 br_62 wl_222 vdd gnd cell_6t
Xbit_r223_c62 bl_62 br_62 wl_223 vdd gnd cell_6t
Xbit_r224_c62 bl_62 br_62 wl_224 vdd gnd cell_6t
Xbit_r225_c62 bl_62 br_62 wl_225 vdd gnd cell_6t
Xbit_r226_c62 bl_62 br_62 wl_226 vdd gnd cell_6t
Xbit_r227_c62 bl_62 br_62 wl_227 vdd gnd cell_6t
Xbit_r228_c62 bl_62 br_62 wl_228 vdd gnd cell_6t
Xbit_r229_c62 bl_62 br_62 wl_229 vdd gnd cell_6t
Xbit_r230_c62 bl_62 br_62 wl_230 vdd gnd cell_6t
Xbit_r231_c62 bl_62 br_62 wl_231 vdd gnd cell_6t
Xbit_r232_c62 bl_62 br_62 wl_232 vdd gnd cell_6t
Xbit_r233_c62 bl_62 br_62 wl_233 vdd gnd cell_6t
Xbit_r234_c62 bl_62 br_62 wl_234 vdd gnd cell_6t
Xbit_r235_c62 bl_62 br_62 wl_235 vdd gnd cell_6t
Xbit_r236_c62 bl_62 br_62 wl_236 vdd gnd cell_6t
Xbit_r237_c62 bl_62 br_62 wl_237 vdd gnd cell_6t
Xbit_r238_c62 bl_62 br_62 wl_238 vdd gnd cell_6t
Xbit_r239_c62 bl_62 br_62 wl_239 vdd gnd cell_6t
Xbit_r240_c62 bl_62 br_62 wl_240 vdd gnd cell_6t
Xbit_r241_c62 bl_62 br_62 wl_241 vdd gnd cell_6t
Xbit_r242_c62 bl_62 br_62 wl_242 vdd gnd cell_6t
Xbit_r243_c62 bl_62 br_62 wl_243 vdd gnd cell_6t
Xbit_r244_c62 bl_62 br_62 wl_244 vdd gnd cell_6t
Xbit_r245_c62 bl_62 br_62 wl_245 vdd gnd cell_6t
Xbit_r246_c62 bl_62 br_62 wl_246 vdd gnd cell_6t
Xbit_r247_c62 bl_62 br_62 wl_247 vdd gnd cell_6t
Xbit_r248_c62 bl_62 br_62 wl_248 vdd gnd cell_6t
Xbit_r249_c62 bl_62 br_62 wl_249 vdd gnd cell_6t
Xbit_r250_c62 bl_62 br_62 wl_250 vdd gnd cell_6t
Xbit_r251_c62 bl_62 br_62 wl_251 vdd gnd cell_6t
Xbit_r252_c62 bl_62 br_62 wl_252 vdd gnd cell_6t
Xbit_r253_c62 bl_62 br_62 wl_253 vdd gnd cell_6t
Xbit_r254_c62 bl_62 br_62 wl_254 vdd gnd cell_6t
Xbit_r255_c62 bl_62 br_62 wl_255 vdd gnd cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd cell_6t
Xbit_r1_c63 bl_63 br_63 wl_1 vdd gnd cell_6t
Xbit_r2_c63 bl_63 br_63 wl_2 vdd gnd cell_6t
Xbit_r3_c63 bl_63 br_63 wl_3 vdd gnd cell_6t
Xbit_r4_c63 bl_63 br_63 wl_4 vdd gnd cell_6t
Xbit_r5_c63 bl_63 br_63 wl_5 vdd gnd cell_6t
Xbit_r6_c63 bl_63 br_63 wl_6 vdd gnd cell_6t
Xbit_r7_c63 bl_63 br_63 wl_7 vdd gnd cell_6t
Xbit_r8_c63 bl_63 br_63 wl_8 vdd gnd cell_6t
Xbit_r9_c63 bl_63 br_63 wl_9 vdd gnd cell_6t
Xbit_r10_c63 bl_63 br_63 wl_10 vdd gnd cell_6t
Xbit_r11_c63 bl_63 br_63 wl_11 vdd gnd cell_6t
Xbit_r12_c63 bl_63 br_63 wl_12 vdd gnd cell_6t
Xbit_r13_c63 bl_63 br_63 wl_13 vdd gnd cell_6t
Xbit_r14_c63 bl_63 br_63 wl_14 vdd gnd cell_6t
Xbit_r15_c63 bl_63 br_63 wl_15 vdd gnd cell_6t
Xbit_r16_c63 bl_63 br_63 wl_16 vdd gnd cell_6t
Xbit_r17_c63 bl_63 br_63 wl_17 vdd gnd cell_6t
Xbit_r18_c63 bl_63 br_63 wl_18 vdd gnd cell_6t
Xbit_r19_c63 bl_63 br_63 wl_19 vdd gnd cell_6t
Xbit_r20_c63 bl_63 br_63 wl_20 vdd gnd cell_6t
Xbit_r21_c63 bl_63 br_63 wl_21 vdd gnd cell_6t
Xbit_r22_c63 bl_63 br_63 wl_22 vdd gnd cell_6t
Xbit_r23_c63 bl_63 br_63 wl_23 vdd gnd cell_6t
Xbit_r24_c63 bl_63 br_63 wl_24 vdd gnd cell_6t
Xbit_r25_c63 bl_63 br_63 wl_25 vdd gnd cell_6t
Xbit_r26_c63 bl_63 br_63 wl_26 vdd gnd cell_6t
Xbit_r27_c63 bl_63 br_63 wl_27 vdd gnd cell_6t
Xbit_r28_c63 bl_63 br_63 wl_28 vdd gnd cell_6t
Xbit_r29_c63 bl_63 br_63 wl_29 vdd gnd cell_6t
Xbit_r30_c63 bl_63 br_63 wl_30 vdd gnd cell_6t
Xbit_r31_c63 bl_63 br_63 wl_31 vdd gnd cell_6t
Xbit_r32_c63 bl_63 br_63 wl_32 vdd gnd cell_6t
Xbit_r33_c63 bl_63 br_63 wl_33 vdd gnd cell_6t
Xbit_r34_c63 bl_63 br_63 wl_34 vdd gnd cell_6t
Xbit_r35_c63 bl_63 br_63 wl_35 vdd gnd cell_6t
Xbit_r36_c63 bl_63 br_63 wl_36 vdd gnd cell_6t
Xbit_r37_c63 bl_63 br_63 wl_37 vdd gnd cell_6t
Xbit_r38_c63 bl_63 br_63 wl_38 vdd gnd cell_6t
Xbit_r39_c63 bl_63 br_63 wl_39 vdd gnd cell_6t
Xbit_r40_c63 bl_63 br_63 wl_40 vdd gnd cell_6t
Xbit_r41_c63 bl_63 br_63 wl_41 vdd gnd cell_6t
Xbit_r42_c63 bl_63 br_63 wl_42 vdd gnd cell_6t
Xbit_r43_c63 bl_63 br_63 wl_43 vdd gnd cell_6t
Xbit_r44_c63 bl_63 br_63 wl_44 vdd gnd cell_6t
Xbit_r45_c63 bl_63 br_63 wl_45 vdd gnd cell_6t
Xbit_r46_c63 bl_63 br_63 wl_46 vdd gnd cell_6t
Xbit_r47_c63 bl_63 br_63 wl_47 vdd gnd cell_6t
Xbit_r48_c63 bl_63 br_63 wl_48 vdd gnd cell_6t
Xbit_r49_c63 bl_63 br_63 wl_49 vdd gnd cell_6t
Xbit_r50_c63 bl_63 br_63 wl_50 vdd gnd cell_6t
Xbit_r51_c63 bl_63 br_63 wl_51 vdd gnd cell_6t
Xbit_r52_c63 bl_63 br_63 wl_52 vdd gnd cell_6t
Xbit_r53_c63 bl_63 br_63 wl_53 vdd gnd cell_6t
Xbit_r54_c63 bl_63 br_63 wl_54 vdd gnd cell_6t
Xbit_r55_c63 bl_63 br_63 wl_55 vdd gnd cell_6t
Xbit_r56_c63 bl_63 br_63 wl_56 vdd gnd cell_6t
Xbit_r57_c63 bl_63 br_63 wl_57 vdd gnd cell_6t
Xbit_r58_c63 bl_63 br_63 wl_58 vdd gnd cell_6t
Xbit_r59_c63 bl_63 br_63 wl_59 vdd gnd cell_6t
Xbit_r60_c63 bl_63 br_63 wl_60 vdd gnd cell_6t
Xbit_r61_c63 bl_63 br_63 wl_61 vdd gnd cell_6t
Xbit_r62_c63 bl_63 br_63 wl_62 vdd gnd cell_6t
Xbit_r63_c63 bl_63 br_63 wl_63 vdd gnd cell_6t
Xbit_r64_c63 bl_63 br_63 wl_64 vdd gnd cell_6t
Xbit_r65_c63 bl_63 br_63 wl_65 vdd gnd cell_6t
Xbit_r66_c63 bl_63 br_63 wl_66 vdd gnd cell_6t
Xbit_r67_c63 bl_63 br_63 wl_67 vdd gnd cell_6t
Xbit_r68_c63 bl_63 br_63 wl_68 vdd gnd cell_6t
Xbit_r69_c63 bl_63 br_63 wl_69 vdd gnd cell_6t
Xbit_r70_c63 bl_63 br_63 wl_70 vdd gnd cell_6t
Xbit_r71_c63 bl_63 br_63 wl_71 vdd gnd cell_6t
Xbit_r72_c63 bl_63 br_63 wl_72 vdd gnd cell_6t
Xbit_r73_c63 bl_63 br_63 wl_73 vdd gnd cell_6t
Xbit_r74_c63 bl_63 br_63 wl_74 vdd gnd cell_6t
Xbit_r75_c63 bl_63 br_63 wl_75 vdd gnd cell_6t
Xbit_r76_c63 bl_63 br_63 wl_76 vdd gnd cell_6t
Xbit_r77_c63 bl_63 br_63 wl_77 vdd gnd cell_6t
Xbit_r78_c63 bl_63 br_63 wl_78 vdd gnd cell_6t
Xbit_r79_c63 bl_63 br_63 wl_79 vdd gnd cell_6t
Xbit_r80_c63 bl_63 br_63 wl_80 vdd gnd cell_6t
Xbit_r81_c63 bl_63 br_63 wl_81 vdd gnd cell_6t
Xbit_r82_c63 bl_63 br_63 wl_82 vdd gnd cell_6t
Xbit_r83_c63 bl_63 br_63 wl_83 vdd gnd cell_6t
Xbit_r84_c63 bl_63 br_63 wl_84 vdd gnd cell_6t
Xbit_r85_c63 bl_63 br_63 wl_85 vdd gnd cell_6t
Xbit_r86_c63 bl_63 br_63 wl_86 vdd gnd cell_6t
Xbit_r87_c63 bl_63 br_63 wl_87 vdd gnd cell_6t
Xbit_r88_c63 bl_63 br_63 wl_88 vdd gnd cell_6t
Xbit_r89_c63 bl_63 br_63 wl_89 vdd gnd cell_6t
Xbit_r90_c63 bl_63 br_63 wl_90 vdd gnd cell_6t
Xbit_r91_c63 bl_63 br_63 wl_91 vdd gnd cell_6t
Xbit_r92_c63 bl_63 br_63 wl_92 vdd gnd cell_6t
Xbit_r93_c63 bl_63 br_63 wl_93 vdd gnd cell_6t
Xbit_r94_c63 bl_63 br_63 wl_94 vdd gnd cell_6t
Xbit_r95_c63 bl_63 br_63 wl_95 vdd gnd cell_6t
Xbit_r96_c63 bl_63 br_63 wl_96 vdd gnd cell_6t
Xbit_r97_c63 bl_63 br_63 wl_97 vdd gnd cell_6t
Xbit_r98_c63 bl_63 br_63 wl_98 vdd gnd cell_6t
Xbit_r99_c63 bl_63 br_63 wl_99 vdd gnd cell_6t
Xbit_r100_c63 bl_63 br_63 wl_100 vdd gnd cell_6t
Xbit_r101_c63 bl_63 br_63 wl_101 vdd gnd cell_6t
Xbit_r102_c63 bl_63 br_63 wl_102 vdd gnd cell_6t
Xbit_r103_c63 bl_63 br_63 wl_103 vdd gnd cell_6t
Xbit_r104_c63 bl_63 br_63 wl_104 vdd gnd cell_6t
Xbit_r105_c63 bl_63 br_63 wl_105 vdd gnd cell_6t
Xbit_r106_c63 bl_63 br_63 wl_106 vdd gnd cell_6t
Xbit_r107_c63 bl_63 br_63 wl_107 vdd gnd cell_6t
Xbit_r108_c63 bl_63 br_63 wl_108 vdd gnd cell_6t
Xbit_r109_c63 bl_63 br_63 wl_109 vdd gnd cell_6t
Xbit_r110_c63 bl_63 br_63 wl_110 vdd gnd cell_6t
Xbit_r111_c63 bl_63 br_63 wl_111 vdd gnd cell_6t
Xbit_r112_c63 bl_63 br_63 wl_112 vdd gnd cell_6t
Xbit_r113_c63 bl_63 br_63 wl_113 vdd gnd cell_6t
Xbit_r114_c63 bl_63 br_63 wl_114 vdd gnd cell_6t
Xbit_r115_c63 bl_63 br_63 wl_115 vdd gnd cell_6t
Xbit_r116_c63 bl_63 br_63 wl_116 vdd gnd cell_6t
Xbit_r117_c63 bl_63 br_63 wl_117 vdd gnd cell_6t
Xbit_r118_c63 bl_63 br_63 wl_118 vdd gnd cell_6t
Xbit_r119_c63 bl_63 br_63 wl_119 vdd gnd cell_6t
Xbit_r120_c63 bl_63 br_63 wl_120 vdd gnd cell_6t
Xbit_r121_c63 bl_63 br_63 wl_121 vdd gnd cell_6t
Xbit_r122_c63 bl_63 br_63 wl_122 vdd gnd cell_6t
Xbit_r123_c63 bl_63 br_63 wl_123 vdd gnd cell_6t
Xbit_r124_c63 bl_63 br_63 wl_124 vdd gnd cell_6t
Xbit_r125_c63 bl_63 br_63 wl_125 vdd gnd cell_6t
Xbit_r126_c63 bl_63 br_63 wl_126 vdd gnd cell_6t
Xbit_r127_c63 bl_63 br_63 wl_127 vdd gnd cell_6t
Xbit_r128_c63 bl_63 br_63 wl_128 vdd gnd cell_6t
Xbit_r129_c63 bl_63 br_63 wl_129 vdd gnd cell_6t
Xbit_r130_c63 bl_63 br_63 wl_130 vdd gnd cell_6t
Xbit_r131_c63 bl_63 br_63 wl_131 vdd gnd cell_6t
Xbit_r132_c63 bl_63 br_63 wl_132 vdd gnd cell_6t
Xbit_r133_c63 bl_63 br_63 wl_133 vdd gnd cell_6t
Xbit_r134_c63 bl_63 br_63 wl_134 vdd gnd cell_6t
Xbit_r135_c63 bl_63 br_63 wl_135 vdd gnd cell_6t
Xbit_r136_c63 bl_63 br_63 wl_136 vdd gnd cell_6t
Xbit_r137_c63 bl_63 br_63 wl_137 vdd gnd cell_6t
Xbit_r138_c63 bl_63 br_63 wl_138 vdd gnd cell_6t
Xbit_r139_c63 bl_63 br_63 wl_139 vdd gnd cell_6t
Xbit_r140_c63 bl_63 br_63 wl_140 vdd gnd cell_6t
Xbit_r141_c63 bl_63 br_63 wl_141 vdd gnd cell_6t
Xbit_r142_c63 bl_63 br_63 wl_142 vdd gnd cell_6t
Xbit_r143_c63 bl_63 br_63 wl_143 vdd gnd cell_6t
Xbit_r144_c63 bl_63 br_63 wl_144 vdd gnd cell_6t
Xbit_r145_c63 bl_63 br_63 wl_145 vdd gnd cell_6t
Xbit_r146_c63 bl_63 br_63 wl_146 vdd gnd cell_6t
Xbit_r147_c63 bl_63 br_63 wl_147 vdd gnd cell_6t
Xbit_r148_c63 bl_63 br_63 wl_148 vdd gnd cell_6t
Xbit_r149_c63 bl_63 br_63 wl_149 vdd gnd cell_6t
Xbit_r150_c63 bl_63 br_63 wl_150 vdd gnd cell_6t
Xbit_r151_c63 bl_63 br_63 wl_151 vdd gnd cell_6t
Xbit_r152_c63 bl_63 br_63 wl_152 vdd gnd cell_6t
Xbit_r153_c63 bl_63 br_63 wl_153 vdd gnd cell_6t
Xbit_r154_c63 bl_63 br_63 wl_154 vdd gnd cell_6t
Xbit_r155_c63 bl_63 br_63 wl_155 vdd gnd cell_6t
Xbit_r156_c63 bl_63 br_63 wl_156 vdd gnd cell_6t
Xbit_r157_c63 bl_63 br_63 wl_157 vdd gnd cell_6t
Xbit_r158_c63 bl_63 br_63 wl_158 vdd gnd cell_6t
Xbit_r159_c63 bl_63 br_63 wl_159 vdd gnd cell_6t
Xbit_r160_c63 bl_63 br_63 wl_160 vdd gnd cell_6t
Xbit_r161_c63 bl_63 br_63 wl_161 vdd gnd cell_6t
Xbit_r162_c63 bl_63 br_63 wl_162 vdd gnd cell_6t
Xbit_r163_c63 bl_63 br_63 wl_163 vdd gnd cell_6t
Xbit_r164_c63 bl_63 br_63 wl_164 vdd gnd cell_6t
Xbit_r165_c63 bl_63 br_63 wl_165 vdd gnd cell_6t
Xbit_r166_c63 bl_63 br_63 wl_166 vdd gnd cell_6t
Xbit_r167_c63 bl_63 br_63 wl_167 vdd gnd cell_6t
Xbit_r168_c63 bl_63 br_63 wl_168 vdd gnd cell_6t
Xbit_r169_c63 bl_63 br_63 wl_169 vdd gnd cell_6t
Xbit_r170_c63 bl_63 br_63 wl_170 vdd gnd cell_6t
Xbit_r171_c63 bl_63 br_63 wl_171 vdd gnd cell_6t
Xbit_r172_c63 bl_63 br_63 wl_172 vdd gnd cell_6t
Xbit_r173_c63 bl_63 br_63 wl_173 vdd gnd cell_6t
Xbit_r174_c63 bl_63 br_63 wl_174 vdd gnd cell_6t
Xbit_r175_c63 bl_63 br_63 wl_175 vdd gnd cell_6t
Xbit_r176_c63 bl_63 br_63 wl_176 vdd gnd cell_6t
Xbit_r177_c63 bl_63 br_63 wl_177 vdd gnd cell_6t
Xbit_r178_c63 bl_63 br_63 wl_178 vdd gnd cell_6t
Xbit_r179_c63 bl_63 br_63 wl_179 vdd gnd cell_6t
Xbit_r180_c63 bl_63 br_63 wl_180 vdd gnd cell_6t
Xbit_r181_c63 bl_63 br_63 wl_181 vdd gnd cell_6t
Xbit_r182_c63 bl_63 br_63 wl_182 vdd gnd cell_6t
Xbit_r183_c63 bl_63 br_63 wl_183 vdd gnd cell_6t
Xbit_r184_c63 bl_63 br_63 wl_184 vdd gnd cell_6t
Xbit_r185_c63 bl_63 br_63 wl_185 vdd gnd cell_6t
Xbit_r186_c63 bl_63 br_63 wl_186 vdd gnd cell_6t
Xbit_r187_c63 bl_63 br_63 wl_187 vdd gnd cell_6t
Xbit_r188_c63 bl_63 br_63 wl_188 vdd gnd cell_6t
Xbit_r189_c63 bl_63 br_63 wl_189 vdd gnd cell_6t
Xbit_r190_c63 bl_63 br_63 wl_190 vdd gnd cell_6t
Xbit_r191_c63 bl_63 br_63 wl_191 vdd gnd cell_6t
Xbit_r192_c63 bl_63 br_63 wl_192 vdd gnd cell_6t
Xbit_r193_c63 bl_63 br_63 wl_193 vdd gnd cell_6t
Xbit_r194_c63 bl_63 br_63 wl_194 vdd gnd cell_6t
Xbit_r195_c63 bl_63 br_63 wl_195 vdd gnd cell_6t
Xbit_r196_c63 bl_63 br_63 wl_196 vdd gnd cell_6t
Xbit_r197_c63 bl_63 br_63 wl_197 vdd gnd cell_6t
Xbit_r198_c63 bl_63 br_63 wl_198 vdd gnd cell_6t
Xbit_r199_c63 bl_63 br_63 wl_199 vdd gnd cell_6t
Xbit_r200_c63 bl_63 br_63 wl_200 vdd gnd cell_6t
Xbit_r201_c63 bl_63 br_63 wl_201 vdd gnd cell_6t
Xbit_r202_c63 bl_63 br_63 wl_202 vdd gnd cell_6t
Xbit_r203_c63 bl_63 br_63 wl_203 vdd gnd cell_6t
Xbit_r204_c63 bl_63 br_63 wl_204 vdd gnd cell_6t
Xbit_r205_c63 bl_63 br_63 wl_205 vdd gnd cell_6t
Xbit_r206_c63 bl_63 br_63 wl_206 vdd gnd cell_6t
Xbit_r207_c63 bl_63 br_63 wl_207 vdd gnd cell_6t
Xbit_r208_c63 bl_63 br_63 wl_208 vdd gnd cell_6t
Xbit_r209_c63 bl_63 br_63 wl_209 vdd gnd cell_6t
Xbit_r210_c63 bl_63 br_63 wl_210 vdd gnd cell_6t
Xbit_r211_c63 bl_63 br_63 wl_211 vdd gnd cell_6t
Xbit_r212_c63 bl_63 br_63 wl_212 vdd gnd cell_6t
Xbit_r213_c63 bl_63 br_63 wl_213 vdd gnd cell_6t
Xbit_r214_c63 bl_63 br_63 wl_214 vdd gnd cell_6t
Xbit_r215_c63 bl_63 br_63 wl_215 vdd gnd cell_6t
Xbit_r216_c63 bl_63 br_63 wl_216 vdd gnd cell_6t
Xbit_r217_c63 bl_63 br_63 wl_217 vdd gnd cell_6t
Xbit_r218_c63 bl_63 br_63 wl_218 vdd gnd cell_6t
Xbit_r219_c63 bl_63 br_63 wl_219 vdd gnd cell_6t
Xbit_r220_c63 bl_63 br_63 wl_220 vdd gnd cell_6t
Xbit_r221_c63 bl_63 br_63 wl_221 vdd gnd cell_6t
Xbit_r222_c63 bl_63 br_63 wl_222 vdd gnd cell_6t
Xbit_r223_c63 bl_63 br_63 wl_223 vdd gnd cell_6t
Xbit_r224_c63 bl_63 br_63 wl_224 vdd gnd cell_6t
Xbit_r225_c63 bl_63 br_63 wl_225 vdd gnd cell_6t
Xbit_r226_c63 bl_63 br_63 wl_226 vdd gnd cell_6t
Xbit_r227_c63 bl_63 br_63 wl_227 vdd gnd cell_6t
Xbit_r228_c63 bl_63 br_63 wl_228 vdd gnd cell_6t
Xbit_r229_c63 bl_63 br_63 wl_229 vdd gnd cell_6t
Xbit_r230_c63 bl_63 br_63 wl_230 vdd gnd cell_6t
Xbit_r231_c63 bl_63 br_63 wl_231 vdd gnd cell_6t
Xbit_r232_c63 bl_63 br_63 wl_232 vdd gnd cell_6t
Xbit_r233_c63 bl_63 br_63 wl_233 vdd gnd cell_6t
Xbit_r234_c63 bl_63 br_63 wl_234 vdd gnd cell_6t
Xbit_r235_c63 bl_63 br_63 wl_235 vdd gnd cell_6t
Xbit_r236_c63 bl_63 br_63 wl_236 vdd gnd cell_6t
Xbit_r237_c63 bl_63 br_63 wl_237 vdd gnd cell_6t
Xbit_r238_c63 bl_63 br_63 wl_238 vdd gnd cell_6t
Xbit_r239_c63 bl_63 br_63 wl_239 vdd gnd cell_6t
Xbit_r240_c63 bl_63 br_63 wl_240 vdd gnd cell_6t
Xbit_r241_c63 bl_63 br_63 wl_241 vdd gnd cell_6t
Xbit_r242_c63 bl_63 br_63 wl_242 vdd gnd cell_6t
Xbit_r243_c63 bl_63 br_63 wl_243 vdd gnd cell_6t
Xbit_r244_c63 bl_63 br_63 wl_244 vdd gnd cell_6t
Xbit_r245_c63 bl_63 br_63 wl_245 vdd gnd cell_6t
Xbit_r246_c63 bl_63 br_63 wl_246 vdd gnd cell_6t
Xbit_r247_c63 bl_63 br_63 wl_247 vdd gnd cell_6t
Xbit_r248_c63 bl_63 br_63 wl_248 vdd gnd cell_6t
Xbit_r249_c63 bl_63 br_63 wl_249 vdd gnd cell_6t
Xbit_r250_c63 bl_63 br_63 wl_250 vdd gnd cell_6t
Xbit_r251_c63 bl_63 br_63 wl_251 vdd gnd cell_6t
Xbit_r252_c63 bl_63 br_63 wl_252 vdd gnd cell_6t
Xbit_r253_c63 bl_63 br_63 wl_253 vdd gnd cell_6t
Xbit_r254_c63 bl_63 br_63 wl_254 vdd gnd cell_6t
Xbit_r255_c63 bl_63 br_63 wl_255 vdd gnd cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd cell_6t
Xbit_r1_c64 bl_64 br_64 wl_1 vdd gnd cell_6t
Xbit_r2_c64 bl_64 br_64 wl_2 vdd gnd cell_6t
Xbit_r3_c64 bl_64 br_64 wl_3 vdd gnd cell_6t
Xbit_r4_c64 bl_64 br_64 wl_4 vdd gnd cell_6t
Xbit_r5_c64 bl_64 br_64 wl_5 vdd gnd cell_6t
Xbit_r6_c64 bl_64 br_64 wl_6 vdd gnd cell_6t
Xbit_r7_c64 bl_64 br_64 wl_7 vdd gnd cell_6t
Xbit_r8_c64 bl_64 br_64 wl_8 vdd gnd cell_6t
Xbit_r9_c64 bl_64 br_64 wl_9 vdd gnd cell_6t
Xbit_r10_c64 bl_64 br_64 wl_10 vdd gnd cell_6t
Xbit_r11_c64 bl_64 br_64 wl_11 vdd gnd cell_6t
Xbit_r12_c64 bl_64 br_64 wl_12 vdd gnd cell_6t
Xbit_r13_c64 bl_64 br_64 wl_13 vdd gnd cell_6t
Xbit_r14_c64 bl_64 br_64 wl_14 vdd gnd cell_6t
Xbit_r15_c64 bl_64 br_64 wl_15 vdd gnd cell_6t
Xbit_r16_c64 bl_64 br_64 wl_16 vdd gnd cell_6t
Xbit_r17_c64 bl_64 br_64 wl_17 vdd gnd cell_6t
Xbit_r18_c64 bl_64 br_64 wl_18 vdd gnd cell_6t
Xbit_r19_c64 bl_64 br_64 wl_19 vdd gnd cell_6t
Xbit_r20_c64 bl_64 br_64 wl_20 vdd gnd cell_6t
Xbit_r21_c64 bl_64 br_64 wl_21 vdd gnd cell_6t
Xbit_r22_c64 bl_64 br_64 wl_22 vdd gnd cell_6t
Xbit_r23_c64 bl_64 br_64 wl_23 vdd gnd cell_6t
Xbit_r24_c64 bl_64 br_64 wl_24 vdd gnd cell_6t
Xbit_r25_c64 bl_64 br_64 wl_25 vdd gnd cell_6t
Xbit_r26_c64 bl_64 br_64 wl_26 vdd gnd cell_6t
Xbit_r27_c64 bl_64 br_64 wl_27 vdd gnd cell_6t
Xbit_r28_c64 bl_64 br_64 wl_28 vdd gnd cell_6t
Xbit_r29_c64 bl_64 br_64 wl_29 vdd gnd cell_6t
Xbit_r30_c64 bl_64 br_64 wl_30 vdd gnd cell_6t
Xbit_r31_c64 bl_64 br_64 wl_31 vdd gnd cell_6t
Xbit_r32_c64 bl_64 br_64 wl_32 vdd gnd cell_6t
Xbit_r33_c64 bl_64 br_64 wl_33 vdd gnd cell_6t
Xbit_r34_c64 bl_64 br_64 wl_34 vdd gnd cell_6t
Xbit_r35_c64 bl_64 br_64 wl_35 vdd gnd cell_6t
Xbit_r36_c64 bl_64 br_64 wl_36 vdd gnd cell_6t
Xbit_r37_c64 bl_64 br_64 wl_37 vdd gnd cell_6t
Xbit_r38_c64 bl_64 br_64 wl_38 vdd gnd cell_6t
Xbit_r39_c64 bl_64 br_64 wl_39 vdd gnd cell_6t
Xbit_r40_c64 bl_64 br_64 wl_40 vdd gnd cell_6t
Xbit_r41_c64 bl_64 br_64 wl_41 vdd gnd cell_6t
Xbit_r42_c64 bl_64 br_64 wl_42 vdd gnd cell_6t
Xbit_r43_c64 bl_64 br_64 wl_43 vdd gnd cell_6t
Xbit_r44_c64 bl_64 br_64 wl_44 vdd gnd cell_6t
Xbit_r45_c64 bl_64 br_64 wl_45 vdd gnd cell_6t
Xbit_r46_c64 bl_64 br_64 wl_46 vdd gnd cell_6t
Xbit_r47_c64 bl_64 br_64 wl_47 vdd gnd cell_6t
Xbit_r48_c64 bl_64 br_64 wl_48 vdd gnd cell_6t
Xbit_r49_c64 bl_64 br_64 wl_49 vdd gnd cell_6t
Xbit_r50_c64 bl_64 br_64 wl_50 vdd gnd cell_6t
Xbit_r51_c64 bl_64 br_64 wl_51 vdd gnd cell_6t
Xbit_r52_c64 bl_64 br_64 wl_52 vdd gnd cell_6t
Xbit_r53_c64 bl_64 br_64 wl_53 vdd gnd cell_6t
Xbit_r54_c64 bl_64 br_64 wl_54 vdd gnd cell_6t
Xbit_r55_c64 bl_64 br_64 wl_55 vdd gnd cell_6t
Xbit_r56_c64 bl_64 br_64 wl_56 vdd gnd cell_6t
Xbit_r57_c64 bl_64 br_64 wl_57 vdd gnd cell_6t
Xbit_r58_c64 bl_64 br_64 wl_58 vdd gnd cell_6t
Xbit_r59_c64 bl_64 br_64 wl_59 vdd gnd cell_6t
Xbit_r60_c64 bl_64 br_64 wl_60 vdd gnd cell_6t
Xbit_r61_c64 bl_64 br_64 wl_61 vdd gnd cell_6t
Xbit_r62_c64 bl_64 br_64 wl_62 vdd gnd cell_6t
Xbit_r63_c64 bl_64 br_64 wl_63 vdd gnd cell_6t
Xbit_r64_c64 bl_64 br_64 wl_64 vdd gnd cell_6t
Xbit_r65_c64 bl_64 br_64 wl_65 vdd gnd cell_6t
Xbit_r66_c64 bl_64 br_64 wl_66 vdd gnd cell_6t
Xbit_r67_c64 bl_64 br_64 wl_67 vdd gnd cell_6t
Xbit_r68_c64 bl_64 br_64 wl_68 vdd gnd cell_6t
Xbit_r69_c64 bl_64 br_64 wl_69 vdd gnd cell_6t
Xbit_r70_c64 bl_64 br_64 wl_70 vdd gnd cell_6t
Xbit_r71_c64 bl_64 br_64 wl_71 vdd gnd cell_6t
Xbit_r72_c64 bl_64 br_64 wl_72 vdd gnd cell_6t
Xbit_r73_c64 bl_64 br_64 wl_73 vdd gnd cell_6t
Xbit_r74_c64 bl_64 br_64 wl_74 vdd gnd cell_6t
Xbit_r75_c64 bl_64 br_64 wl_75 vdd gnd cell_6t
Xbit_r76_c64 bl_64 br_64 wl_76 vdd gnd cell_6t
Xbit_r77_c64 bl_64 br_64 wl_77 vdd gnd cell_6t
Xbit_r78_c64 bl_64 br_64 wl_78 vdd gnd cell_6t
Xbit_r79_c64 bl_64 br_64 wl_79 vdd gnd cell_6t
Xbit_r80_c64 bl_64 br_64 wl_80 vdd gnd cell_6t
Xbit_r81_c64 bl_64 br_64 wl_81 vdd gnd cell_6t
Xbit_r82_c64 bl_64 br_64 wl_82 vdd gnd cell_6t
Xbit_r83_c64 bl_64 br_64 wl_83 vdd gnd cell_6t
Xbit_r84_c64 bl_64 br_64 wl_84 vdd gnd cell_6t
Xbit_r85_c64 bl_64 br_64 wl_85 vdd gnd cell_6t
Xbit_r86_c64 bl_64 br_64 wl_86 vdd gnd cell_6t
Xbit_r87_c64 bl_64 br_64 wl_87 vdd gnd cell_6t
Xbit_r88_c64 bl_64 br_64 wl_88 vdd gnd cell_6t
Xbit_r89_c64 bl_64 br_64 wl_89 vdd gnd cell_6t
Xbit_r90_c64 bl_64 br_64 wl_90 vdd gnd cell_6t
Xbit_r91_c64 bl_64 br_64 wl_91 vdd gnd cell_6t
Xbit_r92_c64 bl_64 br_64 wl_92 vdd gnd cell_6t
Xbit_r93_c64 bl_64 br_64 wl_93 vdd gnd cell_6t
Xbit_r94_c64 bl_64 br_64 wl_94 vdd gnd cell_6t
Xbit_r95_c64 bl_64 br_64 wl_95 vdd gnd cell_6t
Xbit_r96_c64 bl_64 br_64 wl_96 vdd gnd cell_6t
Xbit_r97_c64 bl_64 br_64 wl_97 vdd gnd cell_6t
Xbit_r98_c64 bl_64 br_64 wl_98 vdd gnd cell_6t
Xbit_r99_c64 bl_64 br_64 wl_99 vdd gnd cell_6t
Xbit_r100_c64 bl_64 br_64 wl_100 vdd gnd cell_6t
Xbit_r101_c64 bl_64 br_64 wl_101 vdd gnd cell_6t
Xbit_r102_c64 bl_64 br_64 wl_102 vdd gnd cell_6t
Xbit_r103_c64 bl_64 br_64 wl_103 vdd gnd cell_6t
Xbit_r104_c64 bl_64 br_64 wl_104 vdd gnd cell_6t
Xbit_r105_c64 bl_64 br_64 wl_105 vdd gnd cell_6t
Xbit_r106_c64 bl_64 br_64 wl_106 vdd gnd cell_6t
Xbit_r107_c64 bl_64 br_64 wl_107 vdd gnd cell_6t
Xbit_r108_c64 bl_64 br_64 wl_108 vdd gnd cell_6t
Xbit_r109_c64 bl_64 br_64 wl_109 vdd gnd cell_6t
Xbit_r110_c64 bl_64 br_64 wl_110 vdd gnd cell_6t
Xbit_r111_c64 bl_64 br_64 wl_111 vdd gnd cell_6t
Xbit_r112_c64 bl_64 br_64 wl_112 vdd gnd cell_6t
Xbit_r113_c64 bl_64 br_64 wl_113 vdd gnd cell_6t
Xbit_r114_c64 bl_64 br_64 wl_114 vdd gnd cell_6t
Xbit_r115_c64 bl_64 br_64 wl_115 vdd gnd cell_6t
Xbit_r116_c64 bl_64 br_64 wl_116 vdd gnd cell_6t
Xbit_r117_c64 bl_64 br_64 wl_117 vdd gnd cell_6t
Xbit_r118_c64 bl_64 br_64 wl_118 vdd gnd cell_6t
Xbit_r119_c64 bl_64 br_64 wl_119 vdd gnd cell_6t
Xbit_r120_c64 bl_64 br_64 wl_120 vdd gnd cell_6t
Xbit_r121_c64 bl_64 br_64 wl_121 vdd gnd cell_6t
Xbit_r122_c64 bl_64 br_64 wl_122 vdd gnd cell_6t
Xbit_r123_c64 bl_64 br_64 wl_123 vdd gnd cell_6t
Xbit_r124_c64 bl_64 br_64 wl_124 vdd gnd cell_6t
Xbit_r125_c64 bl_64 br_64 wl_125 vdd gnd cell_6t
Xbit_r126_c64 bl_64 br_64 wl_126 vdd gnd cell_6t
Xbit_r127_c64 bl_64 br_64 wl_127 vdd gnd cell_6t
Xbit_r128_c64 bl_64 br_64 wl_128 vdd gnd cell_6t
Xbit_r129_c64 bl_64 br_64 wl_129 vdd gnd cell_6t
Xbit_r130_c64 bl_64 br_64 wl_130 vdd gnd cell_6t
Xbit_r131_c64 bl_64 br_64 wl_131 vdd gnd cell_6t
Xbit_r132_c64 bl_64 br_64 wl_132 vdd gnd cell_6t
Xbit_r133_c64 bl_64 br_64 wl_133 vdd gnd cell_6t
Xbit_r134_c64 bl_64 br_64 wl_134 vdd gnd cell_6t
Xbit_r135_c64 bl_64 br_64 wl_135 vdd gnd cell_6t
Xbit_r136_c64 bl_64 br_64 wl_136 vdd gnd cell_6t
Xbit_r137_c64 bl_64 br_64 wl_137 vdd gnd cell_6t
Xbit_r138_c64 bl_64 br_64 wl_138 vdd gnd cell_6t
Xbit_r139_c64 bl_64 br_64 wl_139 vdd gnd cell_6t
Xbit_r140_c64 bl_64 br_64 wl_140 vdd gnd cell_6t
Xbit_r141_c64 bl_64 br_64 wl_141 vdd gnd cell_6t
Xbit_r142_c64 bl_64 br_64 wl_142 vdd gnd cell_6t
Xbit_r143_c64 bl_64 br_64 wl_143 vdd gnd cell_6t
Xbit_r144_c64 bl_64 br_64 wl_144 vdd gnd cell_6t
Xbit_r145_c64 bl_64 br_64 wl_145 vdd gnd cell_6t
Xbit_r146_c64 bl_64 br_64 wl_146 vdd gnd cell_6t
Xbit_r147_c64 bl_64 br_64 wl_147 vdd gnd cell_6t
Xbit_r148_c64 bl_64 br_64 wl_148 vdd gnd cell_6t
Xbit_r149_c64 bl_64 br_64 wl_149 vdd gnd cell_6t
Xbit_r150_c64 bl_64 br_64 wl_150 vdd gnd cell_6t
Xbit_r151_c64 bl_64 br_64 wl_151 vdd gnd cell_6t
Xbit_r152_c64 bl_64 br_64 wl_152 vdd gnd cell_6t
Xbit_r153_c64 bl_64 br_64 wl_153 vdd gnd cell_6t
Xbit_r154_c64 bl_64 br_64 wl_154 vdd gnd cell_6t
Xbit_r155_c64 bl_64 br_64 wl_155 vdd gnd cell_6t
Xbit_r156_c64 bl_64 br_64 wl_156 vdd gnd cell_6t
Xbit_r157_c64 bl_64 br_64 wl_157 vdd gnd cell_6t
Xbit_r158_c64 bl_64 br_64 wl_158 vdd gnd cell_6t
Xbit_r159_c64 bl_64 br_64 wl_159 vdd gnd cell_6t
Xbit_r160_c64 bl_64 br_64 wl_160 vdd gnd cell_6t
Xbit_r161_c64 bl_64 br_64 wl_161 vdd gnd cell_6t
Xbit_r162_c64 bl_64 br_64 wl_162 vdd gnd cell_6t
Xbit_r163_c64 bl_64 br_64 wl_163 vdd gnd cell_6t
Xbit_r164_c64 bl_64 br_64 wl_164 vdd gnd cell_6t
Xbit_r165_c64 bl_64 br_64 wl_165 vdd gnd cell_6t
Xbit_r166_c64 bl_64 br_64 wl_166 vdd gnd cell_6t
Xbit_r167_c64 bl_64 br_64 wl_167 vdd gnd cell_6t
Xbit_r168_c64 bl_64 br_64 wl_168 vdd gnd cell_6t
Xbit_r169_c64 bl_64 br_64 wl_169 vdd gnd cell_6t
Xbit_r170_c64 bl_64 br_64 wl_170 vdd gnd cell_6t
Xbit_r171_c64 bl_64 br_64 wl_171 vdd gnd cell_6t
Xbit_r172_c64 bl_64 br_64 wl_172 vdd gnd cell_6t
Xbit_r173_c64 bl_64 br_64 wl_173 vdd gnd cell_6t
Xbit_r174_c64 bl_64 br_64 wl_174 vdd gnd cell_6t
Xbit_r175_c64 bl_64 br_64 wl_175 vdd gnd cell_6t
Xbit_r176_c64 bl_64 br_64 wl_176 vdd gnd cell_6t
Xbit_r177_c64 bl_64 br_64 wl_177 vdd gnd cell_6t
Xbit_r178_c64 bl_64 br_64 wl_178 vdd gnd cell_6t
Xbit_r179_c64 bl_64 br_64 wl_179 vdd gnd cell_6t
Xbit_r180_c64 bl_64 br_64 wl_180 vdd gnd cell_6t
Xbit_r181_c64 bl_64 br_64 wl_181 vdd gnd cell_6t
Xbit_r182_c64 bl_64 br_64 wl_182 vdd gnd cell_6t
Xbit_r183_c64 bl_64 br_64 wl_183 vdd gnd cell_6t
Xbit_r184_c64 bl_64 br_64 wl_184 vdd gnd cell_6t
Xbit_r185_c64 bl_64 br_64 wl_185 vdd gnd cell_6t
Xbit_r186_c64 bl_64 br_64 wl_186 vdd gnd cell_6t
Xbit_r187_c64 bl_64 br_64 wl_187 vdd gnd cell_6t
Xbit_r188_c64 bl_64 br_64 wl_188 vdd gnd cell_6t
Xbit_r189_c64 bl_64 br_64 wl_189 vdd gnd cell_6t
Xbit_r190_c64 bl_64 br_64 wl_190 vdd gnd cell_6t
Xbit_r191_c64 bl_64 br_64 wl_191 vdd gnd cell_6t
Xbit_r192_c64 bl_64 br_64 wl_192 vdd gnd cell_6t
Xbit_r193_c64 bl_64 br_64 wl_193 vdd gnd cell_6t
Xbit_r194_c64 bl_64 br_64 wl_194 vdd gnd cell_6t
Xbit_r195_c64 bl_64 br_64 wl_195 vdd gnd cell_6t
Xbit_r196_c64 bl_64 br_64 wl_196 vdd gnd cell_6t
Xbit_r197_c64 bl_64 br_64 wl_197 vdd gnd cell_6t
Xbit_r198_c64 bl_64 br_64 wl_198 vdd gnd cell_6t
Xbit_r199_c64 bl_64 br_64 wl_199 vdd gnd cell_6t
Xbit_r200_c64 bl_64 br_64 wl_200 vdd gnd cell_6t
Xbit_r201_c64 bl_64 br_64 wl_201 vdd gnd cell_6t
Xbit_r202_c64 bl_64 br_64 wl_202 vdd gnd cell_6t
Xbit_r203_c64 bl_64 br_64 wl_203 vdd gnd cell_6t
Xbit_r204_c64 bl_64 br_64 wl_204 vdd gnd cell_6t
Xbit_r205_c64 bl_64 br_64 wl_205 vdd gnd cell_6t
Xbit_r206_c64 bl_64 br_64 wl_206 vdd gnd cell_6t
Xbit_r207_c64 bl_64 br_64 wl_207 vdd gnd cell_6t
Xbit_r208_c64 bl_64 br_64 wl_208 vdd gnd cell_6t
Xbit_r209_c64 bl_64 br_64 wl_209 vdd gnd cell_6t
Xbit_r210_c64 bl_64 br_64 wl_210 vdd gnd cell_6t
Xbit_r211_c64 bl_64 br_64 wl_211 vdd gnd cell_6t
Xbit_r212_c64 bl_64 br_64 wl_212 vdd gnd cell_6t
Xbit_r213_c64 bl_64 br_64 wl_213 vdd gnd cell_6t
Xbit_r214_c64 bl_64 br_64 wl_214 vdd gnd cell_6t
Xbit_r215_c64 bl_64 br_64 wl_215 vdd gnd cell_6t
Xbit_r216_c64 bl_64 br_64 wl_216 vdd gnd cell_6t
Xbit_r217_c64 bl_64 br_64 wl_217 vdd gnd cell_6t
Xbit_r218_c64 bl_64 br_64 wl_218 vdd gnd cell_6t
Xbit_r219_c64 bl_64 br_64 wl_219 vdd gnd cell_6t
Xbit_r220_c64 bl_64 br_64 wl_220 vdd gnd cell_6t
Xbit_r221_c64 bl_64 br_64 wl_221 vdd gnd cell_6t
Xbit_r222_c64 bl_64 br_64 wl_222 vdd gnd cell_6t
Xbit_r223_c64 bl_64 br_64 wl_223 vdd gnd cell_6t
Xbit_r224_c64 bl_64 br_64 wl_224 vdd gnd cell_6t
Xbit_r225_c64 bl_64 br_64 wl_225 vdd gnd cell_6t
Xbit_r226_c64 bl_64 br_64 wl_226 vdd gnd cell_6t
Xbit_r227_c64 bl_64 br_64 wl_227 vdd gnd cell_6t
Xbit_r228_c64 bl_64 br_64 wl_228 vdd gnd cell_6t
Xbit_r229_c64 bl_64 br_64 wl_229 vdd gnd cell_6t
Xbit_r230_c64 bl_64 br_64 wl_230 vdd gnd cell_6t
Xbit_r231_c64 bl_64 br_64 wl_231 vdd gnd cell_6t
Xbit_r232_c64 bl_64 br_64 wl_232 vdd gnd cell_6t
Xbit_r233_c64 bl_64 br_64 wl_233 vdd gnd cell_6t
Xbit_r234_c64 bl_64 br_64 wl_234 vdd gnd cell_6t
Xbit_r235_c64 bl_64 br_64 wl_235 vdd gnd cell_6t
Xbit_r236_c64 bl_64 br_64 wl_236 vdd gnd cell_6t
Xbit_r237_c64 bl_64 br_64 wl_237 vdd gnd cell_6t
Xbit_r238_c64 bl_64 br_64 wl_238 vdd gnd cell_6t
Xbit_r239_c64 bl_64 br_64 wl_239 vdd gnd cell_6t
Xbit_r240_c64 bl_64 br_64 wl_240 vdd gnd cell_6t
Xbit_r241_c64 bl_64 br_64 wl_241 vdd gnd cell_6t
Xbit_r242_c64 bl_64 br_64 wl_242 vdd gnd cell_6t
Xbit_r243_c64 bl_64 br_64 wl_243 vdd gnd cell_6t
Xbit_r244_c64 bl_64 br_64 wl_244 vdd gnd cell_6t
Xbit_r245_c64 bl_64 br_64 wl_245 vdd gnd cell_6t
Xbit_r246_c64 bl_64 br_64 wl_246 vdd gnd cell_6t
Xbit_r247_c64 bl_64 br_64 wl_247 vdd gnd cell_6t
Xbit_r248_c64 bl_64 br_64 wl_248 vdd gnd cell_6t
Xbit_r249_c64 bl_64 br_64 wl_249 vdd gnd cell_6t
Xbit_r250_c64 bl_64 br_64 wl_250 vdd gnd cell_6t
Xbit_r251_c64 bl_64 br_64 wl_251 vdd gnd cell_6t
Xbit_r252_c64 bl_64 br_64 wl_252 vdd gnd cell_6t
Xbit_r253_c64 bl_64 br_64 wl_253 vdd gnd cell_6t
Xbit_r254_c64 bl_64 br_64 wl_254 vdd gnd cell_6t
Xbit_r255_c64 bl_64 br_64 wl_255 vdd gnd cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd cell_6t
Xbit_r1_c65 bl_65 br_65 wl_1 vdd gnd cell_6t
Xbit_r2_c65 bl_65 br_65 wl_2 vdd gnd cell_6t
Xbit_r3_c65 bl_65 br_65 wl_3 vdd gnd cell_6t
Xbit_r4_c65 bl_65 br_65 wl_4 vdd gnd cell_6t
Xbit_r5_c65 bl_65 br_65 wl_5 vdd gnd cell_6t
Xbit_r6_c65 bl_65 br_65 wl_6 vdd gnd cell_6t
Xbit_r7_c65 bl_65 br_65 wl_7 vdd gnd cell_6t
Xbit_r8_c65 bl_65 br_65 wl_8 vdd gnd cell_6t
Xbit_r9_c65 bl_65 br_65 wl_9 vdd gnd cell_6t
Xbit_r10_c65 bl_65 br_65 wl_10 vdd gnd cell_6t
Xbit_r11_c65 bl_65 br_65 wl_11 vdd gnd cell_6t
Xbit_r12_c65 bl_65 br_65 wl_12 vdd gnd cell_6t
Xbit_r13_c65 bl_65 br_65 wl_13 vdd gnd cell_6t
Xbit_r14_c65 bl_65 br_65 wl_14 vdd gnd cell_6t
Xbit_r15_c65 bl_65 br_65 wl_15 vdd gnd cell_6t
Xbit_r16_c65 bl_65 br_65 wl_16 vdd gnd cell_6t
Xbit_r17_c65 bl_65 br_65 wl_17 vdd gnd cell_6t
Xbit_r18_c65 bl_65 br_65 wl_18 vdd gnd cell_6t
Xbit_r19_c65 bl_65 br_65 wl_19 vdd gnd cell_6t
Xbit_r20_c65 bl_65 br_65 wl_20 vdd gnd cell_6t
Xbit_r21_c65 bl_65 br_65 wl_21 vdd gnd cell_6t
Xbit_r22_c65 bl_65 br_65 wl_22 vdd gnd cell_6t
Xbit_r23_c65 bl_65 br_65 wl_23 vdd gnd cell_6t
Xbit_r24_c65 bl_65 br_65 wl_24 vdd gnd cell_6t
Xbit_r25_c65 bl_65 br_65 wl_25 vdd gnd cell_6t
Xbit_r26_c65 bl_65 br_65 wl_26 vdd gnd cell_6t
Xbit_r27_c65 bl_65 br_65 wl_27 vdd gnd cell_6t
Xbit_r28_c65 bl_65 br_65 wl_28 vdd gnd cell_6t
Xbit_r29_c65 bl_65 br_65 wl_29 vdd gnd cell_6t
Xbit_r30_c65 bl_65 br_65 wl_30 vdd gnd cell_6t
Xbit_r31_c65 bl_65 br_65 wl_31 vdd gnd cell_6t
Xbit_r32_c65 bl_65 br_65 wl_32 vdd gnd cell_6t
Xbit_r33_c65 bl_65 br_65 wl_33 vdd gnd cell_6t
Xbit_r34_c65 bl_65 br_65 wl_34 vdd gnd cell_6t
Xbit_r35_c65 bl_65 br_65 wl_35 vdd gnd cell_6t
Xbit_r36_c65 bl_65 br_65 wl_36 vdd gnd cell_6t
Xbit_r37_c65 bl_65 br_65 wl_37 vdd gnd cell_6t
Xbit_r38_c65 bl_65 br_65 wl_38 vdd gnd cell_6t
Xbit_r39_c65 bl_65 br_65 wl_39 vdd gnd cell_6t
Xbit_r40_c65 bl_65 br_65 wl_40 vdd gnd cell_6t
Xbit_r41_c65 bl_65 br_65 wl_41 vdd gnd cell_6t
Xbit_r42_c65 bl_65 br_65 wl_42 vdd gnd cell_6t
Xbit_r43_c65 bl_65 br_65 wl_43 vdd gnd cell_6t
Xbit_r44_c65 bl_65 br_65 wl_44 vdd gnd cell_6t
Xbit_r45_c65 bl_65 br_65 wl_45 vdd gnd cell_6t
Xbit_r46_c65 bl_65 br_65 wl_46 vdd gnd cell_6t
Xbit_r47_c65 bl_65 br_65 wl_47 vdd gnd cell_6t
Xbit_r48_c65 bl_65 br_65 wl_48 vdd gnd cell_6t
Xbit_r49_c65 bl_65 br_65 wl_49 vdd gnd cell_6t
Xbit_r50_c65 bl_65 br_65 wl_50 vdd gnd cell_6t
Xbit_r51_c65 bl_65 br_65 wl_51 vdd gnd cell_6t
Xbit_r52_c65 bl_65 br_65 wl_52 vdd gnd cell_6t
Xbit_r53_c65 bl_65 br_65 wl_53 vdd gnd cell_6t
Xbit_r54_c65 bl_65 br_65 wl_54 vdd gnd cell_6t
Xbit_r55_c65 bl_65 br_65 wl_55 vdd gnd cell_6t
Xbit_r56_c65 bl_65 br_65 wl_56 vdd gnd cell_6t
Xbit_r57_c65 bl_65 br_65 wl_57 vdd gnd cell_6t
Xbit_r58_c65 bl_65 br_65 wl_58 vdd gnd cell_6t
Xbit_r59_c65 bl_65 br_65 wl_59 vdd gnd cell_6t
Xbit_r60_c65 bl_65 br_65 wl_60 vdd gnd cell_6t
Xbit_r61_c65 bl_65 br_65 wl_61 vdd gnd cell_6t
Xbit_r62_c65 bl_65 br_65 wl_62 vdd gnd cell_6t
Xbit_r63_c65 bl_65 br_65 wl_63 vdd gnd cell_6t
Xbit_r64_c65 bl_65 br_65 wl_64 vdd gnd cell_6t
Xbit_r65_c65 bl_65 br_65 wl_65 vdd gnd cell_6t
Xbit_r66_c65 bl_65 br_65 wl_66 vdd gnd cell_6t
Xbit_r67_c65 bl_65 br_65 wl_67 vdd gnd cell_6t
Xbit_r68_c65 bl_65 br_65 wl_68 vdd gnd cell_6t
Xbit_r69_c65 bl_65 br_65 wl_69 vdd gnd cell_6t
Xbit_r70_c65 bl_65 br_65 wl_70 vdd gnd cell_6t
Xbit_r71_c65 bl_65 br_65 wl_71 vdd gnd cell_6t
Xbit_r72_c65 bl_65 br_65 wl_72 vdd gnd cell_6t
Xbit_r73_c65 bl_65 br_65 wl_73 vdd gnd cell_6t
Xbit_r74_c65 bl_65 br_65 wl_74 vdd gnd cell_6t
Xbit_r75_c65 bl_65 br_65 wl_75 vdd gnd cell_6t
Xbit_r76_c65 bl_65 br_65 wl_76 vdd gnd cell_6t
Xbit_r77_c65 bl_65 br_65 wl_77 vdd gnd cell_6t
Xbit_r78_c65 bl_65 br_65 wl_78 vdd gnd cell_6t
Xbit_r79_c65 bl_65 br_65 wl_79 vdd gnd cell_6t
Xbit_r80_c65 bl_65 br_65 wl_80 vdd gnd cell_6t
Xbit_r81_c65 bl_65 br_65 wl_81 vdd gnd cell_6t
Xbit_r82_c65 bl_65 br_65 wl_82 vdd gnd cell_6t
Xbit_r83_c65 bl_65 br_65 wl_83 vdd gnd cell_6t
Xbit_r84_c65 bl_65 br_65 wl_84 vdd gnd cell_6t
Xbit_r85_c65 bl_65 br_65 wl_85 vdd gnd cell_6t
Xbit_r86_c65 bl_65 br_65 wl_86 vdd gnd cell_6t
Xbit_r87_c65 bl_65 br_65 wl_87 vdd gnd cell_6t
Xbit_r88_c65 bl_65 br_65 wl_88 vdd gnd cell_6t
Xbit_r89_c65 bl_65 br_65 wl_89 vdd gnd cell_6t
Xbit_r90_c65 bl_65 br_65 wl_90 vdd gnd cell_6t
Xbit_r91_c65 bl_65 br_65 wl_91 vdd gnd cell_6t
Xbit_r92_c65 bl_65 br_65 wl_92 vdd gnd cell_6t
Xbit_r93_c65 bl_65 br_65 wl_93 vdd gnd cell_6t
Xbit_r94_c65 bl_65 br_65 wl_94 vdd gnd cell_6t
Xbit_r95_c65 bl_65 br_65 wl_95 vdd gnd cell_6t
Xbit_r96_c65 bl_65 br_65 wl_96 vdd gnd cell_6t
Xbit_r97_c65 bl_65 br_65 wl_97 vdd gnd cell_6t
Xbit_r98_c65 bl_65 br_65 wl_98 vdd gnd cell_6t
Xbit_r99_c65 bl_65 br_65 wl_99 vdd gnd cell_6t
Xbit_r100_c65 bl_65 br_65 wl_100 vdd gnd cell_6t
Xbit_r101_c65 bl_65 br_65 wl_101 vdd gnd cell_6t
Xbit_r102_c65 bl_65 br_65 wl_102 vdd gnd cell_6t
Xbit_r103_c65 bl_65 br_65 wl_103 vdd gnd cell_6t
Xbit_r104_c65 bl_65 br_65 wl_104 vdd gnd cell_6t
Xbit_r105_c65 bl_65 br_65 wl_105 vdd gnd cell_6t
Xbit_r106_c65 bl_65 br_65 wl_106 vdd gnd cell_6t
Xbit_r107_c65 bl_65 br_65 wl_107 vdd gnd cell_6t
Xbit_r108_c65 bl_65 br_65 wl_108 vdd gnd cell_6t
Xbit_r109_c65 bl_65 br_65 wl_109 vdd gnd cell_6t
Xbit_r110_c65 bl_65 br_65 wl_110 vdd gnd cell_6t
Xbit_r111_c65 bl_65 br_65 wl_111 vdd gnd cell_6t
Xbit_r112_c65 bl_65 br_65 wl_112 vdd gnd cell_6t
Xbit_r113_c65 bl_65 br_65 wl_113 vdd gnd cell_6t
Xbit_r114_c65 bl_65 br_65 wl_114 vdd gnd cell_6t
Xbit_r115_c65 bl_65 br_65 wl_115 vdd gnd cell_6t
Xbit_r116_c65 bl_65 br_65 wl_116 vdd gnd cell_6t
Xbit_r117_c65 bl_65 br_65 wl_117 vdd gnd cell_6t
Xbit_r118_c65 bl_65 br_65 wl_118 vdd gnd cell_6t
Xbit_r119_c65 bl_65 br_65 wl_119 vdd gnd cell_6t
Xbit_r120_c65 bl_65 br_65 wl_120 vdd gnd cell_6t
Xbit_r121_c65 bl_65 br_65 wl_121 vdd gnd cell_6t
Xbit_r122_c65 bl_65 br_65 wl_122 vdd gnd cell_6t
Xbit_r123_c65 bl_65 br_65 wl_123 vdd gnd cell_6t
Xbit_r124_c65 bl_65 br_65 wl_124 vdd gnd cell_6t
Xbit_r125_c65 bl_65 br_65 wl_125 vdd gnd cell_6t
Xbit_r126_c65 bl_65 br_65 wl_126 vdd gnd cell_6t
Xbit_r127_c65 bl_65 br_65 wl_127 vdd gnd cell_6t
Xbit_r128_c65 bl_65 br_65 wl_128 vdd gnd cell_6t
Xbit_r129_c65 bl_65 br_65 wl_129 vdd gnd cell_6t
Xbit_r130_c65 bl_65 br_65 wl_130 vdd gnd cell_6t
Xbit_r131_c65 bl_65 br_65 wl_131 vdd gnd cell_6t
Xbit_r132_c65 bl_65 br_65 wl_132 vdd gnd cell_6t
Xbit_r133_c65 bl_65 br_65 wl_133 vdd gnd cell_6t
Xbit_r134_c65 bl_65 br_65 wl_134 vdd gnd cell_6t
Xbit_r135_c65 bl_65 br_65 wl_135 vdd gnd cell_6t
Xbit_r136_c65 bl_65 br_65 wl_136 vdd gnd cell_6t
Xbit_r137_c65 bl_65 br_65 wl_137 vdd gnd cell_6t
Xbit_r138_c65 bl_65 br_65 wl_138 vdd gnd cell_6t
Xbit_r139_c65 bl_65 br_65 wl_139 vdd gnd cell_6t
Xbit_r140_c65 bl_65 br_65 wl_140 vdd gnd cell_6t
Xbit_r141_c65 bl_65 br_65 wl_141 vdd gnd cell_6t
Xbit_r142_c65 bl_65 br_65 wl_142 vdd gnd cell_6t
Xbit_r143_c65 bl_65 br_65 wl_143 vdd gnd cell_6t
Xbit_r144_c65 bl_65 br_65 wl_144 vdd gnd cell_6t
Xbit_r145_c65 bl_65 br_65 wl_145 vdd gnd cell_6t
Xbit_r146_c65 bl_65 br_65 wl_146 vdd gnd cell_6t
Xbit_r147_c65 bl_65 br_65 wl_147 vdd gnd cell_6t
Xbit_r148_c65 bl_65 br_65 wl_148 vdd gnd cell_6t
Xbit_r149_c65 bl_65 br_65 wl_149 vdd gnd cell_6t
Xbit_r150_c65 bl_65 br_65 wl_150 vdd gnd cell_6t
Xbit_r151_c65 bl_65 br_65 wl_151 vdd gnd cell_6t
Xbit_r152_c65 bl_65 br_65 wl_152 vdd gnd cell_6t
Xbit_r153_c65 bl_65 br_65 wl_153 vdd gnd cell_6t
Xbit_r154_c65 bl_65 br_65 wl_154 vdd gnd cell_6t
Xbit_r155_c65 bl_65 br_65 wl_155 vdd gnd cell_6t
Xbit_r156_c65 bl_65 br_65 wl_156 vdd gnd cell_6t
Xbit_r157_c65 bl_65 br_65 wl_157 vdd gnd cell_6t
Xbit_r158_c65 bl_65 br_65 wl_158 vdd gnd cell_6t
Xbit_r159_c65 bl_65 br_65 wl_159 vdd gnd cell_6t
Xbit_r160_c65 bl_65 br_65 wl_160 vdd gnd cell_6t
Xbit_r161_c65 bl_65 br_65 wl_161 vdd gnd cell_6t
Xbit_r162_c65 bl_65 br_65 wl_162 vdd gnd cell_6t
Xbit_r163_c65 bl_65 br_65 wl_163 vdd gnd cell_6t
Xbit_r164_c65 bl_65 br_65 wl_164 vdd gnd cell_6t
Xbit_r165_c65 bl_65 br_65 wl_165 vdd gnd cell_6t
Xbit_r166_c65 bl_65 br_65 wl_166 vdd gnd cell_6t
Xbit_r167_c65 bl_65 br_65 wl_167 vdd gnd cell_6t
Xbit_r168_c65 bl_65 br_65 wl_168 vdd gnd cell_6t
Xbit_r169_c65 bl_65 br_65 wl_169 vdd gnd cell_6t
Xbit_r170_c65 bl_65 br_65 wl_170 vdd gnd cell_6t
Xbit_r171_c65 bl_65 br_65 wl_171 vdd gnd cell_6t
Xbit_r172_c65 bl_65 br_65 wl_172 vdd gnd cell_6t
Xbit_r173_c65 bl_65 br_65 wl_173 vdd gnd cell_6t
Xbit_r174_c65 bl_65 br_65 wl_174 vdd gnd cell_6t
Xbit_r175_c65 bl_65 br_65 wl_175 vdd gnd cell_6t
Xbit_r176_c65 bl_65 br_65 wl_176 vdd gnd cell_6t
Xbit_r177_c65 bl_65 br_65 wl_177 vdd gnd cell_6t
Xbit_r178_c65 bl_65 br_65 wl_178 vdd gnd cell_6t
Xbit_r179_c65 bl_65 br_65 wl_179 vdd gnd cell_6t
Xbit_r180_c65 bl_65 br_65 wl_180 vdd gnd cell_6t
Xbit_r181_c65 bl_65 br_65 wl_181 vdd gnd cell_6t
Xbit_r182_c65 bl_65 br_65 wl_182 vdd gnd cell_6t
Xbit_r183_c65 bl_65 br_65 wl_183 vdd gnd cell_6t
Xbit_r184_c65 bl_65 br_65 wl_184 vdd gnd cell_6t
Xbit_r185_c65 bl_65 br_65 wl_185 vdd gnd cell_6t
Xbit_r186_c65 bl_65 br_65 wl_186 vdd gnd cell_6t
Xbit_r187_c65 bl_65 br_65 wl_187 vdd gnd cell_6t
Xbit_r188_c65 bl_65 br_65 wl_188 vdd gnd cell_6t
Xbit_r189_c65 bl_65 br_65 wl_189 vdd gnd cell_6t
Xbit_r190_c65 bl_65 br_65 wl_190 vdd gnd cell_6t
Xbit_r191_c65 bl_65 br_65 wl_191 vdd gnd cell_6t
Xbit_r192_c65 bl_65 br_65 wl_192 vdd gnd cell_6t
Xbit_r193_c65 bl_65 br_65 wl_193 vdd gnd cell_6t
Xbit_r194_c65 bl_65 br_65 wl_194 vdd gnd cell_6t
Xbit_r195_c65 bl_65 br_65 wl_195 vdd gnd cell_6t
Xbit_r196_c65 bl_65 br_65 wl_196 vdd gnd cell_6t
Xbit_r197_c65 bl_65 br_65 wl_197 vdd gnd cell_6t
Xbit_r198_c65 bl_65 br_65 wl_198 vdd gnd cell_6t
Xbit_r199_c65 bl_65 br_65 wl_199 vdd gnd cell_6t
Xbit_r200_c65 bl_65 br_65 wl_200 vdd gnd cell_6t
Xbit_r201_c65 bl_65 br_65 wl_201 vdd gnd cell_6t
Xbit_r202_c65 bl_65 br_65 wl_202 vdd gnd cell_6t
Xbit_r203_c65 bl_65 br_65 wl_203 vdd gnd cell_6t
Xbit_r204_c65 bl_65 br_65 wl_204 vdd gnd cell_6t
Xbit_r205_c65 bl_65 br_65 wl_205 vdd gnd cell_6t
Xbit_r206_c65 bl_65 br_65 wl_206 vdd gnd cell_6t
Xbit_r207_c65 bl_65 br_65 wl_207 vdd gnd cell_6t
Xbit_r208_c65 bl_65 br_65 wl_208 vdd gnd cell_6t
Xbit_r209_c65 bl_65 br_65 wl_209 vdd gnd cell_6t
Xbit_r210_c65 bl_65 br_65 wl_210 vdd gnd cell_6t
Xbit_r211_c65 bl_65 br_65 wl_211 vdd gnd cell_6t
Xbit_r212_c65 bl_65 br_65 wl_212 vdd gnd cell_6t
Xbit_r213_c65 bl_65 br_65 wl_213 vdd gnd cell_6t
Xbit_r214_c65 bl_65 br_65 wl_214 vdd gnd cell_6t
Xbit_r215_c65 bl_65 br_65 wl_215 vdd gnd cell_6t
Xbit_r216_c65 bl_65 br_65 wl_216 vdd gnd cell_6t
Xbit_r217_c65 bl_65 br_65 wl_217 vdd gnd cell_6t
Xbit_r218_c65 bl_65 br_65 wl_218 vdd gnd cell_6t
Xbit_r219_c65 bl_65 br_65 wl_219 vdd gnd cell_6t
Xbit_r220_c65 bl_65 br_65 wl_220 vdd gnd cell_6t
Xbit_r221_c65 bl_65 br_65 wl_221 vdd gnd cell_6t
Xbit_r222_c65 bl_65 br_65 wl_222 vdd gnd cell_6t
Xbit_r223_c65 bl_65 br_65 wl_223 vdd gnd cell_6t
Xbit_r224_c65 bl_65 br_65 wl_224 vdd gnd cell_6t
Xbit_r225_c65 bl_65 br_65 wl_225 vdd gnd cell_6t
Xbit_r226_c65 bl_65 br_65 wl_226 vdd gnd cell_6t
Xbit_r227_c65 bl_65 br_65 wl_227 vdd gnd cell_6t
Xbit_r228_c65 bl_65 br_65 wl_228 vdd gnd cell_6t
Xbit_r229_c65 bl_65 br_65 wl_229 vdd gnd cell_6t
Xbit_r230_c65 bl_65 br_65 wl_230 vdd gnd cell_6t
Xbit_r231_c65 bl_65 br_65 wl_231 vdd gnd cell_6t
Xbit_r232_c65 bl_65 br_65 wl_232 vdd gnd cell_6t
Xbit_r233_c65 bl_65 br_65 wl_233 vdd gnd cell_6t
Xbit_r234_c65 bl_65 br_65 wl_234 vdd gnd cell_6t
Xbit_r235_c65 bl_65 br_65 wl_235 vdd gnd cell_6t
Xbit_r236_c65 bl_65 br_65 wl_236 vdd gnd cell_6t
Xbit_r237_c65 bl_65 br_65 wl_237 vdd gnd cell_6t
Xbit_r238_c65 bl_65 br_65 wl_238 vdd gnd cell_6t
Xbit_r239_c65 bl_65 br_65 wl_239 vdd gnd cell_6t
Xbit_r240_c65 bl_65 br_65 wl_240 vdd gnd cell_6t
Xbit_r241_c65 bl_65 br_65 wl_241 vdd gnd cell_6t
Xbit_r242_c65 bl_65 br_65 wl_242 vdd gnd cell_6t
Xbit_r243_c65 bl_65 br_65 wl_243 vdd gnd cell_6t
Xbit_r244_c65 bl_65 br_65 wl_244 vdd gnd cell_6t
Xbit_r245_c65 bl_65 br_65 wl_245 vdd gnd cell_6t
Xbit_r246_c65 bl_65 br_65 wl_246 vdd gnd cell_6t
Xbit_r247_c65 bl_65 br_65 wl_247 vdd gnd cell_6t
Xbit_r248_c65 bl_65 br_65 wl_248 vdd gnd cell_6t
Xbit_r249_c65 bl_65 br_65 wl_249 vdd gnd cell_6t
Xbit_r250_c65 bl_65 br_65 wl_250 vdd gnd cell_6t
Xbit_r251_c65 bl_65 br_65 wl_251 vdd gnd cell_6t
Xbit_r252_c65 bl_65 br_65 wl_252 vdd gnd cell_6t
Xbit_r253_c65 bl_65 br_65 wl_253 vdd gnd cell_6t
Xbit_r254_c65 bl_65 br_65 wl_254 vdd gnd cell_6t
Xbit_r255_c65 bl_65 br_65 wl_255 vdd gnd cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd cell_6t
Xbit_r1_c66 bl_66 br_66 wl_1 vdd gnd cell_6t
Xbit_r2_c66 bl_66 br_66 wl_2 vdd gnd cell_6t
Xbit_r3_c66 bl_66 br_66 wl_3 vdd gnd cell_6t
Xbit_r4_c66 bl_66 br_66 wl_4 vdd gnd cell_6t
Xbit_r5_c66 bl_66 br_66 wl_5 vdd gnd cell_6t
Xbit_r6_c66 bl_66 br_66 wl_6 vdd gnd cell_6t
Xbit_r7_c66 bl_66 br_66 wl_7 vdd gnd cell_6t
Xbit_r8_c66 bl_66 br_66 wl_8 vdd gnd cell_6t
Xbit_r9_c66 bl_66 br_66 wl_9 vdd gnd cell_6t
Xbit_r10_c66 bl_66 br_66 wl_10 vdd gnd cell_6t
Xbit_r11_c66 bl_66 br_66 wl_11 vdd gnd cell_6t
Xbit_r12_c66 bl_66 br_66 wl_12 vdd gnd cell_6t
Xbit_r13_c66 bl_66 br_66 wl_13 vdd gnd cell_6t
Xbit_r14_c66 bl_66 br_66 wl_14 vdd gnd cell_6t
Xbit_r15_c66 bl_66 br_66 wl_15 vdd gnd cell_6t
Xbit_r16_c66 bl_66 br_66 wl_16 vdd gnd cell_6t
Xbit_r17_c66 bl_66 br_66 wl_17 vdd gnd cell_6t
Xbit_r18_c66 bl_66 br_66 wl_18 vdd gnd cell_6t
Xbit_r19_c66 bl_66 br_66 wl_19 vdd gnd cell_6t
Xbit_r20_c66 bl_66 br_66 wl_20 vdd gnd cell_6t
Xbit_r21_c66 bl_66 br_66 wl_21 vdd gnd cell_6t
Xbit_r22_c66 bl_66 br_66 wl_22 vdd gnd cell_6t
Xbit_r23_c66 bl_66 br_66 wl_23 vdd gnd cell_6t
Xbit_r24_c66 bl_66 br_66 wl_24 vdd gnd cell_6t
Xbit_r25_c66 bl_66 br_66 wl_25 vdd gnd cell_6t
Xbit_r26_c66 bl_66 br_66 wl_26 vdd gnd cell_6t
Xbit_r27_c66 bl_66 br_66 wl_27 vdd gnd cell_6t
Xbit_r28_c66 bl_66 br_66 wl_28 vdd gnd cell_6t
Xbit_r29_c66 bl_66 br_66 wl_29 vdd gnd cell_6t
Xbit_r30_c66 bl_66 br_66 wl_30 vdd gnd cell_6t
Xbit_r31_c66 bl_66 br_66 wl_31 vdd gnd cell_6t
Xbit_r32_c66 bl_66 br_66 wl_32 vdd gnd cell_6t
Xbit_r33_c66 bl_66 br_66 wl_33 vdd gnd cell_6t
Xbit_r34_c66 bl_66 br_66 wl_34 vdd gnd cell_6t
Xbit_r35_c66 bl_66 br_66 wl_35 vdd gnd cell_6t
Xbit_r36_c66 bl_66 br_66 wl_36 vdd gnd cell_6t
Xbit_r37_c66 bl_66 br_66 wl_37 vdd gnd cell_6t
Xbit_r38_c66 bl_66 br_66 wl_38 vdd gnd cell_6t
Xbit_r39_c66 bl_66 br_66 wl_39 vdd gnd cell_6t
Xbit_r40_c66 bl_66 br_66 wl_40 vdd gnd cell_6t
Xbit_r41_c66 bl_66 br_66 wl_41 vdd gnd cell_6t
Xbit_r42_c66 bl_66 br_66 wl_42 vdd gnd cell_6t
Xbit_r43_c66 bl_66 br_66 wl_43 vdd gnd cell_6t
Xbit_r44_c66 bl_66 br_66 wl_44 vdd gnd cell_6t
Xbit_r45_c66 bl_66 br_66 wl_45 vdd gnd cell_6t
Xbit_r46_c66 bl_66 br_66 wl_46 vdd gnd cell_6t
Xbit_r47_c66 bl_66 br_66 wl_47 vdd gnd cell_6t
Xbit_r48_c66 bl_66 br_66 wl_48 vdd gnd cell_6t
Xbit_r49_c66 bl_66 br_66 wl_49 vdd gnd cell_6t
Xbit_r50_c66 bl_66 br_66 wl_50 vdd gnd cell_6t
Xbit_r51_c66 bl_66 br_66 wl_51 vdd gnd cell_6t
Xbit_r52_c66 bl_66 br_66 wl_52 vdd gnd cell_6t
Xbit_r53_c66 bl_66 br_66 wl_53 vdd gnd cell_6t
Xbit_r54_c66 bl_66 br_66 wl_54 vdd gnd cell_6t
Xbit_r55_c66 bl_66 br_66 wl_55 vdd gnd cell_6t
Xbit_r56_c66 bl_66 br_66 wl_56 vdd gnd cell_6t
Xbit_r57_c66 bl_66 br_66 wl_57 vdd gnd cell_6t
Xbit_r58_c66 bl_66 br_66 wl_58 vdd gnd cell_6t
Xbit_r59_c66 bl_66 br_66 wl_59 vdd gnd cell_6t
Xbit_r60_c66 bl_66 br_66 wl_60 vdd gnd cell_6t
Xbit_r61_c66 bl_66 br_66 wl_61 vdd gnd cell_6t
Xbit_r62_c66 bl_66 br_66 wl_62 vdd gnd cell_6t
Xbit_r63_c66 bl_66 br_66 wl_63 vdd gnd cell_6t
Xbit_r64_c66 bl_66 br_66 wl_64 vdd gnd cell_6t
Xbit_r65_c66 bl_66 br_66 wl_65 vdd gnd cell_6t
Xbit_r66_c66 bl_66 br_66 wl_66 vdd gnd cell_6t
Xbit_r67_c66 bl_66 br_66 wl_67 vdd gnd cell_6t
Xbit_r68_c66 bl_66 br_66 wl_68 vdd gnd cell_6t
Xbit_r69_c66 bl_66 br_66 wl_69 vdd gnd cell_6t
Xbit_r70_c66 bl_66 br_66 wl_70 vdd gnd cell_6t
Xbit_r71_c66 bl_66 br_66 wl_71 vdd gnd cell_6t
Xbit_r72_c66 bl_66 br_66 wl_72 vdd gnd cell_6t
Xbit_r73_c66 bl_66 br_66 wl_73 vdd gnd cell_6t
Xbit_r74_c66 bl_66 br_66 wl_74 vdd gnd cell_6t
Xbit_r75_c66 bl_66 br_66 wl_75 vdd gnd cell_6t
Xbit_r76_c66 bl_66 br_66 wl_76 vdd gnd cell_6t
Xbit_r77_c66 bl_66 br_66 wl_77 vdd gnd cell_6t
Xbit_r78_c66 bl_66 br_66 wl_78 vdd gnd cell_6t
Xbit_r79_c66 bl_66 br_66 wl_79 vdd gnd cell_6t
Xbit_r80_c66 bl_66 br_66 wl_80 vdd gnd cell_6t
Xbit_r81_c66 bl_66 br_66 wl_81 vdd gnd cell_6t
Xbit_r82_c66 bl_66 br_66 wl_82 vdd gnd cell_6t
Xbit_r83_c66 bl_66 br_66 wl_83 vdd gnd cell_6t
Xbit_r84_c66 bl_66 br_66 wl_84 vdd gnd cell_6t
Xbit_r85_c66 bl_66 br_66 wl_85 vdd gnd cell_6t
Xbit_r86_c66 bl_66 br_66 wl_86 vdd gnd cell_6t
Xbit_r87_c66 bl_66 br_66 wl_87 vdd gnd cell_6t
Xbit_r88_c66 bl_66 br_66 wl_88 vdd gnd cell_6t
Xbit_r89_c66 bl_66 br_66 wl_89 vdd gnd cell_6t
Xbit_r90_c66 bl_66 br_66 wl_90 vdd gnd cell_6t
Xbit_r91_c66 bl_66 br_66 wl_91 vdd gnd cell_6t
Xbit_r92_c66 bl_66 br_66 wl_92 vdd gnd cell_6t
Xbit_r93_c66 bl_66 br_66 wl_93 vdd gnd cell_6t
Xbit_r94_c66 bl_66 br_66 wl_94 vdd gnd cell_6t
Xbit_r95_c66 bl_66 br_66 wl_95 vdd gnd cell_6t
Xbit_r96_c66 bl_66 br_66 wl_96 vdd gnd cell_6t
Xbit_r97_c66 bl_66 br_66 wl_97 vdd gnd cell_6t
Xbit_r98_c66 bl_66 br_66 wl_98 vdd gnd cell_6t
Xbit_r99_c66 bl_66 br_66 wl_99 vdd gnd cell_6t
Xbit_r100_c66 bl_66 br_66 wl_100 vdd gnd cell_6t
Xbit_r101_c66 bl_66 br_66 wl_101 vdd gnd cell_6t
Xbit_r102_c66 bl_66 br_66 wl_102 vdd gnd cell_6t
Xbit_r103_c66 bl_66 br_66 wl_103 vdd gnd cell_6t
Xbit_r104_c66 bl_66 br_66 wl_104 vdd gnd cell_6t
Xbit_r105_c66 bl_66 br_66 wl_105 vdd gnd cell_6t
Xbit_r106_c66 bl_66 br_66 wl_106 vdd gnd cell_6t
Xbit_r107_c66 bl_66 br_66 wl_107 vdd gnd cell_6t
Xbit_r108_c66 bl_66 br_66 wl_108 vdd gnd cell_6t
Xbit_r109_c66 bl_66 br_66 wl_109 vdd gnd cell_6t
Xbit_r110_c66 bl_66 br_66 wl_110 vdd gnd cell_6t
Xbit_r111_c66 bl_66 br_66 wl_111 vdd gnd cell_6t
Xbit_r112_c66 bl_66 br_66 wl_112 vdd gnd cell_6t
Xbit_r113_c66 bl_66 br_66 wl_113 vdd gnd cell_6t
Xbit_r114_c66 bl_66 br_66 wl_114 vdd gnd cell_6t
Xbit_r115_c66 bl_66 br_66 wl_115 vdd gnd cell_6t
Xbit_r116_c66 bl_66 br_66 wl_116 vdd gnd cell_6t
Xbit_r117_c66 bl_66 br_66 wl_117 vdd gnd cell_6t
Xbit_r118_c66 bl_66 br_66 wl_118 vdd gnd cell_6t
Xbit_r119_c66 bl_66 br_66 wl_119 vdd gnd cell_6t
Xbit_r120_c66 bl_66 br_66 wl_120 vdd gnd cell_6t
Xbit_r121_c66 bl_66 br_66 wl_121 vdd gnd cell_6t
Xbit_r122_c66 bl_66 br_66 wl_122 vdd gnd cell_6t
Xbit_r123_c66 bl_66 br_66 wl_123 vdd gnd cell_6t
Xbit_r124_c66 bl_66 br_66 wl_124 vdd gnd cell_6t
Xbit_r125_c66 bl_66 br_66 wl_125 vdd gnd cell_6t
Xbit_r126_c66 bl_66 br_66 wl_126 vdd gnd cell_6t
Xbit_r127_c66 bl_66 br_66 wl_127 vdd gnd cell_6t
Xbit_r128_c66 bl_66 br_66 wl_128 vdd gnd cell_6t
Xbit_r129_c66 bl_66 br_66 wl_129 vdd gnd cell_6t
Xbit_r130_c66 bl_66 br_66 wl_130 vdd gnd cell_6t
Xbit_r131_c66 bl_66 br_66 wl_131 vdd gnd cell_6t
Xbit_r132_c66 bl_66 br_66 wl_132 vdd gnd cell_6t
Xbit_r133_c66 bl_66 br_66 wl_133 vdd gnd cell_6t
Xbit_r134_c66 bl_66 br_66 wl_134 vdd gnd cell_6t
Xbit_r135_c66 bl_66 br_66 wl_135 vdd gnd cell_6t
Xbit_r136_c66 bl_66 br_66 wl_136 vdd gnd cell_6t
Xbit_r137_c66 bl_66 br_66 wl_137 vdd gnd cell_6t
Xbit_r138_c66 bl_66 br_66 wl_138 vdd gnd cell_6t
Xbit_r139_c66 bl_66 br_66 wl_139 vdd gnd cell_6t
Xbit_r140_c66 bl_66 br_66 wl_140 vdd gnd cell_6t
Xbit_r141_c66 bl_66 br_66 wl_141 vdd gnd cell_6t
Xbit_r142_c66 bl_66 br_66 wl_142 vdd gnd cell_6t
Xbit_r143_c66 bl_66 br_66 wl_143 vdd gnd cell_6t
Xbit_r144_c66 bl_66 br_66 wl_144 vdd gnd cell_6t
Xbit_r145_c66 bl_66 br_66 wl_145 vdd gnd cell_6t
Xbit_r146_c66 bl_66 br_66 wl_146 vdd gnd cell_6t
Xbit_r147_c66 bl_66 br_66 wl_147 vdd gnd cell_6t
Xbit_r148_c66 bl_66 br_66 wl_148 vdd gnd cell_6t
Xbit_r149_c66 bl_66 br_66 wl_149 vdd gnd cell_6t
Xbit_r150_c66 bl_66 br_66 wl_150 vdd gnd cell_6t
Xbit_r151_c66 bl_66 br_66 wl_151 vdd gnd cell_6t
Xbit_r152_c66 bl_66 br_66 wl_152 vdd gnd cell_6t
Xbit_r153_c66 bl_66 br_66 wl_153 vdd gnd cell_6t
Xbit_r154_c66 bl_66 br_66 wl_154 vdd gnd cell_6t
Xbit_r155_c66 bl_66 br_66 wl_155 vdd gnd cell_6t
Xbit_r156_c66 bl_66 br_66 wl_156 vdd gnd cell_6t
Xbit_r157_c66 bl_66 br_66 wl_157 vdd gnd cell_6t
Xbit_r158_c66 bl_66 br_66 wl_158 vdd gnd cell_6t
Xbit_r159_c66 bl_66 br_66 wl_159 vdd gnd cell_6t
Xbit_r160_c66 bl_66 br_66 wl_160 vdd gnd cell_6t
Xbit_r161_c66 bl_66 br_66 wl_161 vdd gnd cell_6t
Xbit_r162_c66 bl_66 br_66 wl_162 vdd gnd cell_6t
Xbit_r163_c66 bl_66 br_66 wl_163 vdd gnd cell_6t
Xbit_r164_c66 bl_66 br_66 wl_164 vdd gnd cell_6t
Xbit_r165_c66 bl_66 br_66 wl_165 vdd gnd cell_6t
Xbit_r166_c66 bl_66 br_66 wl_166 vdd gnd cell_6t
Xbit_r167_c66 bl_66 br_66 wl_167 vdd gnd cell_6t
Xbit_r168_c66 bl_66 br_66 wl_168 vdd gnd cell_6t
Xbit_r169_c66 bl_66 br_66 wl_169 vdd gnd cell_6t
Xbit_r170_c66 bl_66 br_66 wl_170 vdd gnd cell_6t
Xbit_r171_c66 bl_66 br_66 wl_171 vdd gnd cell_6t
Xbit_r172_c66 bl_66 br_66 wl_172 vdd gnd cell_6t
Xbit_r173_c66 bl_66 br_66 wl_173 vdd gnd cell_6t
Xbit_r174_c66 bl_66 br_66 wl_174 vdd gnd cell_6t
Xbit_r175_c66 bl_66 br_66 wl_175 vdd gnd cell_6t
Xbit_r176_c66 bl_66 br_66 wl_176 vdd gnd cell_6t
Xbit_r177_c66 bl_66 br_66 wl_177 vdd gnd cell_6t
Xbit_r178_c66 bl_66 br_66 wl_178 vdd gnd cell_6t
Xbit_r179_c66 bl_66 br_66 wl_179 vdd gnd cell_6t
Xbit_r180_c66 bl_66 br_66 wl_180 vdd gnd cell_6t
Xbit_r181_c66 bl_66 br_66 wl_181 vdd gnd cell_6t
Xbit_r182_c66 bl_66 br_66 wl_182 vdd gnd cell_6t
Xbit_r183_c66 bl_66 br_66 wl_183 vdd gnd cell_6t
Xbit_r184_c66 bl_66 br_66 wl_184 vdd gnd cell_6t
Xbit_r185_c66 bl_66 br_66 wl_185 vdd gnd cell_6t
Xbit_r186_c66 bl_66 br_66 wl_186 vdd gnd cell_6t
Xbit_r187_c66 bl_66 br_66 wl_187 vdd gnd cell_6t
Xbit_r188_c66 bl_66 br_66 wl_188 vdd gnd cell_6t
Xbit_r189_c66 bl_66 br_66 wl_189 vdd gnd cell_6t
Xbit_r190_c66 bl_66 br_66 wl_190 vdd gnd cell_6t
Xbit_r191_c66 bl_66 br_66 wl_191 vdd gnd cell_6t
Xbit_r192_c66 bl_66 br_66 wl_192 vdd gnd cell_6t
Xbit_r193_c66 bl_66 br_66 wl_193 vdd gnd cell_6t
Xbit_r194_c66 bl_66 br_66 wl_194 vdd gnd cell_6t
Xbit_r195_c66 bl_66 br_66 wl_195 vdd gnd cell_6t
Xbit_r196_c66 bl_66 br_66 wl_196 vdd gnd cell_6t
Xbit_r197_c66 bl_66 br_66 wl_197 vdd gnd cell_6t
Xbit_r198_c66 bl_66 br_66 wl_198 vdd gnd cell_6t
Xbit_r199_c66 bl_66 br_66 wl_199 vdd gnd cell_6t
Xbit_r200_c66 bl_66 br_66 wl_200 vdd gnd cell_6t
Xbit_r201_c66 bl_66 br_66 wl_201 vdd gnd cell_6t
Xbit_r202_c66 bl_66 br_66 wl_202 vdd gnd cell_6t
Xbit_r203_c66 bl_66 br_66 wl_203 vdd gnd cell_6t
Xbit_r204_c66 bl_66 br_66 wl_204 vdd gnd cell_6t
Xbit_r205_c66 bl_66 br_66 wl_205 vdd gnd cell_6t
Xbit_r206_c66 bl_66 br_66 wl_206 vdd gnd cell_6t
Xbit_r207_c66 bl_66 br_66 wl_207 vdd gnd cell_6t
Xbit_r208_c66 bl_66 br_66 wl_208 vdd gnd cell_6t
Xbit_r209_c66 bl_66 br_66 wl_209 vdd gnd cell_6t
Xbit_r210_c66 bl_66 br_66 wl_210 vdd gnd cell_6t
Xbit_r211_c66 bl_66 br_66 wl_211 vdd gnd cell_6t
Xbit_r212_c66 bl_66 br_66 wl_212 vdd gnd cell_6t
Xbit_r213_c66 bl_66 br_66 wl_213 vdd gnd cell_6t
Xbit_r214_c66 bl_66 br_66 wl_214 vdd gnd cell_6t
Xbit_r215_c66 bl_66 br_66 wl_215 vdd gnd cell_6t
Xbit_r216_c66 bl_66 br_66 wl_216 vdd gnd cell_6t
Xbit_r217_c66 bl_66 br_66 wl_217 vdd gnd cell_6t
Xbit_r218_c66 bl_66 br_66 wl_218 vdd gnd cell_6t
Xbit_r219_c66 bl_66 br_66 wl_219 vdd gnd cell_6t
Xbit_r220_c66 bl_66 br_66 wl_220 vdd gnd cell_6t
Xbit_r221_c66 bl_66 br_66 wl_221 vdd gnd cell_6t
Xbit_r222_c66 bl_66 br_66 wl_222 vdd gnd cell_6t
Xbit_r223_c66 bl_66 br_66 wl_223 vdd gnd cell_6t
Xbit_r224_c66 bl_66 br_66 wl_224 vdd gnd cell_6t
Xbit_r225_c66 bl_66 br_66 wl_225 vdd gnd cell_6t
Xbit_r226_c66 bl_66 br_66 wl_226 vdd gnd cell_6t
Xbit_r227_c66 bl_66 br_66 wl_227 vdd gnd cell_6t
Xbit_r228_c66 bl_66 br_66 wl_228 vdd gnd cell_6t
Xbit_r229_c66 bl_66 br_66 wl_229 vdd gnd cell_6t
Xbit_r230_c66 bl_66 br_66 wl_230 vdd gnd cell_6t
Xbit_r231_c66 bl_66 br_66 wl_231 vdd gnd cell_6t
Xbit_r232_c66 bl_66 br_66 wl_232 vdd gnd cell_6t
Xbit_r233_c66 bl_66 br_66 wl_233 vdd gnd cell_6t
Xbit_r234_c66 bl_66 br_66 wl_234 vdd gnd cell_6t
Xbit_r235_c66 bl_66 br_66 wl_235 vdd gnd cell_6t
Xbit_r236_c66 bl_66 br_66 wl_236 vdd gnd cell_6t
Xbit_r237_c66 bl_66 br_66 wl_237 vdd gnd cell_6t
Xbit_r238_c66 bl_66 br_66 wl_238 vdd gnd cell_6t
Xbit_r239_c66 bl_66 br_66 wl_239 vdd gnd cell_6t
Xbit_r240_c66 bl_66 br_66 wl_240 vdd gnd cell_6t
Xbit_r241_c66 bl_66 br_66 wl_241 vdd gnd cell_6t
Xbit_r242_c66 bl_66 br_66 wl_242 vdd gnd cell_6t
Xbit_r243_c66 bl_66 br_66 wl_243 vdd gnd cell_6t
Xbit_r244_c66 bl_66 br_66 wl_244 vdd gnd cell_6t
Xbit_r245_c66 bl_66 br_66 wl_245 vdd gnd cell_6t
Xbit_r246_c66 bl_66 br_66 wl_246 vdd gnd cell_6t
Xbit_r247_c66 bl_66 br_66 wl_247 vdd gnd cell_6t
Xbit_r248_c66 bl_66 br_66 wl_248 vdd gnd cell_6t
Xbit_r249_c66 bl_66 br_66 wl_249 vdd gnd cell_6t
Xbit_r250_c66 bl_66 br_66 wl_250 vdd gnd cell_6t
Xbit_r251_c66 bl_66 br_66 wl_251 vdd gnd cell_6t
Xbit_r252_c66 bl_66 br_66 wl_252 vdd gnd cell_6t
Xbit_r253_c66 bl_66 br_66 wl_253 vdd gnd cell_6t
Xbit_r254_c66 bl_66 br_66 wl_254 vdd gnd cell_6t
Xbit_r255_c66 bl_66 br_66 wl_255 vdd gnd cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd cell_6t
Xbit_r1_c67 bl_67 br_67 wl_1 vdd gnd cell_6t
Xbit_r2_c67 bl_67 br_67 wl_2 vdd gnd cell_6t
Xbit_r3_c67 bl_67 br_67 wl_3 vdd gnd cell_6t
Xbit_r4_c67 bl_67 br_67 wl_4 vdd gnd cell_6t
Xbit_r5_c67 bl_67 br_67 wl_5 vdd gnd cell_6t
Xbit_r6_c67 bl_67 br_67 wl_6 vdd gnd cell_6t
Xbit_r7_c67 bl_67 br_67 wl_7 vdd gnd cell_6t
Xbit_r8_c67 bl_67 br_67 wl_8 vdd gnd cell_6t
Xbit_r9_c67 bl_67 br_67 wl_9 vdd gnd cell_6t
Xbit_r10_c67 bl_67 br_67 wl_10 vdd gnd cell_6t
Xbit_r11_c67 bl_67 br_67 wl_11 vdd gnd cell_6t
Xbit_r12_c67 bl_67 br_67 wl_12 vdd gnd cell_6t
Xbit_r13_c67 bl_67 br_67 wl_13 vdd gnd cell_6t
Xbit_r14_c67 bl_67 br_67 wl_14 vdd gnd cell_6t
Xbit_r15_c67 bl_67 br_67 wl_15 vdd gnd cell_6t
Xbit_r16_c67 bl_67 br_67 wl_16 vdd gnd cell_6t
Xbit_r17_c67 bl_67 br_67 wl_17 vdd gnd cell_6t
Xbit_r18_c67 bl_67 br_67 wl_18 vdd gnd cell_6t
Xbit_r19_c67 bl_67 br_67 wl_19 vdd gnd cell_6t
Xbit_r20_c67 bl_67 br_67 wl_20 vdd gnd cell_6t
Xbit_r21_c67 bl_67 br_67 wl_21 vdd gnd cell_6t
Xbit_r22_c67 bl_67 br_67 wl_22 vdd gnd cell_6t
Xbit_r23_c67 bl_67 br_67 wl_23 vdd gnd cell_6t
Xbit_r24_c67 bl_67 br_67 wl_24 vdd gnd cell_6t
Xbit_r25_c67 bl_67 br_67 wl_25 vdd gnd cell_6t
Xbit_r26_c67 bl_67 br_67 wl_26 vdd gnd cell_6t
Xbit_r27_c67 bl_67 br_67 wl_27 vdd gnd cell_6t
Xbit_r28_c67 bl_67 br_67 wl_28 vdd gnd cell_6t
Xbit_r29_c67 bl_67 br_67 wl_29 vdd gnd cell_6t
Xbit_r30_c67 bl_67 br_67 wl_30 vdd gnd cell_6t
Xbit_r31_c67 bl_67 br_67 wl_31 vdd gnd cell_6t
Xbit_r32_c67 bl_67 br_67 wl_32 vdd gnd cell_6t
Xbit_r33_c67 bl_67 br_67 wl_33 vdd gnd cell_6t
Xbit_r34_c67 bl_67 br_67 wl_34 vdd gnd cell_6t
Xbit_r35_c67 bl_67 br_67 wl_35 vdd gnd cell_6t
Xbit_r36_c67 bl_67 br_67 wl_36 vdd gnd cell_6t
Xbit_r37_c67 bl_67 br_67 wl_37 vdd gnd cell_6t
Xbit_r38_c67 bl_67 br_67 wl_38 vdd gnd cell_6t
Xbit_r39_c67 bl_67 br_67 wl_39 vdd gnd cell_6t
Xbit_r40_c67 bl_67 br_67 wl_40 vdd gnd cell_6t
Xbit_r41_c67 bl_67 br_67 wl_41 vdd gnd cell_6t
Xbit_r42_c67 bl_67 br_67 wl_42 vdd gnd cell_6t
Xbit_r43_c67 bl_67 br_67 wl_43 vdd gnd cell_6t
Xbit_r44_c67 bl_67 br_67 wl_44 vdd gnd cell_6t
Xbit_r45_c67 bl_67 br_67 wl_45 vdd gnd cell_6t
Xbit_r46_c67 bl_67 br_67 wl_46 vdd gnd cell_6t
Xbit_r47_c67 bl_67 br_67 wl_47 vdd gnd cell_6t
Xbit_r48_c67 bl_67 br_67 wl_48 vdd gnd cell_6t
Xbit_r49_c67 bl_67 br_67 wl_49 vdd gnd cell_6t
Xbit_r50_c67 bl_67 br_67 wl_50 vdd gnd cell_6t
Xbit_r51_c67 bl_67 br_67 wl_51 vdd gnd cell_6t
Xbit_r52_c67 bl_67 br_67 wl_52 vdd gnd cell_6t
Xbit_r53_c67 bl_67 br_67 wl_53 vdd gnd cell_6t
Xbit_r54_c67 bl_67 br_67 wl_54 vdd gnd cell_6t
Xbit_r55_c67 bl_67 br_67 wl_55 vdd gnd cell_6t
Xbit_r56_c67 bl_67 br_67 wl_56 vdd gnd cell_6t
Xbit_r57_c67 bl_67 br_67 wl_57 vdd gnd cell_6t
Xbit_r58_c67 bl_67 br_67 wl_58 vdd gnd cell_6t
Xbit_r59_c67 bl_67 br_67 wl_59 vdd gnd cell_6t
Xbit_r60_c67 bl_67 br_67 wl_60 vdd gnd cell_6t
Xbit_r61_c67 bl_67 br_67 wl_61 vdd gnd cell_6t
Xbit_r62_c67 bl_67 br_67 wl_62 vdd gnd cell_6t
Xbit_r63_c67 bl_67 br_67 wl_63 vdd gnd cell_6t
Xbit_r64_c67 bl_67 br_67 wl_64 vdd gnd cell_6t
Xbit_r65_c67 bl_67 br_67 wl_65 vdd gnd cell_6t
Xbit_r66_c67 bl_67 br_67 wl_66 vdd gnd cell_6t
Xbit_r67_c67 bl_67 br_67 wl_67 vdd gnd cell_6t
Xbit_r68_c67 bl_67 br_67 wl_68 vdd gnd cell_6t
Xbit_r69_c67 bl_67 br_67 wl_69 vdd gnd cell_6t
Xbit_r70_c67 bl_67 br_67 wl_70 vdd gnd cell_6t
Xbit_r71_c67 bl_67 br_67 wl_71 vdd gnd cell_6t
Xbit_r72_c67 bl_67 br_67 wl_72 vdd gnd cell_6t
Xbit_r73_c67 bl_67 br_67 wl_73 vdd gnd cell_6t
Xbit_r74_c67 bl_67 br_67 wl_74 vdd gnd cell_6t
Xbit_r75_c67 bl_67 br_67 wl_75 vdd gnd cell_6t
Xbit_r76_c67 bl_67 br_67 wl_76 vdd gnd cell_6t
Xbit_r77_c67 bl_67 br_67 wl_77 vdd gnd cell_6t
Xbit_r78_c67 bl_67 br_67 wl_78 vdd gnd cell_6t
Xbit_r79_c67 bl_67 br_67 wl_79 vdd gnd cell_6t
Xbit_r80_c67 bl_67 br_67 wl_80 vdd gnd cell_6t
Xbit_r81_c67 bl_67 br_67 wl_81 vdd gnd cell_6t
Xbit_r82_c67 bl_67 br_67 wl_82 vdd gnd cell_6t
Xbit_r83_c67 bl_67 br_67 wl_83 vdd gnd cell_6t
Xbit_r84_c67 bl_67 br_67 wl_84 vdd gnd cell_6t
Xbit_r85_c67 bl_67 br_67 wl_85 vdd gnd cell_6t
Xbit_r86_c67 bl_67 br_67 wl_86 vdd gnd cell_6t
Xbit_r87_c67 bl_67 br_67 wl_87 vdd gnd cell_6t
Xbit_r88_c67 bl_67 br_67 wl_88 vdd gnd cell_6t
Xbit_r89_c67 bl_67 br_67 wl_89 vdd gnd cell_6t
Xbit_r90_c67 bl_67 br_67 wl_90 vdd gnd cell_6t
Xbit_r91_c67 bl_67 br_67 wl_91 vdd gnd cell_6t
Xbit_r92_c67 bl_67 br_67 wl_92 vdd gnd cell_6t
Xbit_r93_c67 bl_67 br_67 wl_93 vdd gnd cell_6t
Xbit_r94_c67 bl_67 br_67 wl_94 vdd gnd cell_6t
Xbit_r95_c67 bl_67 br_67 wl_95 vdd gnd cell_6t
Xbit_r96_c67 bl_67 br_67 wl_96 vdd gnd cell_6t
Xbit_r97_c67 bl_67 br_67 wl_97 vdd gnd cell_6t
Xbit_r98_c67 bl_67 br_67 wl_98 vdd gnd cell_6t
Xbit_r99_c67 bl_67 br_67 wl_99 vdd gnd cell_6t
Xbit_r100_c67 bl_67 br_67 wl_100 vdd gnd cell_6t
Xbit_r101_c67 bl_67 br_67 wl_101 vdd gnd cell_6t
Xbit_r102_c67 bl_67 br_67 wl_102 vdd gnd cell_6t
Xbit_r103_c67 bl_67 br_67 wl_103 vdd gnd cell_6t
Xbit_r104_c67 bl_67 br_67 wl_104 vdd gnd cell_6t
Xbit_r105_c67 bl_67 br_67 wl_105 vdd gnd cell_6t
Xbit_r106_c67 bl_67 br_67 wl_106 vdd gnd cell_6t
Xbit_r107_c67 bl_67 br_67 wl_107 vdd gnd cell_6t
Xbit_r108_c67 bl_67 br_67 wl_108 vdd gnd cell_6t
Xbit_r109_c67 bl_67 br_67 wl_109 vdd gnd cell_6t
Xbit_r110_c67 bl_67 br_67 wl_110 vdd gnd cell_6t
Xbit_r111_c67 bl_67 br_67 wl_111 vdd gnd cell_6t
Xbit_r112_c67 bl_67 br_67 wl_112 vdd gnd cell_6t
Xbit_r113_c67 bl_67 br_67 wl_113 vdd gnd cell_6t
Xbit_r114_c67 bl_67 br_67 wl_114 vdd gnd cell_6t
Xbit_r115_c67 bl_67 br_67 wl_115 vdd gnd cell_6t
Xbit_r116_c67 bl_67 br_67 wl_116 vdd gnd cell_6t
Xbit_r117_c67 bl_67 br_67 wl_117 vdd gnd cell_6t
Xbit_r118_c67 bl_67 br_67 wl_118 vdd gnd cell_6t
Xbit_r119_c67 bl_67 br_67 wl_119 vdd gnd cell_6t
Xbit_r120_c67 bl_67 br_67 wl_120 vdd gnd cell_6t
Xbit_r121_c67 bl_67 br_67 wl_121 vdd gnd cell_6t
Xbit_r122_c67 bl_67 br_67 wl_122 vdd gnd cell_6t
Xbit_r123_c67 bl_67 br_67 wl_123 vdd gnd cell_6t
Xbit_r124_c67 bl_67 br_67 wl_124 vdd gnd cell_6t
Xbit_r125_c67 bl_67 br_67 wl_125 vdd gnd cell_6t
Xbit_r126_c67 bl_67 br_67 wl_126 vdd gnd cell_6t
Xbit_r127_c67 bl_67 br_67 wl_127 vdd gnd cell_6t
Xbit_r128_c67 bl_67 br_67 wl_128 vdd gnd cell_6t
Xbit_r129_c67 bl_67 br_67 wl_129 vdd gnd cell_6t
Xbit_r130_c67 bl_67 br_67 wl_130 vdd gnd cell_6t
Xbit_r131_c67 bl_67 br_67 wl_131 vdd gnd cell_6t
Xbit_r132_c67 bl_67 br_67 wl_132 vdd gnd cell_6t
Xbit_r133_c67 bl_67 br_67 wl_133 vdd gnd cell_6t
Xbit_r134_c67 bl_67 br_67 wl_134 vdd gnd cell_6t
Xbit_r135_c67 bl_67 br_67 wl_135 vdd gnd cell_6t
Xbit_r136_c67 bl_67 br_67 wl_136 vdd gnd cell_6t
Xbit_r137_c67 bl_67 br_67 wl_137 vdd gnd cell_6t
Xbit_r138_c67 bl_67 br_67 wl_138 vdd gnd cell_6t
Xbit_r139_c67 bl_67 br_67 wl_139 vdd gnd cell_6t
Xbit_r140_c67 bl_67 br_67 wl_140 vdd gnd cell_6t
Xbit_r141_c67 bl_67 br_67 wl_141 vdd gnd cell_6t
Xbit_r142_c67 bl_67 br_67 wl_142 vdd gnd cell_6t
Xbit_r143_c67 bl_67 br_67 wl_143 vdd gnd cell_6t
Xbit_r144_c67 bl_67 br_67 wl_144 vdd gnd cell_6t
Xbit_r145_c67 bl_67 br_67 wl_145 vdd gnd cell_6t
Xbit_r146_c67 bl_67 br_67 wl_146 vdd gnd cell_6t
Xbit_r147_c67 bl_67 br_67 wl_147 vdd gnd cell_6t
Xbit_r148_c67 bl_67 br_67 wl_148 vdd gnd cell_6t
Xbit_r149_c67 bl_67 br_67 wl_149 vdd gnd cell_6t
Xbit_r150_c67 bl_67 br_67 wl_150 vdd gnd cell_6t
Xbit_r151_c67 bl_67 br_67 wl_151 vdd gnd cell_6t
Xbit_r152_c67 bl_67 br_67 wl_152 vdd gnd cell_6t
Xbit_r153_c67 bl_67 br_67 wl_153 vdd gnd cell_6t
Xbit_r154_c67 bl_67 br_67 wl_154 vdd gnd cell_6t
Xbit_r155_c67 bl_67 br_67 wl_155 vdd gnd cell_6t
Xbit_r156_c67 bl_67 br_67 wl_156 vdd gnd cell_6t
Xbit_r157_c67 bl_67 br_67 wl_157 vdd gnd cell_6t
Xbit_r158_c67 bl_67 br_67 wl_158 vdd gnd cell_6t
Xbit_r159_c67 bl_67 br_67 wl_159 vdd gnd cell_6t
Xbit_r160_c67 bl_67 br_67 wl_160 vdd gnd cell_6t
Xbit_r161_c67 bl_67 br_67 wl_161 vdd gnd cell_6t
Xbit_r162_c67 bl_67 br_67 wl_162 vdd gnd cell_6t
Xbit_r163_c67 bl_67 br_67 wl_163 vdd gnd cell_6t
Xbit_r164_c67 bl_67 br_67 wl_164 vdd gnd cell_6t
Xbit_r165_c67 bl_67 br_67 wl_165 vdd gnd cell_6t
Xbit_r166_c67 bl_67 br_67 wl_166 vdd gnd cell_6t
Xbit_r167_c67 bl_67 br_67 wl_167 vdd gnd cell_6t
Xbit_r168_c67 bl_67 br_67 wl_168 vdd gnd cell_6t
Xbit_r169_c67 bl_67 br_67 wl_169 vdd gnd cell_6t
Xbit_r170_c67 bl_67 br_67 wl_170 vdd gnd cell_6t
Xbit_r171_c67 bl_67 br_67 wl_171 vdd gnd cell_6t
Xbit_r172_c67 bl_67 br_67 wl_172 vdd gnd cell_6t
Xbit_r173_c67 bl_67 br_67 wl_173 vdd gnd cell_6t
Xbit_r174_c67 bl_67 br_67 wl_174 vdd gnd cell_6t
Xbit_r175_c67 bl_67 br_67 wl_175 vdd gnd cell_6t
Xbit_r176_c67 bl_67 br_67 wl_176 vdd gnd cell_6t
Xbit_r177_c67 bl_67 br_67 wl_177 vdd gnd cell_6t
Xbit_r178_c67 bl_67 br_67 wl_178 vdd gnd cell_6t
Xbit_r179_c67 bl_67 br_67 wl_179 vdd gnd cell_6t
Xbit_r180_c67 bl_67 br_67 wl_180 vdd gnd cell_6t
Xbit_r181_c67 bl_67 br_67 wl_181 vdd gnd cell_6t
Xbit_r182_c67 bl_67 br_67 wl_182 vdd gnd cell_6t
Xbit_r183_c67 bl_67 br_67 wl_183 vdd gnd cell_6t
Xbit_r184_c67 bl_67 br_67 wl_184 vdd gnd cell_6t
Xbit_r185_c67 bl_67 br_67 wl_185 vdd gnd cell_6t
Xbit_r186_c67 bl_67 br_67 wl_186 vdd gnd cell_6t
Xbit_r187_c67 bl_67 br_67 wl_187 vdd gnd cell_6t
Xbit_r188_c67 bl_67 br_67 wl_188 vdd gnd cell_6t
Xbit_r189_c67 bl_67 br_67 wl_189 vdd gnd cell_6t
Xbit_r190_c67 bl_67 br_67 wl_190 vdd gnd cell_6t
Xbit_r191_c67 bl_67 br_67 wl_191 vdd gnd cell_6t
Xbit_r192_c67 bl_67 br_67 wl_192 vdd gnd cell_6t
Xbit_r193_c67 bl_67 br_67 wl_193 vdd gnd cell_6t
Xbit_r194_c67 bl_67 br_67 wl_194 vdd gnd cell_6t
Xbit_r195_c67 bl_67 br_67 wl_195 vdd gnd cell_6t
Xbit_r196_c67 bl_67 br_67 wl_196 vdd gnd cell_6t
Xbit_r197_c67 bl_67 br_67 wl_197 vdd gnd cell_6t
Xbit_r198_c67 bl_67 br_67 wl_198 vdd gnd cell_6t
Xbit_r199_c67 bl_67 br_67 wl_199 vdd gnd cell_6t
Xbit_r200_c67 bl_67 br_67 wl_200 vdd gnd cell_6t
Xbit_r201_c67 bl_67 br_67 wl_201 vdd gnd cell_6t
Xbit_r202_c67 bl_67 br_67 wl_202 vdd gnd cell_6t
Xbit_r203_c67 bl_67 br_67 wl_203 vdd gnd cell_6t
Xbit_r204_c67 bl_67 br_67 wl_204 vdd gnd cell_6t
Xbit_r205_c67 bl_67 br_67 wl_205 vdd gnd cell_6t
Xbit_r206_c67 bl_67 br_67 wl_206 vdd gnd cell_6t
Xbit_r207_c67 bl_67 br_67 wl_207 vdd gnd cell_6t
Xbit_r208_c67 bl_67 br_67 wl_208 vdd gnd cell_6t
Xbit_r209_c67 bl_67 br_67 wl_209 vdd gnd cell_6t
Xbit_r210_c67 bl_67 br_67 wl_210 vdd gnd cell_6t
Xbit_r211_c67 bl_67 br_67 wl_211 vdd gnd cell_6t
Xbit_r212_c67 bl_67 br_67 wl_212 vdd gnd cell_6t
Xbit_r213_c67 bl_67 br_67 wl_213 vdd gnd cell_6t
Xbit_r214_c67 bl_67 br_67 wl_214 vdd gnd cell_6t
Xbit_r215_c67 bl_67 br_67 wl_215 vdd gnd cell_6t
Xbit_r216_c67 bl_67 br_67 wl_216 vdd gnd cell_6t
Xbit_r217_c67 bl_67 br_67 wl_217 vdd gnd cell_6t
Xbit_r218_c67 bl_67 br_67 wl_218 vdd gnd cell_6t
Xbit_r219_c67 bl_67 br_67 wl_219 vdd gnd cell_6t
Xbit_r220_c67 bl_67 br_67 wl_220 vdd gnd cell_6t
Xbit_r221_c67 bl_67 br_67 wl_221 vdd gnd cell_6t
Xbit_r222_c67 bl_67 br_67 wl_222 vdd gnd cell_6t
Xbit_r223_c67 bl_67 br_67 wl_223 vdd gnd cell_6t
Xbit_r224_c67 bl_67 br_67 wl_224 vdd gnd cell_6t
Xbit_r225_c67 bl_67 br_67 wl_225 vdd gnd cell_6t
Xbit_r226_c67 bl_67 br_67 wl_226 vdd gnd cell_6t
Xbit_r227_c67 bl_67 br_67 wl_227 vdd gnd cell_6t
Xbit_r228_c67 bl_67 br_67 wl_228 vdd gnd cell_6t
Xbit_r229_c67 bl_67 br_67 wl_229 vdd gnd cell_6t
Xbit_r230_c67 bl_67 br_67 wl_230 vdd gnd cell_6t
Xbit_r231_c67 bl_67 br_67 wl_231 vdd gnd cell_6t
Xbit_r232_c67 bl_67 br_67 wl_232 vdd gnd cell_6t
Xbit_r233_c67 bl_67 br_67 wl_233 vdd gnd cell_6t
Xbit_r234_c67 bl_67 br_67 wl_234 vdd gnd cell_6t
Xbit_r235_c67 bl_67 br_67 wl_235 vdd gnd cell_6t
Xbit_r236_c67 bl_67 br_67 wl_236 vdd gnd cell_6t
Xbit_r237_c67 bl_67 br_67 wl_237 vdd gnd cell_6t
Xbit_r238_c67 bl_67 br_67 wl_238 vdd gnd cell_6t
Xbit_r239_c67 bl_67 br_67 wl_239 vdd gnd cell_6t
Xbit_r240_c67 bl_67 br_67 wl_240 vdd gnd cell_6t
Xbit_r241_c67 bl_67 br_67 wl_241 vdd gnd cell_6t
Xbit_r242_c67 bl_67 br_67 wl_242 vdd gnd cell_6t
Xbit_r243_c67 bl_67 br_67 wl_243 vdd gnd cell_6t
Xbit_r244_c67 bl_67 br_67 wl_244 vdd gnd cell_6t
Xbit_r245_c67 bl_67 br_67 wl_245 vdd gnd cell_6t
Xbit_r246_c67 bl_67 br_67 wl_246 vdd gnd cell_6t
Xbit_r247_c67 bl_67 br_67 wl_247 vdd gnd cell_6t
Xbit_r248_c67 bl_67 br_67 wl_248 vdd gnd cell_6t
Xbit_r249_c67 bl_67 br_67 wl_249 vdd gnd cell_6t
Xbit_r250_c67 bl_67 br_67 wl_250 vdd gnd cell_6t
Xbit_r251_c67 bl_67 br_67 wl_251 vdd gnd cell_6t
Xbit_r252_c67 bl_67 br_67 wl_252 vdd gnd cell_6t
Xbit_r253_c67 bl_67 br_67 wl_253 vdd gnd cell_6t
Xbit_r254_c67 bl_67 br_67 wl_254 vdd gnd cell_6t
Xbit_r255_c67 bl_67 br_67 wl_255 vdd gnd cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd cell_6t
Xbit_r1_c68 bl_68 br_68 wl_1 vdd gnd cell_6t
Xbit_r2_c68 bl_68 br_68 wl_2 vdd gnd cell_6t
Xbit_r3_c68 bl_68 br_68 wl_3 vdd gnd cell_6t
Xbit_r4_c68 bl_68 br_68 wl_4 vdd gnd cell_6t
Xbit_r5_c68 bl_68 br_68 wl_5 vdd gnd cell_6t
Xbit_r6_c68 bl_68 br_68 wl_6 vdd gnd cell_6t
Xbit_r7_c68 bl_68 br_68 wl_7 vdd gnd cell_6t
Xbit_r8_c68 bl_68 br_68 wl_8 vdd gnd cell_6t
Xbit_r9_c68 bl_68 br_68 wl_9 vdd gnd cell_6t
Xbit_r10_c68 bl_68 br_68 wl_10 vdd gnd cell_6t
Xbit_r11_c68 bl_68 br_68 wl_11 vdd gnd cell_6t
Xbit_r12_c68 bl_68 br_68 wl_12 vdd gnd cell_6t
Xbit_r13_c68 bl_68 br_68 wl_13 vdd gnd cell_6t
Xbit_r14_c68 bl_68 br_68 wl_14 vdd gnd cell_6t
Xbit_r15_c68 bl_68 br_68 wl_15 vdd gnd cell_6t
Xbit_r16_c68 bl_68 br_68 wl_16 vdd gnd cell_6t
Xbit_r17_c68 bl_68 br_68 wl_17 vdd gnd cell_6t
Xbit_r18_c68 bl_68 br_68 wl_18 vdd gnd cell_6t
Xbit_r19_c68 bl_68 br_68 wl_19 vdd gnd cell_6t
Xbit_r20_c68 bl_68 br_68 wl_20 vdd gnd cell_6t
Xbit_r21_c68 bl_68 br_68 wl_21 vdd gnd cell_6t
Xbit_r22_c68 bl_68 br_68 wl_22 vdd gnd cell_6t
Xbit_r23_c68 bl_68 br_68 wl_23 vdd gnd cell_6t
Xbit_r24_c68 bl_68 br_68 wl_24 vdd gnd cell_6t
Xbit_r25_c68 bl_68 br_68 wl_25 vdd gnd cell_6t
Xbit_r26_c68 bl_68 br_68 wl_26 vdd gnd cell_6t
Xbit_r27_c68 bl_68 br_68 wl_27 vdd gnd cell_6t
Xbit_r28_c68 bl_68 br_68 wl_28 vdd gnd cell_6t
Xbit_r29_c68 bl_68 br_68 wl_29 vdd gnd cell_6t
Xbit_r30_c68 bl_68 br_68 wl_30 vdd gnd cell_6t
Xbit_r31_c68 bl_68 br_68 wl_31 vdd gnd cell_6t
Xbit_r32_c68 bl_68 br_68 wl_32 vdd gnd cell_6t
Xbit_r33_c68 bl_68 br_68 wl_33 vdd gnd cell_6t
Xbit_r34_c68 bl_68 br_68 wl_34 vdd gnd cell_6t
Xbit_r35_c68 bl_68 br_68 wl_35 vdd gnd cell_6t
Xbit_r36_c68 bl_68 br_68 wl_36 vdd gnd cell_6t
Xbit_r37_c68 bl_68 br_68 wl_37 vdd gnd cell_6t
Xbit_r38_c68 bl_68 br_68 wl_38 vdd gnd cell_6t
Xbit_r39_c68 bl_68 br_68 wl_39 vdd gnd cell_6t
Xbit_r40_c68 bl_68 br_68 wl_40 vdd gnd cell_6t
Xbit_r41_c68 bl_68 br_68 wl_41 vdd gnd cell_6t
Xbit_r42_c68 bl_68 br_68 wl_42 vdd gnd cell_6t
Xbit_r43_c68 bl_68 br_68 wl_43 vdd gnd cell_6t
Xbit_r44_c68 bl_68 br_68 wl_44 vdd gnd cell_6t
Xbit_r45_c68 bl_68 br_68 wl_45 vdd gnd cell_6t
Xbit_r46_c68 bl_68 br_68 wl_46 vdd gnd cell_6t
Xbit_r47_c68 bl_68 br_68 wl_47 vdd gnd cell_6t
Xbit_r48_c68 bl_68 br_68 wl_48 vdd gnd cell_6t
Xbit_r49_c68 bl_68 br_68 wl_49 vdd gnd cell_6t
Xbit_r50_c68 bl_68 br_68 wl_50 vdd gnd cell_6t
Xbit_r51_c68 bl_68 br_68 wl_51 vdd gnd cell_6t
Xbit_r52_c68 bl_68 br_68 wl_52 vdd gnd cell_6t
Xbit_r53_c68 bl_68 br_68 wl_53 vdd gnd cell_6t
Xbit_r54_c68 bl_68 br_68 wl_54 vdd gnd cell_6t
Xbit_r55_c68 bl_68 br_68 wl_55 vdd gnd cell_6t
Xbit_r56_c68 bl_68 br_68 wl_56 vdd gnd cell_6t
Xbit_r57_c68 bl_68 br_68 wl_57 vdd gnd cell_6t
Xbit_r58_c68 bl_68 br_68 wl_58 vdd gnd cell_6t
Xbit_r59_c68 bl_68 br_68 wl_59 vdd gnd cell_6t
Xbit_r60_c68 bl_68 br_68 wl_60 vdd gnd cell_6t
Xbit_r61_c68 bl_68 br_68 wl_61 vdd gnd cell_6t
Xbit_r62_c68 bl_68 br_68 wl_62 vdd gnd cell_6t
Xbit_r63_c68 bl_68 br_68 wl_63 vdd gnd cell_6t
Xbit_r64_c68 bl_68 br_68 wl_64 vdd gnd cell_6t
Xbit_r65_c68 bl_68 br_68 wl_65 vdd gnd cell_6t
Xbit_r66_c68 bl_68 br_68 wl_66 vdd gnd cell_6t
Xbit_r67_c68 bl_68 br_68 wl_67 vdd gnd cell_6t
Xbit_r68_c68 bl_68 br_68 wl_68 vdd gnd cell_6t
Xbit_r69_c68 bl_68 br_68 wl_69 vdd gnd cell_6t
Xbit_r70_c68 bl_68 br_68 wl_70 vdd gnd cell_6t
Xbit_r71_c68 bl_68 br_68 wl_71 vdd gnd cell_6t
Xbit_r72_c68 bl_68 br_68 wl_72 vdd gnd cell_6t
Xbit_r73_c68 bl_68 br_68 wl_73 vdd gnd cell_6t
Xbit_r74_c68 bl_68 br_68 wl_74 vdd gnd cell_6t
Xbit_r75_c68 bl_68 br_68 wl_75 vdd gnd cell_6t
Xbit_r76_c68 bl_68 br_68 wl_76 vdd gnd cell_6t
Xbit_r77_c68 bl_68 br_68 wl_77 vdd gnd cell_6t
Xbit_r78_c68 bl_68 br_68 wl_78 vdd gnd cell_6t
Xbit_r79_c68 bl_68 br_68 wl_79 vdd gnd cell_6t
Xbit_r80_c68 bl_68 br_68 wl_80 vdd gnd cell_6t
Xbit_r81_c68 bl_68 br_68 wl_81 vdd gnd cell_6t
Xbit_r82_c68 bl_68 br_68 wl_82 vdd gnd cell_6t
Xbit_r83_c68 bl_68 br_68 wl_83 vdd gnd cell_6t
Xbit_r84_c68 bl_68 br_68 wl_84 vdd gnd cell_6t
Xbit_r85_c68 bl_68 br_68 wl_85 vdd gnd cell_6t
Xbit_r86_c68 bl_68 br_68 wl_86 vdd gnd cell_6t
Xbit_r87_c68 bl_68 br_68 wl_87 vdd gnd cell_6t
Xbit_r88_c68 bl_68 br_68 wl_88 vdd gnd cell_6t
Xbit_r89_c68 bl_68 br_68 wl_89 vdd gnd cell_6t
Xbit_r90_c68 bl_68 br_68 wl_90 vdd gnd cell_6t
Xbit_r91_c68 bl_68 br_68 wl_91 vdd gnd cell_6t
Xbit_r92_c68 bl_68 br_68 wl_92 vdd gnd cell_6t
Xbit_r93_c68 bl_68 br_68 wl_93 vdd gnd cell_6t
Xbit_r94_c68 bl_68 br_68 wl_94 vdd gnd cell_6t
Xbit_r95_c68 bl_68 br_68 wl_95 vdd gnd cell_6t
Xbit_r96_c68 bl_68 br_68 wl_96 vdd gnd cell_6t
Xbit_r97_c68 bl_68 br_68 wl_97 vdd gnd cell_6t
Xbit_r98_c68 bl_68 br_68 wl_98 vdd gnd cell_6t
Xbit_r99_c68 bl_68 br_68 wl_99 vdd gnd cell_6t
Xbit_r100_c68 bl_68 br_68 wl_100 vdd gnd cell_6t
Xbit_r101_c68 bl_68 br_68 wl_101 vdd gnd cell_6t
Xbit_r102_c68 bl_68 br_68 wl_102 vdd gnd cell_6t
Xbit_r103_c68 bl_68 br_68 wl_103 vdd gnd cell_6t
Xbit_r104_c68 bl_68 br_68 wl_104 vdd gnd cell_6t
Xbit_r105_c68 bl_68 br_68 wl_105 vdd gnd cell_6t
Xbit_r106_c68 bl_68 br_68 wl_106 vdd gnd cell_6t
Xbit_r107_c68 bl_68 br_68 wl_107 vdd gnd cell_6t
Xbit_r108_c68 bl_68 br_68 wl_108 vdd gnd cell_6t
Xbit_r109_c68 bl_68 br_68 wl_109 vdd gnd cell_6t
Xbit_r110_c68 bl_68 br_68 wl_110 vdd gnd cell_6t
Xbit_r111_c68 bl_68 br_68 wl_111 vdd gnd cell_6t
Xbit_r112_c68 bl_68 br_68 wl_112 vdd gnd cell_6t
Xbit_r113_c68 bl_68 br_68 wl_113 vdd gnd cell_6t
Xbit_r114_c68 bl_68 br_68 wl_114 vdd gnd cell_6t
Xbit_r115_c68 bl_68 br_68 wl_115 vdd gnd cell_6t
Xbit_r116_c68 bl_68 br_68 wl_116 vdd gnd cell_6t
Xbit_r117_c68 bl_68 br_68 wl_117 vdd gnd cell_6t
Xbit_r118_c68 bl_68 br_68 wl_118 vdd gnd cell_6t
Xbit_r119_c68 bl_68 br_68 wl_119 vdd gnd cell_6t
Xbit_r120_c68 bl_68 br_68 wl_120 vdd gnd cell_6t
Xbit_r121_c68 bl_68 br_68 wl_121 vdd gnd cell_6t
Xbit_r122_c68 bl_68 br_68 wl_122 vdd gnd cell_6t
Xbit_r123_c68 bl_68 br_68 wl_123 vdd gnd cell_6t
Xbit_r124_c68 bl_68 br_68 wl_124 vdd gnd cell_6t
Xbit_r125_c68 bl_68 br_68 wl_125 vdd gnd cell_6t
Xbit_r126_c68 bl_68 br_68 wl_126 vdd gnd cell_6t
Xbit_r127_c68 bl_68 br_68 wl_127 vdd gnd cell_6t
Xbit_r128_c68 bl_68 br_68 wl_128 vdd gnd cell_6t
Xbit_r129_c68 bl_68 br_68 wl_129 vdd gnd cell_6t
Xbit_r130_c68 bl_68 br_68 wl_130 vdd gnd cell_6t
Xbit_r131_c68 bl_68 br_68 wl_131 vdd gnd cell_6t
Xbit_r132_c68 bl_68 br_68 wl_132 vdd gnd cell_6t
Xbit_r133_c68 bl_68 br_68 wl_133 vdd gnd cell_6t
Xbit_r134_c68 bl_68 br_68 wl_134 vdd gnd cell_6t
Xbit_r135_c68 bl_68 br_68 wl_135 vdd gnd cell_6t
Xbit_r136_c68 bl_68 br_68 wl_136 vdd gnd cell_6t
Xbit_r137_c68 bl_68 br_68 wl_137 vdd gnd cell_6t
Xbit_r138_c68 bl_68 br_68 wl_138 vdd gnd cell_6t
Xbit_r139_c68 bl_68 br_68 wl_139 vdd gnd cell_6t
Xbit_r140_c68 bl_68 br_68 wl_140 vdd gnd cell_6t
Xbit_r141_c68 bl_68 br_68 wl_141 vdd gnd cell_6t
Xbit_r142_c68 bl_68 br_68 wl_142 vdd gnd cell_6t
Xbit_r143_c68 bl_68 br_68 wl_143 vdd gnd cell_6t
Xbit_r144_c68 bl_68 br_68 wl_144 vdd gnd cell_6t
Xbit_r145_c68 bl_68 br_68 wl_145 vdd gnd cell_6t
Xbit_r146_c68 bl_68 br_68 wl_146 vdd gnd cell_6t
Xbit_r147_c68 bl_68 br_68 wl_147 vdd gnd cell_6t
Xbit_r148_c68 bl_68 br_68 wl_148 vdd gnd cell_6t
Xbit_r149_c68 bl_68 br_68 wl_149 vdd gnd cell_6t
Xbit_r150_c68 bl_68 br_68 wl_150 vdd gnd cell_6t
Xbit_r151_c68 bl_68 br_68 wl_151 vdd gnd cell_6t
Xbit_r152_c68 bl_68 br_68 wl_152 vdd gnd cell_6t
Xbit_r153_c68 bl_68 br_68 wl_153 vdd gnd cell_6t
Xbit_r154_c68 bl_68 br_68 wl_154 vdd gnd cell_6t
Xbit_r155_c68 bl_68 br_68 wl_155 vdd gnd cell_6t
Xbit_r156_c68 bl_68 br_68 wl_156 vdd gnd cell_6t
Xbit_r157_c68 bl_68 br_68 wl_157 vdd gnd cell_6t
Xbit_r158_c68 bl_68 br_68 wl_158 vdd gnd cell_6t
Xbit_r159_c68 bl_68 br_68 wl_159 vdd gnd cell_6t
Xbit_r160_c68 bl_68 br_68 wl_160 vdd gnd cell_6t
Xbit_r161_c68 bl_68 br_68 wl_161 vdd gnd cell_6t
Xbit_r162_c68 bl_68 br_68 wl_162 vdd gnd cell_6t
Xbit_r163_c68 bl_68 br_68 wl_163 vdd gnd cell_6t
Xbit_r164_c68 bl_68 br_68 wl_164 vdd gnd cell_6t
Xbit_r165_c68 bl_68 br_68 wl_165 vdd gnd cell_6t
Xbit_r166_c68 bl_68 br_68 wl_166 vdd gnd cell_6t
Xbit_r167_c68 bl_68 br_68 wl_167 vdd gnd cell_6t
Xbit_r168_c68 bl_68 br_68 wl_168 vdd gnd cell_6t
Xbit_r169_c68 bl_68 br_68 wl_169 vdd gnd cell_6t
Xbit_r170_c68 bl_68 br_68 wl_170 vdd gnd cell_6t
Xbit_r171_c68 bl_68 br_68 wl_171 vdd gnd cell_6t
Xbit_r172_c68 bl_68 br_68 wl_172 vdd gnd cell_6t
Xbit_r173_c68 bl_68 br_68 wl_173 vdd gnd cell_6t
Xbit_r174_c68 bl_68 br_68 wl_174 vdd gnd cell_6t
Xbit_r175_c68 bl_68 br_68 wl_175 vdd gnd cell_6t
Xbit_r176_c68 bl_68 br_68 wl_176 vdd gnd cell_6t
Xbit_r177_c68 bl_68 br_68 wl_177 vdd gnd cell_6t
Xbit_r178_c68 bl_68 br_68 wl_178 vdd gnd cell_6t
Xbit_r179_c68 bl_68 br_68 wl_179 vdd gnd cell_6t
Xbit_r180_c68 bl_68 br_68 wl_180 vdd gnd cell_6t
Xbit_r181_c68 bl_68 br_68 wl_181 vdd gnd cell_6t
Xbit_r182_c68 bl_68 br_68 wl_182 vdd gnd cell_6t
Xbit_r183_c68 bl_68 br_68 wl_183 vdd gnd cell_6t
Xbit_r184_c68 bl_68 br_68 wl_184 vdd gnd cell_6t
Xbit_r185_c68 bl_68 br_68 wl_185 vdd gnd cell_6t
Xbit_r186_c68 bl_68 br_68 wl_186 vdd gnd cell_6t
Xbit_r187_c68 bl_68 br_68 wl_187 vdd gnd cell_6t
Xbit_r188_c68 bl_68 br_68 wl_188 vdd gnd cell_6t
Xbit_r189_c68 bl_68 br_68 wl_189 vdd gnd cell_6t
Xbit_r190_c68 bl_68 br_68 wl_190 vdd gnd cell_6t
Xbit_r191_c68 bl_68 br_68 wl_191 vdd gnd cell_6t
Xbit_r192_c68 bl_68 br_68 wl_192 vdd gnd cell_6t
Xbit_r193_c68 bl_68 br_68 wl_193 vdd gnd cell_6t
Xbit_r194_c68 bl_68 br_68 wl_194 vdd gnd cell_6t
Xbit_r195_c68 bl_68 br_68 wl_195 vdd gnd cell_6t
Xbit_r196_c68 bl_68 br_68 wl_196 vdd gnd cell_6t
Xbit_r197_c68 bl_68 br_68 wl_197 vdd gnd cell_6t
Xbit_r198_c68 bl_68 br_68 wl_198 vdd gnd cell_6t
Xbit_r199_c68 bl_68 br_68 wl_199 vdd gnd cell_6t
Xbit_r200_c68 bl_68 br_68 wl_200 vdd gnd cell_6t
Xbit_r201_c68 bl_68 br_68 wl_201 vdd gnd cell_6t
Xbit_r202_c68 bl_68 br_68 wl_202 vdd gnd cell_6t
Xbit_r203_c68 bl_68 br_68 wl_203 vdd gnd cell_6t
Xbit_r204_c68 bl_68 br_68 wl_204 vdd gnd cell_6t
Xbit_r205_c68 bl_68 br_68 wl_205 vdd gnd cell_6t
Xbit_r206_c68 bl_68 br_68 wl_206 vdd gnd cell_6t
Xbit_r207_c68 bl_68 br_68 wl_207 vdd gnd cell_6t
Xbit_r208_c68 bl_68 br_68 wl_208 vdd gnd cell_6t
Xbit_r209_c68 bl_68 br_68 wl_209 vdd gnd cell_6t
Xbit_r210_c68 bl_68 br_68 wl_210 vdd gnd cell_6t
Xbit_r211_c68 bl_68 br_68 wl_211 vdd gnd cell_6t
Xbit_r212_c68 bl_68 br_68 wl_212 vdd gnd cell_6t
Xbit_r213_c68 bl_68 br_68 wl_213 vdd gnd cell_6t
Xbit_r214_c68 bl_68 br_68 wl_214 vdd gnd cell_6t
Xbit_r215_c68 bl_68 br_68 wl_215 vdd gnd cell_6t
Xbit_r216_c68 bl_68 br_68 wl_216 vdd gnd cell_6t
Xbit_r217_c68 bl_68 br_68 wl_217 vdd gnd cell_6t
Xbit_r218_c68 bl_68 br_68 wl_218 vdd gnd cell_6t
Xbit_r219_c68 bl_68 br_68 wl_219 vdd gnd cell_6t
Xbit_r220_c68 bl_68 br_68 wl_220 vdd gnd cell_6t
Xbit_r221_c68 bl_68 br_68 wl_221 vdd gnd cell_6t
Xbit_r222_c68 bl_68 br_68 wl_222 vdd gnd cell_6t
Xbit_r223_c68 bl_68 br_68 wl_223 vdd gnd cell_6t
Xbit_r224_c68 bl_68 br_68 wl_224 vdd gnd cell_6t
Xbit_r225_c68 bl_68 br_68 wl_225 vdd gnd cell_6t
Xbit_r226_c68 bl_68 br_68 wl_226 vdd gnd cell_6t
Xbit_r227_c68 bl_68 br_68 wl_227 vdd gnd cell_6t
Xbit_r228_c68 bl_68 br_68 wl_228 vdd gnd cell_6t
Xbit_r229_c68 bl_68 br_68 wl_229 vdd gnd cell_6t
Xbit_r230_c68 bl_68 br_68 wl_230 vdd gnd cell_6t
Xbit_r231_c68 bl_68 br_68 wl_231 vdd gnd cell_6t
Xbit_r232_c68 bl_68 br_68 wl_232 vdd gnd cell_6t
Xbit_r233_c68 bl_68 br_68 wl_233 vdd gnd cell_6t
Xbit_r234_c68 bl_68 br_68 wl_234 vdd gnd cell_6t
Xbit_r235_c68 bl_68 br_68 wl_235 vdd gnd cell_6t
Xbit_r236_c68 bl_68 br_68 wl_236 vdd gnd cell_6t
Xbit_r237_c68 bl_68 br_68 wl_237 vdd gnd cell_6t
Xbit_r238_c68 bl_68 br_68 wl_238 vdd gnd cell_6t
Xbit_r239_c68 bl_68 br_68 wl_239 vdd gnd cell_6t
Xbit_r240_c68 bl_68 br_68 wl_240 vdd gnd cell_6t
Xbit_r241_c68 bl_68 br_68 wl_241 vdd gnd cell_6t
Xbit_r242_c68 bl_68 br_68 wl_242 vdd gnd cell_6t
Xbit_r243_c68 bl_68 br_68 wl_243 vdd gnd cell_6t
Xbit_r244_c68 bl_68 br_68 wl_244 vdd gnd cell_6t
Xbit_r245_c68 bl_68 br_68 wl_245 vdd gnd cell_6t
Xbit_r246_c68 bl_68 br_68 wl_246 vdd gnd cell_6t
Xbit_r247_c68 bl_68 br_68 wl_247 vdd gnd cell_6t
Xbit_r248_c68 bl_68 br_68 wl_248 vdd gnd cell_6t
Xbit_r249_c68 bl_68 br_68 wl_249 vdd gnd cell_6t
Xbit_r250_c68 bl_68 br_68 wl_250 vdd gnd cell_6t
Xbit_r251_c68 bl_68 br_68 wl_251 vdd gnd cell_6t
Xbit_r252_c68 bl_68 br_68 wl_252 vdd gnd cell_6t
Xbit_r253_c68 bl_68 br_68 wl_253 vdd gnd cell_6t
Xbit_r254_c68 bl_68 br_68 wl_254 vdd gnd cell_6t
Xbit_r255_c68 bl_68 br_68 wl_255 vdd gnd cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd cell_6t
Xbit_r1_c69 bl_69 br_69 wl_1 vdd gnd cell_6t
Xbit_r2_c69 bl_69 br_69 wl_2 vdd gnd cell_6t
Xbit_r3_c69 bl_69 br_69 wl_3 vdd gnd cell_6t
Xbit_r4_c69 bl_69 br_69 wl_4 vdd gnd cell_6t
Xbit_r5_c69 bl_69 br_69 wl_5 vdd gnd cell_6t
Xbit_r6_c69 bl_69 br_69 wl_6 vdd gnd cell_6t
Xbit_r7_c69 bl_69 br_69 wl_7 vdd gnd cell_6t
Xbit_r8_c69 bl_69 br_69 wl_8 vdd gnd cell_6t
Xbit_r9_c69 bl_69 br_69 wl_9 vdd gnd cell_6t
Xbit_r10_c69 bl_69 br_69 wl_10 vdd gnd cell_6t
Xbit_r11_c69 bl_69 br_69 wl_11 vdd gnd cell_6t
Xbit_r12_c69 bl_69 br_69 wl_12 vdd gnd cell_6t
Xbit_r13_c69 bl_69 br_69 wl_13 vdd gnd cell_6t
Xbit_r14_c69 bl_69 br_69 wl_14 vdd gnd cell_6t
Xbit_r15_c69 bl_69 br_69 wl_15 vdd gnd cell_6t
Xbit_r16_c69 bl_69 br_69 wl_16 vdd gnd cell_6t
Xbit_r17_c69 bl_69 br_69 wl_17 vdd gnd cell_6t
Xbit_r18_c69 bl_69 br_69 wl_18 vdd gnd cell_6t
Xbit_r19_c69 bl_69 br_69 wl_19 vdd gnd cell_6t
Xbit_r20_c69 bl_69 br_69 wl_20 vdd gnd cell_6t
Xbit_r21_c69 bl_69 br_69 wl_21 vdd gnd cell_6t
Xbit_r22_c69 bl_69 br_69 wl_22 vdd gnd cell_6t
Xbit_r23_c69 bl_69 br_69 wl_23 vdd gnd cell_6t
Xbit_r24_c69 bl_69 br_69 wl_24 vdd gnd cell_6t
Xbit_r25_c69 bl_69 br_69 wl_25 vdd gnd cell_6t
Xbit_r26_c69 bl_69 br_69 wl_26 vdd gnd cell_6t
Xbit_r27_c69 bl_69 br_69 wl_27 vdd gnd cell_6t
Xbit_r28_c69 bl_69 br_69 wl_28 vdd gnd cell_6t
Xbit_r29_c69 bl_69 br_69 wl_29 vdd gnd cell_6t
Xbit_r30_c69 bl_69 br_69 wl_30 vdd gnd cell_6t
Xbit_r31_c69 bl_69 br_69 wl_31 vdd gnd cell_6t
Xbit_r32_c69 bl_69 br_69 wl_32 vdd gnd cell_6t
Xbit_r33_c69 bl_69 br_69 wl_33 vdd gnd cell_6t
Xbit_r34_c69 bl_69 br_69 wl_34 vdd gnd cell_6t
Xbit_r35_c69 bl_69 br_69 wl_35 vdd gnd cell_6t
Xbit_r36_c69 bl_69 br_69 wl_36 vdd gnd cell_6t
Xbit_r37_c69 bl_69 br_69 wl_37 vdd gnd cell_6t
Xbit_r38_c69 bl_69 br_69 wl_38 vdd gnd cell_6t
Xbit_r39_c69 bl_69 br_69 wl_39 vdd gnd cell_6t
Xbit_r40_c69 bl_69 br_69 wl_40 vdd gnd cell_6t
Xbit_r41_c69 bl_69 br_69 wl_41 vdd gnd cell_6t
Xbit_r42_c69 bl_69 br_69 wl_42 vdd gnd cell_6t
Xbit_r43_c69 bl_69 br_69 wl_43 vdd gnd cell_6t
Xbit_r44_c69 bl_69 br_69 wl_44 vdd gnd cell_6t
Xbit_r45_c69 bl_69 br_69 wl_45 vdd gnd cell_6t
Xbit_r46_c69 bl_69 br_69 wl_46 vdd gnd cell_6t
Xbit_r47_c69 bl_69 br_69 wl_47 vdd gnd cell_6t
Xbit_r48_c69 bl_69 br_69 wl_48 vdd gnd cell_6t
Xbit_r49_c69 bl_69 br_69 wl_49 vdd gnd cell_6t
Xbit_r50_c69 bl_69 br_69 wl_50 vdd gnd cell_6t
Xbit_r51_c69 bl_69 br_69 wl_51 vdd gnd cell_6t
Xbit_r52_c69 bl_69 br_69 wl_52 vdd gnd cell_6t
Xbit_r53_c69 bl_69 br_69 wl_53 vdd gnd cell_6t
Xbit_r54_c69 bl_69 br_69 wl_54 vdd gnd cell_6t
Xbit_r55_c69 bl_69 br_69 wl_55 vdd gnd cell_6t
Xbit_r56_c69 bl_69 br_69 wl_56 vdd gnd cell_6t
Xbit_r57_c69 bl_69 br_69 wl_57 vdd gnd cell_6t
Xbit_r58_c69 bl_69 br_69 wl_58 vdd gnd cell_6t
Xbit_r59_c69 bl_69 br_69 wl_59 vdd gnd cell_6t
Xbit_r60_c69 bl_69 br_69 wl_60 vdd gnd cell_6t
Xbit_r61_c69 bl_69 br_69 wl_61 vdd gnd cell_6t
Xbit_r62_c69 bl_69 br_69 wl_62 vdd gnd cell_6t
Xbit_r63_c69 bl_69 br_69 wl_63 vdd gnd cell_6t
Xbit_r64_c69 bl_69 br_69 wl_64 vdd gnd cell_6t
Xbit_r65_c69 bl_69 br_69 wl_65 vdd gnd cell_6t
Xbit_r66_c69 bl_69 br_69 wl_66 vdd gnd cell_6t
Xbit_r67_c69 bl_69 br_69 wl_67 vdd gnd cell_6t
Xbit_r68_c69 bl_69 br_69 wl_68 vdd gnd cell_6t
Xbit_r69_c69 bl_69 br_69 wl_69 vdd gnd cell_6t
Xbit_r70_c69 bl_69 br_69 wl_70 vdd gnd cell_6t
Xbit_r71_c69 bl_69 br_69 wl_71 vdd gnd cell_6t
Xbit_r72_c69 bl_69 br_69 wl_72 vdd gnd cell_6t
Xbit_r73_c69 bl_69 br_69 wl_73 vdd gnd cell_6t
Xbit_r74_c69 bl_69 br_69 wl_74 vdd gnd cell_6t
Xbit_r75_c69 bl_69 br_69 wl_75 vdd gnd cell_6t
Xbit_r76_c69 bl_69 br_69 wl_76 vdd gnd cell_6t
Xbit_r77_c69 bl_69 br_69 wl_77 vdd gnd cell_6t
Xbit_r78_c69 bl_69 br_69 wl_78 vdd gnd cell_6t
Xbit_r79_c69 bl_69 br_69 wl_79 vdd gnd cell_6t
Xbit_r80_c69 bl_69 br_69 wl_80 vdd gnd cell_6t
Xbit_r81_c69 bl_69 br_69 wl_81 vdd gnd cell_6t
Xbit_r82_c69 bl_69 br_69 wl_82 vdd gnd cell_6t
Xbit_r83_c69 bl_69 br_69 wl_83 vdd gnd cell_6t
Xbit_r84_c69 bl_69 br_69 wl_84 vdd gnd cell_6t
Xbit_r85_c69 bl_69 br_69 wl_85 vdd gnd cell_6t
Xbit_r86_c69 bl_69 br_69 wl_86 vdd gnd cell_6t
Xbit_r87_c69 bl_69 br_69 wl_87 vdd gnd cell_6t
Xbit_r88_c69 bl_69 br_69 wl_88 vdd gnd cell_6t
Xbit_r89_c69 bl_69 br_69 wl_89 vdd gnd cell_6t
Xbit_r90_c69 bl_69 br_69 wl_90 vdd gnd cell_6t
Xbit_r91_c69 bl_69 br_69 wl_91 vdd gnd cell_6t
Xbit_r92_c69 bl_69 br_69 wl_92 vdd gnd cell_6t
Xbit_r93_c69 bl_69 br_69 wl_93 vdd gnd cell_6t
Xbit_r94_c69 bl_69 br_69 wl_94 vdd gnd cell_6t
Xbit_r95_c69 bl_69 br_69 wl_95 vdd gnd cell_6t
Xbit_r96_c69 bl_69 br_69 wl_96 vdd gnd cell_6t
Xbit_r97_c69 bl_69 br_69 wl_97 vdd gnd cell_6t
Xbit_r98_c69 bl_69 br_69 wl_98 vdd gnd cell_6t
Xbit_r99_c69 bl_69 br_69 wl_99 vdd gnd cell_6t
Xbit_r100_c69 bl_69 br_69 wl_100 vdd gnd cell_6t
Xbit_r101_c69 bl_69 br_69 wl_101 vdd gnd cell_6t
Xbit_r102_c69 bl_69 br_69 wl_102 vdd gnd cell_6t
Xbit_r103_c69 bl_69 br_69 wl_103 vdd gnd cell_6t
Xbit_r104_c69 bl_69 br_69 wl_104 vdd gnd cell_6t
Xbit_r105_c69 bl_69 br_69 wl_105 vdd gnd cell_6t
Xbit_r106_c69 bl_69 br_69 wl_106 vdd gnd cell_6t
Xbit_r107_c69 bl_69 br_69 wl_107 vdd gnd cell_6t
Xbit_r108_c69 bl_69 br_69 wl_108 vdd gnd cell_6t
Xbit_r109_c69 bl_69 br_69 wl_109 vdd gnd cell_6t
Xbit_r110_c69 bl_69 br_69 wl_110 vdd gnd cell_6t
Xbit_r111_c69 bl_69 br_69 wl_111 vdd gnd cell_6t
Xbit_r112_c69 bl_69 br_69 wl_112 vdd gnd cell_6t
Xbit_r113_c69 bl_69 br_69 wl_113 vdd gnd cell_6t
Xbit_r114_c69 bl_69 br_69 wl_114 vdd gnd cell_6t
Xbit_r115_c69 bl_69 br_69 wl_115 vdd gnd cell_6t
Xbit_r116_c69 bl_69 br_69 wl_116 vdd gnd cell_6t
Xbit_r117_c69 bl_69 br_69 wl_117 vdd gnd cell_6t
Xbit_r118_c69 bl_69 br_69 wl_118 vdd gnd cell_6t
Xbit_r119_c69 bl_69 br_69 wl_119 vdd gnd cell_6t
Xbit_r120_c69 bl_69 br_69 wl_120 vdd gnd cell_6t
Xbit_r121_c69 bl_69 br_69 wl_121 vdd gnd cell_6t
Xbit_r122_c69 bl_69 br_69 wl_122 vdd gnd cell_6t
Xbit_r123_c69 bl_69 br_69 wl_123 vdd gnd cell_6t
Xbit_r124_c69 bl_69 br_69 wl_124 vdd gnd cell_6t
Xbit_r125_c69 bl_69 br_69 wl_125 vdd gnd cell_6t
Xbit_r126_c69 bl_69 br_69 wl_126 vdd gnd cell_6t
Xbit_r127_c69 bl_69 br_69 wl_127 vdd gnd cell_6t
Xbit_r128_c69 bl_69 br_69 wl_128 vdd gnd cell_6t
Xbit_r129_c69 bl_69 br_69 wl_129 vdd gnd cell_6t
Xbit_r130_c69 bl_69 br_69 wl_130 vdd gnd cell_6t
Xbit_r131_c69 bl_69 br_69 wl_131 vdd gnd cell_6t
Xbit_r132_c69 bl_69 br_69 wl_132 vdd gnd cell_6t
Xbit_r133_c69 bl_69 br_69 wl_133 vdd gnd cell_6t
Xbit_r134_c69 bl_69 br_69 wl_134 vdd gnd cell_6t
Xbit_r135_c69 bl_69 br_69 wl_135 vdd gnd cell_6t
Xbit_r136_c69 bl_69 br_69 wl_136 vdd gnd cell_6t
Xbit_r137_c69 bl_69 br_69 wl_137 vdd gnd cell_6t
Xbit_r138_c69 bl_69 br_69 wl_138 vdd gnd cell_6t
Xbit_r139_c69 bl_69 br_69 wl_139 vdd gnd cell_6t
Xbit_r140_c69 bl_69 br_69 wl_140 vdd gnd cell_6t
Xbit_r141_c69 bl_69 br_69 wl_141 vdd gnd cell_6t
Xbit_r142_c69 bl_69 br_69 wl_142 vdd gnd cell_6t
Xbit_r143_c69 bl_69 br_69 wl_143 vdd gnd cell_6t
Xbit_r144_c69 bl_69 br_69 wl_144 vdd gnd cell_6t
Xbit_r145_c69 bl_69 br_69 wl_145 vdd gnd cell_6t
Xbit_r146_c69 bl_69 br_69 wl_146 vdd gnd cell_6t
Xbit_r147_c69 bl_69 br_69 wl_147 vdd gnd cell_6t
Xbit_r148_c69 bl_69 br_69 wl_148 vdd gnd cell_6t
Xbit_r149_c69 bl_69 br_69 wl_149 vdd gnd cell_6t
Xbit_r150_c69 bl_69 br_69 wl_150 vdd gnd cell_6t
Xbit_r151_c69 bl_69 br_69 wl_151 vdd gnd cell_6t
Xbit_r152_c69 bl_69 br_69 wl_152 vdd gnd cell_6t
Xbit_r153_c69 bl_69 br_69 wl_153 vdd gnd cell_6t
Xbit_r154_c69 bl_69 br_69 wl_154 vdd gnd cell_6t
Xbit_r155_c69 bl_69 br_69 wl_155 vdd gnd cell_6t
Xbit_r156_c69 bl_69 br_69 wl_156 vdd gnd cell_6t
Xbit_r157_c69 bl_69 br_69 wl_157 vdd gnd cell_6t
Xbit_r158_c69 bl_69 br_69 wl_158 vdd gnd cell_6t
Xbit_r159_c69 bl_69 br_69 wl_159 vdd gnd cell_6t
Xbit_r160_c69 bl_69 br_69 wl_160 vdd gnd cell_6t
Xbit_r161_c69 bl_69 br_69 wl_161 vdd gnd cell_6t
Xbit_r162_c69 bl_69 br_69 wl_162 vdd gnd cell_6t
Xbit_r163_c69 bl_69 br_69 wl_163 vdd gnd cell_6t
Xbit_r164_c69 bl_69 br_69 wl_164 vdd gnd cell_6t
Xbit_r165_c69 bl_69 br_69 wl_165 vdd gnd cell_6t
Xbit_r166_c69 bl_69 br_69 wl_166 vdd gnd cell_6t
Xbit_r167_c69 bl_69 br_69 wl_167 vdd gnd cell_6t
Xbit_r168_c69 bl_69 br_69 wl_168 vdd gnd cell_6t
Xbit_r169_c69 bl_69 br_69 wl_169 vdd gnd cell_6t
Xbit_r170_c69 bl_69 br_69 wl_170 vdd gnd cell_6t
Xbit_r171_c69 bl_69 br_69 wl_171 vdd gnd cell_6t
Xbit_r172_c69 bl_69 br_69 wl_172 vdd gnd cell_6t
Xbit_r173_c69 bl_69 br_69 wl_173 vdd gnd cell_6t
Xbit_r174_c69 bl_69 br_69 wl_174 vdd gnd cell_6t
Xbit_r175_c69 bl_69 br_69 wl_175 vdd gnd cell_6t
Xbit_r176_c69 bl_69 br_69 wl_176 vdd gnd cell_6t
Xbit_r177_c69 bl_69 br_69 wl_177 vdd gnd cell_6t
Xbit_r178_c69 bl_69 br_69 wl_178 vdd gnd cell_6t
Xbit_r179_c69 bl_69 br_69 wl_179 vdd gnd cell_6t
Xbit_r180_c69 bl_69 br_69 wl_180 vdd gnd cell_6t
Xbit_r181_c69 bl_69 br_69 wl_181 vdd gnd cell_6t
Xbit_r182_c69 bl_69 br_69 wl_182 vdd gnd cell_6t
Xbit_r183_c69 bl_69 br_69 wl_183 vdd gnd cell_6t
Xbit_r184_c69 bl_69 br_69 wl_184 vdd gnd cell_6t
Xbit_r185_c69 bl_69 br_69 wl_185 vdd gnd cell_6t
Xbit_r186_c69 bl_69 br_69 wl_186 vdd gnd cell_6t
Xbit_r187_c69 bl_69 br_69 wl_187 vdd gnd cell_6t
Xbit_r188_c69 bl_69 br_69 wl_188 vdd gnd cell_6t
Xbit_r189_c69 bl_69 br_69 wl_189 vdd gnd cell_6t
Xbit_r190_c69 bl_69 br_69 wl_190 vdd gnd cell_6t
Xbit_r191_c69 bl_69 br_69 wl_191 vdd gnd cell_6t
Xbit_r192_c69 bl_69 br_69 wl_192 vdd gnd cell_6t
Xbit_r193_c69 bl_69 br_69 wl_193 vdd gnd cell_6t
Xbit_r194_c69 bl_69 br_69 wl_194 vdd gnd cell_6t
Xbit_r195_c69 bl_69 br_69 wl_195 vdd gnd cell_6t
Xbit_r196_c69 bl_69 br_69 wl_196 vdd gnd cell_6t
Xbit_r197_c69 bl_69 br_69 wl_197 vdd gnd cell_6t
Xbit_r198_c69 bl_69 br_69 wl_198 vdd gnd cell_6t
Xbit_r199_c69 bl_69 br_69 wl_199 vdd gnd cell_6t
Xbit_r200_c69 bl_69 br_69 wl_200 vdd gnd cell_6t
Xbit_r201_c69 bl_69 br_69 wl_201 vdd gnd cell_6t
Xbit_r202_c69 bl_69 br_69 wl_202 vdd gnd cell_6t
Xbit_r203_c69 bl_69 br_69 wl_203 vdd gnd cell_6t
Xbit_r204_c69 bl_69 br_69 wl_204 vdd gnd cell_6t
Xbit_r205_c69 bl_69 br_69 wl_205 vdd gnd cell_6t
Xbit_r206_c69 bl_69 br_69 wl_206 vdd gnd cell_6t
Xbit_r207_c69 bl_69 br_69 wl_207 vdd gnd cell_6t
Xbit_r208_c69 bl_69 br_69 wl_208 vdd gnd cell_6t
Xbit_r209_c69 bl_69 br_69 wl_209 vdd gnd cell_6t
Xbit_r210_c69 bl_69 br_69 wl_210 vdd gnd cell_6t
Xbit_r211_c69 bl_69 br_69 wl_211 vdd gnd cell_6t
Xbit_r212_c69 bl_69 br_69 wl_212 vdd gnd cell_6t
Xbit_r213_c69 bl_69 br_69 wl_213 vdd gnd cell_6t
Xbit_r214_c69 bl_69 br_69 wl_214 vdd gnd cell_6t
Xbit_r215_c69 bl_69 br_69 wl_215 vdd gnd cell_6t
Xbit_r216_c69 bl_69 br_69 wl_216 vdd gnd cell_6t
Xbit_r217_c69 bl_69 br_69 wl_217 vdd gnd cell_6t
Xbit_r218_c69 bl_69 br_69 wl_218 vdd gnd cell_6t
Xbit_r219_c69 bl_69 br_69 wl_219 vdd gnd cell_6t
Xbit_r220_c69 bl_69 br_69 wl_220 vdd gnd cell_6t
Xbit_r221_c69 bl_69 br_69 wl_221 vdd gnd cell_6t
Xbit_r222_c69 bl_69 br_69 wl_222 vdd gnd cell_6t
Xbit_r223_c69 bl_69 br_69 wl_223 vdd gnd cell_6t
Xbit_r224_c69 bl_69 br_69 wl_224 vdd gnd cell_6t
Xbit_r225_c69 bl_69 br_69 wl_225 vdd gnd cell_6t
Xbit_r226_c69 bl_69 br_69 wl_226 vdd gnd cell_6t
Xbit_r227_c69 bl_69 br_69 wl_227 vdd gnd cell_6t
Xbit_r228_c69 bl_69 br_69 wl_228 vdd gnd cell_6t
Xbit_r229_c69 bl_69 br_69 wl_229 vdd gnd cell_6t
Xbit_r230_c69 bl_69 br_69 wl_230 vdd gnd cell_6t
Xbit_r231_c69 bl_69 br_69 wl_231 vdd gnd cell_6t
Xbit_r232_c69 bl_69 br_69 wl_232 vdd gnd cell_6t
Xbit_r233_c69 bl_69 br_69 wl_233 vdd gnd cell_6t
Xbit_r234_c69 bl_69 br_69 wl_234 vdd gnd cell_6t
Xbit_r235_c69 bl_69 br_69 wl_235 vdd gnd cell_6t
Xbit_r236_c69 bl_69 br_69 wl_236 vdd gnd cell_6t
Xbit_r237_c69 bl_69 br_69 wl_237 vdd gnd cell_6t
Xbit_r238_c69 bl_69 br_69 wl_238 vdd gnd cell_6t
Xbit_r239_c69 bl_69 br_69 wl_239 vdd gnd cell_6t
Xbit_r240_c69 bl_69 br_69 wl_240 vdd gnd cell_6t
Xbit_r241_c69 bl_69 br_69 wl_241 vdd gnd cell_6t
Xbit_r242_c69 bl_69 br_69 wl_242 vdd gnd cell_6t
Xbit_r243_c69 bl_69 br_69 wl_243 vdd gnd cell_6t
Xbit_r244_c69 bl_69 br_69 wl_244 vdd gnd cell_6t
Xbit_r245_c69 bl_69 br_69 wl_245 vdd gnd cell_6t
Xbit_r246_c69 bl_69 br_69 wl_246 vdd gnd cell_6t
Xbit_r247_c69 bl_69 br_69 wl_247 vdd gnd cell_6t
Xbit_r248_c69 bl_69 br_69 wl_248 vdd gnd cell_6t
Xbit_r249_c69 bl_69 br_69 wl_249 vdd gnd cell_6t
Xbit_r250_c69 bl_69 br_69 wl_250 vdd gnd cell_6t
Xbit_r251_c69 bl_69 br_69 wl_251 vdd gnd cell_6t
Xbit_r252_c69 bl_69 br_69 wl_252 vdd gnd cell_6t
Xbit_r253_c69 bl_69 br_69 wl_253 vdd gnd cell_6t
Xbit_r254_c69 bl_69 br_69 wl_254 vdd gnd cell_6t
Xbit_r255_c69 bl_69 br_69 wl_255 vdd gnd cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd cell_6t
Xbit_r1_c70 bl_70 br_70 wl_1 vdd gnd cell_6t
Xbit_r2_c70 bl_70 br_70 wl_2 vdd gnd cell_6t
Xbit_r3_c70 bl_70 br_70 wl_3 vdd gnd cell_6t
Xbit_r4_c70 bl_70 br_70 wl_4 vdd gnd cell_6t
Xbit_r5_c70 bl_70 br_70 wl_5 vdd gnd cell_6t
Xbit_r6_c70 bl_70 br_70 wl_6 vdd gnd cell_6t
Xbit_r7_c70 bl_70 br_70 wl_7 vdd gnd cell_6t
Xbit_r8_c70 bl_70 br_70 wl_8 vdd gnd cell_6t
Xbit_r9_c70 bl_70 br_70 wl_9 vdd gnd cell_6t
Xbit_r10_c70 bl_70 br_70 wl_10 vdd gnd cell_6t
Xbit_r11_c70 bl_70 br_70 wl_11 vdd gnd cell_6t
Xbit_r12_c70 bl_70 br_70 wl_12 vdd gnd cell_6t
Xbit_r13_c70 bl_70 br_70 wl_13 vdd gnd cell_6t
Xbit_r14_c70 bl_70 br_70 wl_14 vdd gnd cell_6t
Xbit_r15_c70 bl_70 br_70 wl_15 vdd gnd cell_6t
Xbit_r16_c70 bl_70 br_70 wl_16 vdd gnd cell_6t
Xbit_r17_c70 bl_70 br_70 wl_17 vdd gnd cell_6t
Xbit_r18_c70 bl_70 br_70 wl_18 vdd gnd cell_6t
Xbit_r19_c70 bl_70 br_70 wl_19 vdd gnd cell_6t
Xbit_r20_c70 bl_70 br_70 wl_20 vdd gnd cell_6t
Xbit_r21_c70 bl_70 br_70 wl_21 vdd gnd cell_6t
Xbit_r22_c70 bl_70 br_70 wl_22 vdd gnd cell_6t
Xbit_r23_c70 bl_70 br_70 wl_23 vdd gnd cell_6t
Xbit_r24_c70 bl_70 br_70 wl_24 vdd gnd cell_6t
Xbit_r25_c70 bl_70 br_70 wl_25 vdd gnd cell_6t
Xbit_r26_c70 bl_70 br_70 wl_26 vdd gnd cell_6t
Xbit_r27_c70 bl_70 br_70 wl_27 vdd gnd cell_6t
Xbit_r28_c70 bl_70 br_70 wl_28 vdd gnd cell_6t
Xbit_r29_c70 bl_70 br_70 wl_29 vdd gnd cell_6t
Xbit_r30_c70 bl_70 br_70 wl_30 vdd gnd cell_6t
Xbit_r31_c70 bl_70 br_70 wl_31 vdd gnd cell_6t
Xbit_r32_c70 bl_70 br_70 wl_32 vdd gnd cell_6t
Xbit_r33_c70 bl_70 br_70 wl_33 vdd gnd cell_6t
Xbit_r34_c70 bl_70 br_70 wl_34 vdd gnd cell_6t
Xbit_r35_c70 bl_70 br_70 wl_35 vdd gnd cell_6t
Xbit_r36_c70 bl_70 br_70 wl_36 vdd gnd cell_6t
Xbit_r37_c70 bl_70 br_70 wl_37 vdd gnd cell_6t
Xbit_r38_c70 bl_70 br_70 wl_38 vdd gnd cell_6t
Xbit_r39_c70 bl_70 br_70 wl_39 vdd gnd cell_6t
Xbit_r40_c70 bl_70 br_70 wl_40 vdd gnd cell_6t
Xbit_r41_c70 bl_70 br_70 wl_41 vdd gnd cell_6t
Xbit_r42_c70 bl_70 br_70 wl_42 vdd gnd cell_6t
Xbit_r43_c70 bl_70 br_70 wl_43 vdd gnd cell_6t
Xbit_r44_c70 bl_70 br_70 wl_44 vdd gnd cell_6t
Xbit_r45_c70 bl_70 br_70 wl_45 vdd gnd cell_6t
Xbit_r46_c70 bl_70 br_70 wl_46 vdd gnd cell_6t
Xbit_r47_c70 bl_70 br_70 wl_47 vdd gnd cell_6t
Xbit_r48_c70 bl_70 br_70 wl_48 vdd gnd cell_6t
Xbit_r49_c70 bl_70 br_70 wl_49 vdd gnd cell_6t
Xbit_r50_c70 bl_70 br_70 wl_50 vdd gnd cell_6t
Xbit_r51_c70 bl_70 br_70 wl_51 vdd gnd cell_6t
Xbit_r52_c70 bl_70 br_70 wl_52 vdd gnd cell_6t
Xbit_r53_c70 bl_70 br_70 wl_53 vdd gnd cell_6t
Xbit_r54_c70 bl_70 br_70 wl_54 vdd gnd cell_6t
Xbit_r55_c70 bl_70 br_70 wl_55 vdd gnd cell_6t
Xbit_r56_c70 bl_70 br_70 wl_56 vdd gnd cell_6t
Xbit_r57_c70 bl_70 br_70 wl_57 vdd gnd cell_6t
Xbit_r58_c70 bl_70 br_70 wl_58 vdd gnd cell_6t
Xbit_r59_c70 bl_70 br_70 wl_59 vdd gnd cell_6t
Xbit_r60_c70 bl_70 br_70 wl_60 vdd gnd cell_6t
Xbit_r61_c70 bl_70 br_70 wl_61 vdd gnd cell_6t
Xbit_r62_c70 bl_70 br_70 wl_62 vdd gnd cell_6t
Xbit_r63_c70 bl_70 br_70 wl_63 vdd gnd cell_6t
Xbit_r64_c70 bl_70 br_70 wl_64 vdd gnd cell_6t
Xbit_r65_c70 bl_70 br_70 wl_65 vdd gnd cell_6t
Xbit_r66_c70 bl_70 br_70 wl_66 vdd gnd cell_6t
Xbit_r67_c70 bl_70 br_70 wl_67 vdd gnd cell_6t
Xbit_r68_c70 bl_70 br_70 wl_68 vdd gnd cell_6t
Xbit_r69_c70 bl_70 br_70 wl_69 vdd gnd cell_6t
Xbit_r70_c70 bl_70 br_70 wl_70 vdd gnd cell_6t
Xbit_r71_c70 bl_70 br_70 wl_71 vdd gnd cell_6t
Xbit_r72_c70 bl_70 br_70 wl_72 vdd gnd cell_6t
Xbit_r73_c70 bl_70 br_70 wl_73 vdd gnd cell_6t
Xbit_r74_c70 bl_70 br_70 wl_74 vdd gnd cell_6t
Xbit_r75_c70 bl_70 br_70 wl_75 vdd gnd cell_6t
Xbit_r76_c70 bl_70 br_70 wl_76 vdd gnd cell_6t
Xbit_r77_c70 bl_70 br_70 wl_77 vdd gnd cell_6t
Xbit_r78_c70 bl_70 br_70 wl_78 vdd gnd cell_6t
Xbit_r79_c70 bl_70 br_70 wl_79 vdd gnd cell_6t
Xbit_r80_c70 bl_70 br_70 wl_80 vdd gnd cell_6t
Xbit_r81_c70 bl_70 br_70 wl_81 vdd gnd cell_6t
Xbit_r82_c70 bl_70 br_70 wl_82 vdd gnd cell_6t
Xbit_r83_c70 bl_70 br_70 wl_83 vdd gnd cell_6t
Xbit_r84_c70 bl_70 br_70 wl_84 vdd gnd cell_6t
Xbit_r85_c70 bl_70 br_70 wl_85 vdd gnd cell_6t
Xbit_r86_c70 bl_70 br_70 wl_86 vdd gnd cell_6t
Xbit_r87_c70 bl_70 br_70 wl_87 vdd gnd cell_6t
Xbit_r88_c70 bl_70 br_70 wl_88 vdd gnd cell_6t
Xbit_r89_c70 bl_70 br_70 wl_89 vdd gnd cell_6t
Xbit_r90_c70 bl_70 br_70 wl_90 vdd gnd cell_6t
Xbit_r91_c70 bl_70 br_70 wl_91 vdd gnd cell_6t
Xbit_r92_c70 bl_70 br_70 wl_92 vdd gnd cell_6t
Xbit_r93_c70 bl_70 br_70 wl_93 vdd gnd cell_6t
Xbit_r94_c70 bl_70 br_70 wl_94 vdd gnd cell_6t
Xbit_r95_c70 bl_70 br_70 wl_95 vdd gnd cell_6t
Xbit_r96_c70 bl_70 br_70 wl_96 vdd gnd cell_6t
Xbit_r97_c70 bl_70 br_70 wl_97 vdd gnd cell_6t
Xbit_r98_c70 bl_70 br_70 wl_98 vdd gnd cell_6t
Xbit_r99_c70 bl_70 br_70 wl_99 vdd gnd cell_6t
Xbit_r100_c70 bl_70 br_70 wl_100 vdd gnd cell_6t
Xbit_r101_c70 bl_70 br_70 wl_101 vdd gnd cell_6t
Xbit_r102_c70 bl_70 br_70 wl_102 vdd gnd cell_6t
Xbit_r103_c70 bl_70 br_70 wl_103 vdd gnd cell_6t
Xbit_r104_c70 bl_70 br_70 wl_104 vdd gnd cell_6t
Xbit_r105_c70 bl_70 br_70 wl_105 vdd gnd cell_6t
Xbit_r106_c70 bl_70 br_70 wl_106 vdd gnd cell_6t
Xbit_r107_c70 bl_70 br_70 wl_107 vdd gnd cell_6t
Xbit_r108_c70 bl_70 br_70 wl_108 vdd gnd cell_6t
Xbit_r109_c70 bl_70 br_70 wl_109 vdd gnd cell_6t
Xbit_r110_c70 bl_70 br_70 wl_110 vdd gnd cell_6t
Xbit_r111_c70 bl_70 br_70 wl_111 vdd gnd cell_6t
Xbit_r112_c70 bl_70 br_70 wl_112 vdd gnd cell_6t
Xbit_r113_c70 bl_70 br_70 wl_113 vdd gnd cell_6t
Xbit_r114_c70 bl_70 br_70 wl_114 vdd gnd cell_6t
Xbit_r115_c70 bl_70 br_70 wl_115 vdd gnd cell_6t
Xbit_r116_c70 bl_70 br_70 wl_116 vdd gnd cell_6t
Xbit_r117_c70 bl_70 br_70 wl_117 vdd gnd cell_6t
Xbit_r118_c70 bl_70 br_70 wl_118 vdd gnd cell_6t
Xbit_r119_c70 bl_70 br_70 wl_119 vdd gnd cell_6t
Xbit_r120_c70 bl_70 br_70 wl_120 vdd gnd cell_6t
Xbit_r121_c70 bl_70 br_70 wl_121 vdd gnd cell_6t
Xbit_r122_c70 bl_70 br_70 wl_122 vdd gnd cell_6t
Xbit_r123_c70 bl_70 br_70 wl_123 vdd gnd cell_6t
Xbit_r124_c70 bl_70 br_70 wl_124 vdd gnd cell_6t
Xbit_r125_c70 bl_70 br_70 wl_125 vdd gnd cell_6t
Xbit_r126_c70 bl_70 br_70 wl_126 vdd gnd cell_6t
Xbit_r127_c70 bl_70 br_70 wl_127 vdd gnd cell_6t
Xbit_r128_c70 bl_70 br_70 wl_128 vdd gnd cell_6t
Xbit_r129_c70 bl_70 br_70 wl_129 vdd gnd cell_6t
Xbit_r130_c70 bl_70 br_70 wl_130 vdd gnd cell_6t
Xbit_r131_c70 bl_70 br_70 wl_131 vdd gnd cell_6t
Xbit_r132_c70 bl_70 br_70 wl_132 vdd gnd cell_6t
Xbit_r133_c70 bl_70 br_70 wl_133 vdd gnd cell_6t
Xbit_r134_c70 bl_70 br_70 wl_134 vdd gnd cell_6t
Xbit_r135_c70 bl_70 br_70 wl_135 vdd gnd cell_6t
Xbit_r136_c70 bl_70 br_70 wl_136 vdd gnd cell_6t
Xbit_r137_c70 bl_70 br_70 wl_137 vdd gnd cell_6t
Xbit_r138_c70 bl_70 br_70 wl_138 vdd gnd cell_6t
Xbit_r139_c70 bl_70 br_70 wl_139 vdd gnd cell_6t
Xbit_r140_c70 bl_70 br_70 wl_140 vdd gnd cell_6t
Xbit_r141_c70 bl_70 br_70 wl_141 vdd gnd cell_6t
Xbit_r142_c70 bl_70 br_70 wl_142 vdd gnd cell_6t
Xbit_r143_c70 bl_70 br_70 wl_143 vdd gnd cell_6t
Xbit_r144_c70 bl_70 br_70 wl_144 vdd gnd cell_6t
Xbit_r145_c70 bl_70 br_70 wl_145 vdd gnd cell_6t
Xbit_r146_c70 bl_70 br_70 wl_146 vdd gnd cell_6t
Xbit_r147_c70 bl_70 br_70 wl_147 vdd gnd cell_6t
Xbit_r148_c70 bl_70 br_70 wl_148 vdd gnd cell_6t
Xbit_r149_c70 bl_70 br_70 wl_149 vdd gnd cell_6t
Xbit_r150_c70 bl_70 br_70 wl_150 vdd gnd cell_6t
Xbit_r151_c70 bl_70 br_70 wl_151 vdd gnd cell_6t
Xbit_r152_c70 bl_70 br_70 wl_152 vdd gnd cell_6t
Xbit_r153_c70 bl_70 br_70 wl_153 vdd gnd cell_6t
Xbit_r154_c70 bl_70 br_70 wl_154 vdd gnd cell_6t
Xbit_r155_c70 bl_70 br_70 wl_155 vdd gnd cell_6t
Xbit_r156_c70 bl_70 br_70 wl_156 vdd gnd cell_6t
Xbit_r157_c70 bl_70 br_70 wl_157 vdd gnd cell_6t
Xbit_r158_c70 bl_70 br_70 wl_158 vdd gnd cell_6t
Xbit_r159_c70 bl_70 br_70 wl_159 vdd gnd cell_6t
Xbit_r160_c70 bl_70 br_70 wl_160 vdd gnd cell_6t
Xbit_r161_c70 bl_70 br_70 wl_161 vdd gnd cell_6t
Xbit_r162_c70 bl_70 br_70 wl_162 vdd gnd cell_6t
Xbit_r163_c70 bl_70 br_70 wl_163 vdd gnd cell_6t
Xbit_r164_c70 bl_70 br_70 wl_164 vdd gnd cell_6t
Xbit_r165_c70 bl_70 br_70 wl_165 vdd gnd cell_6t
Xbit_r166_c70 bl_70 br_70 wl_166 vdd gnd cell_6t
Xbit_r167_c70 bl_70 br_70 wl_167 vdd gnd cell_6t
Xbit_r168_c70 bl_70 br_70 wl_168 vdd gnd cell_6t
Xbit_r169_c70 bl_70 br_70 wl_169 vdd gnd cell_6t
Xbit_r170_c70 bl_70 br_70 wl_170 vdd gnd cell_6t
Xbit_r171_c70 bl_70 br_70 wl_171 vdd gnd cell_6t
Xbit_r172_c70 bl_70 br_70 wl_172 vdd gnd cell_6t
Xbit_r173_c70 bl_70 br_70 wl_173 vdd gnd cell_6t
Xbit_r174_c70 bl_70 br_70 wl_174 vdd gnd cell_6t
Xbit_r175_c70 bl_70 br_70 wl_175 vdd gnd cell_6t
Xbit_r176_c70 bl_70 br_70 wl_176 vdd gnd cell_6t
Xbit_r177_c70 bl_70 br_70 wl_177 vdd gnd cell_6t
Xbit_r178_c70 bl_70 br_70 wl_178 vdd gnd cell_6t
Xbit_r179_c70 bl_70 br_70 wl_179 vdd gnd cell_6t
Xbit_r180_c70 bl_70 br_70 wl_180 vdd gnd cell_6t
Xbit_r181_c70 bl_70 br_70 wl_181 vdd gnd cell_6t
Xbit_r182_c70 bl_70 br_70 wl_182 vdd gnd cell_6t
Xbit_r183_c70 bl_70 br_70 wl_183 vdd gnd cell_6t
Xbit_r184_c70 bl_70 br_70 wl_184 vdd gnd cell_6t
Xbit_r185_c70 bl_70 br_70 wl_185 vdd gnd cell_6t
Xbit_r186_c70 bl_70 br_70 wl_186 vdd gnd cell_6t
Xbit_r187_c70 bl_70 br_70 wl_187 vdd gnd cell_6t
Xbit_r188_c70 bl_70 br_70 wl_188 vdd gnd cell_6t
Xbit_r189_c70 bl_70 br_70 wl_189 vdd gnd cell_6t
Xbit_r190_c70 bl_70 br_70 wl_190 vdd gnd cell_6t
Xbit_r191_c70 bl_70 br_70 wl_191 vdd gnd cell_6t
Xbit_r192_c70 bl_70 br_70 wl_192 vdd gnd cell_6t
Xbit_r193_c70 bl_70 br_70 wl_193 vdd gnd cell_6t
Xbit_r194_c70 bl_70 br_70 wl_194 vdd gnd cell_6t
Xbit_r195_c70 bl_70 br_70 wl_195 vdd gnd cell_6t
Xbit_r196_c70 bl_70 br_70 wl_196 vdd gnd cell_6t
Xbit_r197_c70 bl_70 br_70 wl_197 vdd gnd cell_6t
Xbit_r198_c70 bl_70 br_70 wl_198 vdd gnd cell_6t
Xbit_r199_c70 bl_70 br_70 wl_199 vdd gnd cell_6t
Xbit_r200_c70 bl_70 br_70 wl_200 vdd gnd cell_6t
Xbit_r201_c70 bl_70 br_70 wl_201 vdd gnd cell_6t
Xbit_r202_c70 bl_70 br_70 wl_202 vdd gnd cell_6t
Xbit_r203_c70 bl_70 br_70 wl_203 vdd gnd cell_6t
Xbit_r204_c70 bl_70 br_70 wl_204 vdd gnd cell_6t
Xbit_r205_c70 bl_70 br_70 wl_205 vdd gnd cell_6t
Xbit_r206_c70 bl_70 br_70 wl_206 vdd gnd cell_6t
Xbit_r207_c70 bl_70 br_70 wl_207 vdd gnd cell_6t
Xbit_r208_c70 bl_70 br_70 wl_208 vdd gnd cell_6t
Xbit_r209_c70 bl_70 br_70 wl_209 vdd gnd cell_6t
Xbit_r210_c70 bl_70 br_70 wl_210 vdd gnd cell_6t
Xbit_r211_c70 bl_70 br_70 wl_211 vdd gnd cell_6t
Xbit_r212_c70 bl_70 br_70 wl_212 vdd gnd cell_6t
Xbit_r213_c70 bl_70 br_70 wl_213 vdd gnd cell_6t
Xbit_r214_c70 bl_70 br_70 wl_214 vdd gnd cell_6t
Xbit_r215_c70 bl_70 br_70 wl_215 vdd gnd cell_6t
Xbit_r216_c70 bl_70 br_70 wl_216 vdd gnd cell_6t
Xbit_r217_c70 bl_70 br_70 wl_217 vdd gnd cell_6t
Xbit_r218_c70 bl_70 br_70 wl_218 vdd gnd cell_6t
Xbit_r219_c70 bl_70 br_70 wl_219 vdd gnd cell_6t
Xbit_r220_c70 bl_70 br_70 wl_220 vdd gnd cell_6t
Xbit_r221_c70 bl_70 br_70 wl_221 vdd gnd cell_6t
Xbit_r222_c70 bl_70 br_70 wl_222 vdd gnd cell_6t
Xbit_r223_c70 bl_70 br_70 wl_223 vdd gnd cell_6t
Xbit_r224_c70 bl_70 br_70 wl_224 vdd gnd cell_6t
Xbit_r225_c70 bl_70 br_70 wl_225 vdd gnd cell_6t
Xbit_r226_c70 bl_70 br_70 wl_226 vdd gnd cell_6t
Xbit_r227_c70 bl_70 br_70 wl_227 vdd gnd cell_6t
Xbit_r228_c70 bl_70 br_70 wl_228 vdd gnd cell_6t
Xbit_r229_c70 bl_70 br_70 wl_229 vdd gnd cell_6t
Xbit_r230_c70 bl_70 br_70 wl_230 vdd gnd cell_6t
Xbit_r231_c70 bl_70 br_70 wl_231 vdd gnd cell_6t
Xbit_r232_c70 bl_70 br_70 wl_232 vdd gnd cell_6t
Xbit_r233_c70 bl_70 br_70 wl_233 vdd gnd cell_6t
Xbit_r234_c70 bl_70 br_70 wl_234 vdd gnd cell_6t
Xbit_r235_c70 bl_70 br_70 wl_235 vdd gnd cell_6t
Xbit_r236_c70 bl_70 br_70 wl_236 vdd gnd cell_6t
Xbit_r237_c70 bl_70 br_70 wl_237 vdd gnd cell_6t
Xbit_r238_c70 bl_70 br_70 wl_238 vdd gnd cell_6t
Xbit_r239_c70 bl_70 br_70 wl_239 vdd gnd cell_6t
Xbit_r240_c70 bl_70 br_70 wl_240 vdd gnd cell_6t
Xbit_r241_c70 bl_70 br_70 wl_241 vdd gnd cell_6t
Xbit_r242_c70 bl_70 br_70 wl_242 vdd gnd cell_6t
Xbit_r243_c70 bl_70 br_70 wl_243 vdd gnd cell_6t
Xbit_r244_c70 bl_70 br_70 wl_244 vdd gnd cell_6t
Xbit_r245_c70 bl_70 br_70 wl_245 vdd gnd cell_6t
Xbit_r246_c70 bl_70 br_70 wl_246 vdd gnd cell_6t
Xbit_r247_c70 bl_70 br_70 wl_247 vdd gnd cell_6t
Xbit_r248_c70 bl_70 br_70 wl_248 vdd gnd cell_6t
Xbit_r249_c70 bl_70 br_70 wl_249 vdd gnd cell_6t
Xbit_r250_c70 bl_70 br_70 wl_250 vdd gnd cell_6t
Xbit_r251_c70 bl_70 br_70 wl_251 vdd gnd cell_6t
Xbit_r252_c70 bl_70 br_70 wl_252 vdd gnd cell_6t
Xbit_r253_c70 bl_70 br_70 wl_253 vdd gnd cell_6t
Xbit_r254_c70 bl_70 br_70 wl_254 vdd gnd cell_6t
Xbit_r255_c70 bl_70 br_70 wl_255 vdd gnd cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd cell_6t
Xbit_r1_c71 bl_71 br_71 wl_1 vdd gnd cell_6t
Xbit_r2_c71 bl_71 br_71 wl_2 vdd gnd cell_6t
Xbit_r3_c71 bl_71 br_71 wl_3 vdd gnd cell_6t
Xbit_r4_c71 bl_71 br_71 wl_4 vdd gnd cell_6t
Xbit_r5_c71 bl_71 br_71 wl_5 vdd gnd cell_6t
Xbit_r6_c71 bl_71 br_71 wl_6 vdd gnd cell_6t
Xbit_r7_c71 bl_71 br_71 wl_7 vdd gnd cell_6t
Xbit_r8_c71 bl_71 br_71 wl_8 vdd gnd cell_6t
Xbit_r9_c71 bl_71 br_71 wl_9 vdd gnd cell_6t
Xbit_r10_c71 bl_71 br_71 wl_10 vdd gnd cell_6t
Xbit_r11_c71 bl_71 br_71 wl_11 vdd gnd cell_6t
Xbit_r12_c71 bl_71 br_71 wl_12 vdd gnd cell_6t
Xbit_r13_c71 bl_71 br_71 wl_13 vdd gnd cell_6t
Xbit_r14_c71 bl_71 br_71 wl_14 vdd gnd cell_6t
Xbit_r15_c71 bl_71 br_71 wl_15 vdd gnd cell_6t
Xbit_r16_c71 bl_71 br_71 wl_16 vdd gnd cell_6t
Xbit_r17_c71 bl_71 br_71 wl_17 vdd gnd cell_6t
Xbit_r18_c71 bl_71 br_71 wl_18 vdd gnd cell_6t
Xbit_r19_c71 bl_71 br_71 wl_19 vdd gnd cell_6t
Xbit_r20_c71 bl_71 br_71 wl_20 vdd gnd cell_6t
Xbit_r21_c71 bl_71 br_71 wl_21 vdd gnd cell_6t
Xbit_r22_c71 bl_71 br_71 wl_22 vdd gnd cell_6t
Xbit_r23_c71 bl_71 br_71 wl_23 vdd gnd cell_6t
Xbit_r24_c71 bl_71 br_71 wl_24 vdd gnd cell_6t
Xbit_r25_c71 bl_71 br_71 wl_25 vdd gnd cell_6t
Xbit_r26_c71 bl_71 br_71 wl_26 vdd gnd cell_6t
Xbit_r27_c71 bl_71 br_71 wl_27 vdd gnd cell_6t
Xbit_r28_c71 bl_71 br_71 wl_28 vdd gnd cell_6t
Xbit_r29_c71 bl_71 br_71 wl_29 vdd gnd cell_6t
Xbit_r30_c71 bl_71 br_71 wl_30 vdd gnd cell_6t
Xbit_r31_c71 bl_71 br_71 wl_31 vdd gnd cell_6t
Xbit_r32_c71 bl_71 br_71 wl_32 vdd gnd cell_6t
Xbit_r33_c71 bl_71 br_71 wl_33 vdd gnd cell_6t
Xbit_r34_c71 bl_71 br_71 wl_34 vdd gnd cell_6t
Xbit_r35_c71 bl_71 br_71 wl_35 vdd gnd cell_6t
Xbit_r36_c71 bl_71 br_71 wl_36 vdd gnd cell_6t
Xbit_r37_c71 bl_71 br_71 wl_37 vdd gnd cell_6t
Xbit_r38_c71 bl_71 br_71 wl_38 vdd gnd cell_6t
Xbit_r39_c71 bl_71 br_71 wl_39 vdd gnd cell_6t
Xbit_r40_c71 bl_71 br_71 wl_40 vdd gnd cell_6t
Xbit_r41_c71 bl_71 br_71 wl_41 vdd gnd cell_6t
Xbit_r42_c71 bl_71 br_71 wl_42 vdd gnd cell_6t
Xbit_r43_c71 bl_71 br_71 wl_43 vdd gnd cell_6t
Xbit_r44_c71 bl_71 br_71 wl_44 vdd gnd cell_6t
Xbit_r45_c71 bl_71 br_71 wl_45 vdd gnd cell_6t
Xbit_r46_c71 bl_71 br_71 wl_46 vdd gnd cell_6t
Xbit_r47_c71 bl_71 br_71 wl_47 vdd gnd cell_6t
Xbit_r48_c71 bl_71 br_71 wl_48 vdd gnd cell_6t
Xbit_r49_c71 bl_71 br_71 wl_49 vdd gnd cell_6t
Xbit_r50_c71 bl_71 br_71 wl_50 vdd gnd cell_6t
Xbit_r51_c71 bl_71 br_71 wl_51 vdd gnd cell_6t
Xbit_r52_c71 bl_71 br_71 wl_52 vdd gnd cell_6t
Xbit_r53_c71 bl_71 br_71 wl_53 vdd gnd cell_6t
Xbit_r54_c71 bl_71 br_71 wl_54 vdd gnd cell_6t
Xbit_r55_c71 bl_71 br_71 wl_55 vdd gnd cell_6t
Xbit_r56_c71 bl_71 br_71 wl_56 vdd gnd cell_6t
Xbit_r57_c71 bl_71 br_71 wl_57 vdd gnd cell_6t
Xbit_r58_c71 bl_71 br_71 wl_58 vdd gnd cell_6t
Xbit_r59_c71 bl_71 br_71 wl_59 vdd gnd cell_6t
Xbit_r60_c71 bl_71 br_71 wl_60 vdd gnd cell_6t
Xbit_r61_c71 bl_71 br_71 wl_61 vdd gnd cell_6t
Xbit_r62_c71 bl_71 br_71 wl_62 vdd gnd cell_6t
Xbit_r63_c71 bl_71 br_71 wl_63 vdd gnd cell_6t
Xbit_r64_c71 bl_71 br_71 wl_64 vdd gnd cell_6t
Xbit_r65_c71 bl_71 br_71 wl_65 vdd gnd cell_6t
Xbit_r66_c71 bl_71 br_71 wl_66 vdd gnd cell_6t
Xbit_r67_c71 bl_71 br_71 wl_67 vdd gnd cell_6t
Xbit_r68_c71 bl_71 br_71 wl_68 vdd gnd cell_6t
Xbit_r69_c71 bl_71 br_71 wl_69 vdd gnd cell_6t
Xbit_r70_c71 bl_71 br_71 wl_70 vdd gnd cell_6t
Xbit_r71_c71 bl_71 br_71 wl_71 vdd gnd cell_6t
Xbit_r72_c71 bl_71 br_71 wl_72 vdd gnd cell_6t
Xbit_r73_c71 bl_71 br_71 wl_73 vdd gnd cell_6t
Xbit_r74_c71 bl_71 br_71 wl_74 vdd gnd cell_6t
Xbit_r75_c71 bl_71 br_71 wl_75 vdd gnd cell_6t
Xbit_r76_c71 bl_71 br_71 wl_76 vdd gnd cell_6t
Xbit_r77_c71 bl_71 br_71 wl_77 vdd gnd cell_6t
Xbit_r78_c71 bl_71 br_71 wl_78 vdd gnd cell_6t
Xbit_r79_c71 bl_71 br_71 wl_79 vdd gnd cell_6t
Xbit_r80_c71 bl_71 br_71 wl_80 vdd gnd cell_6t
Xbit_r81_c71 bl_71 br_71 wl_81 vdd gnd cell_6t
Xbit_r82_c71 bl_71 br_71 wl_82 vdd gnd cell_6t
Xbit_r83_c71 bl_71 br_71 wl_83 vdd gnd cell_6t
Xbit_r84_c71 bl_71 br_71 wl_84 vdd gnd cell_6t
Xbit_r85_c71 bl_71 br_71 wl_85 vdd gnd cell_6t
Xbit_r86_c71 bl_71 br_71 wl_86 vdd gnd cell_6t
Xbit_r87_c71 bl_71 br_71 wl_87 vdd gnd cell_6t
Xbit_r88_c71 bl_71 br_71 wl_88 vdd gnd cell_6t
Xbit_r89_c71 bl_71 br_71 wl_89 vdd gnd cell_6t
Xbit_r90_c71 bl_71 br_71 wl_90 vdd gnd cell_6t
Xbit_r91_c71 bl_71 br_71 wl_91 vdd gnd cell_6t
Xbit_r92_c71 bl_71 br_71 wl_92 vdd gnd cell_6t
Xbit_r93_c71 bl_71 br_71 wl_93 vdd gnd cell_6t
Xbit_r94_c71 bl_71 br_71 wl_94 vdd gnd cell_6t
Xbit_r95_c71 bl_71 br_71 wl_95 vdd gnd cell_6t
Xbit_r96_c71 bl_71 br_71 wl_96 vdd gnd cell_6t
Xbit_r97_c71 bl_71 br_71 wl_97 vdd gnd cell_6t
Xbit_r98_c71 bl_71 br_71 wl_98 vdd gnd cell_6t
Xbit_r99_c71 bl_71 br_71 wl_99 vdd gnd cell_6t
Xbit_r100_c71 bl_71 br_71 wl_100 vdd gnd cell_6t
Xbit_r101_c71 bl_71 br_71 wl_101 vdd gnd cell_6t
Xbit_r102_c71 bl_71 br_71 wl_102 vdd gnd cell_6t
Xbit_r103_c71 bl_71 br_71 wl_103 vdd gnd cell_6t
Xbit_r104_c71 bl_71 br_71 wl_104 vdd gnd cell_6t
Xbit_r105_c71 bl_71 br_71 wl_105 vdd gnd cell_6t
Xbit_r106_c71 bl_71 br_71 wl_106 vdd gnd cell_6t
Xbit_r107_c71 bl_71 br_71 wl_107 vdd gnd cell_6t
Xbit_r108_c71 bl_71 br_71 wl_108 vdd gnd cell_6t
Xbit_r109_c71 bl_71 br_71 wl_109 vdd gnd cell_6t
Xbit_r110_c71 bl_71 br_71 wl_110 vdd gnd cell_6t
Xbit_r111_c71 bl_71 br_71 wl_111 vdd gnd cell_6t
Xbit_r112_c71 bl_71 br_71 wl_112 vdd gnd cell_6t
Xbit_r113_c71 bl_71 br_71 wl_113 vdd gnd cell_6t
Xbit_r114_c71 bl_71 br_71 wl_114 vdd gnd cell_6t
Xbit_r115_c71 bl_71 br_71 wl_115 vdd gnd cell_6t
Xbit_r116_c71 bl_71 br_71 wl_116 vdd gnd cell_6t
Xbit_r117_c71 bl_71 br_71 wl_117 vdd gnd cell_6t
Xbit_r118_c71 bl_71 br_71 wl_118 vdd gnd cell_6t
Xbit_r119_c71 bl_71 br_71 wl_119 vdd gnd cell_6t
Xbit_r120_c71 bl_71 br_71 wl_120 vdd gnd cell_6t
Xbit_r121_c71 bl_71 br_71 wl_121 vdd gnd cell_6t
Xbit_r122_c71 bl_71 br_71 wl_122 vdd gnd cell_6t
Xbit_r123_c71 bl_71 br_71 wl_123 vdd gnd cell_6t
Xbit_r124_c71 bl_71 br_71 wl_124 vdd gnd cell_6t
Xbit_r125_c71 bl_71 br_71 wl_125 vdd gnd cell_6t
Xbit_r126_c71 bl_71 br_71 wl_126 vdd gnd cell_6t
Xbit_r127_c71 bl_71 br_71 wl_127 vdd gnd cell_6t
Xbit_r128_c71 bl_71 br_71 wl_128 vdd gnd cell_6t
Xbit_r129_c71 bl_71 br_71 wl_129 vdd gnd cell_6t
Xbit_r130_c71 bl_71 br_71 wl_130 vdd gnd cell_6t
Xbit_r131_c71 bl_71 br_71 wl_131 vdd gnd cell_6t
Xbit_r132_c71 bl_71 br_71 wl_132 vdd gnd cell_6t
Xbit_r133_c71 bl_71 br_71 wl_133 vdd gnd cell_6t
Xbit_r134_c71 bl_71 br_71 wl_134 vdd gnd cell_6t
Xbit_r135_c71 bl_71 br_71 wl_135 vdd gnd cell_6t
Xbit_r136_c71 bl_71 br_71 wl_136 vdd gnd cell_6t
Xbit_r137_c71 bl_71 br_71 wl_137 vdd gnd cell_6t
Xbit_r138_c71 bl_71 br_71 wl_138 vdd gnd cell_6t
Xbit_r139_c71 bl_71 br_71 wl_139 vdd gnd cell_6t
Xbit_r140_c71 bl_71 br_71 wl_140 vdd gnd cell_6t
Xbit_r141_c71 bl_71 br_71 wl_141 vdd gnd cell_6t
Xbit_r142_c71 bl_71 br_71 wl_142 vdd gnd cell_6t
Xbit_r143_c71 bl_71 br_71 wl_143 vdd gnd cell_6t
Xbit_r144_c71 bl_71 br_71 wl_144 vdd gnd cell_6t
Xbit_r145_c71 bl_71 br_71 wl_145 vdd gnd cell_6t
Xbit_r146_c71 bl_71 br_71 wl_146 vdd gnd cell_6t
Xbit_r147_c71 bl_71 br_71 wl_147 vdd gnd cell_6t
Xbit_r148_c71 bl_71 br_71 wl_148 vdd gnd cell_6t
Xbit_r149_c71 bl_71 br_71 wl_149 vdd gnd cell_6t
Xbit_r150_c71 bl_71 br_71 wl_150 vdd gnd cell_6t
Xbit_r151_c71 bl_71 br_71 wl_151 vdd gnd cell_6t
Xbit_r152_c71 bl_71 br_71 wl_152 vdd gnd cell_6t
Xbit_r153_c71 bl_71 br_71 wl_153 vdd gnd cell_6t
Xbit_r154_c71 bl_71 br_71 wl_154 vdd gnd cell_6t
Xbit_r155_c71 bl_71 br_71 wl_155 vdd gnd cell_6t
Xbit_r156_c71 bl_71 br_71 wl_156 vdd gnd cell_6t
Xbit_r157_c71 bl_71 br_71 wl_157 vdd gnd cell_6t
Xbit_r158_c71 bl_71 br_71 wl_158 vdd gnd cell_6t
Xbit_r159_c71 bl_71 br_71 wl_159 vdd gnd cell_6t
Xbit_r160_c71 bl_71 br_71 wl_160 vdd gnd cell_6t
Xbit_r161_c71 bl_71 br_71 wl_161 vdd gnd cell_6t
Xbit_r162_c71 bl_71 br_71 wl_162 vdd gnd cell_6t
Xbit_r163_c71 bl_71 br_71 wl_163 vdd gnd cell_6t
Xbit_r164_c71 bl_71 br_71 wl_164 vdd gnd cell_6t
Xbit_r165_c71 bl_71 br_71 wl_165 vdd gnd cell_6t
Xbit_r166_c71 bl_71 br_71 wl_166 vdd gnd cell_6t
Xbit_r167_c71 bl_71 br_71 wl_167 vdd gnd cell_6t
Xbit_r168_c71 bl_71 br_71 wl_168 vdd gnd cell_6t
Xbit_r169_c71 bl_71 br_71 wl_169 vdd gnd cell_6t
Xbit_r170_c71 bl_71 br_71 wl_170 vdd gnd cell_6t
Xbit_r171_c71 bl_71 br_71 wl_171 vdd gnd cell_6t
Xbit_r172_c71 bl_71 br_71 wl_172 vdd gnd cell_6t
Xbit_r173_c71 bl_71 br_71 wl_173 vdd gnd cell_6t
Xbit_r174_c71 bl_71 br_71 wl_174 vdd gnd cell_6t
Xbit_r175_c71 bl_71 br_71 wl_175 vdd gnd cell_6t
Xbit_r176_c71 bl_71 br_71 wl_176 vdd gnd cell_6t
Xbit_r177_c71 bl_71 br_71 wl_177 vdd gnd cell_6t
Xbit_r178_c71 bl_71 br_71 wl_178 vdd gnd cell_6t
Xbit_r179_c71 bl_71 br_71 wl_179 vdd gnd cell_6t
Xbit_r180_c71 bl_71 br_71 wl_180 vdd gnd cell_6t
Xbit_r181_c71 bl_71 br_71 wl_181 vdd gnd cell_6t
Xbit_r182_c71 bl_71 br_71 wl_182 vdd gnd cell_6t
Xbit_r183_c71 bl_71 br_71 wl_183 vdd gnd cell_6t
Xbit_r184_c71 bl_71 br_71 wl_184 vdd gnd cell_6t
Xbit_r185_c71 bl_71 br_71 wl_185 vdd gnd cell_6t
Xbit_r186_c71 bl_71 br_71 wl_186 vdd gnd cell_6t
Xbit_r187_c71 bl_71 br_71 wl_187 vdd gnd cell_6t
Xbit_r188_c71 bl_71 br_71 wl_188 vdd gnd cell_6t
Xbit_r189_c71 bl_71 br_71 wl_189 vdd gnd cell_6t
Xbit_r190_c71 bl_71 br_71 wl_190 vdd gnd cell_6t
Xbit_r191_c71 bl_71 br_71 wl_191 vdd gnd cell_6t
Xbit_r192_c71 bl_71 br_71 wl_192 vdd gnd cell_6t
Xbit_r193_c71 bl_71 br_71 wl_193 vdd gnd cell_6t
Xbit_r194_c71 bl_71 br_71 wl_194 vdd gnd cell_6t
Xbit_r195_c71 bl_71 br_71 wl_195 vdd gnd cell_6t
Xbit_r196_c71 bl_71 br_71 wl_196 vdd gnd cell_6t
Xbit_r197_c71 bl_71 br_71 wl_197 vdd gnd cell_6t
Xbit_r198_c71 bl_71 br_71 wl_198 vdd gnd cell_6t
Xbit_r199_c71 bl_71 br_71 wl_199 vdd gnd cell_6t
Xbit_r200_c71 bl_71 br_71 wl_200 vdd gnd cell_6t
Xbit_r201_c71 bl_71 br_71 wl_201 vdd gnd cell_6t
Xbit_r202_c71 bl_71 br_71 wl_202 vdd gnd cell_6t
Xbit_r203_c71 bl_71 br_71 wl_203 vdd gnd cell_6t
Xbit_r204_c71 bl_71 br_71 wl_204 vdd gnd cell_6t
Xbit_r205_c71 bl_71 br_71 wl_205 vdd gnd cell_6t
Xbit_r206_c71 bl_71 br_71 wl_206 vdd gnd cell_6t
Xbit_r207_c71 bl_71 br_71 wl_207 vdd gnd cell_6t
Xbit_r208_c71 bl_71 br_71 wl_208 vdd gnd cell_6t
Xbit_r209_c71 bl_71 br_71 wl_209 vdd gnd cell_6t
Xbit_r210_c71 bl_71 br_71 wl_210 vdd gnd cell_6t
Xbit_r211_c71 bl_71 br_71 wl_211 vdd gnd cell_6t
Xbit_r212_c71 bl_71 br_71 wl_212 vdd gnd cell_6t
Xbit_r213_c71 bl_71 br_71 wl_213 vdd gnd cell_6t
Xbit_r214_c71 bl_71 br_71 wl_214 vdd gnd cell_6t
Xbit_r215_c71 bl_71 br_71 wl_215 vdd gnd cell_6t
Xbit_r216_c71 bl_71 br_71 wl_216 vdd gnd cell_6t
Xbit_r217_c71 bl_71 br_71 wl_217 vdd gnd cell_6t
Xbit_r218_c71 bl_71 br_71 wl_218 vdd gnd cell_6t
Xbit_r219_c71 bl_71 br_71 wl_219 vdd gnd cell_6t
Xbit_r220_c71 bl_71 br_71 wl_220 vdd gnd cell_6t
Xbit_r221_c71 bl_71 br_71 wl_221 vdd gnd cell_6t
Xbit_r222_c71 bl_71 br_71 wl_222 vdd gnd cell_6t
Xbit_r223_c71 bl_71 br_71 wl_223 vdd gnd cell_6t
Xbit_r224_c71 bl_71 br_71 wl_224 vdd gnd cell_6t
Xbit_r225_c71 bl_71 br_71 wl_225 vdd gnd cell_6t
Xbit_r226_c71 bl_71 br_71 wl_226 vdd gnd cell_6t
Xbit_r227_c71 bl_71 br_71 wl_227 vdd gnd cell_6t
Xbit_r228_c71 bl_71 br_71 wl_228 vdd gnd cell_6t
Xbit_r229_c71 bl_71 br_71 wl_229 vdd gnd cell_6t
Xbit_r230_c71 bl_71 br_71 wl_230 vdd gnd cell_6t
Xbit_r231_c71 bl_71 br_71 wl_231 vdd gnd cell_6t
Xbit_r232_c71 bl_71 br_71 wl_232 vdd gnd cell_6t
Xbit_r233_c71 bl_71 br_71 wl_233 vdd gnd cell_6t
Xbit_r234_c71 bl_71 br_71 wl_234 vdd gnd cell_6t
Xbit_r235_c71 bl_71 br_71 wl_235 vdd gnd cell_6t
Xbit_r236_c71 bl_71 br_71 wl_236 vdd gnd cell_6t
Xbit_r237_c71 bl_71 br_71 wl_237 vdd gnd cell_6t
Xbit_r238_c71 bl_71 br_71 wl_238 vdd gnd cell_6t
Xbit_r239_c71 bl_71 br_71 wl_239 vdd gnd cell_6t
Xbit_r240_c71 bl_71 br_71 wl_240 vdd gnd cell_6t
Xbit_r241_c71 bl_71 br_71 wl_241 vdd gnd cell_6t
Xbit_r242_c71 bl_71 br_71 wl_242 vdd gnd cell_6t
Xbit_r243_c71 bl_71 br_71 wl_243 vdd gnd cell_6t
Xbit_r244_c71 bl_71 br_71 wl_244 vdd gnd cell_6t
Xbit_r245_c71 bl_71 br_71 wl_245 vdd gnd cell_6t
Xbit_r246_c71 bl_71 br_71 wl_246 vdd gnd cell_6t
Xbit_r247_c71 bl_71 br_71 wl_247 vdd gnd cell_6t
Xbit_r248_c71 bl_71 br_71 wl_248 vdd gnd cell_6t
Xbit_r249_c71 bl_71 br_71 wl_249 vdd gnd cell_6t
Xbit_r250_c71 bl_71 br_71 wl_250 vdd gnd cell_6t
Xbit_r251_c71 bl_71 br_71 wl_251 vdd gnd cell_6t
Xbit_r252_c71 bl_71 br_71 wl_252 vdd gnd cell_6t
Xbit_r253_c71 bl_71 br_71 wl_253 vdd gnd cell_6t
Xbit_r254_c71 bl_71 br_71 wl_254 vdd gnd cell_6t
Xbit_r255_c71 bl_71 br_71 wl_255 vdd gnd cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd cell_6t
Xbit_r1_c72 bl_72 br_72 wl_1 vdd gnd cell_6t
Xbit_r2_c72 bl_72 br_72 wl_2 vdd gnd cell_6t
Xbit_r3_c72 bl_72 br_72 wl_3 vdd gnd cell_6t
Xbit_r4_c72 bl_72 br_72 wl_4 vdd gnd cell_6t
Xbit_r5_c72 bl_72 br_72 wl_5 vdd gnd cell_6t
Xbit_r6_c72 bl_72 br_72 wl_6 vdd gnd cell_6t
Xbit_r7_c72 bl_72 br_72 wl_7 vdd gnd cell_6t
Xbit_r8_c72 bl_72 br_72 wl_8 vdd gnd cell_6t
Xbit_r9_c72 bl_72 br_72 wl_9 vdd gnd cell_6t
Xbit_r10_c72 bl_72 br_72 wl_10 vdd gnd cell_6t
Xbit_r11_c72 bl_72 br_72 wl_11 vdd gnd cell_6t
Xbit_r12_c72 bl_72 br_72 wl_12 vdd gnd cell_6t
Xbit_r13_c72 bl_72 br_72 wl_13 vdd gnd cell_6t
Xbit_r14_c72 bl_72 br_72 wl_14 vdd gnd cell_6t
Xbit_r15_c72 bl_72 br_72 wl_15 vdd gnd cell_6t
Xbit_r16_c72 bl_72 br_72 wl_16 vdd gnd cell_6t
Xbit_r17_c72 bl_72 br_72 wl_17 vdd gnd cell_6t
Xbit_r18_c72 bl_72 br_72 wl_18 vdd gnd cell_6t
Xbit_r19_c72 bl_72 br_72 wl_19 vdd gnd cell_6t
Xbit_r20_c72 bl_72 br_72 wl_20 vdd gnd cell_6t
Xbit_r21_c72 bl_72 br_72 wl_21 vdd gnd cell_6t
Xbit_r22_c72 bl_72 br_72 wl_22 vdd gnd cell_6t
Xbit_r23_c72 bl_72 br_72 wl_23 vdd gnd cell_6t
Xbit_r24_c72 bl_72 br_72 wl_24 vdd gnd cell_6t
Xbit_r25_c72 bl_72 br_72 wl_25 vdd gnd cell_6t
Xbit_r26_c72 bl_72 br_72 wl_26 vdd gnd cell_6t
Xbit_r27_c72 bl_72 br_72 wl_27 vdd gnd cell_6t
Xbit_r28_c72 bl_72 br_72 wl_28 vdd gnd cell_6t
Xbit_r29_c72 bl_72 br_72 wl_29 vdd gnd cell_6t
Xbit_r30_c72 bl_72 br_72 wl_30 vdd gnd cell_6t
Xbit_r31_c72 bl_72 br_72 wl_31 vdd gnd cell_6t
Xbit_r32_c72 bl_72 br_72 wl_32 vdd gnd cell_6t
Xbit_r33_c72 bl_72 br_72 wl_33 vdd gnd cell_6t
Xbit_r34_c72 bl_72 br_72 wl_34 vdd gnd cell_6t
Xbit_r35_c72 bl_72 br_72 wl_35 vdd gnd cell_6t
Xbit_r36_c72 bl_72 br_72 wl_36 vdd gnd cell_6t
Xbit_r37_c72 bl_72 br_72 wl_37 vdd gnd cell_6t
Xbit_r38_c72 bl_72 br_72 wl_38 vdd gnd cell_6t
Xbit_r39_c72 bl_72 br_72 wl_39 vdd gnd cell_6t
Xbit_r40_c72 bl_72 br_72 wl_40 vdd gnd cell_6t
Xbit_r41_c72 bl_72 br_72 wl_41 vdd gnd cell_6t
Xbit_r42_c72 bl_72 br_72 wl_42 vdd gnd cell_6t
Xbit_r43_c72 bl_72 br_72 wl_43 vdd gnd cell_6t
Xbit_r44_c72 bl_72 br_72 wl_44 vdd gnd cell_6t
Xbit_r45_c72 bl_72 br_72 wl_45 vdd gnd cell_6t
Xbit_r46_c72 bl_72 br_72 wl_46 vdd gnd cell_6t
Xbit_r47_c72 bl_72 br_72 wl_47 vdd gnd cell_6t
Xbit_r48_c72 bl_72 br_72 wl_48 vdd gnd cell_6t
Xbit_r49_c72 bl_72 br_72 wl_49 vdd gnd cell_6t
Xbit_r50_c72 bl_72 br_72 wl_50 vdd gnd cell_6t
Xbit_r51_c72 bl_72 br_72 wl_51 vdd gnd cell_6t
Xbit_r52_c72 bl_72 br_72 wl_52 vdd gnd cell_6t
Xbit_r53_c72 bl_72 br_72 wl_53 vdd gnd cell_6t
Xbit_r54_c72 bl_72 br_72 wl_54 vdd gnd cell_6t
Xbit_r55_c72 bl_72 br_72 wl_55 vdd gnd cell_6t
Xbit_r56_c72 bl_72 br_72 wl_56 vdd gnd cell_6t
Xbit_r57_c72 bl_72 br_72 wl_57 vdd gnd cell_6t
Xbit_r58_c72 bl_72 br_72 wl_58 vdd gnd cell_6t
Xbit_r59_c72 bl_72 br_72 wl_59 vdd gnd cell_6t
Xbit_r60_c72 bl_72 br_72 wl_60 vdd gnd cell_6t
Xbit_r61_c72 bl_72 br_72 wl_61 vdd gnd cell_6t
Xbit_r62_c72 bl_72 br_72 wl_62 vdd gnd cell_6t
Xbit_r63_c72 bl_72 br_72 wl_63 vdd gnd cell_6t
Xbit_r64_c72 bl_72 br_72 wl_64 vdd gnd cell_6t
Xbit_r65_c72 bl_72 br_72 wl_65 vdd gnd cell_6t
Xbit_r66_c72 bl_72 br_72 wl_66 vdd gnd cell_6t
Xbit_r67_c72 bl_72 br_72 wl_67 vdd gnd cell_6t
Xbit_r68_c72 bl_72 br_72 wl_68 vdd gnd cell_6t
Xbit_r69_c72 bl_72 br_72 wl_69 vdd gnd cell_6t
Xbit_r70_c72 bl_72 br_72 wl_70 vdd gnd cell_6t
Xbit_r71_c72 bl_72 br_72 wl_71 vdd gnd cell_6t
Xbit_r72_c72 bl_72 br_72 wl_72 vdd gnd cell_6t
Xbit_r73_c72 bl_72 br_72 wl_73 vdd gnd cell_6t
Xbit_r74_c72 bl_72 br_72 wl_74 vdd gnd cell_6t
Xbit_r75_c72 bl_72 br_72 wl_75 vdd gnd cell_6t
Xbit_r76_c72 bl_72 br_72 wl_76 vdd gnd cell_6t
Xbit_r77_c72 bl_72 br_72 wl_77 vdd gnd cell_6t
Xbit_r78_c72 bl_72 br_72 wl_78 vdd gnd cell_6t
Xbit_r79_c72 bl_72 br_72 wl_79 vdd gnd cell_6t
Xbit_r80_c72 bl_72 br_72 wl_80 vdd gnd cell_6t
Xbit_r81_c72 bl_72 br_72 wl_81 vdd gnd cell_6t
Xbit_r82_c72 bl_72 br_72 wl_82 vdd gnd cell_6t
Xbit_r83_c72 bl_72 br_72 wl_83 vdd gnd cell_6t
Xbit_r84_c72 bl_72 br_72 wl_84 vdd gnd cell_6t
Xbit_r85_c72 bl_72 br_72 wl_85 vdd gnd cell_6t
Xbit_r86_c72 bl_72 br_72 wl_86 vdd gnd cell_6t
Xbit_r87_c72 bl_72 br_72 wl_87 vdd gnd cell_6t
Xbit_r88_c72 bl_72 br_72 wl_88 vdd gnd cell_6t
Xbit_r89_c72 bl_72 br_72 wl_89 vdd gnd cell_6t
Xbit_r90_c72 bl_72 br_72 wl_90 vdd gnd cell_6t
Xbit_r91_c72 bl_72 br_72 wl_91 vdd gnd cell_6t
Xbit_r92_c72 bl_72 br_72 wl_92 vdd gnd cell_6t
Xbit_r93_c72 bl_72 br_72 wl_93 vdd gnd cell_6t
Xbit_r94_c72 bl_72 br_72 wl_94 vdd gnd cell_6t
Xbit_r95_c72 bl_72 br_72 wl_95 vdd gnd cell_6t
Xbit_r96_c72 bl_72 br_72 wl_96 vdd gnd cell_6t
Xbit_r97_c72 bl_72 br_72 wl_97 vdd gnd cell_6t
Xbit_r98_c72 bl_72 br_72 wl_98 vdd gnd cell_6t
Xbit_r99_c72 bl_72 br_72 wl_99 vdd gnd cell_6t
Xbit_r100_c72 bl_72 br_72 wl_100 vdd gnd cell_6t
Xbit_r101_c72 bl_72 br_72 wl_101 vdd gnd cell_6t
Xbit_r102_c72 bl_72 br_72 wl_102 vdd gnd cell_6t
Xbit_r103_c72 bl_72 br_72 wl_103 vdd gnd cell_6t
Xbit_r104_c72 bl_72 br_72 wl_104 vdd gnd cell_6t
Xbit_r105_c72 bl_72 br_72 wl_105 vdd gnd cell_6t
Xbit_r106_c72 bl_72 br_72 wl_106 vdd gnd cell_6t
Xbit_r107_c72 bl_72 br_72 wl_107 vdd gnd cell_6t
Xbit_r108_c72 bl_72 br_72 wl_108 vdd gnd cell_6t
Xbit_r109_c72 bl_72 br_72 wl_109 vdd gnd cell_6t
Xbit_r110_c72 bl_72 br_72 wl_110 vdd gnd cell_6t
Xbit_r111_c72 bl_72 br_72 wl_111 vdd gnd cell_6t
Xbit_r112_c72 bl_72 br_72 wl_112 vdd gnd cell_6t
Xbit_r113_c72 bl_72 br_72 wl_113 vdd gnd cell_6t
Xbit_r114_c72 bl_72 br_72 wl_114 vdd gnd cell_6t
Xbit_r115_c72 bl_72 br_72 wl_115 vdd gnd cell_6t
Xbit_r116_c72 bl_72 br_72 wl_116 vdd gnd cell_6t
Xbit_r117_c72 bl_72 br_72 wl_117 vdd gnd cell_6t
Xbit_r118_c72 bl_72 br_72 wl_118 vdd gnd cell_6t
Xbit_r119_c72 bl_72 br_72 wl_119 vdd gnd cell_6t
Xbit_r120_c72 bl_72 br_72 wl_120 vdd gnd cell_6t
Xbit_r121_c72 bl_72 br_72 wl_121 vdd gnd cell_6t
Xbit_r122_c72 bl_72 br_72 wl_122 vdd gnd cell_6t
Xbit_r123_c72 bl_72 br_72 wl_123 vdd gnd cell_6t
Xbit_r124_c72 bl_72 br_72 wl_124 vdd gnd cell_6t
Xbit_r125_c72 bl_72 br_72 wl_125 vdd gnd cell_6t
Xbit_r126_c72 bl_72 br_72 wl_126 vdd gnd cell_6t
Xbit_r127_c72 bl_72 br_72 wl_127 vdd gnd cell_6t
Xbit_r128_c72 bl_72 br_72 wl_128 vdd gnd cell_6t
Xbit_r129_c72 bl_72 br_72 wl_129 vdd gnd cell_6t
Xbit_r130_c72 bl_72 br_72 wl_130 vdd gnd cell_6t
Xbit_r131_c72 bl_72 br_72 wl_131 vdd gnd cell_6t
Xbit_r132_c72 bl_72 br_72 wl_132 vdd gnd cell_6t
Xbit_r133_c72 bl_72 br_72 wl_133 vdd gnd cell_6t
Xbit_r134_c72 bl_72 br_72 wl_134 vdd gnd cell_6t
Xbit_r135_c72 bl_72 br_72 wl_135 vdd gnd cell_6t
Xbit_r136_c72 bl_72 br_72 wl_136 vdd gnd cell_6t
Xbit_r137_c72 bl_72 br_72 wl_137 vdd gnd cell_6t
Xbit_r138_c72 bl_72 br_72 wl_138 vdd gnd cell_6t
Xbit_r139_c72 bl_72 br_72 wl_139 vdd gnd cell_6t
Xbit_r140_c72 bl_72 br_72 wl_140 vdd gnd cell_6t
Xbit_r141_c72 bl_72 br_72 wl_141 vdd gnd cell_6t
Xbit_r142_c72 bl_72 br_72 wl_142 vdd gnd cell_6t
Xbit_r143_c72 bl_72 br_72 wl_143 vdd gnd cell_6t
Xbit_r144_c72 bl_72 br_72 wl_144 vdd gnd cell_6t
Xbit_r145_c72 bl_72 br_72 wl_145 vdd gnd cell_6t
Xbit_r146_c72 bl_72 br_72 wl_146 vdd gnd cell_6t
Xbit_r147_c72 bl_72 br_72 wl_147 vdd gnd cell_6t
Xbit_r148_c72 bl_72 br_72 wl_148 vdd gnd cell_6t
Xbit_r149_c72 bl_72 br_72 wl_149 vdd gnd cell_6t
Xbit_r150_c72 bl_72 br_72 wl_150 vdd gnd cell_6t
Xbit_r151_c72 bl_72 br_72 wl_151 vdd gnd cell_6t
Xbit_r152_c72 bl_72 br_72 wl_152 vdd gnd cell_6t
Xbit_r153_c72 bl_72 br_72 wl_153 vdd gnd cell_6t
Xbit_r154_c72 bl_72 br_72 wl_154 vdd gnd cell_6t
Xbit_r155_c72 bl_72 br_72 wl_155 vdd gnd cell_6t
Xbit_r156_c72 bl_72 br_72 wl_156 vdd gnd cell_6t
Xbit_r157_c72 bl_72 br_72 wl_157 vdd gnd cell_6t
Xbit_r158_c72 bl_72 br_72 wl_158 vdd gnd cell_6t
Xbit_r159_c72 bl_72 br_72 wl_159 vdd gnd cell_6t
Xbit_r160_c72 bl_72 br_72 wl_160 vdd gnd cell_6t
Xbit_r161_c72 bl_72 br_72 wl_161 vdd gnd cell_6t
Xbit_r162_c72 bl_72 br_72 wl_162 vdd gnd cell_6t
Xbit_r163_c72 bl_72 br_72 wl_163 vdd gnd cell_6t
Xbit_r164_c72 bl_72 br_72 wl_164 vdd gnd cell_6t
Xbit_r165_c72 bl_72 br_72 wl_165 vdd gnd cell_6t
Xbit_r166_c72 bl_72 br_72 wl_166 vdd gnd cell_6t
Xbit_r167_c72 bl_72 br_72 wl_167 vdd gnd cell_6t
Xbit_r168_c72 bl_72 br_72 wl_168 vdd gnd cell_6t
Xbit_r169_c72 bl_72 br_72 wl_169 vdd gnd cell_6t
Xbit_r170_c72 bl_72 br_72 wl_170 vdd gnd cell_6t
Xbit_r171_c72 bl_72 br_72 wl_171 vdd gnd cell_6t
Xbit_r172_c72 bl_72 br_72 wl_172 vdd gnd cell_6t
Xbit_r173_c72 bl_72 br_72 wl_173 vdd gnd cell_6t
Xbit_r174_c72 bl_72 br_72 wl_174 vdd gnd cell_6t
Xbit_r175_c72 bl_72 br_72 wl_175 vdd gnd cell_6t
Xbit_r176_c72 bl_72 br_72 wl_176 vdd gnd cell_6t
Xbit_r177_c72 bl_72 br_72 wl_177 vdd gnd cell_6t
Xbit_r178_c72 bl_72 br_72 wl_178 vdd gnd cell_6t
Xbit_r179_c72 bl_72 br_72 wl_179 vdd gnd cell_6t
Xbit_r180_c72 bl_72 br_72 wl_180 vdd gnd cell_6t
Xbit_r181_c72 bl_72 br_72 wl_181 vdd gnd cell_6t
Xbit_r182_c72 bl_72 br_72 wl_182 vdd gnd cell_6t
Xbit_r183_c72 bl_72 br_72 wl_183 vdd gnd cell_6t
Xbit_r184_c72 bl_72 br_72 wl_184 vdd gnd cell_6t
Xbit_r185_c72 bl_72 br_72 wl_185 vdd gnd cell_6t
Xbit_r186_c72 bl_72 br_72 wl_186 vdd gnd cell_6t
Xbit_r187_c72 bl_72 br_72 wl_187 vdd gnd cell_6t
Xbit_r188_c72 bl_72 br_72 wl_188 vdd gnd cell_6t
Xbit_r189_c72 bl_72 br_72 wl_189 vdd gnd cell_6t
Xbit_r190_c72 bl_72 br_72 wl_190 vdd gnd cell_6t
Xbit_r191_c72 bl_72 br_72 wl_191 vdd gnd cell_6t
Xbit_r192_c72 bl_72 br_72 wl_192 vdd gnd cell_6t
Xbit_r193_c72 bl_72 br_72 wl_193 vdd gnd cell_6t
Xbit_r194_c72 bl_72 br_72 wl_194 vdd gnd cell_6t
Xbit_r195_c72 bl_72 br_72 wl_195 vdd gnd cell_6t
Xbit_r196_c72 bl_72 br_72 wl_196 vdd gnd cell_6t
Xbit_r197_c72 bl_72 br_72 wl_197 vdd gnd cell_6t
Xbit_r198_c72 bl_72 br_72 wl_198 vdd gnd cell_6t
Xbit_r199_c72 bl_72 br_72 wl_199 vdd gnd cell_6t
Xbit_r200_c72 bl_72 br_72 wl_200 vdd gnd cell_6t
Xbit_r201_c72 bl_72 br_72 wl_201 vdd gnd cell_6t
Xbit_r202_c72 bl_72 br_72 wl_202 vdd gnd cell_6t
Xbit_r203_c72 bl_72 br_72 wl_203 vdd gnd cell_6t
Xbit_r204_c72 bl_72 br_72 wl_204 vdd gnd cell_6t
Xbit_r205_c72 bl_72 br_72 wl_205 vdd gnd cell_6t
Xbit_r206_c72 bl_72 br_72 wl_206 vdd gnd cell_6t
Xbit_r207_c72 bl_72 br_72 wl_207 vdd gnd cell_6t
Xbit_r208_c72 bl_72 br_72 wl_208 vdd gnd cell_6t
Xbit_r209_c72 bl_72 br_72 wl_209 vdd gnd cell_6t
Xbit_r210_c72 bl_72 br_72 wl_210 vdd gnd cell_6t
Xbit_r211_c72 bl_72 br_72 wl_211 vdd gnd cell_6t
Xbit_r212_c72 bl_72 br_72 wl_212 vdd gnd cell_6t
Xbit_r213_c72 bl_72 br_72 wl_213 vdd gnd cell_6t
Xbit_r214_c72 bl_72 br_72 wl_214 vdd gnd cell_6t
Xbit_r215_c72 bl_72 br_72 wl_215 vdd gnd cell_6t
Xbit_r216_c72 bl_72 br_72 wl_216 vdd gnd cell_6t
Xbit_r217_c72 bl_72 br_72 wl_217 vdd gnd cell_6t
Xbit_r218_c72 bl_72 br_72 wl_218 vdd gnd cell_6t
Xbit_r219_c72 bl_72 br_72 wl_219 vdd gnd cell_6t
Xbit_r220_c72 bl_72 br_72 wl_220 vdd gnd cell_6t
Xbit_r221_c72 bl_72 br_72 wl_221 vdd gnd cell_6t
Xbit_r222_c72 bl_72 br_72 wl_222 vdd gnd cell_6t
Xbit_r223_c72 bl_72 br_72 wl_223 vdd gnd cell_6t
Xbit_r224_c72 bl_72 br_72 wl_224 vdd gnd cell_6t
Xbit_r225_c72 bl_72 br_72 wl_225 vdd gnd cell_6t
Xbit_r226_c72 bl_72 br_72 wl_226 vdd gnd cell_6t
Xbit_r227_c72 bl_72 br_72 wl_227 vdd gnd cell_6t
Xbit_r228_c72 bl_72 br_72 wl_228 vdd gnd cell_6t
Xbit_r229_c72 bl_72 br_72 wl_229 vdd gnd cell_6t
Xbit_r230_c72 bl_72 br_72 wl_230 vdd gnd cell_6t
Xbit_r231_c72 bl_72 br_72 wl_231 vdd gnd cell_6t
Xbit_r232_c72 bl_72 br_72 wl_232 vdd gnd cell_6t
Xbit_r233_c72 bl_72 br_72 wl_233 vdd gnd cell_6t
Xbit_r234_c72 bl_72 br_72 wl_234 vdd gnd cell_6t
Xbit_r235_c72 bl_72 br_72 wl_235 vdd gnd cell_6t
Xbit_r236_c72 bl_72 br_72 wl_236 vdd gnd cell_6t
Xbit_r237_c72 bl_72 br_72 wl_237 vdd gnd cell_6t
Xbit_r238_c72 bl_72 br_72 wl_238 vdd gnd cell_6t
Xbit_r239_c72 bl_72 br_72 wl_239 vdd gnd cell_6t
Xbit_r240_c72 bl_72 br_72 wl_240 vdd gnd cell_6t
Xbit_r241_c72 bl_72 br_72 wl_241 vdd gnd cell_6t
Xbit_r242_c72 bl_72 br_72 wl_242 vdd gnd cell_6t
Xbit_r243_c72 bl_72 br_72 wl_243 vdd gnd cell_6t
Xbit_r244_c72 bl_72 br_72 wl_244 vdd gnd cell_6t
Xbit_r245_c72 bl_72 br_72 wl_245 vdd gnd cell_6t
Xbit_r246_c72 bl_72 br_72 wl_246 vdd gnd cell_6t
Xbit_r247_c72 bl_72 br_72 wl_247 vdd gnd cell_6t
Xbit_r248_c72 bl_72 br_72 wl_248 vdd gnd cell_6t
Xbit_r249_c72 bl_72 br_72 wl_249 vdd gnd cell_6t
Xbit_r250_c72 bl_72 br_72 wl_250 vdd gnd cell_6t
Xbit_r251_c72 bl_72 br_72 wl_251 vdd gnd cell_6t
Xbit_r252_c72 bl_72 br_72 wl_252 vdd gnd cell_6t
Xbit_r253_c72 bl_72 br_72 wl_253 vdd gnd cell_6t
Xbit_r254_c72 bl_72 br_72 wl_254 vdd gnd cell_6t
Xbit_r255_c72 bl_72 br_72 wl_255 vdd gnd cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd cell_6t
Xbit_r1_c73 bl_73 br_73 wl_1 vdd gnd cell_6t
Xbit_r2_c73 bl_73 br_73 wl_2 vdd gnd cell_6t
Xbit_r3_c73 bl_73 br_73 wl_3 vdd gnd cell_6t
Xbit_r4_c73 bl_73 br_73 wl_4 vdd gnd cell_6t
Xbit_r5_c73 bl_73 br_73 wl_5 vdd gnd cell_6t
Xbit_r6_c73 bl_73 br_73 wl_6 vdd gnd cell_6t
Xbit_r7_c73 bl_73 br_73 wl_7 vdd gnd cell_6t
Xbit_r8_c73 bl_73 br_73 wl_8 vdd gnd cell_6t
Xbit_r9_c73 bl_73 br_73 wl_9 vdd gnd cell_6t
Xbit_r10_c73 bl_73 br_73 wl_10 vdd gnd cell_6t
Xbit_r11_c73 bl_73 br_73 wl_11 vdd gnd cell_6t
Xbit_r12_c73 bl_73 br_73 wl_12 vdd gnd cell_6t
Xbit_r13_c73 bl_73 br_73 wl_13 vdd gnd cell_6t
Xbit_r14_c73 bl_73 br_73 wl_14 vdd gnd cell_6t
Xbit_r15_c73 bl_73 br_73 wl_15 vdd gnd cell_6t
Xbit_r16_c73 bl_73 br_73 wl_16 vdd gnd cell_6t
Xbit_r17_c73 bl_73 br_73 wl_17 vdd gnd cell_6t
Xbit_r18_c73 bl_73 br_73 wl_18 vdd gnd cell_6t
Xbit_r19_c73 bl_73 br_73 wl_19 vdd gnd cell_6t
Xbit_r20_c73 bl_73 br_73 wl_20 vdd gnd cell_6t
Xbit_r21_c73 bl_73 br_73 wl_21 vdd gnd cell_6t
Xbit_r22_c73 bl_73 br_73 wl_22 vdd gnd cell_6t
Xbit_r23_c73 bl_73 br_73 wl_23 vdd gnd cell_6t
Xbit_r24_c73 bl_73 br_73 wl_24 vdd gnd cell_6t
Xbit_r25_c73 bl_73 br_73 wl_25 vdd gnd cell_6t
Xbit_r26_c73 bl_73 br_73 wl_26 vdd gnd cell_6t
Xbit_r27_c73 bl_73 br_73 wl_27 vdd gnd cell_6t
Xbit_r28_c73 bl_73 br_73 wl_28 vdd gnd cell_6t
Xbit_r29_c73 bl_73 br_73 wl_29 vdd gnd cell_6t
Xbit_r30_c73 bl_73 br_73 wl_30 vdd gnd cell_6t
Xbit_r31_c73 bl_73 br_73 wl_31 vdd gnd cell_6t
Xbit_r32_c73 bl_73 br_73 wl_32 vdd gnd cell_6t
Xbit_r33_c73 bl_73 br_73 wl_33 vdd gnd cell_6t
Xbit_r34_c73 bl_73 br_73 wl_34 vdd gnd cell_6t
Xbit_r35_c73 bl_73 br_73 wl_35 vdd gnd cell_6t
Xbit_r36_c73 bl_73 br_73 wl_36 vdd gnd cell_6t
Xbit_r37_c73 bl_73 br_73 wl_37 vdd gnd cell_6t
Xbit_r38_c73 bl_73 br_73 wl_38 vdd gnd cell_6t
Xbit_r39_c73 bl_73 br_73 wl_39 vdd gnd cell_6t
Xbit_r40_c73 bl_73 br_73 wl_40 vdd gnd cell_6t
Xbit_r41_c73 bl_73 br_73 wl_41 vdd gnd cell_6t
Xbit_r42_c73 bl_73 br_73 wl_42 vdd gnd cell_6t
Xbit_r43_c73 bl_73 br_73 wl_43 vdd gnd cell_6t
Xbit_r44_c73 bl_73 br_73 wl_44 vdd gnd cell_6t
Xbit_r45_c73 bl_73 br_73 wl_45 vdd gnd cell_6t
Xbit_r46_c73 bl_73 br_73 wl_46 vdd gnd cell_6t
Xbit_r47_c73 bl_73 br_73 wl_47 vdd gnd cell_6t
Xbit_r48_c73 bl_73 br_73 wl_48 vdd gnd cell_6t
Xbit_r49_c73 bl_73 br_73 wl_49 vdd gnd cell_6t
Xbit_r50_c73 bl_73 br_73 wl_50 vdd gnd cell_6t
Xbit_r51_c73 bl_73 br_73 wl_51 vdd gnd cell_6t
Xbit_r52_c73 bl_73 br_73 wl_52 vdd gnd cell_6t
Xbit_r53_c73 bl_73 br_73 wl_53 vdd gnd cell_6t
Xbit_r54_c73 bl_73 br_73 wl_54 vdd gnd cell_6t
Xbit_r55_c73 bl_73 br_73 wl_55 vdd gnd cell_6t
Xbit_r56_c73 bl_73 br_73 wl_56 vdd gnd cell_6t
Xbit_r57_c73 bl_73 br_73 wl_57 vdd gnd cell_6t
Xbit_r58_c73 bl_73 br_73 wl_58 vdd gnd cell_6t
Xbit_r59_c73 bl_73 br_73 wl_59 vdd gnd cell_6t
Xbit_r60_c73 bl_73 br_73 wl_60 vdd gnd cell_6t
Xbit_r61_c73 bl_73 br_73 wl_61 vdd gnd cell_6t
Xbit_r62_c73 bl_73 br_73 wl_62 vdd gnd cell_6t
Xbit_r63_c73 bl_73 br_73 wl_63 vdd gnd cell_6t
Xbit_r64_c73 bl_73 br_73 wl_64 vdd gnd cell_6t
Xbit_r65_c73 bl_73 br_73 wl_65 vdd gnd cell_6t
Xbit_r66_c73 bl_73 br_73 wl_66 vdd gnd cell_6t
Xbit_r67_c73 bl_73 br_73 wl_67 vdd gnd cell_6t
Xbit_r68_c73 bl_73 br_73 wl_68 vdd gnd cell_6t
Xbit_r69_c73 bl_73 br_73 wl_69 vdd gnd cell_6t
Xbit_r70_c73 bl_73 br_73 wl_70 vdd gnd cell_6t
Xbit_r71_c73 bl_73 br_73 wl_71 vdd gnd cell_6t
Xbit_r72_c73 bl_73 br_73 wl_72 vdd gnd cell_6t
Xbit_r73_c73 bl_73 br_73 wl_73 vdd gnd cell_6t
Xbit_r74_c73 bl_73 br_73 wl_74 vdd gnd cell_6t
Xbit_r75_c73 bl_73 br_73 wl_75 vdd gnd cell_6t
Xbit_r76_c73 bl_73 br_73 wl_76 vdd gnd cell_6t
Xbit_r77_c73 bl_73 br_73 wl_77 vdd gnd cell_6t
Xbit_r78_c73 bl_73 br_73 wl_78 vdd gnd cell_6t
Xbit_r79_c73 bl_73 br_73 wl_79 vdd gnd cell_6t
Xbit_r80_c73 bl_73 br_73 wl_80 vdd gnd cell_6t
Xbit_r81_c73 bl_73 br_73 wl_81 vdd gnd cell_6t
Xbit_r82_c73 bl_73 br_73 wl_82 vdd gnd cell_6t
Xbit_r83_c73 bl_73 br_73 wl_83 vdd gnd cell_6t
Xbit_r84_c73 bl_73 br_73 wl_84 vdd gnd cell_6t
Xbit_r85_c73 bl_73 br_73 wl_85 vdd gnd cell_6t
Xbit_r86_c73 bl_73 br_73 wl_86 vdd gnd cell_6t
Xbit_r87_c73 bl_73 br_73 wl_87 vdd gnd cell_6t
Xbit_r88_c73 bl_73 br_73 wl_88 vdd gnd cell_6t
Xbit_r89_c73 bl_73 br_73 wl_89 vdd gnd cell_6t
Xbit_r90_c73 bl_73 br_73 wl_90 vdd gnd cell_6t
Xbit_r91_c73 bl_73 br_73 wl_91 vdd gnd cell_6t
Xbit_r92_c73 bl_73 br_73 wl_92 vdd gnd cell_6t
Xbit_r93_c73 bl_73 br_73 wl_93 vdd gnd cell_6t
Xbit_r94_c73 bl_73 br_73 wl_94 vdd gnd cell_6t
Xbit_r95_c73 bl_73 br_73 wl_95 vdd gnd cell_6t
Xbit_r96_c73 bl_73 br_73 wl_96 vdd gnd cell_6t
Xbit_r97_c73 bl_73 br_73 wl_97 vdd gnd cell_6t
Xbit_r98_c73 bl_73 br_73 wl_98 vdd gnd cell_6t
Xbit_r99_c73 bl_73 br_73 wl_99 vdd gnd cell_6t
Xbit_r100_c73 bl_73 br_73 wl_100 vdd gnd cell_6t
Xbit_r101_c73 bl_73 br_73 wl_101 vdd gnd cell_6t
Xbit_r102_c73 bl_73 br_73 wl_102 vdd gnd cell_6t
Xbit_r103_c73 bl_73 br_73 wl_103 vdd gnd cell_6t
Xbit_r104_c73 bl_73 br_73 wl_104 vdd gnd cell_6t
Xbit_r105_c73 bl_73 br_73 wl_105 vdd gnd cell_6t
Xbit_r106_c73 bl_73 br_73 wl_106 vdd gnd cell_6t
Xbit_r107_c73 bl_73 br_73 wl_107 vdd gnd cell_6t
Xbit_r108_c73 bl_73 br_73 wl_108 vdd gnd cell_6t
Xbit_r109_c73 bl_73 br_73 wl_109 vdd gnd cell_6t
Xbit_r110_c73 bl_73 br_73 wl_110 vdd gnd cell_6t
Xbit_r111_c73 bl_73 br_73 wl_111 vdd gnd cell_6t
Xbit_r112_c73 bl_73 br_73 wl_112 vdd gnd cell_6t
Xbit_r113_c73 bl_73 br_73 wl_113 vdd gnd cell_6t
Xbit_r114_c73 bl_73 br_73 wl_114 vdd gnd cell_6t
Xbit_r115_c73 bl_73 br_73 wl_115 vdd gnd cell_6t
Xbit_r116_c73 bl_73 br_73 wl_116 vdd gnd cell_6t
Xbit_r117_c73 bl_73 br_73 wl_117 vdd gnd cell_6t
Xbit_r118_c73 bl_73 br_73 wl_118 vdd gnd cell_6t
Xbit_r119_c73 bl_73 br_73 wl_119 vdd gnd cell_6t
Xbit_r120_c73 bl_73 br_73 wl_120 vdd gnd cell_6t
Xbit_r121_c73 bl_73 br_73 wl_121 vdd gnd cell_6t
Xbit_r122_c73 bl_73 br_73 wl_122 vdd gnd cell_6t
Xbit_r123_c73 bl_73 br_73 wl_123 vdd gnd cell_6t
Xbit_r124_c73 bl_73 br_73 wl_124 vdd gnd cell_6t
Xbit_r125_c73 bl_73 br_73 wl_125 vdd gnd cell_6t
Xbit_r126_c73 bl_73 br_73 wl_126 vdd gnd cell_6t
Xbit_r127_c73 bl_73 br_73 wl_127 vdd gnd cell_6t
Xbit_r128_c73 bl_73 br_73 wl_128 vdd gnd cell_6t
Xbit_r129_c73 bl_73 br_73 wl_129 vdd gnd cell_6t
Xbit_r130_c73 bl_73 br_73 wl_130 vdd gnd cell_6t
Xbit_r131_c73 bl_73 br_73 wl_131 vdd gnd cell_6t
Xbit_r132_c73 bl_73 br_73 wl_132 vdd gnd cell_6t
Xbit_r133_c73 bl_73 br_73 wl_133 vdd gnd cell_6t
Xbit_r134_c73 bl_73 br_73 wl_134 vdd gnd cell_6t
Xbit_r135_c73 bl_73 br_73 wl_135 vdd gnd cell_6t
Xbit_r136_c73 bl_73 br_73 wl_136 vdd gnd cell_6t
Xbit_r137_c73 bl_73 br_73 wl_137 vdd gnd cell_6t
Xbit_r138_c73 bl_73 br_73 wl_138 vdd gnd cell_6t
Xbit_r139_c73 bl_73 br_73 wl_139 vdd gnd cell_6t
Xbit_r140_c73 bl_73 br_73 wl_140 vdd gnd cell_6t
Xbit_r141_c73 bl_73 br_73 wl_141 vdd gnd cell_6t
Xbit_r142_c73 bl_73 br_73 wl_142 vdd gnd cell_6t
Xbit_r143_c73 bl_73 br_73 wl_143 vdd gnd cell_6t
Xbit_r144_c73 bl_73 br_73 wl_144 vdd gnd cell_6t
Xbit_r145_c73 bl_73 br_73 wl_145 vdd gnd cell_6t
Xbit_r146_c73 bl_73 br_73 wl_146 vdd gnd cell_6t
Xbit_r147_c73 bl_73 br_73 wl_147 vdd gnd cell_6t
Xbit_r148_c73 bl_73 br_73 wl_148 vdd gnd cell_6t
Xbit_r149_c73 bl_73 br_73 wl_149 vdd gnd cell_6t
Xbit_r150_c73 bl_73 br_73 wl_150 vdd gnd cell_6t
Xbit_r151_c73 bl_73 br_73 wl_151 vdd gnd cell_6t
Xbit_r152_c73 bl_73 br_73 wl_152 vdd gnd cell_6t
Xbit_r153_c73 bl_73 br_73 wl_153 vdd gnd cell_6t
Xbit_r154_c73 bl_73 br_73 wl_154 vdd gnd cell_6t
Xbit_r155_c73 bl_73 br_73 wl_155 vdd gnd cell_6t
Xbit_r156_c73 bl_73 br_73 wl_156 vdd gnd cell_6t
Xbit_r157_c73 bl_73 br_73 wl_157 vdd gnd cell_6t
Xbit_r158_c73 bl_73 br_73 wl_158 vdd gnd cell_6t
Xbit_r159_c73 bl_73 br_73 wl_159 vdd gnd cell_6t
Xbit_r160_c73 bl_73 br_73 wl_160 vdd gnd cell_6t
Xbit_r161_c73 bl_73 br_73 wl_161 vdd gnd cell_6t
Xbit_r162_c73 bl_73 br_73 wl_162 vdd gnd cell_6t
Xbit_r163_c73 bl_73 br_73 wl_163 vdd gnd cell_6t
Xbit_r164_c73 bl_73 br_73 wl_164 vdd gnd cell_6t
Xbit_r165_c73 bl_73 br_73 wl_165 vdd gnd cell_6t
Xbit_r166_c73 bl_73 br_73 wl_166 vdd gnd cell_6t
Xbit_r167_c73 bl_73 br_73 wl_167 vdd gnd cell_6t
Xbit_r168_c73 bl_73 br_73 wl_168 vdd gnd cell_6t
Xbit_r169_c73 bl_73 br_73 wl_169 vdd gnd cell_6t
Xbit_r170_c73 bl_73 br_73 wl_170 vdd gnd cell_6t
Xbit_r171_c73 bl_73 br_73 wl_171 vdd gnd cell_6t
Xbit_r172_c73 bl_73 br_73 wl_172 vdd gnd cell_6t
Xbit_r173_c73 bl_73 br_73 wl_173 vdd gnd cell_6t
Xbit_r174_c73 bl_73 br_73 wl_174 vdd gnd cell_6t
Xbit_r175_c73 bl_73 br_73 wl_175 vdd gnd cell_6t
Xbit_r176_c73 bl_73 br_73 wl_176 vdd gnd cell_6t
Xbit_r177_c73 bl_73 br_73 wl_177 vdd gnd cell_6t
Xbit_r178_c73 bl_73 br_73 wl_178 vdd gnd cell_6t
Xbit_r179_c73 bl_73 br_73 wl_179 vdd gnd cell_6t
Xbit_r180_c73 bl_73 br_73 wl_180 vdd gnd cell_6t
Xbit_r181_c73 bl_73 br_73 wl_181 vdd gnd cell_6t
Xbit_r182_c73 bl_73 br_73 wl_182 vdd gnd cell_6t
Xbit_r183_c73 bl_73 br_73 wl_183 vdd gnd cell_6t
Xbit_r184_c73 bl_73 br_73 wl_184 vdd gnd cell_6t
Xbit_r185_c73 bl_73 br_73 wl_185 vdd gnd cell_6t
Xbit_r186_c73 bl_73 br_73 wl_186 vdd gnd cell_6t
Xbit_r187_c73 bl_73 br_73 wl_187 vdd gnd cell_6t
Xbit_r188_c73 bl_73 br_73 wl_188 vdd gnd cell_6t
Xbit_r189_c73 bl_73 br_73 wl_189 vdd gnd cell_6t
Xbit_r190_c73 bl_73 br_73 wl_190 vdd gnd cell_6t
Xbit_r191_c73 bl_73 br_73 wl_191 vdd gnd cell_6t
Xbit_r192_c73 bl_73 br_73 wl_192 vdd gnd cell_6t
Xbit_r193_c73 bl_73 br_73 wl_193 vdd gnd cell_6t
Xbit_r194_c73 bl_73 br_73 wl_194 vdd gnd cell_6t
Xbit_r195_c73 bl_73 br_73 wl_195 vdd gnd cell_6t
Xbit_r196_c73 bl_73 br_73 wl_196 vdd gnd cell_6t
Xbit_r197_c73 bl_73 br_73 wl_197 vdd gnd cell_6t
Xbit_r198_c73 bl_73 br_73 wl_198 vdd gnd cell_6t
Xbit_r199_c73 bl_73 br_73 wl_199 vdd gnd cell_6t
Xbit_r200_c73 bl_73 br_73 wl_200 vdd gnd cell_6t
Xbit_r201_c73 bl_73 br_73 wl_201 vdd gnd cell_6t
Xbit_r202_c73 bl_73 br_73 wl_202 vdd gnd cell_6t
Xbit_r203_c73 bl_73 br_73 wl_203 vdd gnd cell_6t
Xbit_r204_c73 bl_73 br_73 wl_204 vdd gnd cell_6t
Xbit_r205_c73 bl_73 br_73 wl_205 vdd gnd cell_6t
Xbit_r206_c73 bl_73 br_73 wl_206 vdd gnd cell_6t
Xbit_r207_c73 bl_73 br_73 wl_207 vdd gnd cell_6t
Xbit_r208_c73 bl_73 br_73 wl_208 vdd gnd cell_6t
Xbit_r209_c73 bl_73 br_73 wl_209 vdd gnd cell_6t
Xbit_r210_c73 bl_73 br_73 wl_210 vdd gnd cell_6t
Xbit_r211_c73 bl_73 br_73 wl_211 vdd gnd cell_6t
Xbit_r212_c73 bl_73 br_73 wl_212 vdd gnd cell_6t
Xbit_r213_c73 bl_73 br_73 wl_213 vdd gnd cell_6t
Xbit_r214_c73 bl_73 br_73 wl_214 vdd gnd cell_6t
Xbit_r215_c73 bl_73 br_73 wl_215 vdd gnd cell_6t
Xbit_r216_c73 bl_73 br_73 wl_216 vdd gnd cell_6t
Xbit_r217_c73 bl_73 br_73 wl_217 vdd gnd cell_6t
Xbit_r218_c73 bl_73 br_73 wl_218 vdd gnd cell_6t
Xbit_r219_c73 bl_73 br_73 wl_219 vdd gnd cell_6t
Xbit_r220_c73 bl_73 br_73 wl_220 vdd gnd cell_6t
Xbit_r221_c73 bl_73 br_73 wl_221 vdd gnd cell_6t
Xbit_r222_c73 bl_73 br_73 wl_222 vdd gnd cell_6t
Xbit_r223_c73 bl_73 br_73 wl_223 vdd gnd cell_6t
Xbit_r224_c73 bl_73 br_73 wl_224 vdd gnd cell_6t
Xbit_r225_c73 bl_73 br_73 wl_225 vdd gnd cell_6t
Xbit_r226_c73 bl_73 br_73 wl_226 vdd gnd cell_6t
Xbit_r227_c73 bl_73 br_73 wl_227 vdd gnd cell_6t
Xbit_r228_c73 bl_73 br_73 wl_228 vdd gnd cell_6t
Xbit_r229_c73 bl_73 br_73 wl_229 vdd gnd cell_6t
Xbit_r230_c73 bl_73 br_73 wl_230 vdd gnd cell_6t
Xbit_r231_c73 bl_73 br_73 wl_231 vdd gnd cell_6t
Xbit_r232_c73 bl_73 br_73 wl_232 vdd gnd cell_6t
Xbit_r233_c73 bl_73 br_73 wl_233 vdd gnd cell_6t
Xbit_r234_c73 bl_73 br_73 wl_234 vdd gnd cell_6t
Xbit_r235_c73 bl_73 br_73 wl_235 vdd gnd cell_6t
Xbit_r236_c73 bl_73 br_73 wl_236 vdd gnd cell_6t
Xbit_r237_c73 bl_73 br_73 wl_237 vdd gnd cell_6t
Xbit_r238_c73 bl_73 br_73 wl_238 vdd gnd cell_6t
Xbit_r239_c73 bl_73 br_73 wl_239 vdd gnd cell_6t
Xbit_r240_c73 bl_73 br_73 wl_240 vdd gnd cell_6t
Xbit_r241_c73 bl_73 br_73 wl_241 vdd gnd cell_6t
Xbit_r242_c73 bl_73 br_73 wl_242 vdd gnd cell_6t
Xbit_r243_c73 bl_73 br_73 wl_243 vdd gnd cell_6t
Xbit_r244_c73 bl_73 br_73 wl_244 vdd gnd cell_6t
Xbit_r245_c73 bl_73 br_73 wl_245 vdd gnd cell_6t
Xbit_r246_c73 bl_73 br_73 wl_246 vdd gnd cell_6t
Xbit_r247_c73 bl_73 br_73 wl_247 vdd gnd cell_6t
Xbit_r248_c73 bl_73 br_73 wl_248 vdd gnd cell_6t
Xbit_r249_c73 bl_73 br_73 wl_249 vdd gnd cell_6t
Xbit_r250_c73 bl_73 br_73 wl_250 vdd gnd cell_6t
Xbit_r251_c73 bl_73 br_73 wl_251 vdd gnd cell_6t
Xbit_r252_c73 bl_73 br_73 wl_252 vdd gnd cell_6t
Xbit_r253_c73 bl_73 br_73 wl_253 vdd gnd cell_6t
Xbit_r254_c73 bl_73 br_73 wl_254 vdd gnd cell_6t
Xbit_r255_c73 bl_73 br_73 wl_255 vdd gnd cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd cell_6t
Xbit_r1_c74 bl_74 br_74 wl_1 vdd gnd cell_6t
Xbit_r2_c74 bl_74 br_74 wl_2 vdd gnd cell_6t
Xbit_r3_c74 bl_74 br_74 wl_3 vdd gnd cell_6t
Xbit_r4_c74 bl_74 br_74 wl_4 vdd gnd cell_6t
Xbit_r5_c74 bl_74 br_74 wl_5 vdd gnd cell_6t
Xbit_r6_c74 bl_74 br_74 wl_6 vdd gnd cell_6t
Xbit_r7_c74 bl_74 br_74 wl_7 vdd gnd cell_6t
Xbit_r8_c74 bl_74 br_74 wl_8 vdd gnd cell_6t
Xbit_r9_c74 bl_74 br_74 wl_9 vdd gnd cell_6t
Xbit_r10_c74 bl_74 br_74 wl_10 vdd gnd cell_6t
Xbit_r11_c74 bl_74 br_74 wl_11 vdd gnd cell_6t
Xbit_r12_c74 bl_74 br_74 wl_12 vdd gnd cell_6t
Xbit_r13_c74 bl_74 br_74 wl_13 vdd gnd cell_6t
Xbit_r14_c74 bl_74 br_74 wl_14 vdd gnd cell_6t
Xbit_r15_c74 bl_74 br_74 wl_15 vdd gnd cell_6t
Xbit_r16_c74 bl_74 br_74 wl_16 vdd gnd cell_6t
Xbit_r17_c74 bl_74 br_74 wl_17 vdd gnd cell_6t
Xbit_r18_c74 bl_74 br_74 wl_18 vdd gnd cell_6t
Xbit_r19_c74 bl_74 br_74 wl_19 vdd gnd cell_6t
Xbit_r20_c74 bl_74 br_74 wl_20 vdd gnd cell_6t
Xbit_r21_c74 bl_74 br_74 wl_21 vdd gnd cell_6t
Xbit_r22_c74 bl_74 br_74 wl_22 vdd gnd cell_6t
Xbit_r23_c74 bl_74 br_74 wl_23 vdd gnd cell_6t
Xbit_r24_c74 bl_74 br_74 wl_24 vdd gnd cell_6t
Xbit_r25_c74 bl_74 br_74 wl_25 vdd gnd cell_6t
Xbit_r26_c74 bl_74 br_74 wl_26 vdd gnd cell_6t
Xbit_r27_c74 bl_74 br_74 wl_27 vdd gnd cell_6t
Xbit_r28_c74 bl_74 br_74 wl_28 vdd gnd cell_6t
Xbit_r29_c74 bl_74 br_74 wl_29 vdd gnd cell_6t
Xbit_r30_c74 bl_74 br_74 wl_30 vdd gnd cell_6t
Xbit_r31_c74 bl_74 br_74 wl_31 vdd gnd cell_6t
Xbit_r32_c74 bl_74 br_74 wl_32 vdd gnd cell_6t
Xbit_r33_c74 bl_74 br_74 wl_33 vdd gnd cell_6t
Xbit_r34_c74 bl_74 br_74 wl_34 vdd gnd cell_6t
Xbit_r35_c74 bl_74 br_74 wl_35 vdd gnd cell_6t
Xbit_r36_c74 bl_74 br_74 wl_36 vdd gnd cell_6t
Xbit_r37_c74 bl_74 br_74 wl_37 vdd gnd cell_6t
Xbit_r38_c74 bl_74 br_74 wl_38 vdd gnd cell_6t
Xbit_r39_c74 bl_74 br_74 wl_39 vdd gnd cell_6t
Xbit_r40_c74 bl_74 br_74 wl_40 vdd gnd cell_6t
Xbit_r41_c74 bl_74 br_74 wl_41 vdd gnd cell_6t
Xbit_r42_c74 bl_74 br_74 wl_42 vdd gnd cell_6t
Xbit_r43_c74 bl_74 br_74 wl_43 vdd gnd cell_6t
Xbit_r44_c74 bl_74 br_74 wl_44 vdd gnd cell_6t
Xbit_r45_c74 bl_74 br_74 wl_45 vdd gnd cell_6t
Xbit_r46_c74 bl_74 br_74 wl_46 vdd gnd cell_6t
Xbit_r47_c74 bl_74 br_74 wl_47 vdd gnd cell_6t
Xbit_r48_c74 bl_74 br_74 wl_48 vdd gnd cell_6t
Xbit_r49_c74 bl_74 br_74 wl_49 vdd gnd cell_6t
Xbit_r50_c74 bl_74 br_74 wl_50 vdd gnd cell_6t
Xbit_r51_c74 bl_74 br_74 wl_51 vdd gnd cell_6t
Xbit_r52_c74 bl_74 br_74 wl_52 vdd gnd cell_6t
Xbit_r53_c74 bl_74 br_74 wl_53 vdd gnd cell_6t
Xbit_r54_c74 bl_74 br_74 wl_54 vdd gnd cell_6t
Xbit_r55_c74 bl_74 br_74 wl_55 vdd gnd cell_6t
Xbit_r56_c74 bl_74 br_74 wl_56 vdd gnd cell_6t
Xbit_r57_c74 bl_74 br_74 wl_57 vdd gnd cell_6t
Xbit_r58_c74 bl_74 br_74 wl_58 vdd gnd cell_6t
Xbit_r59_c74 bl_74 br_74 wl_59 vdd gnd cell_6t
Xbit_r60_c74 bl_74 br_74 wl_60 vdd gnd cell_6t
Xbit_r61_c74 bl_74 br_74 wl_61 vdd gnd cell_6t
Xbit_r62_c74 bl_74 br_74 wl_62 vdd gnd cell_6t
Xbit_r63_c74 bl_74 br_74 wl_63 vdd gnd cell_6t
Xbit_r64_c74 bl_74 br_74 wl_64 vdd gnd cell_6t
Xbit_r65_c74 bl_74 br_74 wl_65 vdd gnd cell_6t
Xbit_r66_c74 bl_74 br_74 wl_66 vdd gnd cell_6t
Xbit_r67_c74 bl_74 br_74 wl_67 vdd gnd cell_6t
Xbit_r68_c74 bl_74 br_74 wl_68 vdd gnd cell_6t
Xbit_r69_c74 bl_74 br_74 wl_69 vdd gnd cell_6t
Xbit_r70_c74 bl_74 br_74 wl_70 vdd gnd cell_6t
Xbit_r71_c74 bl_74 br_74 wl_71 vdd gnd cell_6t
Xbit_r72_c74 bl_74 br_74 wl_72 vdd gnd cell_6t
Xbit_r73_c74 bl_74 br_74 wl_73 vdd gnd cell_6t
Xbit_r74_c74 bl_74 br_74 wl_74 vdd gnd cell_6t
Xbit_r75_c74 bl_74 br_74 wl_75 vdd gnd cell_6t
Xbit_r76_c74 bl_74 br_74 wl_76 vdd gnd cell_6t
Xbit_r77_c74 bl_74 br_74 wl_77 vdd gnd cell_6t
Xbit_r78_c74 bl_74 br_74 wl_78 vdd gnd cell_6t
Xbit_r79_c74 bl_74 br_74 wl_79 vdd gnd cell_6t
Xbit_r80_c74 bl_74 br_74 wl_80 vdd gnd cell_6t
Xbit_r81_c74 bl_74 br_74 wl_81 vdd gnd cell_6t
Xbit_r82_c74 bl_74 br_74 wl_82 vdd gnd cell_6t
Xbit_r83_c74 bl_74 br_74 wl_83 vdd gnd cell_6t
Xbit_r84_c74 bl_74 br_74 wl_84 vdd gnd cell_6t
Xbit_r85_c74 bl_74 br_74 wl_85 vdd gnd cell_6t
Xbit_r86_c74 bl_74 br_74 wl_86 vdd gnd cell_6t
Xbit_r87_c74 bl_74 br_74 wl_87 vdd gnd cell_6t
Xbit_r88_c74 bl_74 br_74 wl_88 vdd gnd cell_6t
Xbit_r89_c74 bl_74 br_74 wl_89 vdd gnd cell_6t
Xbit_r90_c74 bl_74 br_74 wl_90 vdd gnd cell_6t
Xbit_r91_c74 bl_74 br_74 wl_91 vdd gnd cell_6t
Xbit_r92_c74 bl_74 br_74 wl_92 vdd gnd cell_6t
Xbit_r93_c74 bl_74 br_74 wl_93 vdd gnd cell_6t
Xbit_r94_c74 bl_74 br_74 wl_94 vdd gnd cell_6t
Xbit_r95_c74 bl_74 br_74 wl_95 vdd gnd cell_6t
Xbit_r96_c74 bl_74 br_74 wl_96 vdd gnd cell_6t
Xbit_r97_c74 bl_74 br_74 wl_97 vdd gnd cell_6t
Xbit_r98_c74 bl_74 br_74 wl_98 vdd gnd cell_6t
Xbit_r99_c74 bl_74 br_74 wl_99 vdd gnd cell_6t
Xbit_r100_c74 bl_74 br_74 wl_100 vdd gnd cell_6t
Xbit_r101_c74 bl_74 br_74 wl_101 vdd gnd cell_6t
Xbit_r102_c74 bl_74 br_74 wl_102 vdd gnd cell_6t
Xbit_r103_c74 bl_74 br_74 wl_103 vdd gnd cell_6t
Xbit_r104_c74 bl_74 br_74 wl_104 vdd gnd cell_6t
Xbit_r105_c74 bl_74 br_74 wl_105 vdd gnd cell_6t
Xbit_r106_c74 bl_74 br_74 wl_106 vdd gnd cell_6t
Xbit_r107_c74 bl_74 br_74 wl_107 vdd gnd cell_6t
Xbit_r108_c74 bl_74 br_74 wl_108 vdd gnd cell_6t
Xbit_r109_c74 bl_74 br_74 wl_109 vdd gnd cell_6t
Xbit_r110_c74 bl_74 br_74 wl_110 vdd gnd cell_6t
Xbit_r111_c74 bl_74 br_74 wl_111 vdd gnd cell_6t
Xbit_r112_c74 bl_74 br_74 wl_112 vdd gnd cell_6t
Xbit_r113_c74 bl_74 br_74 wl_113 vdd gnd cell_6t
Xbit_r114_c74 bl_74 br_74 wl_114 vdd gnd cell_6t
Xbit_r115_c74 bl_74 br_74 wl_115 vdd gnd cell_6t
Xbit_r116_c74 bl_74 br_74 wl_116 vdd gnd cell_6t
Xbit_r117_c74 bl_74 br_74 wl_117 vdd gnd cell_6t
Xbit_r118_c74 bl_74 br_74 wl_118 vdd gnd cell_6t
Xbit_r119_c74 bl_74 br_74 wl_119 vdd gnd cell_6t
Xbit_r120_c74 bl_74 br_74 wl_120 vdd gnd cell_6t
Xbit_r121_c74 bl_74 br_74 wl_121 vdd gnd cell_6t
Xbit_r122_c74 bl_74 br_74 wl_122 vdd gnd cell_6t
Xbit_r123_c74 bl_74 br_74 wl_123 vdd gnd cell_6t
Xbit_r124_c74 bl_74 br_74 wl_124 vdd gnd cell_6t
Xbit_r125_c74 bl_74 br_74 wl_125 vdd gnd cell_6t
Xbit_r126_c74 bl_74 br_74 wl_126 vdd gnd cell_6t
Xbit_r127_c74 bl_74 br_74 wl_127 vdd gnd cell_6t
Xbit_r128_c74 bl_74 br_74 wl_128 vdd gnd cell_6t
Xbit_r129_c74 bl_74 br_74 wl_129 vdd gnd cell_6t
Xbit_r130_c74 bl_74 br_74 wl_130 vdd gnd cell_6t
Xbit_r131_c74 bl_74 br_74 wl_131 vdd gnd cell_6t
Xbit_r132_c74 bl_74 br_74 wl_132 vdd gnd cell_6t
Xbit_r133_c74 bl_74 br_74 wl_133 vdd gnd cell_6t
Xbit_r134_c74 bl_74 br_74 wl_134 vdd gnd cell_6t
Xbit_r135_c74 bl_74 br_74 wl_135 vdd gnd cell_6t
Xbit_r136_c74 bl_74 br_74 wl_136 vdd gnd cell_6t
Xbit_r137_c74 bl_74 br_74 wl_137 vdd gnd cell_6t
Xbit_r138_c74 bl_74 br_74 wl_138 vdd gnd cell_6t
Xbit_r139_c74 bl_74 br_74 wl_139 vdd gnd cell_6t
Xbit_r140_c74 bl_74 br_74 wl_140 vdd gnd cell_6t
Xbit_r141_c74 bl_74 br_74 wl_141 vdd gnd cell_6t
Xbit_r142_c74 bl_74 br_74 wl_142 vdd gnd cell_6t
Xbit_r143_c74 bl_74 br_74 wl_143 vdd gnd cell_6t
Xbit_r144_c74 bl_74 br_74 wl_144 vdd gnd cell_6t
Xbit_r145_c74 bl_74 br_74 wl_145 vdd gnd cell_6t
Xbit_r146_c74 bl_74 br_74 wl_146 vdd gnd cell_6t
Xbit_r147_c74 bl_74 br_74 wl_147 vdd gnd cell_6t
Xbit_r148_c74 bl_74 br_74 wl_148 vdd gnd cell_6t
Xbit_r149_c74 bl_74 br_74 wl_149 vdd gnd cell_6t
Xbit_r150_c74 bl_74 br_74 wl_150 vdd gnd cell_6t
Xbit_r151_c74 bl_74 br_74 wl_151 vdd gnd cell_6t
Xbit_r152_c74 bl_74 br_74 wl_152 vdd gnd cell_6t
Xbit_r153_c74 bl_74 br_74 wl_153 vdd gnd cell_6t
Xbit_r154_c74 bl_74 br_74 wl_154 vdd gnd cell_6t
Xbit_r155_c74 bl_74 br_74 wl_155 vdd gnd cell_6t
Xbit_r156_c74 bl_74 br_74 wl_156 vdd gnd cell_6t
Xbit_r157_c74 bl_74 br_74 wl_157 vdd gnd cell_6t
Xbit_r158_c74 bl_74 br_74 wl_158 vdd gnd cell_6t
Xbit_r159_c74 bl_74 br_74 wl_159 vdd gnd cell_6t
Xbit_r160_c74 bl_74 br_74 wl_160 vdd gnd cell_6t
Xbit_r161_c74 bl_74 br_74 wl_161 vdd gnd cell_6t
Xbit_r162_c74 bl_74 br_74 wl_162 vdd gnd cell_6t
Xbit_r163_c74 bl_74 br_74 wl_163 vdd gnd cell_6t
Xbit_r164_c74 bl_74 br_74 wl_164 vdd gnd cell_6t
Xbit_r165_c74 bl_74 br_74 wl_165 vdd gnd cell_6t
Xbit_r166_c74 bl_74 br_74 wl_166 vdd gnd cell_6t
Xbit_r167_c74 bl_74 br_74 wl_167 vdd gnd cell_6t
Xbit_r168_c74 bl_74 br_74 wl_168 vdd gnd cell_6t
Xbit_r169_c74 bl_74 br_74 wl_169 vdd gnd cell_6t
Xbit_r170_c74 bl_74 br_74 wl_170 vdd gnd cell_6t
Xbit_r171_c74 bl_74 br_74 wl_171 vdd gnd cell_6t
Xbit_r172_c74 bl_74 br_74 wl_172 vdd gnd cell_6t
Xbit_r173_c74 bl_74 br_74 wl_173 vdd gnd cell_6t
Xbit_r174_c74 bl_74 br_74 wl_174 vdd gnd cell_6t
Xbit_r175_c74 bl_74 br_74 wl_175 vdd gnd cell_6t
Xbit_r176_c74 bl_74 br_74 wl_176 vdd gnd cell_6t
Xbit_r177_c74 bl_74 br_74 wl_177 vdd gnd cell_6t
Xbit_r178_c74 bl_74 br_74 wl_178 vdd gnd cell_6t
Xbit_r179_c74 bl_74 br_74 wl_179 vdd gnd cell_6t
Xbit_r180_c74 bl_74 br_74 wl_180 vdd gnd cell_6t
Xbit_r181_c74 bl_74 br_74 wl_181 vdd gnd cell_6t
Xbit_r182_c74 bl_74 br_74 wl_182 vdd gnd cell_6t
Xbit_r183_c74 bl_74 br_74 wl_183 vdd gnd cell_6t
Xbit_r184_c74 bl_74 br_74 wl_184 vdd gnd cell_6t
Xbit_r185_c74 bl_74 br_74 wl_185 vdd gnd cell_6t
Xbit_r186_c74 bl_74 br_74 wl_186 vdd gnd cell_6t
Xbit_r187_c74 bl_74 br_74 wl_187 vdd gnd cell_6t
Xbit_r188_c74 bl_74 br_74 wl_188 vdd gnd cell_6t
Xbit_r189_c74 bl_74 br_74 wl_189 vdd gnd cell_6t
Xbit_r190_c74 bl_74 br_74 wl_190 vdd gnd cell_6t
Xbit_r191_c74 bl_74 br_74 wl_191 vdd gnd cell_6t
Xbit_r192_c74 bl_74 br_74 wl_192 vdd gnd cell_6t
Xbit_r193_c74 bl_74 br_74 wl_193 vdd gnd cell_6t
Xbit_r194_c74 bl_74 br_74 wl_194 vdd gnd cell_6t
Xbit_r195_c74 bl_74 br_74 wl_195 vdd gnd cell_6t
Xbit_r196_c74 bl_74 br_74 wl_196 vdd gnd cell_6t
Xbit_r197_c74 bl_74 br_74 wl_197 vdd gnd cell_6t
Xbit_r198_c74 bl_74 br_74 wl_198 vdd gnd cell_6t
Xbit_r199_c74 bl_74 br_74 wl_199 vdd gnd cell_6t
Xbit_r200_c74 bl_74 br_74 wl_200 vdd gnd cell_6t
Xbit_r201_c74 bl_74 br_74 wl_201 vdd gnd cell_6t
Xbit_r202_c74 bl_74 br_74 wl_202 vdd gnd cell_6t
Xbit_r203_c74 bl_74 br_74 wl_203 vdd gnd cell_6t
Xbit_r204_c74 bl_74 br_74 wl_204 vdd gnd cell_6t
Xbit_r205_c74 bl_74 br_74 wl_205 vdd gnd cell_6t
Xbit_r206_c74 bl_74 br_74 wl_206 vdd gnd cell_6t
Xbit_r207_c74 bl_74 br_74 wl_207 vdd gnd cell_6t
Xbit_r208_c74 bl_74 br_74 wl_208 vdd gnd cell_6t
Xbit_r209_c74 bl_74 br_74 wl_209 vdd gnd cell_6t
Xbit_r210_c74 bl_74 br_74 wl_210 vdd gnd cell_6t
Xbit_r211_c74 bl_74 br_74 wl_211 vdd gnd cell_6t
Xbit_r212_c74 bl_74 br_74 wl_212 vdd gnd cell_6t
Xbit_r213_c74 bl_74 br_74 wl_213 vdd gnd cell_6t
Xbit_r214_c74 bl_74 br_74 wl_214 vdd gnd cell_6t
Xbit_r215_c74 bl_74 br_74 wl_215 vdd gnd cell_6t
Xbit_r216_c74 bl_74 br_74 wl_216 vdd gnd cell_6t
Xbit_r217_c74 bl_74 br_74 wl_217 vdd gnd cell_6t
Xbit_r218_c74 bl_74 br_74 wl_218 vdd gnd cell_6t
Xbit_r219_c74 bl_74 br_74 wl_219 vdd gnd cell_6t
Xbit_r220_c74 bl_74 br_74 wl_220 vdd gnd cell_6t
Xbit_r221_c74 bl_74 br_74 wl_221 vdd gnd cell_6t
Xbit_r222_c74 bl_74 br_74 wl_222 vdd gnd cell_6t
Xbit_r223_c74 bl_74 br_74 wl_223 vdd gnd cell_6t
Xbit_r224_c74 bl_74 br_74 wl_224 vdd gnd cell_6t
Xbit_r225_c74 bl_74 br_74 wl_225 vdd gnd cell_6t
Xbit_r226_c74 bl_74 br_74 wl_226 vdd gnd cell_6t
Xbit_r227_c74 bl_74 br_74 wl_227 vdd gnd cell_6t
Xbit_r228_c74 bl_74 br_74 wl_228 vdd gnd cell_6t
Xbit_r229_c74 bl_74 br_74 wl_229 vdd gnd cell_6t
Xbit_r230_c74 bl_74 br_74 wl_230 vdd gnd cell_6t
Xbit_r231_c74 bl_74 br_74 wl_231 vdd gnd cell_6t
Xbit_r232_c74 bl_74 br_74 wl_232 vdd gnd cell_6t
Xbit_r233_c74 bl_74 br_74 wl_233 vdd gnd cell_6t
Xbit_r234_c74 bl_74 br_74 wl_234 vdd gnd cell_6t
Xbit_r235_c74 bl_74 br_74 wl_235 vdd gnd cell_6t
Xbit_r236_c74 bl_74 br_74 wl_236 vdd gnd cell_6t
Xbit_r237_c74 bl_74 br_74 wl_237 vdd gnd cell_6t
Xbit_r238_c74 bl_74 br_74 wl_238 vdd gnd cell_6t
Xbit_r239_c74 bl_74 br_74 wl_239 vdd gnd cell_6t
Xbit_r240_c74 bl_74 br_74 wl_240 vdd gnd cell_6t
Xbit_r241_c74 bl_74 br_74 wl_241 vdd gnd cell_6t
Xbit_r242_c74 bl_74 br_74 wl_242 vdd gnd cell_6t
Xbit_r243_c74 bl_74 br_74 wl_243 vdd gnd cell_6t
Xbit_r244_c74 bl_74 br_74 wl_244 vdd gnd cell_6t
Xbit_r245_c74 bl_74 br_74 wl_245 vdd gnd cell_6t
Xbit_r246_c74 bl_74 br_74 wl_246 vdd gnd cell_6t
Xbit_r247_c74 bl_74 br_74 wl_247 vdd gnd cell_6t
Xbit_r248_c74 bl_74 br_74 wl_248 vdd gnd cell_6t
Xbit_r249_c74 bl_74 br_74 wl_249 vdd gnd cell_6t
Xbit_r250_c74 bl_74 br_74 wl_250 vdd gnd cell_6t
Xbit_r251_c74 bl_74 br_74 wl_251 vdd gnd cell_6t
Xbit_r252_c74 bl_74 br_74 wl_252 vdd gnd cell_6t
Xbit_r253_c74 bl_74 br_74 wl_253 vdd gnd cell_6t
Xbit_r254_c74 bl_74 br_74 wl_254 vdd gnd cell_6t
Xbit_r255_c74 bl_74 br_74 wl_255 vdd gnd cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd cell_6t
Xbit_r1_c75 bl_75 br_75 wl_1 vdd gnd cell_6t
Xbit_r2_c75 bl_75 br_75 wl_2 vdd gnd cell_6t
Xbit_r3_c75 bl_75 br_75 wl_3 vdd gnd cell_6t
Xbit_r4_c75 bl_75 br_75 wl_4 vdd gnd cell_6t
Xbit_r5_c75 bl_75 br_75 wl_5 vdd gnd cell_6t
Xbit_r6_c75 bl_75 br_75 wl_6 vdd gnd cell_6t
Xbit_r7_c75 bl_75 br_75 wl_7 vdd gnd cell_6t
Xbit_r8_c75 bl_75 br_75 wl_8 vdd gnd cell_6t
Xbit_r9_c75 bl_75 br_75 wl_9 vdd gnd cell_6t
Xbit_r10_c75 bl_75 br_75 wl_10 vdd gnd cell_6t
Xbit_r11_c75 bl_75 br_75 wl_11 vdd gnd cell_6t
Xbit_r12_c75 bl_75 br_75 wl_12 vdd gnd cell_6t
Xbit_r13_c75 bl_75 br_75 wl_13 vdd gnd cell_6t
Xbit_r14_c75 bl_75 br_75 wl_14 vdd gnd cell_6t
Xbit_r15_c75 bl_75 br_75 wl_15 vdd gnd cell_6t
Xbit_r16_c75 bl_75 br_75 wl_16 vdd gnd cell_6t
Xbit_r17_c75 bl_75 br_75 wl_17 vdd gnd cell_6t
Xbit_r18_c75 bl_75 br_75 wl_18 vdd gnd cell_6t
Xbit_r19_c75 bl_75 br_75 wl_19 vdd gnd cell_6t
Xbit_r20_c75 bl_75 br_75 wl_20 vdd gnd cell_6t
Xbit_r21_c75 bl_75 br_75 wl_21 vdd gnd cell_6t
Xbit_r22_c75 bl_75 br_75 wl_22 vdd gnd cell_6t
Xbit_r23_c75 bl_75 br_75 wl_23 vdd gnd cell_6t
Xbit_r24_c75 bl_75 br_75 wl_24 vdd gnd cell_6t
Xbit_r25_c75 bl_75 br_75 wl_25 vdd gnd cell_6t
Xbit_r26_c75 bl_75 br_75 wl_26 vdd gnd cell_6t
Xbit_r27_c75 bl_75 br_75 wl_27 vdd gnd cell_6t
Xbit_r28_c75 bl_75 br_75 wl_28 vdd gnd cell_6t
Xbit_r29_c75 bl_75 br_75 wl_29 vdd gnd cell_6t
Xbit_r30_c75 bl_75 br_75 wl_30 vdd gnd cell_6t
Xbit_r31_c75 bl_75 br_75 wl_31 vdd gnd cell_6t
Xbit_r32_c75 bl_75 br_75 wl_32 vdd gnd cell_6t
Xbit_r33_c75 bl_75 br_75 wl_33 vdd gnd cell_6t
Xbit_r34_c75 bl_75 br_75 wl_34 vdd gnd cell_6t
Xbit_r35_c75 bl_75 br_75 wl_35 vdd gnd cell_6t
Xbit_r36_c75 bl_75 br_75 wl_36 vdd gnd cell_6t
Xbit_r37_c75 bl_75 br_75 wl_37 vdd gnd cell_6t
Xbit_r38_c75 bl_75 br_75 wl_38 vdd gnd cell_6t
Xbit_r39_c75 bl_75 br_75 wl_39 vdd gnd cell_6t
Xbit_r40_c75 bl_75 br_75 wl_40 vdd gnd cell_6t
Xbit_r41_c75 bl_75 br_75 wl_41 vdd gnd cell_6t
Xbit_r42_c75 bl_75 br_75 wl_42 vdd gnd cell_6t
Xbit_r43_c75 bl_75 br_75 wl_43 vdd gnd cell_6t
Xbit_r44_c75 bl_75 br_75 wl_44 vdd gnd cell_6t
Xbit_r45_c75 bl_75 br_75 wl_45 vdd gnd cell_6t
Xbit_r46_c75 bl_75 br_75 wl_46 vdd gnd cell_6t
Xbit_r47_c75 bl_75 br_75 wl_47 vdd gnd cell_6t
Xbit_r48_c75 bl_75 br_75 wl_48 vdd gnd cell_6t
Xbit_r49_c75 bl_75 br_75 wl_49 vdd gnd cell_6t
Xbit_r50_c75 bl_75 br_75 wl_50 vdd gnd cell_6t
Xbit_r51_c75 bl_75 br_75 wl_51 vdd gnd cell_6t
Xbit_r52_c75 bl_75 br_75 wl_52 vdd gnd cell_6t
Xbit_r53_c75 bl_75 br_75 wl_53 vdd gnd cell_6t
Xbit_r54_c75 bl_75 br_75 wl_54 vdd gnd cell_6t
Xbit_r55_c75 bl_75 br_75 wl_55 vdd gnd cell_6t
Xbit_r56_c75 bl_75 br_75 wl_56 vdd gnd cell_6t
Xbit_r57_c75 bl_75 br_75 wl_57 vdd gnd cell_6t
Xbit_r58_c75 bl_75 br_75 wl_58 vdd gnd cell_6t
Xbit_r59_c75 bl_75 br_75 wl_59 vdd gnd cell_6t
Xbit_r60_c75 bl_75 br_75 wl_60 vdd gnd cell_6t
Xbit_r61_c75 bl_75 br_75 wl_61 vdd gnd cell_6t
Xbit_r62_c75 bl_75 br_75 wl_62 vdd gnd cell_6t
Xbit_r63_c75 bl_75 br_75 wl_63 vdd gnd cell_6t
Xbit_r64_c75 bl_75 br_75 wl_64 vdd gnd cell_6t
Xbit_r65_c75 bl_75 br_75 wl_65 vdd gnd cell_6t
Xbit_r66_c75 bl_75 br_75 wl_66 vdd gnd cell_6t
Xbit_r67_c75 bl_75 br_75 wl_67 vdd gnd cell_6t
Xbit_r68_c75 bl_75 br_75 wl_68 vdd gnd cell_6t
Xbit_r69_c75 bl_75 br_75 wl_69 vdd gnd cell_6t
Xbit_r70_c75 bl_75 br_75 wl_70 vdd gnd cell_6t
Xbit_r71_c75 bl_75 br_75 wl_71 vdd gnd cell_6t
Xbit_r72_c75 bl_75 br_75 wl_72 vdd gnd cell_6t
Xbit_r73_c75 bl_75 br_75 wl_73 vdd gnd cell_6t
Xbit_r74_c75 bl_75 br_75 wl_74 vdd gnd cell_6t
Xbit_r75_c75 bl_75 br_75 wl_75 vdd gnd cell_6t
Xbit_r76_c75 bl_75 br_75 wl_76 vdd gnd cell_6t
Xbit_r77_c75 bl_75 br_75 wl_77 vdd gnd cell_6t
Xbit_r78_c75 bl_75 br_75 wl_78 vdd gnd cell_6t
Xbit_r79_c75 bl_75 br_75 wl_79 vdd gnd cell_6t
Xbit_r80_c75 bl_75 br_75 wl_80 vdd gnd cell_6t
Xbit_r81_c75 bl_75 br_75 wl_81 vdd gnd cell_6t
Xbit_r82_c75 bl_75 br_75 wl_82 vdd gnd cell_6t
Xbit_r83_c75 bl_75 br_75 wl_83 vdd gnd cell_6t
Xbit_r84_c75 bl_75 br_75 wl_84 vdd gnd cell_6t
Xbit_r85_c75 bl_75 br_75 wl_85 vdd gnd cell_6t
Xbit_r86_c75 bl_75 br_75 wl_86 vdd gnd cell_6t
Xbit_r87_c75 bl_75 br_75 wl_87 vdd gnd cell_6t
Xbit_r88_c75 bl_75 br_75 wl_88 vdd gnd cell_6t
Xbit_r89_c75 bl_75 br_75 wl_89 vdd gnd cell_6t
Xbit_r90_c75 bl_75 br_75 wl_90 vdd gnd cell_6t
Xbit_r91_c75 bl_75 br_75 wl_91 vdd gnd cell_6t
Xbit_r92_c75 bl_75 br_75 wl_92 vdd gnd cell_6t
Xbit_r93_c75 bl_75 br_75 wl_93 vdd gnd cell_6t
Xbit_r94_c75 bl_75 br_75 wl_94 vdd gnd cell_6t
Xbit_r95_c75 bl_75 br_75 wl_95 vdd gnd cell_6t
Xbit_r96_c75 bl_75 br_75 wl_96 vdd gnd cell_6t
Xbit_r97_c75 bl_75 br_75 wl_97 vdd gnd cell_6t
Xbit_r98_c75 bl_75 br_75 wl_98 vdd gnd cell_6t
Xbit_r99_c75 bl_75 br_75 wl_99 vdd gnd cell_6t
Xbit_r100_c75 bl_75 br_75 wl_100 vdd gnd cell_6t
Xbit_r101_c75 bl_75 br_75 wl_101 vdd gnd cell_6t
Xbit_r102_c75 bl_75 br_75 wl_102 vdd gnd cell_6t
Xbit_r103_c75 bl_75 br_75 wl_103 vdd gnd cell_6t
Xbit_r104_c75 bl_75 br_75 wl_104 vdd gnd cell_6t
Xbit_r105_c75 bl_75 br_75 wl_105 vdd gnd cell_6t
Xbit_r106_c75 bl_75 br_75 wl_106 vdd gnd cell_6t
Xbit_r107_c75 bl_75 br_75 wl_107 vdd gnd cell_6t
Xbit_r108_c75 bl_75 br_75 wl_108 vdd gnd cell_6t
Xbit_r109_c75 bl_75 br_75 wl_109 vdd gnd cell_6t
Xbit_r110_c75 bl_75 br_75 wl_110 vdd gnd cell_6t
Xbit_r111_c75 bl_75 br_75 wl_111 vdd gnd cell_6t
Xbit_r112_c75 bl_75 br_75 wl_112 vdd gnd cell_6t
Xbit_r113_c75 bl_75 br_75 wl_113 vdd gnd cell_6t
Xbit_r114_c75 bl_75 br_75 wl_114 vdd gnd cell_6t
Xbit_r115_c75 bl_75 br_75 wl_115 vdd gnd cell_6t
Xbit_r116_c75 bl_75 br_75 wl_116 vdd gnd cell_6t
Xbit_r117_c75 bl_75 br_75 wl_117 vdd gnd cell_6t
Xbit_r118_c75 bl_75 br_75 wl_118 vdd gnd cell_6t
Xbit_r119_c75 bl_75 br_75 wl_119 vdd gnd cell_6t
Xbit_r120_c75 bl_75 br_75 wl_120 vdd gnd cell_6t
Xbit_r121_c75 bl_75 br_75 wl_121 vdd gnd cell_6t
Xbit_r122_c75 bl_75 br_75 wl_122 vdd gnd cell_6t
Xbit_r123_c75 bl_75 br_75 wl_123 vdd gnd cell_6t
Xbit_r124_c75 bl_75 br_75 wl_124 vdd gnd cell_6t
Xbit_r125_c75 bl_75 br_75 wl_125 vdd gnd cell_6t
Xbit_r126_c75 bl_75 br_75 wl_126 vdd gnd cell_6t
Xbit_r127_c75 bl_75 br_75 wl_127 vdd gnd cell_6t
Xbit_r128_c75 bl_75 br_75 wl_128 vdd gnd cell_6t
Xbit_r129_c75 bl_75 br_75 wl_129 vdd gnd cell_6t
Xbit_r130_c75 bl_75 br_75 wl_130 vdd gnd cell_6t
Xbit_r131_c75 bl_75 br_75 wl_131 vdd gnd cell_6t
Xbit_r132_c75 bl_75 br_75 wl_132 vdd gnd cell_6t
Xbit_r133_c75 bl_75 br_75 wl_133 vdd gnd cell_6t
Xbit_r134_c75 bl_75 br_75 wl_134 vdd gnd cell_6t
Xbit_r135_c75 bl_75 br_75 wl_135 vdd gnd cell_6t
Xbit_r136_c75 bl_75 br_75 wl_136 vdd gnd cell_6t
Xbit_r137_c75 bl_75 br_75 wl_137 vdd gnd cell_6t
Xbit_r138_c75 bl_75 br_75 wl_138 vdd gnd cell_6t
Xbit_r139_c75 bl_75 br_75 wl_139 vdd gnd cell_6t
Xbit_r140_c75 bl_75 br_75 wl_140 vdd gnd cell_6t
Xbit_r141_c75 bl_75 br_75 wl_141 vdd gnd cell_6t
Xbit_r142_c75 bl_75 br_75 wl_142 vdd gnd cell_6t
Xbit_r143_c75 bl_75 br_75 wl_143 vdd gnd cell_6t
Xbit_r144_c75 bl_75 br_75 wl_144 vdd gnd cell_6t
Xbit_r145_c75 bl_75 br_75 wl_145 vdd gnd cell_6t
Xbit_r146_c75 bl_75 br_75 wl_146 vdd gnd cell_6t
Xbit_r147_c75 bl_75 br_75 wl_147 vdd gnd cell_6t
Xbit_r148_c75 bl_75 br_75 wl_148 vdd gnd cell_6t
Xbit_r149_c75 bl_75 br_75 wl_149 vdd gnd cell_6t
Xbit_r150_c75 bl_75 br_75 wl_150 vdd gnd cell_6t
Xbit_r151_c75 bl_75 br_75 wl_151 vdd gnd cell_6t
Xbit_r152_c75 bl_75 br_75 wl_152 vdd gnd cell_6t
Xbit_r153_c75 bl_75 br_75 wl_153 vdd gnd cell_6t
Xbit_r154_c75 bl_75 br_75 wl_154 vdd gnd cell_6t
Xbit_r155_c75 bl_75 br_75 wl_155 vdd gnd cell_6t
Xbit_r156_c75 bl_75 br_75 wl_156 vdd gnd cell_6t
Xbit_r157_c75 bl_75 br_75 wl_157 vdd gnd cell_6t
Xbit_r158_c75 bl_75 br_75 wl_158 vdd gnd cell_6t
Xbit_r159_c75 bl_75 br_75 wl_159 vdd gnd cell_6t
Xbit_r160_c75 bl_75 br_75 wl_160 vdd gnd cell_6t
Xbit_r161_c75 bl_75 br_75 wl_161 vdd gnd cell_6t
Xbit_r162_c75 bl_75 br_75 wl_162 vdd gnd cell_6t
Xbit_r163_c75 bl_75 br_75 wl_163 vdd gnd cell_6t
Xbit_r164_c75 bl_75 br_75 wl_164 vdd gnd cell_6t
Xbit_r165_c75 bl_75 br_75 wl_165 vdd gnd cell_6t
Xbit_r166_c75 bl_75 br_75 wl_166 vdd gnd cell_6t
Xbit_r167_c75 bl_75 br_75 wl_167 vdd gnd cell_6t
Xbit_r168_c75 bl_75 br_75 wl_168 vdd gnd cell_6t
Xbit_r169_c75 bl_75 br_75 wl_169 vdd gnd cell_6t
Xbit_r170_c75 bl_75 br_75 wl_170 vdd gnd cell_6t
Xbit_r171_c75 bl_75 br_75 wl_171 vdd gnd cell_6t
Xbit_r172_c75 bl_75 br_75 wl_172 vdd gnd cell_6t
Xbit_r173_c75 bl_75 br_75 wl_173 vdd gnd cell_6t
Xbit_r174_c75 bl_75 br_75 wl_174 vdd gnd cell_6t
Xbit_r175_c75 bl_75 br_75 wl_175 vdd gnd cell_6t
Xbit_r176_c75 bl_75 br_75 wl_176 vdd gnd cell_6t
Xbit_r177_c75 bl_75 br_75 wl_177 vdd gnd cell_6t
Xbit_r178_c75 bl_75 br_75 wl_178 vdd gnd cell_6t
Xbit_r179_c75 bl_75 br_75 wl_179 vdd gnd cell_6t
Xbit_r180_c75 bl_75 br_75 wl_180 vdd gnd cell_6t
Xbit_r181_c75 bl_75 br_75 wl_181 vdd gnd cell_6t
Xbit_r182_c75 bl_75 br_75 wl_182 vdd gnd cell_6t
Xbit_r183_c75 bl_75 br_75 wl_183 vdd gnd cell_6t
Xbit_r184_c75 bl_75 br_75 wl_184 vdd gnd cell_6t
Xbit_r185_c75 bl_75 br_75 wl_185 vdd gnd cell_6t
Xbit_r186_c75 bl_75 br_75 wl_186 vdd gnd cell_6t
Xbit_r187_c75 bl_75 br_75 wl_187 vdd gnd cell_6t
Xbit_r188_c75 bl_75 br_75 wl_188 vdd gnd cell_6t
Xbit_r189_c75 bl_75 br_75 wl_189 vdd gnd cell_6t
Xbit_r190_c75 bl_75 br_75 wl_190 vdd gnd cell_6t
Xbit_r191_c75 bl_75 br_75 wl_191 vdd gnd cell_6t
Xbit_r192_c75 bl_75 br_75 wl_192 vdd gnd cell_6t
Xbit_r193_c75 bl_75 br_75 wl_193 vdd gnd cell_6t
Xbit_r194_c75 bl_75 br_75 wl_194 vdd gnd cell_6t
Xbit_r195_c75 bl_75 br_75 wl_195 vdd gnd cell_6t
Xbit_r196_c75 bl_75 br_75 wl_196 vdd gnd cell_6t
Xbit_r197_c75 bl_75 br_75 wl_197 vdd gnd cell_6t
Xbit_r198_c75 bl_75 br_75 wl_198 vdd gnd cell_6t
Xbit_r199_c75 bl_75 br_75 wl_199 vdd gnd cell_6t
Xbit_r200_c75 bl_75 br_75 wl_200 vdd gnd cell_6t
Xbit_r201_c75 bl_75 br_75 wl_201 vdd gnd cell_6t
Xbit_r202_c75 bl_75 br_75 wl_202 vdd gnd cell_6t
Xbit_r203_c75 bl_75 br_75 wl_203 vdd gnd cell_6t
Xbit_r204_c75 bl_75 br_75 wl_204 vdd gnd cell_6t
Xbit_r205_c75 bl_75 br_75 wl_205 vdd gnd cell_6t
Xbit_r206_c75 bl_75 br_75 wl_206 vdd gnd cell_6t
Xbit_r207_c75 bl_75 br_75 wl_207 vdd gnd cell_6t
Xbit_r208_c75 bl_75 br_75 wl_208 vdd gnd cell_6t
Xbit_r209_c75 bl_75 br_75 wl_209 vdd gnd cell_6t
Xbit_r210_c75 bl_75 br_75 wl_210 vdd gnd cell_6t
Xbit_r211_c75 bl_75 br_75 wl_211 vdd gnd cell_6t
Xbit_r212_c75 bl_75 br_75 wl_212 vdd gnd cell_6t
Xbit_r213_c75 bl_75 br_75 wl_213 vdd gnd cell_6t
Xbit_r214_c75 bl_75 br_75 wl_214 vdd gnd cell_6t
Xbit_r215_c75 bl_75 br_75 wl_215 vdd gnd cell_6t
Xbit_r216_c75 bl_75 br_75 wl_216 vdd gnd cell_6t
Xbit_r217_c75 bl_75 br_75 wl_217 vdd gnd cell_6t
Xbit_r218_c75 bl_75 br_75 wl_218 vdd gnd cell_6t
Xbit_r219_c75 bl_75 br_75 wl_219 vdd gnd cell_6t
Xbit_r220_c75 bl_75 br_75 wl_220 vdd gnd cell_6t
Xbit_r221_c75 bl_75 br_75 wl_221 vdd gnd cell_6t
Xbit_r222_c75 bl_75 br_75 wl_222 vdd gnd cell_6t
Xbit_r223_c75 bl_75 br_75 wl_223 vdd gnd cell_6t
Xbit_r224_c75 bl_75 br_75 wl_224 vdd gnd cell_6t
Xbit_r225_c75 bl_75 br_75 wl_225 vdd gnd cell_6t
Xbit_r226_c75 bl_75 br_75 wl_226 vdd gnd cell_6t
Xbit_r227_c75 bl_75 br_75 wl_227 vdd gnd cell_6t
Xbit_r228_c75 bl_75 br_75 wl_228 vdd gnd cell_6t
Xbit_r229_c75 bl_75 br_75 wl_229 vdd gnd cell_6t
Xbit_r230_c75 bl_75 br_75 wl_230 vdd gnd cell_6t
Xbit_r231_c75 bl_75 br_75 wl_231 vdd gnd cell_6t
Xbit_r232_c75 bl_75 br_75 wl_232 vdd gnd cell_6t
Xbit_r233_c75 bl_75 br_75 wl_233 vdd gnd cell_6t
Xbit_r234_c75 bl_75 br_75 wl_234 vdd gnd cell_6t
Xbit_r235_c75 bl_75 br_75 wl_235 vdd gnd cell_6t
Xbit_r236_c75 bl_75 br_75 wl_236 vdd gnd cell_6t
Xbit_r237_c75 bl_75 br_75 wl_237 vdd gnd cell_6t
Xbit_r238_c75 bl_75 br_75 wl_238 vdd gnd cell_6t
Xbit_r239_c75 bl_75 br_75 wl_239 vdd gnd cell_6t
Xbit_r240_c75 bl_75 br_75 wl_240 vdd gnd cell_6t
Xbit_r241_c75 bl_75 br_75 wl_241 vdd gnd cell_6t
Xbit_r242_c75 bl_75 br_75 wl_242 vdd gnd cell_6t
Xbit_r243_c75 bl_75 br_75 wl_243 vdd gnd cell_6t
Xbit_r244_c75 bl_75 br_75 wl_244 vdd gnd cell_6t
Xbit_r245_c75 bl_75 br_75 wl_245 vdd gnd cell_6t
Xbit_r246_c75 bl_75 br_75 wl_246 vdd gnd cell_6t
Xbit_r247_c75 bl_75 br_75 wl_247 vdd gnd cell_6t
Xbit_r248_c75 bl_75 br_75 wl_248 vdd gnd cell_6t
Xbit_r249_c75 bl_75 br_75 wl_249 vdd gnd cell_6t
Xbit_r250_c75 bl_75 br_75 wl_250 vdd gnd cell_6t
Xbit_r251_c75 bl_75 br_75 wl_251 vdd gnd cell_6t
Xbit_r252_c75 bl_75 br_75 wl_252 vdd gnd cell_6t
Xbit_r253_c75 bl_75 br_75 wl_253 vdd gnd cell_6t
Xbit_r254_c75 bl_75 br_75 wl_254 vdd gnd cell_6t
Xbit_r255_c75 bl_75 br_75 wl_255 vdd gnd cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd cell_6t
Xbit_r1_c76 bl_76 br_76 wl_1 vdd gnd cell_6t
Xbit_r2_c76 bl_76 br_76 wl_2 vdd gnd cell_6t
Xbit_r3_c76 bl_76 br_76 wl_3 vdd gnd cell_6t
Xbit_r4_c76 bl_76 br_76 wl_4 vdd gnd cell_6t
Xbit_r5_c76 bl_76 br_76 wl_5 vdd gnd cell_6t
Xbit_r6_c76 bl_76 br_76 wl_6 vdd gnd cell_6t
Xbit_r7_c76 bl_76 br_76 wl_7 vdd gnd cell_6t
Xbit_r8_c76 bl_76 br_76 wl_8 vdd gnd cell_6t
Xbit_r9_c76 bl_76 br_76 wl_9 vdd gnd cell_6t
Xbit_r10_c76 bl_76 br_76 wl_10 vdd gnd cell_6t
Xbit_r11_c76 bl_76 br_76 wl_11 vdd gnd cell_6t
Xbit_r12_c76 bl_76 br_76 wl_12 vdd gnd cell_6t
Xbit_r13_c76 bl_76 br_76 wl_13 vdd gnd cell_6t
Xbit_r14_c76 bl_76 br_76 wl_14 vdd gnd cell_6t
Xbit_r15_c76 bl_76 br_76 wl_15 vdd gnd cell_6t
Xbit_r16_c76 bl_76 br_76 wl_16 vdd gnd cell_6t
Xbit_r17_c76 bl_76 br_76 wl_17 vdd gnd cell_6t
Xbit_r18_c76 bl_76 br_76 wl_18 vdd gnd cell_6t
Xbit_r19_c76 bl_76 br_76 wl_19 vdd gnd cell_6t
Xbit_r20_c76 bl_76 br_76 wl_20 vdd gnd cell_6t
Xbit_r21_c76 bl_76 br_76 wl_21 vdd gnd cell_6t
Xbit_r22_c76 bl_76 br_76 wl_22 vdd gnd cell_6t
Xbit_r23_c76 bl_76 br_76 wl_23 vdd gnd cell_6t
Xbit_r24_c76 bl_76 br_76 wl_24 vdd gnd cell_6t
Xbit_r25_c76 bl_76 br_76 wl_25 vdd gnd cell_6t
Xbit_r26_c76 bl_76 br_76 wl_26 vdd gnd cell_6t
Xbit_r27_c76 bl_76 br_76 wl_27 vdd gnd cell_6t
Xbit_r28_c76 bl_76 br_76 wl_28 vdd gnd cell_6t
Xbit_r29_c76 bl_76 br_76 wl_29 vdd gnd cell_6t
Xbit_r30_c76 bl_76 br_76 wl_30 vdd gnd cell_6t
Xbit_r31_c76 bl_76 br_76 wl_31 vdd gnd cell_6t
Xbit_r32_c76 bl_76 br_76 wl_32 vdd gnd cell_6t
Xbit_r33_c76 bl_76 br_76 wl_33 vdd gnd cell_6t
Xbit_r34_c76 bl_76 br_76 wl_34 vdd gnd cell_6t
Xbit_r35_c76 bl_76 br_76 wl_35 vdd gnd cell_6t
Xbit_r36_c76 bl_76 br_76 wl_36 vdd gnd cell_6t
Xbit_r37_c76 bl_76 br_76 wl_37 vdd gnd cell_6t
Xbit_r38_c76 bl_76 br_76 wl_38 vdd gnd cell_6t
Xbit_r39_c76 bl_76 br_76 wl_39 vdd gnd cell_6t
Xbit_r40_c76 bl_76 br_76 wl_40 vdd gnd cell_6t
Xbit_r41_c76 bl_76 br_76 wl_41 vdd gnd cell_6t
Xbit_r42_c76 bl_76 br_76 wl_42 vdd gnd cell_6t
Xbit_r43_c76 bl_76 br_76 wl_43 vdd gnd cell_6t
Xbit_r44_c76 bl_76 br_76 wl_44 vdd gnd cell_6t
Xbit_r45_c76 bl_76 br_76 wl_45 vdd gnd cell_6t
Xbit_r46_c76 bl_76 br_76 wl_46 vdd gnd cell_6t
Xbit_r47_c76 bl_76 br_76 wl_47 vdd gnd cell_6t
Xbit_r48_c76 bl_76 br_76 wl_48 vdd gnd cell_6t
Xbit_r49_c76 bl_76 br_76 wl_49 vdd gnd cell_6t
Xbit_r50_c76 bl_76 br_76 wl_50 vdd gnd cell_6t
Xbit_r51_c76 bl_76 br_76 wl_51 vdd gnd cell_6t
Xbit_r52_c76 bl_76 br_76 wl_52 vdd gnd cell_6t
Xbit_r53_c76 bl_76 br_76 wl_53 vdd gnd cell_6t
Xbit_r54_c76 bl_76 br_76 wl_54 vdd gnd cell_6t
Xbit_r55_c76 bl_76 br_76 wl_55 vdd gnd cell_6t
Xbit_r56_c76 bl_76 br_76 wl_56 vdd gnd cell_6t
Xbit_r57_c76 bl_76 br_76 wl_57 vdd gnd cell_6t
Xbit_r58_c76 bl_76 br_76 wl_58 vdd gnd cell_6t
Xbit_r59_c76 bl_76 br_76 wl_59 vdd gnd cell_6t
Xbit_r60_c76 bl_76 br_76 wl_60 vdd gnd cell_6t
Xbit_r61_c76 bl_76 br_76 wl_61 vdd gnd cell_6t
Xbit_r62_c76 bl_76 br_76 wl_62 vdd gnd cell_6t
Xbit_r63_c76 bl_76 br_76 wl_63 vdd gnd cell_6t
Xbit_r64_c76 bl_76 br_76 wl_64 vdd gnd cell_6t
Xbit_r65_c76 bl_76 br_76 wl_65 vdd gnd cell_6t
Xbit_r66_c76 bl_76 br_76 wl_66 vdd gnd cell_6t
Xbit_r67_c76 bl_76 br_76 wl_67 vdd gnd cell_6t
Xbit_r68_c76 bl_76 br_76 wl_68 vdd gnd cell_6t
Xbit_r69_c76 bl_76 br_76 wl_69 vdd gnd cell_6t
Xbit_r70_c76 bl_76 br_76 wl_70 vdd gnd cell_6t
Xbit_r71_c76 bl_76 br_76 wl_71 vdd gnd cell_6t
Xbit_r72_c76 bl_76 br_76 wl_72 vdd gnd cell_6t
Xbit_r73_c76 bl_76 br_76 wl_73 vdd gnd cell_6t
Xbit_r74_c76 bl_76 br_76 wl_74 vdd gnd cell_6t
Xbit_r75_c76 bl_76 br_76 wl_75 vdd gnd cell_6t
Xbit_r76_c76 bl_76 br_76 wl_76 vdd gnd cell_6t
Xbit_r77_c76 bl_76 br_76 wl_77 vdd gnd cell_6t
Xbit_r78_c76 bl_76 br_76 wl_78 vdd gnd cell_6t
Xbit_r79_c76 bl_76 br_76 wl_79 vdd gnd cell_6t
Xbit_r80_c76 bl_76 br_76 wl_80 vdd gnd cell_6t
Xbit_r81_c76 bl_76 br_76 wl_81 vdd gnd cell_6t
Xbit_r82_c76 bl_76 br_76 wl_82 vdd gnd cell_6t
Xbit_r83_c76 bl_76 br_76 wl_83 vdd gnd cell_6t
Xbit_r84_c76 bl_76 br_76 wl_84 vdd gnd cell_6t
Xbit_r85_c76 bl_76 br_76 wl_85 vdd gnd cell_6t
Xbit_r86_c76 bl_76 br_76 wl_86 vdd gnd cell_6t
Xbit_r87_c76 bl_76 br_76 wl_87 vdd gnd cell_6t
Xbit_r88_c76 bl_76 br_76 wl_88 vdd gnd cell_6t
Xbit_r89_c76 bl_76 br_76 wl_89 vdd gnd cell_6t
Xbit_r90_c76 bl_76 br_76 wl_90 vdd gnd cell_6t
Xbit_r91_c76 bl_76 br_76 wl_91 vdd gnd cell_6t
Xbit_r92_c76 bl_76 br_76 wl_92 vdd gnd cell_6t
Xbit_r93_c76 bl_76 br_76 wl_93 vdd gnd cell_6t
Xbit_r94_c76 bl_76 br_76 wl_94 vdd gnd cell_6t
Xbit_r95_c76 bl_76 br_76 wl_95 vdd gnd cell_6t
Xbit_r96_c76 bl_76 br_76 wl_96 vdd gnd cell_6t
Xbit_r97_c76 bl_76 br_76 wl_97 vdd gnd cell_6t
Xbit_r98_c76 bl_76 br_76 wl_98 vdd gnd cell_6t
Xbit_r99_c76 bl_76 br_76 wl_99 vdd gnd cell_6t
Xbit_r100_c76 bl_76 br_76 wl_100 vdd gnd cell_6t
Xbit_r101_c76 bl_76 br_76 wl_101 vdd gnd cell_6t
Xbit_r102_c76 bl_76 br_76 wl_102 vdd gnd cell_6t
Xbit_r103_c76 bl_76 br_76 wl_103 vdd gnd cell_6t
Xbit_r104_c76 bl_76 br_76 wl_104 vdd gnd cell_6t
Xbit_r105_c76 bl_76 br_76 wl_105 vdd gnd cell_6t
Xbit_r106_c76 bl_76 br_76 wl_106 vdd gnd cell_6t
Xbit_r107_c76 bl_76 br_76 wl_107 vdd gnd cell_6t
Xbit_r108_c76 bl_76 br_76 wl_108 vdd gnd cell_6t
Xbit_r109_c76 bl_76 br_76 wl_109 vdd gnd cell_6t
Xbit_r110_c76 bl_76 br_76 wl_110 vdd gnd cell_6t
Xbit_r111_c76 bl_76 br_76 wl_111 vdd gnd cell_6t
Xbit_r112_c76 bl_76 br_76 wl_112 vdd gnd cell_6t
Xbit_r113_c76 bl_76 br_76 wl_113 vdd gnd cell_6t
Xbit_r114_c76 bl_76 br_76 wl_114 vdd gnd cell_6t
Xbit_r115_c76 bl_76 br_76 wl_115 vdd gnd cell_6t
Xbit_r116_c76 bl_76 br_76 wl_116 vdd gnd cell_6t
Xbit_r117_c76 bl_76 br_76 wl_117 vdd gnd cell_6t
Xbit_r118_c76 bl_76 br_76 wl_118 vdd gnd cell_6t
Xbit_r119_c76 bl_76 br_76 wl_119 vdd gnd cell_6t
Xbit_r120_c76 bl_76 br_76 wl_120 vdd gnd cell_6t
Xbit_r121_c76 bl_76 br_76 wl_121 vdd gnd cell_6t
Xbit_r122_c76 bl_76 br_76 wl_122 vdd gnd cell_6t
Xbit_r123_c76 bl_76 br_76 wl_123 vdd gnd cell_6t
Xbit_r124_c76 bl_76 br_76 wl_124 vdd gnd cell_6t
Xbit_r125_c76 bl_76 br_76 wl_125 vdd gnd cell_6t
Xbit_r126_c76 bl_76 br_76 wl_126 vdd gnd cell_6t
Xbit_r127_c76 bl_76 br_76 wl_127 vdd gnd cell_6t
Xbit_r128_c76 bl_76 br_76 wl_128 vdd gnd cell_6t
Xbit_r129_c76 bl_76 br_76 wl_129 vdd gnd cell_6t
Xbit_r130_c76 bl_76 br_76 wl_130 vdd gnd cell_6t
Xbit_r131_c76 bl_76 br_76 wl_131 vdd gnd cell_6t
Xbit_r132_c76 bl_76 br_76 wl_132 vdd gnd cell_6t
Xbit_r133_c76 bl_76 br_76 wl_133 vdd gnd cell_6t
Xbit_r134_c76 bl_76 br_76 wl_134 vdd gnd cell_6t
Xbit_r135_c76 bl_76 br_76 wl_135 vdd gnd cell_6t
Xbit_r136_c76 bl_76 br_76 wl_136 vdd gnd cell_6t
Xbit_r137_c76 bl_76 br_76 wl_137 vdd gnd cell_6t
Xbit_r138_c76 bl_76 br_76 wl_138 vdd gnd cell_6t
Xbit_r139_c76 bl_76 br_76 wl_139 vdd gnd cell_6t
Xbit_r140_c76 bl_76 br_76 wl_140 vdd gnd cell_6t
Xbit_r141_c76 bl_76 br_76 wl_141 vdd gnd cell_6t
Xbit_r142_c76 bl_76 br_76 wl_142 vdd gnd cell_6t
Xbit_r143_c76 bl_76 br_76 wl_143 vdd gnd cell_6t
Xbit_r144_c76 bl_76 br_76 wl_144 vdd gnd cell_6t
Xbit_r145_c76 bl_76 br_76 wl_145 vdd gnd cell_6t
Xbit_r146_c76 bl_76 br_76 wl_146 vdd gnd cell_6t
Xbit_r147_c76 bl_76 br_76 wl_147 vdd gnd cell_6t
Xbit_r148_c76 bl_76 br_76 wl_148 vdd gnd cell_6t
Xbit_r149_c76 bl_76 br_76 wl_149 vdd gnd cell_6t
Xbit_r150_c76 bl_76 br_76 wl_150 vdd gnd cell_6t
Xbit_r151_c76 bl_76 br_76 wl_151 vdd gnd cell_6t
Xbit_r152_c76 bl_76 br_76 wl_152 vdd gnd cell_6t
Xbit_r153_c76 bl_76 br_76 wl_153 vdd gnd cell_6t
Xbit_r154_c76 bl_76 br_76 wl_154 vdd gnd cell_6t
Xbit_r155_c76 bl_76 br_76 wl_155 vdd gnd cell_6t
Xbit_r156_c76 bl_76 br_76 wl_156 vdd gnd cell_6t
Xbit_r157_c76 bl_76 br_76 wl_157 vdd gnd cell_6t
Xbit_r158_c76 bl_76 br_76 wl_158 vdd gnd cell_6t
Xbit_r159_c76 bl_76 br_76 wl_159 vdd gnd cell_6t
Xbit_r160_c76 bl_76 br_76 wl_160 vdd gnd cell_6t
Xbit_r161_c76 bl_76 br_76 wl_161 vdd gnd cell_6t
Xbit_r162_c76 bl_76 br_76 wl_162 vdd gnd cell_6t
Xbit_r163_c76 bl_76 br_76 wl_163 vdd gnd cell_6t
Xbit_r164_c76 bl_76 br_76 wl_164 vdd gnd cell_6t
Xbit_r165_c76 bl_76 br_76 wl_165 vdd gnd cell_6t
Xbit_r166_c76 bl_76 br_76 wl_166 vdd gnd cell_6t
Xbit_r167_c76 bl_76 br_76 wl_167 vdd gnd cell_6t
Xbit_r168_c76 bl_76 br_76 wl_168 vdd gnd cell_6t
Xbit_r169_c76 bl_76 br_76 wl_169 vdd gnd cell_6t
Xbit_r170_c76 bl_76 br_76 wl_170 vdd gnd cell_6t
Xbit_r171_c76 bl_76 br_76 wl_171 vdd gnd cell_6t
Xbit_r172_c76 bl_76 br_76 wl_172 vdd gnd cell_6t
Xbit_r173_c76 bl_76 br_76 wl_173 vdd gnd cell_6t
Xbit_r174_c76 bl_76 br_76 wl_174 vdd gnd cell_6t
Xbit_r175_c76 bl_76 br_76 wl_175 vdd gnd cell_6t
Xbit_r176_c76 bl_76 br_76 wl_176 vdd gnd cell_6t
Xbit_r177_c76 bl_76 br_76 wl_177 vdd gnd cell_6t
Xbit_r178_c76 bl_76 br_76 wl_178 vdd gnd cell_6t
Xbit_r179_c76 bl_76 br_76 wl_179 vdd gnd cell_6t
Xbit_r180_c76 bl_76 br_76 wl_180 vdd gnd cell_6t
Xbit_r181_c76 bl_76 br_76 wl_181 vdd gnd cell_6t
Xbit_r182_c76 bl_76 br_76 wl_182 vdd gnd cell_6t
Xbit_r183_c76 bl_76 br_76 wl_183 vdd gnd cell_6t
Xbit_r184_c76 bl_76 br_76 wl_184 vdd gnd cell_6t
Xbit_r185_c76 bl_76 br_76 wl_185 vdd gnd cell_6t
Xbit_r186_c76 bl_76 br_76 wl_186 vdd gnd cell_6t
Xbit_r187_c76 bl_76 br_76 wl_187 vdd gnd cell_6t
Xbit_r188_c76 bl_76 br_76 wl_188 vdd gnd cell_6t
Xbit_r189_c76 bl_76 br_76 wl_189 vdd gnd cell_6t
Xbit_r190_c76 bl_76 br_76 wl_190 vdd gnd cell_6t
Xbit_r191_c76 bl_76 br_76 wl_191 vdd gnd cell_6t
Xbit_r192_c76 bl_76 br_76 wl_192 vdd gnd cell_6t
Xbit_r193_c76 bl_76 br_76 wl_193 vdd gnd cell_6t
Xbit_r194_c76 bl_76 br_76 wl_194 vdd gnd cell_6t
Xbit_r195_c76 bl_76 br_76 wl_195 vdd gnd cell_6t
Xbit_r196_c76 bl_76 br_76 wl_196 vdd gnd cell_6t
Xbit_r197_c76 bl_76 br_76 wl_197 vdd gnd cell_6t
Xbit_r198_c76 bl_76 br_76 wl_198 vdd gnd cell_6t
Xbit_r199_c76 bl_76 br_76 wl_199 vdd gnd cell_6t
Xbit_r200_c76 bl_76 br_76 wl_200 vdd gnd cell_6t
Xbit_r201_c76 bl_76 br_76 wl_201 vdd gnd cell_6t
Xbit_r202_c76 bl_76 br_76 wl_202 vdd gnd cell_6t
Xbit_r203_c76 bl_76 br_76 wl_203 vdd gnd cell_6t
Xbit_r204_c76 bl_76 br_76 wl_204 vdd gnd cell_6t
Xbit_r205_c76 bl_76 br_76 wl_205 vdd gnd cell_6t
Xbit_r206_c76 bl_76 br_76 wl_206 vdd gnd cell_6t
Xbit_r207_c76 bl_76 br_76 wl_207 vdd gnd cell_6t
Xbit_r208_c76 bl_76 br_76 wl_208 vdd gnd cell_6t
Xbit_r209_c76 bl_76 br_76 wl_209 vdd gnd cell_6t
Xbit_r210_c76 bl_76 br_76 wl_210 vdd gnd cell_6t
Xbit_r211_c76 bl_76 br_76 wl_211 vdd gnd cell_6t
Xbit_r212_c76 bl_76 br_76 wl_212 vdd gnd cell_6t
Xbit_r213_c76 bl_76 br_76 wl_213 vdd gnd cell_6t
Xbit_r214_c76 bl_76 br_76 wl_214 vdd gnd cell_6t
Xbit_r215_c76 bl_76 br_76 wl_215 vdd gnd cell_6t
Xbit_r216_c76 bl_76 br_76 wl_216 vdd gnd cell_6t
Xbit_r217_c76 bl_76 br_76 wl_217 vdd gnd cell_6t
Xbit_r218_c76 bl_76 br_76 wl_218 vdd gnd cell_6t
Xbit_r219_c76 bl_76 br_76 wl_219 vdd gnd cell_6t
Xbit_r220_c76 bl_76 br_76 wl_220 vdd gnd cell_6t
Xbit_r221_c76 bl_76 br_76 wl_221 vdd gnd cell_6t
Xbit_r222_c76 bl_76 br_76 wl_222 vdd gnd cell_6t
Xbit_r223_c76 bl_76 br_76 wl_223 vdd gnd cell_6t
Xbit_r224_c76 bl_76 br_76 wl_224 vdd gnd cell_6t
Xbit_r225_c76 bl_76 br_76 wl_225 vdd gnd cell_6t
Xbit_r226_c76 bl_76 br_76 wl_226 vdd gnd cell_6t
Xbit_r227_c76 bl_76 br_76 wl_227 vdd gnd cell_6t
Xbit_r228_c76 bl_76 br_76 wl_228 vdd gnd cell_6t
Xbit_r229_c76 bl_76 br_76 wl_229 vdd gnd cell_6t
Xbit_r230_c76 bl_76 br_76 wl_230 vdd gnd cell_6t
Xbit_r231_c76 bl_76 br_76 wl_231 vdd gnd cell_6t
Xbit_r232_c76 bl_76 br_76 wl_232 vdd gnd cell_6t
Xbit_r233_c76 bl_76 br_76 wl_233 vdd gnd cell_6t
Xbit_r234_c76 bl_76 br_76 wl_234 vdd gnd cell_6t
Xbit_r235_c76 bl_76 br_76 wl_235 vdd gnd cell_6t
Xbit_r236_c76 bl_76 br_76 wl_236 vdd gnd cell_6t
Xbit_r237_c76 bl_76 br_76 wl_237 vdd gnd cell_6t
Xbit_r238_c76 bl_76 br_76 wl_238 vdd gnd cell_6t
Xbit_r239_c76 bl_76 br_76 wl_239 vdd gnd cell_6t
Xbit_r240_c76 bl_76 br_76 wl_240 vdd gnd cell_6t
Xbit_r241_c76 bl_76 br_76 wl_241 vdd gnd cell_6t
Xbit_r242_c76 bl_76 br_76 wl_242 vdd gnd cell_6t
Xbit_r243_c76 bl_76 br_76 wl_243 vdd gnd cell_6t
Xbit_r244_c76 bl_76 br_76 wl_244 vdd gnd cell_6t
Xbit_r245_c76 bl_76 br_76 wl_245 vdd gnd cell_6t
Xbit_r246_c76 bl_76 br_76 wl_246 vdd gnd cell_6t
Xbit_r247_c76 bl_76 br_76 wl_247 vdd gnd cell_6t
Xbit_r248_c76 bl_76 br_76 wl_248 vdd gnd cell_6t
Xbit_r249_c76 bl_76 br_76 wl_249 vdd gnd cell_6t
Xbit_r250_c76 bl_76 br_76 wl_250 vdd gnd cell_6t
Xbit_r251_c76 bl_76 br_76 wl_251 vdd gnd cell_6t
Xbit_r252_c76 bl_76 br_76 wl_252 vdd gnd cell_6t
Xbit_r253_c76 bl_76 br_76 wl_253 vdd gnd cell_6t
Xbit_r254_c76 bl_76 br_76 wl_254 vdd gnd cell_6t
Xbit_r255_c76 bl_76 br_76 wl_255 vdd gnd cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd cell_6t
Xbit_r1_c77 bl_77 br_77 wl_1 vdd gnd cell_6t
Xbit_r2_c77 bl_77 br_77 wl_2 vdd gnd cell_6t
Xbit_r3_c77 bl_77 br_77 wl_3 vdd gnd cell_6t
Xbit_r4_c77 bl_77 br_77 wl_4 vdd gnd cell_6t
Xbit_r5_c77 bl_77 br_77 wl_5 vdd gnd cell_6t
Xbit_r6_c77 bl_77 br_77 wl_6 vdd gnd cell_6t
Xbit_r7_c77 bl_77 br_77 wl_7 vdd gnd cell_6t
Xbit_r8_c77 bl_77 br_77 wl_8 vdd gnd cell_6t
Xbit_r9_c77 bl_77 br_77 wl_9 vdd gnd cell_6t
Xbit_r10_c77 bl_77 br_77 wl_10 vdd gnd cell_6t
Xbit_r11_c77 bl_77 br_77 wl_11 vdd gnd cell_6t
Xbit_r12_c77 bl_77 br_77 wl_12 vdd gnd cell_6t
Xbit_r13_c77 bl_77 br_77 wl_13 vdd gnd cell_6t
Xbit_r14_c77 bl_77 br_77 wl_14 vdd gnd cell_6t
Xbit_r15_c77 bl_77 br_77 wl_15 vdd gnd cell_6t
Xbit_r16_c77 bl_77 br_77 wl_16 vdd gnd cell_6t
Xbit_r17_c77 bl_77 br_77 wl_17 vdd gnd cell_6t
Xbit_r18_c77 bl_77 br_77 wl_18 vdd gnd cell_6t
Xbit_r19_c77 bl_77 br_77 wl_19 vdd gnd cell_6t
Xbit_r20_c77 bl_77 br_77 wl_20 vdd gnd cell_6t
Xbit_r21_c77 bl_77 br_77 wl_21 vdd gnd cell_6t
Xbit_r22_c77 bl_77 br_77 wl_22 vdd gnd cell_6t
Xbit_r23_c77 bl_77 br_77 wl_23 vdd gnd cell_6t
Xbit_r24_c77 bl_77 br_77 wl_24 vdd gnd cell_6t
Xbit_r25_c77 bl_77 br_77 wl_25 vdd gnd cell_6t
Xbit_r26_c77 bl_77 br_77 wl_26 vdd gnd cell_6t
Xbit_r27_c77 bl_77 br_77 wl_27 vdd gnd cell_6t
Xbit_r28_c77 bl_77 br_77 wl_28 vdd gnd cell_6t
Xbit_r29_c77 bl_77 br_77 wl_29 vdd gnd cell_6t
Xbit_r30_c77 bl_77 br_77 wl_30 vdd gnd cell_6t
Xbit_r31_c77 bl_77 br_77 wl_31 vdd gnd cell_6t
Xbit_r32_c77 bl_77 br_77 wl_32 vdd gnd cell_6t
Xbit_r33_c77 bl_77 br_77 wl_33 vdd gnd cell_6t
Xbit_r34_c77 bl_77 br_77 wl_34 vdd gnd cell_6t
Xbit_r35_c77 bl_77 br_77 wl_35 vdd gnd cell_6t
Xbit_r36_c77 bl_77 br_77 wl_36 vdd gnd cell_6t
Xbit_r37_c77 bl_77 br_77 wl_37 vdd gnd cell_6t
Xbit_r38_c77 bl_77 br_77 wl_38 vdd gnd cell_6t
Xbit_r39_c77 bl_77 br_77 wl_39 vdd gnd cell_6t
Xbit_r40_c77 bl_77 br_77 wl_40 vdd gnd cell_6t
Xbit_r41_c77 bl_77 br_77 wl_41 vdd gnd cell_6t
Xbit_r42_c77 bl_77 br_77 wl_42 vdd gnd cell_6t
Xbit_r43_c77 bl_77 br_77 wl_43 vdd gnd cell_6t
Xbit_r44_c77 bl_77 br_77 wl_44 vdd gnd cell_6t
Xbit_r45_c77 bl_77 br_77 wl_45 vdd gnd cell_6t
Xbit_r46_c77 bl_77 br_77 wl_46 vdd gnd cell_6t
Xbit_r47_c77 bl_77 br_77 wl_47 vdd gnd cell_6t
Xbit_r48_c77 bl_77 br_77 wl_48 vdd gnd cell_6t
Xbit_r49_c77 bl_77 br_77 wl_49 vdd gnd cell_6t
Xbit_r50_c77 bl_77 br_77 wl_50 vdd gnd cell_6t
Xbit_r51_c77 bl_77 br_77 wl_51 vdd gnd cell_6t
Xbit_r52_c77 bl_77 br_77 wl_52 vdd gnd cell_6t
Xbit_r53_c77 bl_77 br_77 wl_53 vdd gnd cell_6t
Xbit_r54_c77 bl_77 br_77 wl_54 vdd gnd cell_6t
Xbit_r55_c77 bl_77 br_77 wl_55 vdd gnd cell_6t
Xbit_r56_c77 bl_77 br_77 wl_56 vdd gnd cell_6t
Xbit_r57_c77 bl_77 br_77 wl_57 vdd gnd cell_6t
Xbit_r58_c77 bl_77 br_77 wl_58 vdd gnd cell_6t
Xbit_r59_c77 bl_77 br_77 wl_59 vdd gnd cell_6t
Xbit_r60_c77 bl_77 br_77 wl_60 vdd gnd cell_6t
Xbit_r61_c77 bl_77 br_77 wl_61 vdd gnd cell_6t
Xbit_r62_c77 bl_77 br_77 wl_62 vdd gnd cell_6t
Xbit_r63_c77 bl_77 br_77 wl_63 vdd gnd cell_6t
Xbit_r64_c77 bl_77 br_77 wl_64 vdd gnd cell_6t
Xbit_r65_c77 bl_77 br_77 wl_65 vdd gnd cell_6t
Xbit_r66_c77 bl_77 br_77 wl_66 vdd gnd cell_6t
Xbit_r67_c77 bl_77 br_77 wl_67 vdd gnd cell_6t
Xbit_r68_c77 bl_77 br_77 wl_68 vdd gnd cell_6t
Xbit_r69_c77 bl_77 br_77 wl_69 vdd gnd cell_6t
Xbit_r70_c77 bl_77 br_77 wl_70 vdd gnd cell_6t
Xbit_r71_c77 bl_77 br_77 wl_71 vdd gnd cell_6t
Xbit_r72_c77 bl_77 br_77 wl_72 vdd gnd cell_6t
Xbit_r73_c77 bl_77 br_77 wl_73 vdd gnd cell_6t
Xbit_r74_c77 bl_77 br_77 wl_74 vdd gnd cell_6t
Xbit_r75_c77 bl_77 br_77 wl_75 vdd gnd cell_6t
Xbit_r76_c77 bl_77 br_77 wl_76 vdd gnd cell_6t
Xbit_r77_c77 bl_77 br_77 wl_77 vdd gnd cell_6t
Xbit_r78_c77 bl_77 br_77 wl_78 vdd gnd cell_6t
Xbit_r79_c77 bl_77 br_77 wl_79 vdd gnd cell_6t
Xbit_r80_c77 bl_77 br_77 wl_80 vdd gnd cell_6t
Xbit_r81_c77 bl_77 br_77 wl_81 vdd gnd cell_6t
Xbit_r82_c77 bl_77 br_77 wl_82 vdd gnd cell_6t
Xbit_r83_c77 bl_77 br_77 wl_83 vdd gnd cell_6t
Xbit_r84_c77 bl_77 br_77 wl_84 vdd gnd cell_6t
Xbit_r85_c77 bl_77 br_77 wl_85 vdd gnd cell_6t
Xbit_r86_c77 bl_77 br_77 wl_86 vdd gnd cell_6t
Xbit_r87_c77 bl_77 br_77 wl_87 vdd gnd cell_6t
Xbit_r88_c77 bl_77 br_77 wl_88 vdd gnd cell_6t
Xbit_r89_c77 bl_77 br_77 wl_89 vdd gnd cell_6t
Xbit_r90_c77 bl_77 br_77 wl_90 vdd gnd cell_6t
Xbit_r91_c77 bl_77 br_77 wl_91 vdd gnd cell_6t
Xbit_r92_c77 bl_77 br_77 wl_92 vdd gnd cell_6t
Xbit_r93_c77 bl_77 br_77 wl_93 vdd gnd cell_6t
Xbit_r94_c77 bl_77 br_77 wl_94 vdd gnd cell_6t
Xbit_r95_c77 bl_77 br_77 wl_95 vdd gnd cell_6t
Xbit_r96_c77 bl_77 br_77 wl_96 vdd gnd cell_6t
Xbit_r97_c77 bl_77 br_77 wl_97 vdd gnd cell_6t
Xbit_r98_c77 bl_77 br_77 wl_98 vdd gnd cell_6t
Xbit_r99_c77 bl_77 br_77 wl_99 vdd gnd cell_6t
Xbit_r100_c77 bl_77 br_77 wl_100 vdd gnd cell_6t
Xbit_r101_c77 bl_77 br_77 wl_101 vdd gnd cell_6t
Xbit_r102_c77 bl_77 br_77 wl_102 vdd gnd cell_6t
Xbit_r103_c77 bl_77 br_77 wl_103 vdd gnd cell_6t
Xbit_r104_c77 bl_77 br_77 wl_104 vdd gnd cell_6t
Xbit_r105_c77 bl_77 br_77 wl_105 vdd gnd cell_6t
Xbit_r106_c77 bl_77 br_77 wl_106 vdd gnd cell_6t
Xbit_r107_c77 bl_77 br_77 wl_107 vdd gnd cell_6t
Xbit_r108_c77 bl_77 br_77 wl_108 vdd gnd cell_6t
Xbit_r109_c77 bl_77 br_77 wl_109 vdd gnd cell_6t
Xbit_r110_c77 bl_77 br_77 wl_110 vdd gnd cell_6t
Xbit_r111_c77 bl_77 br_77 wl_111 vdd gnd cell_6t
Xbit_r112_c77 bl_77 br_77 wl_112 vdd gnd cell_6t
Xbit_r113_c77 bl_77 br_77 wl_113 vdd gnd cell_6t
Xbit_r114_c77 bl_77 br_77 wl_114 vdd gnd cell_6t
Xbit_r115_c77 bl_77 br_77 wl_115 vdd gnd cell_6t
Xbit_r116_c77 bl_77 br_77 wl_116 vdd gnd cell_6t
Xbit_r117_c77 bl_77 br_77 wl_117 vdd gnd cell_6t
Xbit_r118_c77 bl_77 br_77 wl_118 vdd gnd cell_6t
Xbit_r119_c77 bl_77 br_77 wl_119 vdd gnd cell_6t
Xbit_r120_c77 bl_77 br_77 wl_120 vdd gnd cell_6t
Xbit_r121_c77 bl_77 br_77 wl_121 vdd gnd cell_6t
Xbit_r122_c77 bl_77 br_77 wl_122 vdd gnd cell_6t
Xbit_r123_c77 bl_77 br_77 wl_123 vdd gnd cell_6t
Xbit_r124_c77 bl_77 br_77 wl_124 vdd gnd cell_6t
Xbit_r125_c77 bl_77 br_77 wl_125 vdd gnd cell_6t
Xbit_r126_c77 bl_77 br_77 wl_126 vdd gnd cell_6t
Xbit_r127_c77 bl_77 br_77 wl_127 vdd gnd cell_6t
Xbit_r128_c77 bl_77 br_77 wl_128 vdd gnd cell_6t
Xbit_r129_c77 bl_77 br_77 wl_129 vdd gnd cell_6t
Xbit_r130_c77 bl_77 br_77 wl_130 vdd gnd cell_6t
Xbit_r131_c77 bl_77 br_77 wl_131 vdd gnd cell_6t
Xbit_r132_c77 bl_77 br_77 wl_132 vdd gnd cell_6t
Xbit_r133_c77 bl_77 br_77 wl_133 vdd gnd cell_6t
Xbit_r134_c77 bl_77 br_77 wl_134 vdd gnd cell_6t
Xbit_r135_c77 bl_77 br_77 wl_135 vdd gnd cell_6t
Xbit_r136_c77 bl_77 br_77 wl_136 vdd gnd cell_6t
Xbit_r137_c77 bl_77 br_77 wl_137 vdd gnd cell_6t
Xbit_r138_c77 bl_77 br_77 wl_138 vdd gnd cell_6t
Xbit_r139_c77 bl_77 br_77 wl_139 vdd gnd cell_6t
Xbit_r140_c77 bl_77 br_77 wl_140 vdd gnd cell_6t
Xbit_r141_c77 bl_77 br_77 wl_141 vdd gnd cell_6t
Xbit_r142_c77 bl_77 br_77 wl_142 vdd gnd cell_6t
Xbit_r143_c77 bl_77 br_77 wl_143 vdd gnd cell_6t
Xbit_r144_c77 bl_77 br_77 wl_144 vdd gnd cell_6t
Xbit_r145_c77 bl_77 br_77 wl_145 vdd gnd cell_6t
Xbit_r146_c77 bl_77 br_77 wl_146 vdd gnd cell_6t
Xbit_r147_c77 bl_77 br_77 wl_147 vdd gnd cell_6t
Xbit_r148_c77 bl_77 br_77 wl_148 vdd gnd cell_6t
Xbit_r149_c77 bl_77 br_77 wl_149 vdd gnd cell_6t
Xbit_r150_c77 bl_77 br_77 wl_150 vdd gnd cell_6t
Xbit_r151_c77 bl_77 br_77 wl_151 vdd gnd cell_6t
Xbit_r152_c77 bl_77 br_77 wl_152 vdd gnd cell_6t
Xbit_r153_c77 bl_77 br_77 wl_153 vdd gnd cell_6t
Xbit_r154_c77 bl_77 br_77 wl_154 vdd gnd cell_6t
Xbit_r155_c77 bl_77 br_77 wl_155 vdd gnd cell_6t
Xbit_r156_c77 bl_77 br_77 wl_156 vdd gnd cell_6t
Xbit_r157_c77 bl_77 br_77 wl_157 vdd gnd cell_6t
Xbit_r158_c77 bl_77 br_77 wl_158 vdd gnd cell_6t
Xbit_r159_c77 bl_77 br_77 wl_159 vdd gnd cell_6t
Xbit_r160_c77 bl_77 br_77 wl_160 vdd gnd cell_6t
Xbit_r161_c77 bl_77 br_77 wl_161 vdd gnd cell_6t
Xbit_r162_c77 bl_77 br_77 wl_162 vdd gnd cell_6t
Xbit_r163_c77 bl_77 br_77 wl_163 vdd gnd cell_6t
Xbit_r164_c77 bl_77 br_77 wl_164 vdd gnd cell_6t
Xbit_r165_c77 bl_77 br_77 wl_165 vdd gnd cell_6t
Xbit_r166_c77 bl_77 br_77 wl_166 vdd gnd cell_6t
Xbit_r167_c77 bl_77 br_77 wl_167 vdd gnd cell_6t
Xbit_r168_c77 bl_77 br_77 wl_168 vdd gnd cell_6t
Xbit_r169_c77 bl_77 br_77 wl_169 vdd gnd cell_6t
Xbit_r170_c77 bl_77 br_77 wl_170 vdd gnd cell_6t
Xbit_r171_c77 bl_77 br_77 wl_171 vdd gnd cell_6t
Xbit_r172_c77 bl_77 br_77 wl_172 vdd gnd cell_6t
Xbit_r173_c77 bl_77 br_77 wl_173 vdd gnd cell_6t
Xbit_r174_c77 bl_77 br_77 wl_174 vdd gnd cell_6t
Xbit_r175_c77 bl_77 br_77 wl_175 vdd gnd cell_6t
Xbit_r176_c77 bl_77 br_77 wl_176 vdd gnd cell_6t
Xbit_r177_c77 bl_77 br_77 wl_177 vdd gnd cell_6t
Xbit_r178_c77 bl_77 br_77 wl_178 vdd gnd cell_6t
Xbit_r179_c77 bl_77 br_77 wl_179 vdd gnd cell_6t
Xbit_r180_c77 bl_77 br_77 wl_180 vdd gnd cell_6t
Xbit_r181_c77 bl_77 br_77 wl_181 vdd gnd cell_6t
Xbit_r182_c77 bl_77 br_77 wl_182 vdd gnd cell_6t
Xbit_r183_c77 bl_77 br_77 wl_183 vdd gnd cell_6t
Xbit_r184_c77 bl_77 br_77 wl_184 vdd gnd cell_6t
Xbit_r185_c77 bl_77 br_77 wl_185 vdd gnd cell_6t
Xbit_r186_c77 bl_77 br_77 wl_186 vdd gnd cell_6t
Xbit_r187_c77 bl_77 br_77 wl_187 vdd gnd cell_6t
Xbit_r188_c77 bl_77 br_77 wl_188 vdd gnd cell_6t
Xbit_r189_c77 bl_77 br_77 wl_189 vdd gnd cell_6t
Xbit_r190_c77 bl_77 br_77 wl_190 vdd gnd cell_6t
Xbit_r191_c77 bl_77 br_77 wl_191 vdd gnd cell_6t
Xbit_r192_c77 bl_77 br_77 wl_192 vdd gnd cell_6t
Xbit_r193_c77 bl_77 br_77 wl_193 vdd gnd cell_6t
Xbit_r194_c77 bl_77 br_77 wl_194 vdd gnd cell_6t
Xbit_r195_c77 bl_77 br_77 wl_195 vdd gnd cell_6t
Xbit_r196_c77 bl_77 br_77 wl_196 vdd gnd cell_6t
Xbit_r197_c77 bl_77 br_77 wl_197 vdd gnd cell_6t
Xbit_r198_c77 bl_77 br_77 wl_198 vdd gnd cell_6t
Xbit_r199_c77 bl_77 br_77 wl_199 vdd gnd cell_6t
Xbit_r200_c77 bl_77 br_77 wl_200 vdd gnd cell_6t
Xbit_r201_c77 bl_77 br_77 wl_201 vdd gnd cell_6t
Xbit_r202_c77 bl_77 br_77 wl_202 vdd gnd cell_6t
Xbit_r203_c77 bl_77 br_77 wl_203 vdd gnd cell_6t
Xbit_r204_c77 bl_77 br_77 wl_204 vdd gnd cell_6t
Xbit_r205_c77 bl_77 br_77 wl_205 vdd gnd cell_6t
Xbit_r206_c77 bl_77 br_77 wl_206 vdd gnd cell_6t
Xbit_r207_c77 bl_77 br_77 wl_207 vdd gnd cell_6t
Xbit_r208_c77 bl_77 br_77 wl_208 vdd gnd cell_6t
Xbit_r209_c77 bl_77 br_77 wl_209 vdd gnd cell_6t
Xbit_r210_c77 bl_77 br_77 wl_210 vdd gnd cell_6t
Xbit_r211_c77 bl_77 br_77 wl_211 vdd gnd cell_6t
Xbit_r212_c77 bl_77 br_77 wl_212 vdd gnd cell_6t
Xbit_r213_c77 bl_77 br_77 wl_213 vdd gnd cell_6t
Xbit_r214_c77 bl_77 br_77 wl_214 vdd gnd cell_6t
Xbit_r215_c77 bl_77 br_77 wl_215 vdd gnd cell_6t
Xbit_r216_c77 bl_77 br_77 wl_216 vdd gnd cell_6t
Xbit_r217_c77 bl_77 br_77 wl_217 vdd gnd cell_6t
Xbit_r218_c77 bl_77 br_77 wl_218 vdd gnd cell_6t
Xbit_r219_c77 bl_77 br_77 wl_219 vdd gnd cell_6t
Xbit_r220_c77 bl_77 br_77 wl_220 vdd gnd cell_6t
Xbit_r221_c77 bl_77 br_77 wl_221 vdd gnd cell_6t
Xbit_r222_c77 bl_77 br_77 wl_222 vdd gnd cell_6t
Xbit_r223_c77 bl_77 br_77 wl_223 vdd gnd cell_6t
Xbit_r224_c77 bl_77 br_77 wl_224 vdd gnd cell_6t
Xbit_r225_c77 bl_77 br_77 wl_225 vdd gnd cell_6t
Xbit_r226_c77 bl_77 br_77 wl_226 vdd gnd cell_6t
Xbit_r227_c77 bl_77 br_77 wl_227 vdd gnd cell_6t
Xbit_r228_c77 bl_77 br_77 wl_228 vdd gnd cell_6t
Xbit_r229_c77 bl_77 br_77 wl_229 vdd gnd cell_6t
Xbit_r230_c77 bl_77 br_77 wl_230 vdd gnd cell_6t
Xbit_r231_c77 bl_77 br_77 wl_231 vdd gnd cell_6t
Xbit_r232_c77 bl_77 br_77 wl_232 vdd gnd cell_6t
Xbit_r233_c77 bl_77 br_77 wl_233 vdd gnd cell_6t
Xbit_r234_c77 bl_77 br_77 wl_234 vdd gnd cell_6t
Xbit_r235_c77 bl_77 br_77 wl_235 vdd gnd cell_6t
Xbit_r236_c77 bl_77 br_77 wl_236 vdd gnd cell_6t
Xbit_r237_c77 bl_77 br_77 wl_237 vdd gnd cell_6t
Xbit_r238_c77 bl_77 br_77 wl_238 vdd gnd cell_6t
Xbit_r239_c77 bl_77 br_77 wl_239 vdd gnd cell_6t
Xbit_r240_c77 bl_77 br_77 wl_240 vdd gnd cell_6t
Xbit_r241_c77 bl_77 br_77 wl_241 vdd gnd cell_6t
Xbit_r242_c77 bl_77 br_77 wl_242 vdd gnd cell_6t
Xbit_r243_c77 bl_77 br_77 wl_243 vdd gnd cell_6t
Xbit_r244_c77 bl_77 br_77 wl_244 vdd gnd cell_6t
Xbit_r245_c77 bl_77 br_77 wl_245 vdd gnd cell_6t
Xbit_r246_c77 bl_77 br_77 wl_246 vdd gnd cell_6t
Xbit_r247_c77 bl_77 br_77 wl_247 vdd gnd cell_6t
Xbit_r248_c77 bl_77 br_77 wl_248 vdd gnd cell_6t
Xbit_r249_c77 bl_77 br_77 wl_249 vdd gnd cell_6t
Xbit_r250_c77 bl_77 br_77 wl_250 vdd gnd cell_6t
Xbit_r251_c77 bl_77 br_77 wl_251 vdd gnd cell_6t
Xbit_r252_c77 bl_77 br_77 wl_252 vdd gnd cell_6t
Xbit_r253_c77 bl_77 br_77 wl_253 vdd gnd cell_6t
Xbit_r254_c77 bl_77 br_77 wl_254 vdd gnd cell_6t
Xbit_r255_c77 bl_77 br_77 wl_255 vdd gnd cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd cell_6t
Xbit_r1_c78 bl_78 br_78 wl_1 vdd gnd cell_6t
Xbit_r2_c78 bl_78 br_78 wl_2 vdd gnd cell_6t
Xbit_r3_c78 bl_78 br_78 wl_3 vdd gnd cell_6t
Xbit_r4_c78 bl_78 br_78 wl_4 vdd gnd cell_6t
Xbit_r5_c78 bl_78 br_78 wl_5 vdd gnd cell_6t
Xbit_r6_c78 bl_78 br_78 wl_6 vdd gnd cell_6t
Xbit_r7_c78 bl_78 br_78 wl_7 vdd gnd cell_6t
Xbit_r8_c78 bl_78 br_78 wl_8 vdd gnd cell_6t
Xbit_r9_c78 bl_78 br_78 wl_9 vdd gnd cell_6t
Xbit_r10_c78 bl_78 br_78 wl_10 vdd gnd cell_6t
Xbit_r11_c78 bl_78 br_78 wl_11 vdd gnd cell_6t
Xbit_r12_c78 bl_78 br_78 wl_12 vdd gnd cell_6t
Xbit_r13_c78 bl_78 br_78 wl_13 vdd gnd cell_6t
Xbit_r14_c78 bl_78 br_78 wl_14 vdd gnd cell_6t
Xbit_r15_c78 bl_78 br_78 wl_15 vdd gnd cell_6t
Xbit_r16_c78 bl_78 br_78 wl_16 vdd gnd cell_6t
Xbit_r17_c78 bl_78 br_78 wl_17 vdd gnd cell_6t
Xbit_r18_c78 bl_78 br_78 wl_18 vdd gnd cell_6t
Xbit_r19_c78 bl_78 br_78 wl_19 vdd gnd cell_6t
Xbit_r20_c78 bl_78 br_78 wl_20 vdd gnd cell_6t
Xbit_r21_c78 bl_78 br_78 wl_21 vdd gnd cell_6t
Xbit_r22_c78 bl_78 br_78 wl_22 vdd gnd cell_6t
Xbit_r23_c78 bl_78 br_78 wl_23 vdd gnd cell_6t
Xbit_r24_c78 bl_78 br_78 wl_24 vdd gnd cell_6t
Xbit_r25_c78 bl_78 br_78 wl_25 vdd gnd cell_6t
Xbit_r26_c78 bl_78 br_78 wl_26 vdd gnd cell_6t
Xbit_r27_c78 bl_78 br_78 wl_27 vdd gnd cell_6t
Xbit_r28_c78 bl_78 br_78 wl_28 vdd gnd cell_6t
Xbit_r29_c78 bl_78 br_78 wl_29 vdd gnd cell_6t
Xbit_r30_c78 bl_78 br_78 wl_30 vdd gnd cell_6t
Xbit_r31_c78 bl_78 br_78 wl_31 vdd gnd cell_6t
Xbit_r32_c78 bl_78 br_78 wl_32 vdd gnd cell_6t
Xbit_r33_c78 bl_78 br_78 wl_33 vdd gnd cell_6t
Xbit_r34_c78 bl_78 br_78 wl_34 vdd gnd cell_6t
Xbit_r35_c78 bl_78 br_78 wl_35 vdd gnd cell_6t
Xbit_r36_c78 bl_78 br_78 wl_36 vdd gnd cell_6t
Xbit_r37_c78 bl_78 br_78 wl_37 vdd gnd cell_6t
Xbit_r38_c78 bl_78 br_78 wl_38 vdd gnd cell_6t
Xbit_r39_c78 bl_78 br_78 wl_39 vdd gnd cell_6t
Xbit_r40_c78 bl_78 br_78 wl_40 vdd gnd cell_6t
Xbit_r41_c78 bl_78 br_78 wl_41 vdd gnd cell_6t
Xbit_r42_c78 bl_78 br_78 wl_42 vdd gnd cell_6t
Xbit_r43_c78 bl_78 br_78 wl_43 vdd gnd cell_6t
Xbit_r44_c78 bl_78 br_78 wl_44 vdd gnd cell_6t
Xbit_r45_c78 bl_78 br_78 wl_45 vdd gnd cell_6t
Xbit_r46_c78 bl_78 br_78 wl_46 vdd gnd cell_6t
Xbit_r47_c78 bl_78 br_78 wl_47 vdd gnd cell_6t
Xbit_r48_c78 bl_78 br_78 wl_48 vdd gnd cell_6t
Xbit_r49_c78 bl_78 br_78 wl_49 vdd gnd cell_6t
Xbit_r50_c78 bl_78 br_78 wl_50 vdd gnd cell_6t
Xbit_r51_c78 bl_78 br_78 wl_51 vdd gnd cell_6t
Xbit_r52_c78 bl_78 br_78 wl_52 vdd gnd cell_6t
Xbit_r53_c78 bl_78 br_78 wl_53 vdd gnd cell_6t
Xbit_r54_c78 bl_78 br_78 wl_54 vdd gnd cell_6t
Xbit_r55_c78 bl_78 br_78 wl_55 vdd gnd cell_6t
Xbit_r56_c78 bl_78 br_78 wl_56 vdd gnd cell_6t
Xbit_r57_c78 bl_78 br_78 wl_57 vdd gnd cell_6t
Xbit_r58_c78 bl_78 br_78 wl_58 vdd gnd cell_6t
Xbit_r59_c78 bl_78 br_78 wl_59 vdd gnd cell_6t
Xbit_r60_c78 bl_78 br_78 wl_60 vdd gnd cell_6t
Xbit_r61_c78 bl_78 br_78 wl_61 vdd gnd cell_6t
Xbit_r62_c78 bl_78 br_78 wl_62 vdd gnd cell_6t
Xbit_r63_c78 bl_78 br_78 wl_63 vdd gnd cell_6t
Xbit_r64_c78 bl_78 br_78 wl_64 vdd gnd cell_6t
Xbit_r65_c78 bl_78 br_78 wl_65 vdd gnd cell_6t
Xbit_r66_c78 bl_78 br_78 wl_66 vdd gnd cell_6t
Xbit_r67_c78 bl_78 br_78 wl_67 vdd gnd cell_6t
Xbit_r68_c78 bl_78 br_78 wl_68 vdd gnd cell_6t
Xbit_r69_c78 bl_78 br_78 wl_69 vdd gnd cell_6t
Xbit_r70_c78 bl_78 br_78 wl_70 vdd gnd cell_6t
Xbit_r71_c78 bl_78 br_78 wl_71 vdd gnd cell_6t
Xbit_r72_c78 bl_78 br_78 wl_72 vdd gnd cell_6t
Xbit_r73_c78 bl_78 br_78 wl_73 vdd gnd cell_6t
Xbit_r74_c78 bl_78 br_78 wl_74 vdd gnd cell_6t
Xbit_r75_c78 bl_78 br_78 wl_75 vdd gnd cell_6t
Xbit_r76_c78 bl_78 br_78 wl_76 vdd gnd cell_6t
Xbit_r77_c78 bl_78 br_78 wl_77 vdd gnd cell_6t
Xbit_r78_c78 bl_78 br_78 wl_78 vdd gnd cell_6t
Xbit_r79_c78 bl_78 br_78 wl_79 vdd gnd cell_6t
Xbit_r80_c78 bl_78 br_78 wl_80 vdd gnd cell_6t
Xbit_r81_c78 bl_78 br_78 wl_81 vdd gnd cell_6t
Xbit_r82_c78 bl_78 br_78 wl_82 vdd gnd cell_6t
Xbit_r83_c78 bl_78 br_78 wl_83 vdd gnd cell_6t
Xbit_r84_c78 bl_78 br_78 wl_84 vdd gnd cell_6t
Xbit_r85_c78 bl_78 br_78 wl_85 vdd gnd cell_6t
Xbit_r86_c78 bl_78 br_78 wl_86 vdd gnd cell_6t
Xbit_r87_c78 bl_78 br_78 wl_87 vdd gnd cell_6t
Xbit_r88_c78 bl_78 br_78 wl_88 vdd gnd cell_6t
Xbit_r89_c78 bl_78 br_78 wl_89 vdd gnd cell_6t
Xbit_r90_c78 bl_78 br_78 wl_90 vdd gnd cell_6t
Xbit_r91_c78 bl_78 br_78 wl_91 vdd gnd cell_6t
Xbit_r92_c78 bl_78 br_78 wl_92 vdd gnd cell_6t
Xbit_r93_c78 bl_78 br_78 wl_93 vdd gnd cell_6t
Xbit_r94_c78 bl_78 br_78 wl_94 vdd gnd cell_6t
Xbit_r95_c78 bl_78 br_78 wl_95 vdd gnd cell_6t
Xbit_r96_c78 bl_78 br_78 wl_96 vdd gnd cell_6t
Xbit_r97_c78 bl_78 br_78 wl_97 vdd gnd cell_6t
Xbit_r98_c78 bl_78 br_78 wl_98 vdd gnd cell_6t
Xbit_r99_c78 bl_78 br_78 wl_99 vdd gnd cell_6t
Xbit_r100_c78 bl_78 br_78 wl_100 vdd gnd cell_6t
Xbit_r101_c78 bl_78 br_78 wl_101 vdd gnd cell_6t
Xbit_r102_c78 bl_78 br_78 wl_102 vdd gnd cell_6t
Xbit_r103_c78 bl_78 br_78 wl_103 vdd gnd cell_6t
Xbit_r104_c78 bl_78 br_78 wl_104 vdd gnd cell_6t
Xbit_r105_c78 bl_78 br_78 wl_105 vdd gnd cell_6t
Xbit_r106_c78 bl_78 br_78 wl_106 vdd gnd cell_6t
Xbit_r107_c78 bl_78 br_78 wl_107 vdd gnd cell_6t
Xbit_r108_c78 bl_78 br_78 wl_108 vdd gnd cell_6t
Xbit_r109_c78 bl_78 br_78 wl_109 vdd gnd cell_6t
Xbit_r110_c78 bl_78 br_78 wl_110 vdd gnd cell_6t
Xbit_r111_c78 bl_78 br_78 wl_111 vdd gnd cell_6t
Xbit_r112_c78 bl_78 br_78 wl_112 vdd gnd cell_6t
Xbit_r113_c78 bl_78 br_78 wl_113 vdd gnd cell_6t
Xbit_r114_c78 bl_78 br_78 wl_114 vdd gnd cell_6t
Xbit_r115_c78 bl_78 br_78 wl_115 vdd gnd cell_6t
Xbit_r116_c78 bl_78 br_78 wl_116 vdd gnd cell_6t
Xbit_r117_c78 bl_78 br_78 wl_117 vdd gnd cell_6t
Xbit_r118_c78 bl_78 br_78 wl_118 vdd gnd cell_6t
Xbit_r119_c78 bl_78 br_78 wl_119 vdd gnd cell_6t
Xbit_r120_c78 bl_78 br_78 wl_120 vdd gnd cell_6t
Xbit_r121_c78 bl_78 br_78 wl_121 vdd gnd cell_6t
Xbit_r122_c78 bl_78 br_78 wl_122 vdd gnd cell_6t
Xbit_r123_c78 bl_78 br_78 wl_123 vdd gnd cell_6t
Xbit_r124_c78 bl_78 br_78 wl_124 vdd gnd cell_6t
Xbit_r125_c78 bl_78 br_78 wl_125 vdd gnd cell_6t
Xbit_r126_c78 bl_78 br_78 wl_126 vdd gnd cell_6t
Xbit_r127_c78 bl_78 br_78 wl_127 vdd gnd cell_6t
Xbit_r128_c78 bl_78 br_78 wl_128 vdd gnd cell_6t
Xbit_r129_c78 bl_78 br_78 wl_129 vdd gnd cell_6t
Xbit_r130_c78 bl_78 br_78 wl_130 vdd gnd cell_6t
Xbit_r131_c78 bl_78 br_78 wl_131 vdd gnd cell_6t
Xbit_r132_c78 bl_78 br_78 wl_132 vdd gnd cell_6t
Xbit_r133_c78 bl_78 br_78 wl_133 vdd gnd cell_6t
Xbit_r134_c78 bl_78 br_78 wl_134 vdd gnd cell_6t
Xbit_r135_c78 bl_78 br_78 wl_135 vdd gnd cell_6t
Xbit_r136_c78 bl_78 br_78 wl_136 vdd gnd cell_6t
Xbit_r137_c78 bl_78 br_78 wl_137 vdd gnd cell_6t
Xbit_r138_c78 bl_78 br_78 wl_138 vdd gnd cell_6t
Xbit_r139_c78 bl_78 br_78 wl_139 vdd gnd cell_6t
Xbit_r140_c78 bl_78 br_78 wl_140 vdd gnd cell_6t
Xbit_r141_c78 bl_78 br_78 wl_141 vdd gnd cell_6t
Xbit_r142_c78 bl_78 br_78 wl_142 vdd gnd cell_6t
Xbit_r143_c78 bl_78 br_78 wl_143 vdd gnd cell_6t
Xbit_r144_c78 bl_78 br_78 wl_144 vdd gnd cell_6t
Xbit_r145_c78 bl_78 br_78 wl_145 vdd gnd cell_6t
Xbit_r146_c78 bl_78 br_78 wl_146 vdd gnd cell_6t
Xbit_r147_c78 bl_78 br_78 wl_147 vdd gnd cell_6t
Xbit_r148_c78 bl_78 br_78 wl_148 vdd gnd cell_6t
Xbit_r149_c78 bl_78 br_78 wl_149 vdd gnd cell_6t
Xbit_r150_c78 bl_78 br_78 wl_150 vdd gnd cell_6t
Xbit_r151_c78 bl_78 br_78 wl_151 vdd gnd cell_6t
Xbit_r152_c78 bl_78 br_78 wl_152 vdd gnd cell_6t
Xbit_r153_c78 bl_78 br_78 wl_153 vdd gnd cell_6t
Xbit_r154_c78 bl_78 br_78 wl_154 vdd gnd cell_6t
Xbit_r155_c78 bl_78 br_78 wl_155 vdd gnd cell_6t
Xbit_r156_c78 bl_78 br_78 wl_156 vdd gnd cell_6t
Xbit_r157_c78 bl_78 br_78 wl_157 vdd gnd cell_6t
Xbit_r158_c78 bl_78 br_78 wl_158 vdd gnd cell_6t
Xbit_r159_c78 bl_78 br_78 wl_159 vdd gnd cell_6t
Xbit_r160_c78 bl_78 br_78 wl_160 vdd gnd cell_6t
Xbit_r161_c78 bl_78 br_78 wl_161 vdd gnd cell_6t
Xbit_r162_c78 bl_78 br_78 wl_162 vdd gnd cell_6t
Xbit_r163_c78 bl_78 br_78 wl_163 vdd gnd cell_6t
Xbit_r164_c78 bl_78 br_78 wl_164 vdd gnd cell_6t
Xbit_r165_c78 bl_78 br_78 wl_165 vdd gnd cell_6t
Xbit_r166_c78 bl_78 br_78 wl_166 vdd gnd cell_6t
Xbit_r167_c78 bl_78 br_78 wl_167 vdd gnd cell_6t
Xbit_r168_c78 bl_78 br_78 wl_168 vdd gnd cell_6t
Xbit_r169_c78 bl_78 br_78 wl_169 vdd gnd cell_6t
Xbit_r170_c78 bl_78 br_78 wl_170 vdd gnd cell_6t
Xbit_r171_c78 bl_78 br_78 wl_171 vdd gnd cell_6t
Xbit_r172_c78 bl_78 br_78 wl_172 vdd gnd cell_6t
Xbit_r173_c78 bl_78 br_78 wl_173 vdd gnd cell_6t
Xbit_r174_c78 bl_78 br_78 wl_174 vdd gnd cell_6t
Xbit_r175_c78 bl_78 br_78 wl_175 vdd gnd cell_6t
Xbit_r176_c78 bl_78 br_78 wl_176 vdd gnd cell_6t
Xbit_r177_c78 bl_78 br_78 wl_177 vdd gnd cell_6t
Xbit_r178_c78 bl_78 br_78 wl_178 vdd gnd cell_6t
Xbit_r179_c78 bl_78 br_78 wl_179 vdd gnd cell_6t
Xbit_r180_c78 bl_78 br_78 wl_180 vdd gnd cell_6t
Xbit_r181_c78 bl_78 br_78 wl_181 vdd gnd cell_6t
Xbit_r182_c78 bl_78 br_78 wl_182 vdd gnd cell_6t
Xbit_r183_c78 bl_78 br_78 wl_183 vdd gnd cell_6t
Xbit_r184_c78 bl_78 br_78 wl_184 vdd gnd cell_6t
Xbit_r185_c78 bl_78 br_78 wl_185 vdd gnd cell_6t
Xbit_r186_c78 bl_78 br_78 wl_186 vdd gnd cell_6t
Xbit_r187_c78 bl_78 br_78 wl_187 vdd gnd cell_6t
Xbit_r188_c78 bl_78 br_78 wl_188 vdd gnd cell_6t
Xbit_r189_c78 bl_78 br_78 wl_189 vdd gnd cell_6t
Xbit_r190_c78 bl_78 br_78 wl_190 vdd gnd cell_6t
Xbit_r191_c78 bl_78 br_78 wl_191 vdd gnd cell_6t
Xbit_r192_c78 bl_78 br_78 wl_192 vdd gnd cell_6t
Xbit_r193_c78 bl_78 br_78 wl_193 vdd gnd cell_6t
Xbit_r194_c78 bl_78 br_78 wl_194 vdd gnd cell_6t
Xbit_r195_c78 bl_78 br_78 wl_195 vdd gnd cell_6t
Xbit_r196_c78 bl_78 br_78 wl_196 vdd gnd cell_6t
Xbit_r197_c78 bl_78 br_78 wl_197 vdd gnd cell_6t
Xbit_r198_c78 bl_78 br_78 wl_198 vdd gnd cell_6t
Xbit_r199_c78 bl_78 br_78 wl_199 vdd gnd cell_6t
Xbit_r200_c78 bl_78 br_78 wl_200 vdd gnd cell_6t
Xbit_r201_c78 bl_78 br_78 wl_201 vdd gnd cell_6t
Xbit_r202_c78 bl_78 br_78 wl_202 vdd gnd cell_6t
Xbit_r203_c78 bl_78 br_78 wl_203 vdd gnd cell_6t
Xbit_r204_c78 bl_78 br_78 wl_204 vdd gnd cell_6t
Xbit_r205_c78 bl_78 br_78 wl_205 vdd gnd cell_6t
Xbit_r206_c78 bl_78 br_78 wl_206 vdd gnd cell_6t
Xbit_r207_c78 bl_78 br_78 wl_207 vdd gnd cell_6t
Xbit_r208_c78 bl_78 br_78 wl_208 vdd gnd cell_6t
Xbit_r209_c78 bl_78 br_78 wl_209 vdd gnd cell_6t
Xbit_r210_c78 bl_78 br_78 wl_210 vdd gnd cell_6t
Xbit_r211_c78 bl_78 br_78 wl_211 vdd gnd cell_6t
Xbit_r212_c78 bl_78 br_78 wl_212 vdd gnd cell_6t
Xbit_r213_c78 bl_78 br_78 wl_213 vdd gnd cell_6t
Xbit_r214_c78 bl_78 br_78 wl_214 vdd gnd cell_6t
Xbit_r215_c78 bl_78 br_78 wl_215 vdd gnd cell_6t
Xbit_r216_c78 bl_78 br_78 wl_216 vdd gnd cell_6t
Xbit_r217_c78 bl_78 br_78 wl_217 vdd gnd cell_6t
Xbit_r218_c78 bl_78 br_78 wl_218 vdd gnd cell_6t
Xbit_r219_c78 bl_78 br_78 wl_219 vdd gnd cell_6t
Xbit_r220_c78 bl_78 br_78 wl_220 vdd gnd cell_6t
Xbit_r221_c78 bl_78 br_78 wl_221 vdd gnd cell_6t
Xbit_r222_c78 bl_78 br_78 wl_222 vdd gnd cell_6t
Xbit_r223_c78 bl_78 br_78 wl_223 vdd gnd cell_6t
Xbit_r224_c78 bl_78 br_78 wl_224 vdd gnd cell_6t
Xbit_r225_c78 bl_78 br_78 wl_225 vdd gnd cell_6t
Xbit_r226_c78 bl_78 br_78 wl_226 vdd gnd cell_6t
Xbit_r227_c78 bl_78 br_78 wl_227 vdd gnd cell_6t
Xbit_r228_c78 bl_78 br_78 wl_228 vdd gnd cell_6t
Xbit_r229_c78 bl_78 br_78 wl_229 vdd gnd cell_6t
Xbit_r230_c78 bl_78 br_78 wl_230 vdd gnd cell_6t
Xbit_r231_c78 bl_78 br_78 wl_231 vdd gnd cell_6t
Xbit_r232_c78 bl_78 br_78 wl_232 vdd gnd cell_6t
Xbit_r233_c78 bl_78 br_78 wl_233 vdd gnd cell_6t
Xbit_r234_c78 bl_78 br_78 wl_234 vdd gnd cell_6t
Xbit_r235_c78 bl_78 br_78 wl_235 vdd gnd cell_6t
Xbit_r236_c78 bl_78 br_78 wl_236 vdd gnd cell_6t
Xbit_r237_c78 bl_78 br_78 wl_237 vdd gnd cell_6t
Xbit_r238_c78 bl_78 br_78 wl_238 vdd gnd cell_6t
Xbit_r239_c78 bl_78 br_78 wl_239 vdd gnd cell_6t
Xbit_r240_c78 bl_78 br_78 wl_240 vdd gnd cell_6t
Xbit_r241_c78 bl_78 br_78 wl_241 vdd gnd cell_6t
Xbit_r242_c78 bl_78 br_78 wl_242 vdd gnd cell_6t
Xbit_r243_c78 bl_78 br_78 wl_243 vdd gnd cell_6t
Xbit_r244_c78 bl_78 br_78 wl_244 vdd gnd cell_6t
Xbit_r245_c78 bl_78 br_78 wl_245 vdd gnd cell_6t
Xbit_r246_c78 bl_78 br_78 wl_246 vdd gnd cell_6t
Xbit_r247_c78 bl_78 br_78 wl_247 vdd gnd cell_6t
Xbit_r248_c78 bl_78 br_78 wl_248 vdd gnd cell_6t
Xbit_r249_c78 bl_78 br_78 wl_249 vdd gnd cell_6t
Xbit_r250_c78 bl_78 br_78 wl_250 vdd gnd cell_6t
Xbit_r251_c78 bl_78 br_78 wl_251 vdd gnd cell_6t
Xbit_r252_c78 bl_78 br_78 wl_252 vdd gnd cell_6t
Xbit_r253_c78 bl_78 br_78 wl_253 vdd gnd cell_6t
Xbit_r254_c78 bl_78 br_78 wl_254 vdd gnd cell_6t
Xbit_r255_c78 bl_78 br_78 wl_255 vdd gnd cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd cell_6t
Xbit_r1_c79 bl_79 br_79 wl_1 vdd gnd cell_6t
Xbit_r2_c79 bl_79 br_79 wl_2 vdd gnd cell_6t
Xbit_r3_c79 bl_79 br_79 wl_3 vdd gnd cell_6t
Xbit_r4_c79 bl_79 br_79 wl_4 vdd gnd cell_6t
Xbit_r5_c79 bl_79 br_79 wl_5 vdd gnd cell_6t
Xbit_r6_c79 bl_79 br_79 wl_6 vdd gnd cell_6t
Xbit_r7_c79 bl_79 br_79 wl_7 vdd gnd cell_6t
Xbit_r8_c79 bl_79 br_79 wl_8 vdd gnd cell_6t
Xbit_r9_c79 bl_79 br_79 wl_9 vdd gnd cell_6t
Xbit_r10_c79 bl_79 br_79 wl_10 vdd gnd cell_6t
Xbit_r11_c79 bl_79 br_79 wl_11 vdd gnd cell_6t
Xbit_r12_c79 bl_79 br_79 wl_12 vdd gnd cell_6t
Xbit_r13_c79 bl_79 br_79 wl_13 vdd gnd cell_6t
Xbit_r14_c79 bl_79 br_79 wl_14 vdd gnd cell_6t
Xbit_r15_c79 bl_79 br_79 wl_15 vdd gnd cell_6t
Xbit_r16_c79 bl_79 br_79 wl_16 vdd gnd cell_6t
Xbit_r17_c79 bl_79 br_79 wl_17 vdd gnd cell_6t
Xbit_r18_c79 bl_79 br_79 wl_18 vdd gnd cell_6t
Xbit_r19_c79 bl_79 br_79 wl_19 vdd gnd cell_6t
Xbit_r20_c79 bl_79 br_79 wl_20 vdd gnd cell_6t
Xbit_r21_c79 bl_79 br_79 wl_21 vdd gnd cell_6t
Xbit_r22_c79 bl_79 br_79 wl_22 vdd gnd cell_6t
Xbit_r23_c79 bl_79 br_79 wl_23 vdd gnd cell_6t
Xbit_r24_c79 bl_79 br_79 wl_24 vdd gnd cell_6t
Xbit_r25_c79 bl_79 br_79 wl_25 vdd gnd cell_6t
Xbit_r26_c79 bl_79 br_79 wl_26 vdd gnd cell_6t
Xbit_r27_c79 bl_79 br_79 wl_27 vdd gnd cell_6t
Xbit_r28_c79 bl_79 br_79 wl_28 vdd gnd cell_6t
Xbit_r29_c79 bl_79 br_79 wl_29 vdd gnd cell_6t
Xbit_r30_c79 bl_79 br_79 wl_30 vdd gnd cell_6t
Xbit_r31_c79 bl_79 br_79 wl_31 vdd gnd cell_6t
Xbit_r32_c79 bl_79 br_79 wl_32 vdd gnd cell_6t
Xbit_r33_c79 bl_79 br_79 wl_33 vdd gnd cell_6t
Xbit_r34_c79 bl_79 br_79 wl_34 vdd gnd cell_6t
Xbit_r35_c79 bl_79 br_79 wl_35 vdd gnd cell_6t
Xbit_r36_c79 bl_79 br_79 wl_36 vdd gnd cell_6t
Xbit_r37_c79 bl_79 br_79 wl_37 vdd gnd cell_6t
Xbit_r38_c79 bl_79 br_79 wl_38 vdd gnd cell_6t
Xbit_r39_c79 bl_79 br_79 wl_39 vdd gnd cell_6t
Xbit_r40_c79 bl_79 br_79 wl_40 vdd gnd cell_6t
Xbit_r41_c79 bl_79 br_79 wl_41 vdd gnd cell_6t
Xbit_r42_c79 bl_79 br_79 wl_42 vdd gnd cell_6t
Xbit_r43_c79 bl_79 br_79 wl_43 vdd gnd cell_6t
Xbit_r44_c79 bl_79 br_79 wl_44 vdd gnd cell_6t
Xbit_r45_c79 bl_79 br_79 wl_45 vdd gnd cell_6t
Xbit_r46_c79 bl_79 br_79 wl_46 vdd gnd cell_6t
Xbit_r47_c79 bl_79 br_79 wl_47 vdd gnd cell_6t
Xbit_r48_c79 bl_79 br_79 wl_48 vdd gnd cell_6t
Xbit_r49_c79 bl_79 br_79 wl_49 vdd gnd cell_6t
Xbit_r50_c79 bl_79 br_79 wl_50 vdd gnd cell_6t
Xbit_r51_c79 bl_79 br_79 wl_51 vdd gnd cell_6t
Xbit_r52_c79 bl_79 br_79 wl_52 vdd gnd cell_6t
Xbit_r53_c79 bl_79 br_79 wl_53 vdd gnd cell_6t
Xbit_r54_c79 bl_79 br_79 wl_54 vdd gnd cell_6t
Xbit_r55_c79 bl_79 br_79 wl_55 vdd gnd cell_6t
Xbit_r56_c79 bl_79 br_79 wl_56 vdd gnd cell_6t
Xbit_r57_c79 bl_79 br_79 wl_57 vdd gnd cell_6t
Xbit_r58_c79 bl_79 br_79 wl_58 vdd gnd cell_6t
Xbit_r59_c79 bl_79 br_79 wl_59 vdd gnd cell_6t
Xbit_r60_c79 bl_79 br_79 wl_60 vdd gnd cell_6t
Xbit_r61_c79 bl_79 br_79 wl_61 vdd gnd cell_6t
Xbit_r62_c79 bl_79 br_79 wl_62 vdd gnd cell_6t
Xbit_r63_c79 bl_79 br_79 wl_63 vdd gnd cell_6t
Xbit_r64_c79 bl_79 br_79 wl_64 vdd gnd cell_6t
Xbit_r65_c79 bl_79 br_79 wl_65 vdd gnd cell_6t
Xbit_r66_c79 bl_79 br_79 wl_66 vdd gnd cell_6t
Xbit_r67_c79 bl_79 br_79 wl_67 vdd gnd cell_6t
Xbit_r68_c79 bl_79 br_79 wl_68 vdd gnd cell_6t
Xbit_r69_c79 bl_79 br_79 wl_69 vdd gnd cell_6t
Xbit_r70_c79 bl_79 br_79 wl_70 vdd gnd cell_6t
Xbit_r71_c79 bl_79 br_79 wl_71 vdd gnd cell_6t
Xbit_r72_c79 bl_79 br_79 wl_72 vdd gnd cell_6t
Xbit_r73_c79 bl_79 br_79 wl_73 vdd gnd cell_6t
Xbit_r74_c79 bl_79 br_79 wl_74 vdd gnd cell_6t
Xbit_r75_c79 bl_79 br_79 wl_75 vdd gnd cell_6t
Xbit_r76_c79 bl_79 br_79 wl_76 vdd gnd cell_6t
Xbit_r77_c79 bl_79 br_79 wl_77 vdd gnd cell_6t
Xbit_r78_c79 bl_79 br_79 wl_78 vdd gnd cell_6t
Xbit_r79_c79 bl_79 br_79 wl_79 vdd gnd cell_6t
Xbit_r80_c79 bl_79 br_79 wl_80 vdd gnd cell_6t
Xbit_r81_c79 bl_79 br_79 wl_81 vdd gnd cell_6t
Xbit_r82_c79 bl_79 br_79 wl_82 vdd gnd cell_6t
Xbit_r83_c79 bl_79 br_79 wl_83 vdd gnd cell_6t
Xbit_r84_c79 bl_79 br_79 wl_84 vdd gnd cell_6t
Xbit_r85_c79 bl_79 br_79 wl_85 vdd gnd cell_6t
Xbit_r86_c79 bl_79 br_79 wl_86 vdd gnd cell_6t
Xbit_r87_c79 bl_79 br_79 wl_87 vdd gnd cell_6t
Xbit_r88_c79 bl_79 br_79 wl_88 vdd gnd cell_6t
Xbit_r89_c79 bl_79 br_79 wl_89 vdd gnd cell_6t
Xbit_r90_c79 bl_79 br_79 wl_90 vdd gnd cell_6t
Xbit_r91_c79 bl_79 br_79 wl_91 vdd gnd cell_6t
Xbit_r92_c79 bl_79 br_79 wl_92 vdd gnd cell_6t
Xbit_r93_c79 bl_79 br_79 wl_93 vdd gnd cell_6t
Xbit_r94_c79 bl_79 br_79 wl_94 vdd gnd cell_6t
Xbit_r95_c79 bl_79 br_79 wl_95 vdd gnd cell_6t
Xbit_r96_c79 bl_79 br_79 wl_96 vdd gnd cell_6t
Xbit_r97_c79 bl_79 br_79 wl_97 vdd gnd cell_6t
Xbit_r98_c79 bl_79 br_79 wl_98 vdd gnd cell_6t
Xbit_r99_c79 bl_79 br_79 wl_99 vdd gnd cell_6t
Xbit_r100_c79 bl_79 br_79 wl_100 vdd gnd cell_6t
Xbit_r101_c79 bl_79 br_79 wl_101 vdd gnd cell_6t
Xbit_r102_c79 bl_79 br_79 wl_102 vdd gnd cell_6t
Xbit_r103_c79 bl_79 br_79 wl_103 vdd gnd cell_6t
Xbit_r104_c79 bl_79 br_79 wl_104 vdd gnd cell_6t
Xbit_r105_c79 bl_79 br_79 wl_105 vdd gnd cell_6t
Xbit_r106_c79 bl_79 br_79 wl_106 vdd gnd cell_6t
Xbit_r107_c79 bl_79 br_79 wl_107 vdd gnd cell_6t
Xbit_r108_c79 bl_79 br_79 wl_108 vdd gnd cell_6t
Xbit_r109_c79 bl_79 br_79 wl_109 vdd gnd cell_6t
Xbit_r110_c79 bl_79 br_79 wl_110 vdd gnd cell_6t
Xbit_r111_c79 bl_79 br_79 wl_111 vdd gnd cell_6t
Xbit_r112_c79 bl_79 br_79 wl_112 vdd gnd cell_6t
Xbit_r113_c79 bl_79 br_79 wl_113 vdd gnd cell_6t
Xbit_r114_c79 bl_79 br_79 wl_114 vdd gnd cell_6t
Xbit_r115_c79 bl_79 br_79 wl_115 vdd gnd cell_6t
Xbit_r116_c79 bl_79 br_79 wl_116 vdd gnd cell_6t
Xbit_r117_c79 bl_79 br_79 wl_117 vdd gnd cell_6t
Xbit_r118_c79 bl_79 br_79 wl_118 vdd gnd cell_6t
Xbit_r119_c79 bl_79 br_79 wl_119 vdd gnd cell_6t
Xbit_r120_c79 bl_79 br_79 wl_120 vdd gnd cell_6t
Xbit_r121_c79 bl_79 br_79 wl_121 vdd gnd cell_6t
Xbit_r122_c79 bl_79 br_79 wl_122 vdd gnd cell_6t
Xbit_r123_c79 bl_79 br_79 wl_123 vdd gnd cell_6t
Xbit_r124_c79 bl_79 br_79 wl_124 vdd gnd cell_6t
Xbit_r125_c79 bl_79 br_79 wl_125 vdd gnd cell_6t
Xbit_r126_c79 bl_79 br_79 wl_126 vdd gnd cell_6t
Xbit_r127_c79 bl_79 br_79 wl_127 vdd gnd cell_6t
Xbit_r128_c79 bl_79 br_79 wl_128 vdd gnd cell_6t
Xbit_r129_c79 bl_79 br_79 wl_129 vdd gnd cell_6t
Xbit_r130_c79 bl_79 br_79 wl_130 vdd gnd cell_6t
Xbit_r131_c79 bl_79 br_79 wl_131 vdd gnd cell_6t
Xbit_r132_c79 bl_79 br_79 wl_132 vdd gnd cell_6t
Xbit_r133_c79 bl_79 br_79 wl_133 vdd gnd cell_6t
Xbit_r134_c79 bl_79 br_79 wl_134 vdd gnd cell_6t
Xbit_r135_c79 bl_79 br_79 wl_135 vdd gnd cell_6t
Xbit_r136_c79 bl_79 br_79 wl_136 vdd gnd cell_6t
Xbit_r137_c79 bl_79 br_79 wl_137 vdd gnd cell_6t
Xbit_r138_c79 bl_79 br_79 wl_138 vdd gnd cell_6t
Xbit_r139_c79 bl_79 br_79 wl_139 vdd gnd cell_6t
Xbit_r140_c79 bl_79 br_79 wl_140 vdd gnd cell_6t
Xbit_r141_c79 bl_79 br_79 wl_141 vdd gnd cell_6t
Xbit_r142_c79 bl_79 br_79 wl_142 vdd gnd cell_6t
Xbit_r143_c79 bl_79 br_79 wl_143 vdd gnd cell_6t
Xbit_r144_c79 bl_79 br_79 wl_144 vdd gnd cell_6t
Xbit_r145_c79 bl_79 br_79 wl_145 vdd gnd cell_6t
Xbit_r146_c79 bl_79 br_79 wl_146 vdd gnd cell_6t
Xbit_r147_c79 bl_79 br_79 wl_147 vdd gnd cell_6t
Xbit_r148_c79 bl_79 br_79 wl_148 vdd gnd cell_6t
Xbit_r149_c79 bl_79 br_79 wl_149 vdd gnd cell_6t
Xbit_r150_c79 bl_79 br_79 wl_150 vdd gnd cell_6t
Xbit_r151_c79 bl_79 br_79 wl_151 vdd gnd cell_6t
Xbit_r152_c79 bl_79 br_79 wl_152 vdd gnd cell_6t
Xbit_r153_c79 bl_79 br_79 wl_153 vdd gnd cell_6t
Xbit_r154_c79 bl_79 br_79 wl_154 vdd gnd cell_6t
Xbit_r155_c79 bl_79 br_79 wl_155 vdd gnd cell_6t
Xbit_r156_c79 bl_79 br_79 wl_156 vdd gnd cell_6t
Xbit_r157_c79 bl_79 br_79 wl_157 vdd gnd cell_6t
Xbit_r158_c79 bl_79 br_79 wl_158 vdd gnd cell_6t
Xbit_r159_c79 bl_79 br_79 wl_159 vdd gnd cell_6t
Xbit_r160_c79 bl_79 br_79 wl_160 vdd gnd cell_6t
Xbit_r161_c79 bl_79 br_79 wl_161 vdd gnd cell_6t
Xbit_r162_c79 bl_79 br_79 wl_162 vdd gnd cell_6t
Xbit_r163_c79 bl_79 br_79 wl_163 vdd gnd cell_6t
Xbit_r164_c79 bl_79 br_79 wl_164 vdd gnd cell_6t
Xbit_r165_c79 bl_79 br_79 wl_165 vdd gnd cell_6t
Xbit_r166_c79 bl_79 br_79 wl_166 vdd gnd cell_6t
Xbit_r167_c79 bl_79 br_79 wl_167 vdd gnd cell_6t
Xbit_r168_c79 bl_79 br_79 wl_168 vdd gnd cell_6t
Xbit_r169_c79 bl_79 br_79 wl_169 vdd gnd cell_6t
Xbit_r170_c79 bl_79 br_79 wl_170 vdd gnd cell_6t
Xbit_r171_c79 bl_79 br_79 wl_171 vdd gnd cell_6t
Xbit_r172_c79 bl_79 br_79 wl_172 vdd gnd cell_6t
Xbit_r173_c79 bl_79 br_79 wl_173 vdd gnd cell_6t
Xbit_r174_c79 bl_79 br_79 wl_174 vdd gnd cell_6t
Xbit_r175_c79 bl_79 br_79 wl_175 vdd gnd cell_6t
Xbit_r176_c79 bl_79 br_79 wl_176 vdd gnd cell_6t
Xbit_r177_c79 bl_79 br_79 wl_177 vdd gnd cell_6t
Xbit_r178_c79 bl_79 br_79 wl_178 vdd gnd cell_6t
Xbit_r179_c79 bl_79 br_79 wl_179 vdd gnd cell_6t
Xbit_r180_c79 bl_79 br_79 wl_180 vdd gnd cell_6t
Xbit_r181_c79 bl_79 br_79 wl_181 vdd gnd cell_6t
Xbit_r182_c79 bl_79 br_79 wl_182 vdd gnd cell_6t
Xbit_r183_c79 bl_79 br_79 wl_183 vdd gnd cell_6t
Xbit_r184_c79 bl_79 br_79 wl_184 vdd gnd cell_6t
Xbit_r185_c79 bl_79 br_79 wl_185 vdd gnd cell_6t
Xbit_r186_c79 bl_79 br_79 wl_186 vdd gnd cell_6t
Xbit_r187_c79 bl_79 br_79 wl_187 vdd gnd cell_6t
Xbit_r188_c79 bl_79 br_79 wl_188 vdd gnd cell_6t
Xbit_r189_c79 bl_79 br_79 wl_189 vdd gnd cell_6t
Xbit_r190_c79 bl_79 br_79 wl_190 vdd gnd cell_6t
Xbit_r191_c79 bl_79 br_79 wl_191 vdd gnd cell_6t
Xbit_r192_c79 bl_79 br_79 wl_192 vdd gnd cell_6t
Xbit_r193_c79 bl_79 br_79 wl_193 vdd gnd cell_6t
Xbit_r194_c79 bl_79 br_79 wl_194 vdd gnd cell_6t
Xbit_r195_c79 bl_79 br_79 wl_195 vdd gnd cell_6t
Xbit_r196_c79 bl_79 br_79 wl_196 vdd gnd cell_6t
Xbit_r197_c79 bl_79 br_79 wl_197 vdd gnd cell_6t
Xbit_r198_c79 bl_79 br_79 wl_198 vdd gnd cell_6t
Xbit_r199_c79 bl_79 br_79 wl_199 vdd gnd cell_6t
Xbit_r200_c79 bl_79 br_79 wl_200 vdd gnd cell_6t
Xbit_r201_c79 bl_79 br_79 wl_201 vdd gnd cell_6t
Xbit_r202_c79 bl_79 br_79 wl_202 vdd gnd cell_6t
Xbit_r203_c79 bl_79 br_79 wl_203 vdd gnd cell_6t
Xbit_r204_c79 bl_79 br_79 wl_204 vdd gnd cell_6t
Xbit_r205_c79 bl_79 br_79 wl_205 vdd gnd cell_6t
Xbit_r206_c79 bl_79 br_79 wl_206 vdd gnd cell_6t
Xbit_r207_c79 bl_79 br_79 wl_207 vdd gnd cell_6t
Xbit_r208_c79 bl_79 br_79 wl_208 vdd gnd cell_6t
Xbit_r209_c79 bl_79 br_79 wl_209 vdd gnd cell_6t
Xbit_r210_c79 bl_79 br_79 wl_210 vdd gnd cell_6t
Xbit_r211_c79 bl_79 br_79 wl_211 vdd gnd cell_6t
Xbit_r212_c79 bl_79 br_79 wl_212 vdd gnd cell_6t
Xbit_r213_c79 bl_79 br_79 wl_213 vdd gnd cell_6t
Xbit_r214_c79 bl_79 br_79 wl_214 vdd gnd cell_6t
Xbit_r215_c79 bl_79 br_79 wl_215 vdd gnd cell_6t
Xbit_r216_c79 bl_79 br_79 wl_216 vdd gnd cell_6t
Xbit_r217_c79 bl_79 br_79 wl_217 vdd gnd cell_6t
Xbit_r218_c79 bl_79 br_79 wl_218 vdd gnd cell_6t
Xbit_r219_c79 bl_79 br_79 wl_219 vdd gnd cell_6t
Xbit_r220_c79 bl_79 br_79 wl_220 vdd gnd cell_6t
Xbit_r221_c79 bl_79 br_79 wl_221 vdd gnd cell_6t
Xbit_r222_c79 bl_79 br_79 wl_222 vdd gnd cell_6t
Xbit_r223_c79 bl_79 br_79 wl_223 vdd gnd cell_6t
Xbit_r224_c79 bl_79 br_79 wl_224 vdd gnd cell_6t
Xbit_r225_c79 bl_79 br_79 wl_225 vdd gnd cell_6t
Xbit_r226_c79 bl_79 br_79 wl_226 vdd gnd cell_6t
Xbit_r227_c79 bl_79 br_79 wl_227 vdd gnd cell_6t
Xbit_r228_c79 bl_79 br_79 wl_228 vdd gnd cell_6t
Xbit_r229_c79 bl_79 br_79 wl_229 vdd gnd cell_6t
Xbit_r230_c79 bl_79 br_79 wl_230 vdd gnd cell_6t
Xbit_r231_c79 bl_79 br_79 wl_231 vdd gnd cell_6t
Xbit_r232_c79 bl_79 br_79 wl_232 vdd gnd cell_6t
Xbit_r233_c79 bl_79 br_79 wl_233 vdd gnd cell_6t
Xbit_r234_c79 bl_79 br_79 wl_234 vdd gnd cell_6t
Xbit_r235_c79 bl_79 br_79 wl_235 vdd gnd cell_6t
Xbit_r236_c79 bl_79 br_79 wl_236 vdd gnd cell_6t
Xbit_r237_c79 bl_79 br_79 wl_237 vdd gnd cell_6t
Xbit_r238_c79 bl_79 br_79 wl_238 vdd gnd cell_6t
Xbit_r239_c79 bl_79 br_79 wl_239 vdd gnd cell_6t
Xbit_r240_c79 bl_79 br_79 wl_240 vdd gnd cell_6t
Xbit_r241_c79 bl_79 br_79 wl_241 vdd gnd cell_6t
Xbit_r242_c79 bl_79 br_79 wl_242 vdd gnd cell_6t
Xbit_r243_c79 bl_79 br_79 wl_243 vdd gnd cell_6t
Xbit_r244_c79 bl_79 br_79 wl_244 vdd gnd cell_6t
Xbit_r245_c79 bl_79 br_79 wl_245 vdd gnd cell_6t
Xbit_r246_c79 bl_79 br_79 wl_246 vdd gnd cell_6t
Xbit_r247_c79 bl_79 br_79 wl_247 vdd gnd cell_6t
Xbit_r248_c79 bl_79 br_79 wl_248 vdd gnd cell_6t
Xbit_r249_c79 bl_79 br_79 wl_249 vdd gnd cell_6t
Xbit_r250_c79 bl_79 br_79 wl_250 vdd gnd cell_6t
Xbit_r251_c79 bl_79 br_79 wl_251 vdd gnd cell_6t
Xbit_r252_c79 bl_79 br_79 wl_252 vdd gnd cell_6t
Xbit_r253_c79 bl_79 br_79 wl_253 vdd gnd cell_6t
Xbit_r254_c79 bl_79 br_79 wl_254 vdd gnd cell_6t
Xbit_r255_c79 bl_79 br_79 wl_255 vdd gnd cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd cell_6t
Xbit_r1_c80 bl_80 br_80 wl_1 vdd gnd cell_6t
Xbit_r2_c80 bl_80 br_80 wl_2 vdd gnd cell_6t
Xbit_r3_c80 bl_80 br_80 wl_3 vdd gnd cell_6t
Xbit_r4_c80 bl_80 br_80 wl_4 vdd gnd cell_6t
Xbit_r5_c80 bl_80 br_80 wl_5 vdd gnd cell_6t
Xbit_r6_c80 bl_80 br_80 wl_6 vdd gnd cell_6t
Xbit_r7_c80 bl_80 br_80 wl_7 vdd gnd cell_6t
Xbit_r8_c80 bl_80 br_80 wl_8 vdd gnd cell_6t
Xbit_r9_c80 bl_80 br_80 wl_9 vdd gnd cell_6t
Xbit_r10_c80 bl_80 br_80 wl_10 vdd gnd cell_6t
Xbit_r11_c80 bl_80 br_80 wl_11 vdd gnd cell_6t
Xbit_r12_c80 bl_80 br_80 wl_12 vdd gnd cell_6t
Xbit_r13_c80 bl_80 br_80 wl_13 vdd gnd cell_6t
Xbit_r14_c80 bl_80 br_80 wl_14 vdd gnd cell_6t
Xbit_r15_c80 bl_80 br_80 wl_15 vdd gnd cell_6t
Xbit_r16_c80 bl_80 br_80 wl_16 vdd gnd cell_6t
Xbit_r17_c80 bl_80 br_80 wl_17 vdd gnd cell_6t
Xbit_r18_c80 bl_80 br_80 wl_18 vdd gnd cell_6t
Xbit_r19_c80 bl_80 br_80 wl_19 vdd gnd cell_6t
Xbit_r20_c80 bl_80 br_80 wl_20 vdd gnd cell_6t
Xbit_r21_c80 bl_80 br_80 wl_21 vdd gnd cell_6t
Xbit_r22_c80 bl_80 br_80 wl_22 vdd gnd cell_6t
Xbit_r23_c80 bl_80 br_80 wl_23 vdd gnd cell_6t
Xbit_r24_c80 bl_80 br_80 wl_24 vdd gnd cell_6t
Xbit_r25_c80 bl_80 br_80 wl_25 vdd gnd cell_6t
Xbit_r26_c80 bl_80 br_80 wl_26 vdd gnd cell_6t
Xbit_r27_c80 bl_80 br_80 wl_27 vdd gnd cell_6t
Xbit_r28_c80 bl_80 br_80 wl_28 vdd gnd cell_6t
Xbit_r29_c80 bl_80 br_80 wl_29 vdd gnd cell_6t
Xbit_r30_c80 bl_80 br_80 wl_30 vdd gnd cell_6t
Xbit_r31_c80 bl_80 br_80 wl_31 vdd gnd cell_6t
Xbit_r32_c80 bl_80 br_80 wl_32 vdd gnd cell_6t
Xbit_r33_c80 bl_80 br_80 wl_33 vdd gnd cell_6t
Xbit_r34_c80 bl_80 br_80 wl_34 vdd gnd cell_6t
Xbit_r35_c80 bl_80 br_80 wl_35 vdd gnd cell_6t
Xbit_r36_c80 bl_80 br_80 wl_36 vdd gnd cell_6t
Xbit_r37_c80 bl_80 br_80 wl_37 vdd gnd cell_6t
Xbit_r38_c80 bl_80 br_80 wl_38 vdd gnd cell_6t
Xbit_r39_c80 bl_80 br_80 wl_39 vdd gnd cell_6t
Xbit_r40_c80 bl_80 br_80 wl_40 vdd gnd cell_6t
Xbit_r41_c80 bl_80 br_80 wl_41 vdd gnd cell_6t
Xbit_r42_c80 bl_80 br_80 wl_42 vdd gnd cell_6t
Xbit_r43_c80 bl_80 br_80 wl_43 vdd gnd cell_6t
Xbit_r44_c80 bl_80 br_80 wl_44 vdd gnd cell_6t
Xbit_r45_c80 bl_80 br_80 wl_45 vdd gnd cell_6t
Xbit_r46_c80 bl_80 br_80 wl_46 vdd gnd cell_6t
Xbit_r47_c80 bl_80 br_80 wl_47 vdd gnd cell_6t
Xbit_r48_c80 bl_80 br_80 wl_48 vdd gnd cell_6t
Xbit_r49_c80 bl_80 br_80 wl_49 vdd gnd cell_6t
Xbit_r50_c80 bl_80 br_80 wl_50 vdd gnd cell_6t
Xbit_r51_c80 bl_80 br_80 wl_51 vdd gnd cell_6t
Xbit_r52_c80 bl_80 br_80 wl_52 vdd gnd cell_6t
Xbit_r53_c80 bl_80 br_80 wl_53 vdd gnd cell_6t
Xbit_r54_c80 bl_80 br_80 wl_54 vdd gnd cell_6t
Xbit_r55_c80 bl_80 br_80 wl_55 vdd gnd cell_6t
Xbit_r56_c80 bl_80 br_80 wl_56 vdd gnd cell_6t
Xbit_r57_c80 bl_80 br_80 wl_57 vdd gnd cell_6t
Xbit_r58_c80 bl_80 br_80 wl_58 vdd gnd cell_6t
Xbit_r59_c80 bl_80 br_80 wl_59 vdd gnd cell_6t
Xbit_r60_c80 bl_80 br_80 wl_60 vdd gnd cell_6t
Xbit_r61_c80 bl_80 br_80 wl_61 vdd gnd cell_6t
Xbit_r62_c80 bl_80 br_80 wl_62 vdd gnd cell_6t
Xbit_r63_c80 bl_80 br_80 wl_63 vdd gnd cell_6t
Xbit_r64_c80 bl_80 br_80 wl_64 vdd gnd cell_6t
Xbit_r65_c80 bl_80 br_80 wl_65 vdd gnd cell_6t
Xbit_r66_c80 bl_80 br_80 wl_66 vdd gnd cell_6t
Xbit_r67_c80 bl_80 br_80 wl_67 vdd gnd cell_6t
Xbit_r68_c80 bl_80 br_80 wl_68 vdd gnd cell_6t
Xbit_r69_c80 bl_80 br_80 wl_69 vdd gnd cell_6t
Xbit_r70_c80 bl_80 br_80 wl_70 vdd gnd cell_6t
Xbit_r71_c80 bl_80 br_80 wl_71 vdd gnd cell_6t
Xbit_r72_c80 bl_80 br_80 wl_72 vdd gnd cell_6t
Xbit_r73_c80 bl_80 br_80 wl_73 vdd gnd cell_6t
Xbit_r74_c80 bl_80 br_80 wl_74 vdd gnd cell_6t
Xbit_r75_c80 bl_80 br_80 wl_75 vdd gnd cell_6t
Xbit_r76_c80 bl_80 br_80 wl_76 vdd gnd cell_6t
Xbit_r77_c80 bl_80 br_80 wl_77 vdd gnd cell_6t
Xbit_r78_c80 bl_80 br_80 wl_78 vdd gnd cell_6t
Xbit_r79_c80 bl_80 br_80 wl_79 vdd gnd cell_6t
Xbit_r80_c80 bl_80 br_80 wl_80 vdd gnd cell_6t
Xbit_r81_c80 bl_80 br_80 wl_81 vdd gnd cell_6t
Xbit_r82_c80 bl_80 br_80 wl_82 vdd gnd cell_6t
Xbit_r83_c80 bl_80 br_80 wl_83 vdd gnd cell_6t
Xbit_r84_c80 bl_80 br_80 wl_84 vdd gnd cell_6t
Xbit_r85_c80 bl_80 br_80 wl_85 vdd gnd cell_6t
Xbit_r86_c80 bl_80 br_80 wl_86 vdd gnd cell_6t
Xbit_r87_c80 bl_80 br_80 wl_87 vdd gnd cell_6t
Xbit_r88_c80 bl_80 br_80 wl_88 vdd gnd cell_6t
Xbit_r89_c80 bl_80 br_80 wl_89 vdd gnd cell_6t
Xbit_r90_c80 bl_80 br_80 wl_90 vdd gnd cell_6t
Xbit_r91_c80 bl_80 br_80 wl_91 vdd gnd cell_6t
Xbit_r92_c80 bl_80 br_80 wl_92 vdd gnd cell_6t
Xbit_r93_c80 bl_80 br_80 wl_93 vdd gnd cell_6t
Xbit_r94_c80 bl_80 br_80 wl_94 vdd gnd cell_6t
Xbit_r95_c80 bl_80 br_80 wl_95 vdd gnd cell_6t
Xbit_r96_c80 bl_80 br_80 wl_96 vdd gnd cell_6t
Xbit_r97_c80 bl_80 br_80 wl_97 vdd gnd cell_6t
Xbit_r98_c80 bl_80 br_80 wl_98 vdd gnd cell_6t
Xbit_r99_c80 bl_80 br_80 wl_99 vdd gnd cell_6t
Xbit_r100_c80 bl_80 br_80 wl_100 vdd gnd cell_6t
Xbit_r101_c80 bl_80 br_80 wl_101 vdd gnd cell_6t
Xbit_r102_c80 bl_80 br_80 wl_102 vdd gnd cell_6t
Xbit_r103_c80 bl_80 br_80 wl_103 vdd gnd cell_6t
Xbit_r104_c80 bl_80 br_80 wl_104 vdd gnd cell_6t
Xbit_r105_c80 bl_80 br_80 wl_105 vdd gnd cell_6t
Xbit_r106_c80 bl_80 br_80 wl_106 vdd gnd cell_6t
Xbit_r107_c80 bl_80 br_80 wl_107 vdd gnd cell_6t
Xbit_r108_c80 bl_80 br_80 wl_108 vdd gnd cell_6t
Xbit_r109_c80 bl_80 br_80 wl_109 vdd gnd cell_6t
Xbit_r110_c80 bl_80 br_80 wl_110 vdd gnd cell_6t
Xbit_r111_c80 bl_80 br_80 wl_111 vdd gnd cell_6t
Xbit_r112_c80 bl_80 br_80 wl_112 vdd gnd cell_6t
Xbit_r113_c80 bl_80 br_80 wl_113 vdd gnd cell_6t
Xbit_r114_c80 bl_80 br_80 wl_114 vdd gnd cell_6t
Xbit_r115_c80 bl_80 br_80 wl_115 vdd gnd cell_6t
Xbit_r116_c80 bl_80 br_80 wl_116 vdd gnd cell_6t
Xbit_r117_c80 bl_80 br_80 wl_117 vdd gnd cell_6t
Xbit_r118_c80 bl_80 br_80 wl_118 vdd gnd cell_6t
Xbit_r119_c80 bl_80 br_80 wl_119 vdd gnd cell_6t
Xbit_r120_c80 bl_80 br_80 wl_120 vdd gnd cell_6t
Xbit_r121_c80 bl_80 br_80 wl_121 vdd gnd cell_6t
Xbit_r122_c80 bl_80 br_80 wl_122 vdd gnd cell_6t
Xbit_r123_c80 bl_80 br_80 wl_123 vdd gnd cell_6t
Xbit_r124_c80 bl_80 br_80 wl_124 vdd gnd cell_6t
Xbit_r125_c80 bl_80 br_80 wl_125 vdd gnd cell_6t
Xbit_r126_c80 bl_80 br_80 wl_126 vdd gnd cell_6t
Xbit_r127_c80 bl_80 br_80 wl_127 vdd gnd cell_6t
Xbit_r128_c80 bl_80 br_80 wl_128 vdd gnd cell_6t
Xbit_r129_c80 bl_80 br_80 wl_129 vdd gnd cell_6t
Xbit_r130_c80 bl_80 br_80 wl_130 vdd gnd cell_6t
Xbit_r131_c80 bl_80 br_80 wl_131 vdd gnd cell_6t
Xbit_r132_c80 bl_80 br_80 wl_132 vdd gnd cell_6t
Xbit_r133_c80 bl_80 br_80 wl_133 vdd gnd cell_6t
Xbit_r134_c80 bl_80 br_80 wl_134 vdd gnd cell_6t
Xbit_r135_c80 bl_80 br_80 wl_135 vdd gnd cell_6t
Xbit_r136_c80 bl_80 br_80 wl_136 vdd gnd cell_6t
Xbit_r137_c80 bl_80 br_80 wl_137 vdd gnd cell_6t
Xbit_r138_c80 bl_80 br_80 wl_138 vdd gnd cell_6t
Xbit_r139_c80 bl_80 br_80 wl_139 vdd gnd cell_6t
Xbit_r140_c80 bl_80 br_80 wl_140 vdd gnd cell_6t
Xbit_r141_c80 bl_80 br_80 wl_141 vdd gnd cell_6t
Xbit_r142_c80 bl_80 br_80 wl_142 vdd gnd cell_6t
Xbit_r143_c80 bl_80 br_80 wl_143 vdd gnd cell_6t
Xbit_r144_c80 bl_80 br_80 wl_144 vdd gnd cell_6t
Xbit_r145_c80 bl_80 br_80 wl_145 vdd gnd cell_6t
Xbit_r146_c80 bl_80 br_80 wl_146 vdd gnd cell_6t
Xbit_r147_c80 bl_80 br_80 wl_147 vdd gnd cell_6t
Xbit_r148_c80 bl_80 br_80 wl_148 vdd gnd cell_6t
Xbit_r149_c80 bl_80 br_80 wl_149 vdd gnd cell_6t
Xbit_r150_c80 bl_80 br_80 wl_150 vdd gnd cell_6t
Xbit_r151_c80 bl_80 br_80 wl_151 vdd gnd cell_6t
Xbit_r152_c80 bl_80 br_80 wl_152 vdd gnd cell_6t
Xbit_r153_c80 bl_80 br_80 wl_153 vdd gnd cell_6t
Xbit_r154_c80 bl_80 br_80 wl_154 vdd gnd cell_6t
Xbit_r155_c80 bl_80 br_80 wl_155 vdd gnd cell_6t
Xbit_r156_c80 bl_80 br_80 wl_156 vdd gnd cell_6t
Xbit_r157_c80 bl_80 br_80 wl_157 vdd gnd cell_6t
Xbit_r158_c80 bl_80 br_80 wl_158 vdd gnd cell_6t
Xbit_r159_c80 bl_80 br_80 wl_159 vdd gnd cell_6t
Xbit_r160_c80 bl_80 br_80 wl_160 vdd gnd cell_6t
Xbit_r161_c80 bl_80 br_80 wl_161 vdd gnd cell_6t
Xbit_r162_c80 bl_80 br_80 wl_162 vdd gnd cell_6t
Xbit_r163_c80 bl_80 br_80 wl_163 vdd gnd cell_6t
Xbit_r164_c80 bl_80 br_80 wl_164 vdd gnd cell_6t
Xbit_r165_c80 bl_80 br_80 wl_165 vdd gnd cell_6t
Xbit_r166_c80 bl_80 br_80 wl_166 vdd gnd cell_6t
Xbit_r167_c80 bl_80 br_80 wl_167 vdd gnd cell_6t
Xbit_r168_c80 bl_80 br_80 wl_168 vdd gnd cell_6t
Xbit_r169_c80 bl_80 br_80 wl_169 vdd gnd cell_6t
Xbit_r170_c80 bl_80 br_80 wl_170 vdd gnd cell_6t
Xbit_r171_c80 bl_80 br_80 wl_171 vdd gnd cell_6t
Xbit_r172_c80 bl_80 br_80 wl_172 vdd gnd cell_6t
Xbit_r173_c80 bl_80 br_80 wl_173 vdd gnd cell_6t
Xbit_r174_c80 bl_80 br_80 wl_174 vdd gnd cell_6t
Xbit_r175_c80 bl_80 br_80 wl_175 vdd gnd cell_6t
Xbit_r176_c80 bl_80 br_80 wl_176 vdd gnd cell_6t
Xbit_r177_c80 bl_80 br_80 wl_177 vdd gnd cell_6t
Xbit_r178_c80 bl_80 br_80 wl_178 vdd gnd cell_6t
Xbit_r179_c80 bl_80 br_80 wl_179 vdd gnd cell_6t
Xbit_r180_c80 bl_80 br_80 wl_180 vdd gnd cell_6t
Xbit_r181_c80 bl_80 br_80 wl_181 vdd gnd cell_6t
Xbit_r182_c80 bl_80 br_80 wl_182 vdd gnd cell_6t
Xbit_r183_c80 bl_80 br_80 wl_183 vdd gnd cell_6t
Xbit_r184_c80 bl_80 br_80 wl_184 vdd gnd cell_6t
Xbit_r185_c80 bl_80 br_80 wl_185 vdd gnd cell_6t
Xbit_r186_c80 bl_80 br_80 wl_186 vdd gnd cell_6t
Xbit_r187_c80 bl_80 br_80 wl_187 vdd gnd cell_6t
Xbit_r188_c80 bl_80 br_80 wl_188 vdd gnd cell_6t
Xbit_r189_c80 bl_80 br_80 wl_189 vdd gnd cell_6t
Xbit_r190_c80 bl_80 br_80 wl_190 vdd gnd cell_6t
Xbit_r191_c80 bl_80 br_80 wl_191 vdd gnd cell_6t
Xbit_r192_c80 bl_80 br_80 wl_192 vdd gnd cell_6t
Xbit_r193_c80 bl_80 br_80 wl_193 vdd gnd cell_6t
Xbit_r194_c80 bl_80 br_80 wl_194 vdd gnd cell_6t
Xbit_r195_c80 bl_80 br_80 wl_195 vdd gnd cell_6t
Xbit_r196_c80 bl_80 br_80 wl_196 vdd gnd cell_6t
Xbit_r197_c80 bl_80 br_80 wl_197 vdd gnd cell_6t
Xbit_r198_c80 bl_80 br_80 wl_198 vdd gnd cell_6t
Xbit_r199_c80 bl_80 br_80 wl_199 vdd gnd cell_6t
Xbit_r200_c80 bl_80 br_80 wl_200 vdd gnd cell_6t
Xbit_r201_c80 bl_80 br_80 wl_201 vdd gnd cell_6t
Xbit_r202_c80 bl_80 br_80 wl_202 vdd gnd cell_6t
Xbit_r203_c80 bl_80 br_80 wl_203 vdd gnd cell_6t
Xbit_r204_c80 bl_80 br_80 wl_204 vdd gnd cell_6t
Xbit_r205_c80 bl_80 br_80 wl_205 vdd gnd cell_6t
Xbit_r206_c80 bl_80 br_80 wl_206 vdd gnd cell_6t
Xbit_r207_c80 bl_80 br_80 wl_207 vdd gnd cell_6t
Xbit_r208_c80 bl_80 br_80 wl_208 vdd gnd cell_6t
Xbit_r209_c80 bl_80 br_80 wl_209 vdd gnd cell_6t
Xbit_r210_c80 bl_80 br_80 wl_210 vdd gnd cell_6t
Xbit_r211_c80 bl_80 br_80 wl_211 vdd gnd cell_6t
Xbit_r212_c80 bl_80 br_80 wl_212 vdd gnd cell_6t
Xbit_r213_c80 bl_80 br_80 wl_213 vdd gnd cell_6t
Xbit_r214_c80 bl_80 br_80 wl_214 vdd gnd cell_6t
Xbit_r215_c80 bl_80 br_80 wl_215 vdd gnd cell_6t
Xbit_r216_c80 bl_80 br_80 wl_216 vdd gnd cell_6t
Xbit_r217_c80 bl_80 br_80 wl_217 vdd gnd cell_6t
Xbit_r218_c80 bl_80 br_80 wl_218 vdd gnd cell_6t
Xbit_r219_c80 bl_80 br_80 wl_219 vdd gnd cell_6t
Xbit_r220_c80 bl_80 br_80 wl_220 vdd gnd cell_6t
Xbit_r221_c80 bl_80 br_80 wl_221 vdd gnd cell_6t
Xbit_r222_c80 bl_80 br_80 wl_222 vdd gnd cell_6t
Xbit_r223_c80 bl_80 br_80 wl_223 vdd gnd cell_6t
Xbit_r224_c80 bl_80 br_80 wl_224 vdd gnd cell_6t
Xbit_r225_c80 bl_80 br_80 wl_225 vdd gnd cell_6t
Xbit_r226_c80 bl_80 br_80 wl_226 vdd gnd cell_6t
Xbit_r227_c80 bl_80 br_80 wl_227 vdd gnd cell_6t
Xbit_r228_c80 bl_80 br_80 wl_228 vdd gnd cell_6t
Xbit_r229_c80 bl_80 br_80 wl_229 vdd gnd cell_6t
Xbit_r230_c80 bl_80 br_80 wl_230 vdd gnd cell_6t
Xbit_r231_c80 bl_80 br_80 wl_231 vdd gnd cell_6t
Xbit_r232_c80 bl_80 br_80 wl_232 vdd gnd cell_6t
Xbit_r233_c80 bl_80 br_80 wl_233 vdd gnd cell_6t
Xbit_r234_c80 bl_80 br_80 wl_234 vdd gnd cell_6t
Xbit_r235_c80 bl_80 br_80 wl_235 vdd gnd cell_6t
Xbit_r236_c80 bl_80 br_80 wl_236 vdd gnd cell_6t
Xbit_r237_c80 bl_80 br_80 wl_237 vdd gnd cell_6t
Xbit_r238_c80 bl_80 br_80 wl_238 vdd gnd cell_6t
Xbit_r239_c80 bl_80 br_80 wl_239 vdd gnd cell_6t
Xbit_r240_c80 bl_80 br_80 wl_240 vdd gnd cell_6t
Xbit_r241_c80 bl_80 br_80 wl_241 vdd gnd cell_6t
Xbit_r242_c80 bl_80 br_80 wl_242 vdd gnd cell_6t
Xbit_r243_c80 bl_80 br_80 wl_243 vdd gnd cell_6t
Xbit_r244_c80 bl_80 br_80 wl_244 vdd gnd cell_6t
Xbit_r245_c80 bl_80 br_80 wl_245 vdd gnd cell_6t
Xbit_r246_c80 bl_80 br_80 wl_246 vdd gnd cell_6t
Xbit_r247_c80 bl_80 br_80 wl_247 vdd gnd cell_6t
Xbit_r248_c80 bl_80 br_80 wl_248 vdd gnd cell_6t
Xbit_r249_c80 bl_80 br_80 wl_249 vdd gnd cell_6t
Xbit_r250_c80 bl_80 br_80 wl_250 vdd gnd cell_6t
Xbit_r251_c80 bl_80 br_80 wl_251 vdd gnd cell_6t
Xbit_r252_c80 bl_80 br_80 wl_252 vdd gnd cell_6t
Xbit_r253_c80 bl_80 br_80 wl_253 vdd gnd cell_6t
Xbit_r254_c80 bl_80 br_80 wl_254 vdd gnd cell_6t
Xbit_r255_c80 bl_80 br_80 wl_255 vdd gnd cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd cell_6t
Xbit_r1_c81 bl_81 br_81 wl_1 vdd gnd cell_6t
Xbit_r2_c81 bl_81 br_81 wl_2 vdd gnd cell_6t
Xbit_r3_c81 bl_81 br_81 wl_3 vdd gnd cell_6t
Xbit_r4_c81 bl_81 br_81 wl_4 vdd gnd cell_6t
Xbit_r5_c81 bl_81 br_81 wl_5 vdd gnd cell_6t
Xbit_r6_c81 bl_81 br_81 wl_6 vdd gnd cell_6t
Xbit_r7_c81 bl_81 br_81 wl_7 vdd gnd cell_6t
Xbit_r8_c81 bl_81 br_81 wl_8 vdd gnd cell_6t
Xbit_r9_c81 bl_81 br_81 wl_9 vdd gnd cell_6t
Xbit_r10_c81 bl_81 br_81 wl_10 vdd gnd cell_6t
Xbit_r11_c81 bl_81 br_81 wl_11 vdd gnd cell_6t
Xbit_r12_c81 bl_81 br_81 wl_12 vdd gnd cell_6t
Xbit_r13_c81 bl_81 br_81 wl_13 vdd gnd cell_6t
Xbit_r14_c81 bl_81 br_81 wl_14 vdd gnd cell_6t
Xbit_r15_c81 bl_81 br_81 wl_15 vdd gnd cell_6t
Xbit_r16_c81 bl_81 br_81 wl_16 vdd gnd cell_6t
Xbit_r17_c81 bl_81 br_81 wl_17 vdd gnd cell_6t
Xbit_r18_c81 bl_81 br_81 wl_18 vdd gnd cell_6t
Xbit_r19_c81 bl_81 br_81 wl_19 vdd gnd cell_6t
Xbit_r20_c81 bl_81 br_81 wl_20 vdd gnd cell_6t
Xbit_r21_c81 bl_81 br_81 wl_21 vdd gnd cell_6t
Xbit_r22_c81 bl_81 br_81 wl_22 vdd gnd cell_6t
Xbit_r23_c81 bl_81 br_81 wl_23 vdd gnd cell_6t
Xbit_r24_c81 bl_81 br_81 wl_24 vdd gnd cell_6t
Xbit_r25_c81 bl_81 br_81 wl_25 vdd gnd cell_6t
Xbit_r26_c81 bl_81 br_81 wl_26 vdd gnd cell_6t
Xbit_r27_c81 bl_81 br_81 wl_27 vdd gnd cell_6t
Xbit_r28_c81 bl_81 br_81 wl_28 vdd gnd cell_6t
Xbit_r29_c81 bl_81 br_81 wl_29 vdd gnd cell_6t
Xbit_r30_c81 bl_81 br_81 wl_30 vdd gnd cell_6t
Xbit_r31_c81 bl_81 br_81 wl_31 vdd gnd cell_6t
Xbit_r32_c81 bl_81 br_81 wl_32 vdd gnd cell_6t
Xbit_r33_c81 bl_81 br_81 wl_33 vdd gnd cell_6t
Xbit_r34_c81 bl_81 br_81 wl_34 vdd gnd cell_6t
Xbit_r35_c81 bl_81 br_81 wl_35 vdd gnd cell_6t
Xbit_r36_c81 bl_81 br_81 wl_36 vdd gnd cell_6t
Xbit_r37_c81 bl_81 br_81 wl_37 vdd gnd cell_6t
Xbit_r38_c81 bl_81 br_81 wl_38 vdd gnd cell_6t
Xbit_r39_c81 bl_81 br_81 wl_39 vdd gnd cell_6t
Xbit_r40_c81 bl_81 br_81 wl_40 vdd gnd cell_6t
Xbit_r41_c81 bl_81 br_81 wl_41 vdd gnd cell_6t
Xbit_r42_c81 bl_81 br_81 wl_42 vdd gnd cell_6t
Xbit_r43_c81 bl_81 br_81 wl_43 vdd gnd cell_6t
Xbit_r44_c81 bl_81 br_81 wl_44 vdd gnd cell_6t
Xbit_r45_c81 bl_81 br_81 wl_45 vdd gnd cell_6t
Xbit_r46_c81 bl_81 br_81 wl_46 vdd gnd cell_6t
Xbit_r47_c81 bl_81 br_81 wl_47 vdd gnd cell_6t
Xbit_r48_c81 bl_81 br_81 wl_48 vdd gnd cell_6t
Xbit_r49_c81 bl_81 br_81 wl_49 vdd gnd cell_6t
Xbit_r50_c81 bl_81 br_81 wl_50 vdd gnd cell_6t
Xbit_r51_c81 bl_81 br_81 wl_51 vdd gnd cell_6t
Xbit_r52_c81 bl_81 br_81 wl_52 vdd gnd cell_6t
Xbit_r53_c81 bl_81 br_81 wl_53 vdd gnd cell_6t
Xbit_r54_c81 bl_81 br_81 wl_54 vdd gnd cell_6t
Xbit_r55_c81 bl_81 br_81 wl_55 vdd gnd cell_6t
Xbit_r56_c81 bl_81 br_81 wl_56 vdd gnd cell_6t
Xbit_r57_c81 bl_81 br_81 wl_57 vdd gnd cell_6t
Xbit_r58_c81 bl_81 br_81 wl_58 vdd gnd cell_6t
Xbit_r59_c81 bl_81 br_81 wl_59 vdd gnd cell_6t
Xbit_r60_c81 bl_81 br_81 wl_60 vdd gnd cell_6t
Xbit_r61_c81 bl_81 br_81 wl_61 vdd gnd cell_6t
Xbit_r62_c81 bl_81 br_81 wl_62 vdd gnd cell_6t
Xbit_r63_c81 bl_81 br_81 wl_63 vdd gnd cell_6t
Xbit_r64_c81 bl_81 br_81 wl_64 vdd gnd cell_6t
Xbit_r65_c81 bl_81 br_81 wl_65 vdd gnd cell_6t
Xbit_r66_c81 bl_81 br_81 wl_66 vdd gnd cell_6t
Xbit_r67_c81 bl_81 br_81 wl_67 vdd gnd cell_6t
Xbit_r68_c81 bl_81 br_81 wl_68 vdd gnd cell_6t
Xbit_r69_c81 bl_81 br_81 wl_69 vdd gnd cell_6t
Xbit_r70_c81 bl_81 br_81 wl_70 vdd gnd cell_6t
Xbit_r71_c81 bl_81 br_81 wl_71 vdd gnd cell_6t
Xbit_r72_c81 bl_81 br_81 wl_72 vdd gnd cell_6t
Xbit_r73_c81 bl_81 br_81 wl_73 vdd gnd cell_6t
Xbit_r74_c81 bl_81 br_81 wl_74 vdd gnd cell_6t
Xbit_r75_c81 bl_81 br_81 wl_75 vdd gnd cell_6t
Xbit_r76_c81 bl_81 br_81 wl_76 vdd gnd cell_6t
Xbit_r77_c81 bl_81 br_81 wl_77 vdd gnd cell_6t
Xbit_r78_c81 bl_81 br_81 wl_78 vdd gnd cell_6t
Xbit_r79_c81 bl_81 br_81 wl_79 vdd gnd cell_6t
Xbit_r80_c81 bl_81 br_81 wl_80 vdd gnd cell_6t
Xbit_r81_c81 bl_81 br_81 wl_81 vdd gnd cell_6t
Xbit_r82_c81 bl_81 br_81 wl_82 vdd gnd cell_6t
Xbit_r83_c81 bl_81 br_81 wl_83 vdd gnd cell_6t
Xbit_r84_c81 bl_81 br_81 wl_84 vdd gnd cell_6t
Xbit_r85_c81 bl_81 br_81 wl_85 vdd gnd cell_6t
Xbit_r86_c81 bl_81 br_81 wl_86 vdd gnd cell_6t
Xbit_r87_c81 bl_81 br_81 wl_87 vdd gnd cell_6t
Xbit_r88_c81 bl_81 br_81 wl_88 vdd gnd cell_6t
Xbit_r89_c81 bl_81 br_81 wl_89 vdd gnd cell_6t
Xbit_r90_c81 bl_81 br_81 wl_90 vdd gnd cell_6t
Xbit_r91_c81 bl_81 br_81 wl_91 vdd gnd cell_6t
Xbit_r92_c81 bl_81 br_81 wl_92 vdd gnd cell_6t
Xbit_r93_c81 bl_81 br_81 wl_93 vdd gnd cell_6t
Xbit_r94_c81 bl_81 br_81 wl_94 vdd gnd cell_6t
Xbit_r95_c81 bl_81 br_81 wl_95 vdd gnd cell_6t
Xbit_r96_c81 bl_81 br_81 wl_96 vdd gnd cell_6t
Xbit_r97_c81 bl_81 br_81 wl_97 vdd gnd cell_6t
Xbit_r98_c81 bl_81 br_81 wl_98 vdd gnd cell_6t
Xbit_r99_c81 bl_81 br_81 wl_99 vdd gnd cell_6t
Xbit_r100_c81 bl_81 br_81 wl_100 vdd gnd cell_6t
Xbit_r101_c81 bl_81 br_81 wl_101 vdd gnd cell_6t
Xbit_r102_c81 bl_81 br_81 wl_102 vdd gnd cell_6t
Xbit_r103_c81 bl_81 br_81 wl_103 vdd gnd cell_6t
Xbit_r104_c81 bl_81 br_81 wl_104 vdd gnd cell_6t
Xbit_r105_c81 bl_81 br_81 wl_105 vdd gnd cell_6t
Xbit_r106_c81 bl_81 br_81 wl_106 vdd gnd cell_6t
Xbit_r107_c81 bl_81 br_81 wl_107 vdd gnd cell_6t
Xbit_r108_c81 bl_81 br_81 wl_108 vdd gnd cell_6t
Xbit_r109_c81 bl_81 br_81 wl_109 vdd gnd cell_6t
Xbit_r110_c81 bl_81 br_81 wl_110 vdd gnd cell_6t
Xbit_r111_c81 bl_81 br_81 wl_111 vdd gnd cell_6t
Xbit_r112_c81 bl_81 br_81 wl_112 vdd gnd cell_6t
Xbit_r113_c81 bl_81 br_81 wl_113 vdd gnd cell_6t
Xbit_r114_c81 bl_81 br_81 wl_114 vdd gnd cell_6t
Xbit_r115_c81 bl_81 br_81 wl_115 vdd gnd cell_6t
Xbit_r116_c81 bl_81 br_81 wl_116 vdd gnd cell_6t
Xbit_r117_c81 bl_81 br_81 wl_117 vdd gnd cell_6t
Xbit_r118_c81 bl_81 br_81 wl_118 vdd gnd cell_6t
Xbit_r119_c81 bl_81 br_81 wl_119 vdd gnd cell_6t
Xbit_r120_c81 bl_81 br_81 wl_120 vdd gnd cell_6t
Xbit_r121_c81 bl_81 br_81 wl_121 vdd gnd cell_6t
Xbit_r122_c81 bl_81 br_81 wl_122 vdd gnd cell_6t
Xbit_r123_c81 bl_81 br_81 wl_123 vdd gnd cell_6t
Xbit_r124_c81 bl_81 br_81 wl_124 vdd gnd cell_6t
Xbit_r125_c81 bl_81 br_81 wl_125 vdd gnd cell_6t
Xbit_r126_c81 bl_81 br_81 wl_126 vdd gnd cell_6t
Xbit_r127_c81 bl_81 br_81 wl_127 vdd gnd cell_6t
Xbit_r128_c81 bl_81 br_81 wl_128 vdd gnd cell_6t
Xbit_r129_c81 bl_81 br_81 wl_129 vdd gnd cell_6t
Xbit_r130_c81 bl_81 br_81 wl_130 vdd gnd cell_6t
Xbit_r131_c81 bl_81 br_81 wl_131 vdd gnd cell_6t
Xbit_r132_c81 bl_81 br_81 wl_132 vdd gnd cell_6t
Xbit_r133_c81 bl_81 br_81 wl_133 vdd gnd cell_6t
Xbit_r134_c81 bl_81 br_81 wl_134 vdd gnd cell_6t
Xbit_r135_c81 bl_81 br_81 wl_135 vdd gnd cell_6t
Xbit_r136_c81 bl_81 br_81 wl_136 vdd gnd cell_6t
Xbit_r137_c81 bl_81 br_81 wl_137 vdd gnd cell_6t
Xbit_r138_c81 bl_81 br_81 wl_138 vdd gnd cell_6t
Xbit_r139_c81 bl_81 br_81 wl_139 vdd gnd cell_6t
Xbit_r140_c81 bl_81 br_81 wl_140 vdd gnd cell_6t
Xbit_r141_c81 bl_81 br_81 wl_141 vdd gnd cell_6t
Xbit_r142_c81 bl_81 br_81 wl_142 vdd gnd cell_6t
Xbit_r143_c81 bl_81 br_81 wl_143 vdd gnd cell_6t
Xbit_r144_c81 bl_81 br_81 wl_144 vdd gnd cell_6t
Xbit_r145_c81 bl_81 br_81 wl_145 vdd gnd cell_6t
Xbit_r146_c81 bl_81 br_81 wl_146 vdd gnd cell_6t
Xbit_r147_c81 bl_81 br_81 wl_147 vdd gnd cell_6t
Xbit_r148_c81 bl_81 br_81 wl_148 vdd gnd cell_6t
Xbit_r149_c81 bl_81 br_81 wl_149 vdd gnd cell_6t
Xbit_r150_c81 bl_81 br_81 wl_150 vdd gnd cell_6t
Xbit_r151_c81 bl_81 br_81 wl_151 vdd gnd cell_6t
Xbit_r152_c81 bl_81 br_81 wl_152 vdd gnd cell_6t
Xbit_r153_c81 bl_81 br_81 wl_153 vdd gnd cell_6t
Xbit_r154_c81 bl_81 br_81 wl_154 vdd gnd cell_6t
Xbit_r155_c81 bl_81 br_81 wl_155 vdd gnd cell_6t
Xbit_r156_c81 bl_81 br_81 wl_156 vdd gnd cell_6t
Xbit_r157_c81 bl_81 br_81 wl_157 vdd gnd cell_6t
Xbit_r158_c81 bl_81 br_81 wl_158 vdd gnd cell_6t
Xbit_r159_c81 bl_81 br_81 wl_159 vdd gnd cell_6t
Xbit_r160_c81 bl_81 br_81 wl_160 vdd gnd cell_6t
Xbit_r161_c81 bl_81 br_81 wl_161 vdd gnd cell_6t
Xbit_r162_c81 bl_81 br_81 wl_162 vdd gnd cell_6t
Xbit_r163_c81 bl_81 br_81 wl_163 vdd gnd cell_6t
Xbit_r164_c81 bl_81 br_81 wl_164 vdd gnd cell_6t
Xbit_r165_c81 bl_81 br_81 wl_165 vdd gnd cell_6t
Xbit_r166_c81 bl_81 br_81 wl_166 vdd gnd cell_6t
Xbit_r167_c81 bl_81 br_81 wl_167 vdd gnd cell_6t
Xbit_r168_c81 bl_81 br_81 wl_168 vdd gnd cell_6t
Xbit_r169_c81 bl_81 br_81 wl_169 vdd gnd cell_6t
Xbit_r170_c81 bl_81 br_81 wl_170 vdd gnd cell_6t
Xbit_r171_c81 bl_81 br_81 wl_171 vdd gnd cell_6t
Xbit_r172_c81 bl_81 br_81 wl_172 vdd gnd cell_6t
Xbit_r173_c81 bl_81 br_81 wl_173 vdd gnd cell_6t
Xbit_r174_c81 bl_81 br_81 wl_174 vdd gnd cell_6t
Xbit_r175_c81 bl_81 br_81 wl_175 vdd gnd cell_6t
Xbit_r176_c81 bl_81 br_81 wl_176 vdd gnd cell_6t
Xbit_r177_c81 bl_81 br_81 wl_177 vdd gnd cell_6t
Xbit_r178_c81 bl_81 br_81 wl_178 vdd gnd cell_6t
Xbit_r179_c81 bl_81 br_81 wl_179 vdd gnd cell_6t
Xbit_r180_c81 bl_81 br_81 wl_180 vdd gnd cell_6t
Xbit_r181_c81 bl_81 br_81 wl_181 vdd gnd cell_6t
Xbit_r182_c81 bl_81 br_81 wl_182 vdd gnd cell_6t
Xbit_r183_c81 bl_81 br_81 wl_183 vdd gnd cell_6t
Xbit_r184_c81 bl_81 br_81 wl_184 vdd gnd cell_6t
Xbit_r185_c81 bl_81 br_81 wl_185 vdd gnd cell_6t
Xbit_r186_c81 bl_81 br_81 wl_186 vdd gnd cell_6t
Xbit_r187_c81 bl_81 br_81 wl_187 vdd gnd cell_6t
Xbit_r188_c81 bl_81 br_81 wl_188 vdd gnd cell_6t
Xbit_r189_c81 bl_81 br_81 wl_189 vdd gnd cell_6t
Xbit_r190_c81 bl_81 br_81 wl_190 vdd gnd cell_6t
Xbit_r191_c81 bl_81 br_81 wl_191 vdd gnd cell_6t
Xbit_r192_c81 bl_81 br_81 wl_192 vdd gnd cell_6t
Xbit_r193_c81 bl_81 br_81 wl_193 vdd gnd cell_6t
Xbit_r194_c81 bl_81 br_81 wl_194 vdd gnd cell_6t
Xbit_r195_c81 bl_81 br_81 wl_195 vdd gnd cell_6t
Xbit_r196_c81 bl_81 br_81 wl_196 vdd gnd cell_6t
Xbit_r197_c81 bl_81 br_81 wl_197 vdd gnd cell_6t
Xbit_r198_c81 bl_81 br_81 wl_198 vdd gnd cell_6t
Xbit_r199_c81 bl_81 br_81 wl_199 vdd gnd cell_6t
Xbit_r200_c81 bl_81 br_81 wl_200 vdd gnd cell_6t
Xbit_r201_c81 bl_81 br_81 wl_201 vdd gnd cell_6t
Xbit_r202_c81 bl_81 br_81 wl_202 vdd gnd cell_6t
Xbit_r203_c81 bl_81 br_81 wl_203 vdd gnd cell_6t
Xbit_r204_c81 bl_81 br_81 wl_204 vdd gnd cell_6t
Xbit_r205_c81 bl_81 br_81 wl_205 vdd gnd cell_6t
Xbit_r206_c81 bl_81 br_81 wl_206 vdd gnd cell_6t
Xbit_r207_c81 bl_81 br_81 wl_207 vdd gnd cell_6t
Xbit_r208_c81 bl_81 br_81 wl_208 vdd gnd cell_6t
Xbit_r209_c81 bl_81 br_81 wl_209 vdd gnd cell_6t
Xbit_r210_c81 bl_81 br_81 wl_210 vdd gnd cell_6t
Xbit_r211_c81 bl_81 br_81 wl_211 vdd gnd cell_6t
Xbit_r212_c81 bl_81 br_81 wl_212 vdd gnd cell_6t
Xbit_r213_c81 bl_81 br_81 wl_213 vdd gnd cell_6t
Xbit_r214_c81 bl_81 br_81 wl_214 vdd gnd cell_6t
Xbit_r215_c81 bl_81 br_81 wl_215 vdd gnd cell_6t
Xbit_r216_c81 bl_81 br_81 wl_216 vdd gnd cell_6t
Xbit_r217_c81 bl_81 br_81 wl_217 vdd gnd cell_6t
Xbit_r218_c81 bl_81 br_81 wl_218 vdd gnd cell_6t
Xbit_r219_c81 bl_81 br_81 wl_219 vdd gnd cell_6t
Xbit_r220_c81 bl_81 br_81 wl_220 vdd gnd cell_6t
Xbit_r221_c81 bl_81 br_81 wl_221 vdd gnd cell_6t
Xbit_r222_c81 bl_81 br_81 wl_222 vdd gnd cell_6t
Xbit_r223_c81 bl_81 br_81 wl_223 vdd gnd cell_6t
Xbit_r224_c81 bl_81 br_81 wl_224 vdd gnd cell_6t
Xbit_r225_c81 bl_81 br_81 wl_225 vdd gnd cell_6t
Xbit_r226_c81 bl_81 br_81 wl_226 vdd gnd cell_6t
Xbit_r227_c81 bl_81 br_81 wl_227 vdd gnd cell_6t
Xbit_r228_c81 bl_81 br_81 wl_228 vdd gnd cell_6t
Xbit_r229_c81 bl_81 br_81 wl_229 vdd gnd cell_6t
Xbit_r230_c81 bl_81 br_81 wl_230 vdd gnd cell_6t
Xbit_r231_c81 bl_81 br_81 wl_231 vdd gnd cell_6t
Xbit_r232_c81 bl_81 br_81 wl_232 vdd gnd cell_6t
Xbit_r233_c81 bl_81 br_81 wl_233 vdd gnd cell_6t
Xbit_r234_c81 bl_81 br_81 wl_234 vdd gnd cell_6t
Xbit_r235_c81 bl_81 br_81 wl_235 vdd gnd cell_6t
Xbit_r236_c81 bl_81 br_81 wl_236 vdd gnd cell_6t
Xbit_r237_c81 bl_81 br_81 wl_237 vdd gnd cell_6t
Xbit_r238_c81 bl_81 br_81 wl_238 vdd gnd cell_6t
Xbit_r239_c81 bl_81 br_81 wl_239 vdd gnd cell_6t
Xbit_r240_c81 bl_81 br_81 wl_240 vdd gnd cell_6t
Xbit_r241_c81 bl_81 br_81 wl_241 vdd gnd cell_6t
Xbit_r242_c81 bl_81 br_81 wl_242 vdd gnd cell_6t
Xbit_r243_c81 bl_81 br_81 wl_243 vdd gnd cell_6t
Xbit_r244_c81 bl_81 br_81 wl_244 vdd gnd cell_6t
Xbit_r245_c81 bl_81 br_81 wl_245 vdd gnd cell_6t
Xbit_r246_c81 bl_81 br_81 wl_246 vdd gnd cell_6t
Xbit_r247_c81 bl_81 br_81 wl_247 vdd gnd cell_6t
Xbit_r248_c81 bl_81 br_81 wl_248 vdd gnd cell_6t
Xbit_r249_c81 bl_81 br_81 wl_249 vdd gnd cell_6t
Xbit_r250_c81 bl_81 br_81 wl_250 vdd gnd cell_6t
Xbit_r251_c81 bl_81 br_81 wl_251 vdd gnd cell_6t
Xbit_r252_c81 bl_81 br_81 wl_252 vdd gnd cell_6t
Xbit_r253_c81 bl_81 br_81 wl_253 vdd gnd cell_6t
Xbit_r254_c81 bl_81 br_81 wl_254 vdd gnd cell_6t
Xbit_r255_c81 bl_81 br_81 wl_255 vdd gnd cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd cell_6t
Xbit_r1_c82 bl_82 br_82 wl_1 vdd gnd cell_6t
Xbit_r2_c82 bl_82 br_82 wl_2 vdd gnd cell_6t
Xbit_r3_c82 bl_82 br_82 wl_3 vdd gnd cell_6t
Xbit_r4_c82 bl_82 br_82 wl_4 vdd gnd cell_6t
Xbit_r5_c82 bl_82 br_82 wl_5 vdd gnd cell_6t
Xbit_r6_c82 bl_82 br_82 wl_6 vdd gnd cell_6t
Xbit_r7_c82 bl_82 br_82 wl_7 vdd gnd cell_6t
Xbit_r8_c82 bl_82 br_82 wl_8 vdd gnd cell_6t
Xbit_r9_c82 bl_82 br_82 wl_9 vdd gnd cell_6t
Xbit_r10_c82 bl_82 br_82 wl_10 vdd gnd cell_6t
Xbit_r11_c82 bl_82 br_82 wl_11 vdd gnd cell_6t
Xbit_r12_c82 bl_82 br_82 wl_12 vdd gnd cell_6t
Xbit_r13_c82 bl_82 br_82 wl_13 vdd gnd cell_6t
Xbit_r14_c82 bl_82 br_82 wl_14 vdd gnd cell_6t
Xbit_r15_c82 bl_82 br_82 wl_15 vdd gnd cell_6t
Xbit_r16_c82 bl_82 br_82 wl_16 vdd gnd cell_6t
Xbit_r17_c82 bl_82 br_82 wl_17 vdd gnd cell_6t
Xbit_r18_c82 bl_82 br_82 wl_18 vdd gnd cell_6t
Xbit_r19_c82 bl_82 br_82 wl_19 vdd gnd cell_6t
Xbit_r20_c82 bl_82 br_82 wl_20 vdd gnd cell_6t
Xbit_r21_c82 bl_82 br_82 wl_21 vdd gnd cell_6t
Xbit_r22_c82 bl_82 br_82 wl_22 vdd gnd cell_6t
Xbit_r23_c82 bl_82 br_82 wl_23 vdd gnd cell_6t
Xbit_r24_c82 bl_82 br_82 wl_24 vdd gnd cell_6t
Xbit_r25_c82 bl_82 br_82 wl_25 vdd gnd cell_6t
Xbit_r26_c82 bl_82 br_82 wl_26 vdd gnd cell_6t
Xbit_r27_c82 bl_82 br_82 wl_27 vdd gnd cell_6t
Xbit_r28_c82 bl_82 br_82 wl_28 vdd gnd cell_6t
Xbit_r29_c82 bl_82 br_82 wl_29 vdd gnd cell_6t
Xbit_r30_c82 bl_82 br_82 wl_30 vdd gnd cell_6t
Xbit_r31_c82 bl_82 br_82 wl_31 vdd gnd cell_6t
Xbit_r32_c82 bl_82 br_82 wl_32 vdd gnd cell_6t
Xbit_r33_c82 bl_82 br_82 wl_33 vdd gnd cell_6t
Xbit_r34_c82 bl_82 br_82 wl_34 vdd gnd cell_6t
Xbit_r35_c82 bl_82 br_82 wl_35 vdd gnd cell_6t
Xbit_r36_c82 bl_82 br_82 wl_36 vdd gnd cell_6t
Xbit_r37_c82 bl_82 br_82 wl_37 vdd gnd cell_6t
Xbit_r38_c82 bl_82 br_82 wl_38 vdd gnd cell_6t
Xbit_r39_c82 bl_82 br_82 wl_39 vdd gnd cell_6t
Xbit_r40_c82 bl_82 br_82 wl_40 vdd gnd cell_6t
Xbit_r41_c82 bl_82 br_82 wl_41 vdd gnd cell_6t
Xbit_r42_c82 bl_82 br_82 wl_42 vdd gnd cell_6t
Xbit_r43_c82 bl_82 br_82 wl_43 vdd gnd cell_6t
Xbit_r44_c82 bl_82 br_82 wl_44 vdd gnd cell_6t
Xbit_r45_c82 bl_82 br_82 wl_45 vdd gnd cell_6t
Xbit_r46_c82 bl_82 br_82 wl_46 vdd gnd cell_6t
Xbit_r47_c82 bl_82 br_82 wl_47 vdd gnd cell_6t
Xbit_r48_c82 bl_82 br_82 wl_48 vdd gnd cell_6t
Xbit_r49_c82 bl_82 br_82 wl_49 vdd gnd cell_6t
Xbit_r50_c82 bl_82 br_82 wl_50 vdd gnd cell_6t
Xbit_r51_c82 bl_82 br_82 wl_51 vdd gnd cell_6t
Xbit_r52_c82 bl_82 br_82 wl_52 vdd gnd cell_6t
Xbit_r53_c82 bl_82 br_82 wl_53 vdd gnd cell_6t
Xbit_r54_c82 bl_82 br_82 wl_54 vdd gnd cell_6t
Xbit_r55_c82 bl_82 br_82 wl_55 vdd gnd cell_6t
Xbit_r56_c82 bl_82 br_82 wl_56 vdd gnd cell_6t
Xbit_r57_c82 bl_82 br_82 wl_57 vdd gnd cell_6t
Xbit_r58_c82 bl_82 br_82 wl_58 vdd gnd cell_6t
Xbit_r59_c82 bl_82 br_82 wl_59 vdd gnd cell_6t
Xbit_r60_c82 bl_82 br_82 wl_60 vdd gnd cell_6t
Xbit_r61_c82 bl_82 br_82 wl_61 vdd gnd cell_6t
Xbit_r62_c82 bl_82 br_82 wl_62 vdd gnd cell_6t
Xbit_r63_c82 bl_82 br_82 wl_63 vdd gnd cell_6t
Xbit_r64_c82 bl_82 br_82 wl_64 vdd gnd cell_6t
Xbit_r65_c82 bl_82 br_82 wl_65 vdd gnd cell_6t
Xbit_r66_c82 bl_82 br_82 wl_66 vdd gnd cell_6t
Xbit_r67_c82 bl_82 br_82 wl_67 vdd gnd cell_6t
Xbit_r68_c82 bl_82 br_82 wl_68 vdd gnd cell_6t
Xbit_r69_c82 bl_82 br_82 wl_69 vdd gnd cell_6t
Xbit_r70_c82 bl_82 br_82 wl_70 vdd gnd cell_6t
Xbit_r71_c82 bl_82 br_82 wl_71 vdd gnd cell_6t
Xbit_r72_c82 bl_82 br_82 wl_72 vdd gnd cell_6t
Xbit_r73_c82 bl_82 br_82 wl_73 vdd gnd cell_6t
Xbit_r74_c82 bl_82 br_82 wl_74 vdd gnd cell_6t
Xbit_r75_c82 bl_82 br_82 wl_75 vdd gnd cell_6t
Xbit_r76_c82 bl_82 br_82 wl_76 vdd gnd cell_6t
Xbit_r77_c82 bl_82 br_82 wl_77 vdd gnd cell_6t
Xbit_r78_c82 bl_82 br_82 wl_78 vdd gnd cell_6t
Xbit_r79_c82 bl_82 br_82 wl_79 vdd gnd cell_6t
Xbit_r80_c82 bl_82 br_82 wl_80 vdd gnd cell_6t
Xbit_r81_c82 bl_82 br_82 wl_81 vdd gnd cell_6t
Xbit_r82_c82 bl_82 br_82 wl_82 vdd gnd cell_6t
Xbit_r83_c82 bl_82 br_82 wl_83 vdd gnd cell_6t
Xbit_r84_c82 bl_82 br_82 wl_84 vdd gnd cell_6t
Xbit_r85_c82 bl_82 br_82 wl_85 vdd gnd cell_6t
Xbit_r86_c82 bl_82 br_82 wl_86 vdd gnd cell_6t
Xbit_r87_c82 bl_82 br_82 wl_87 vdd gnd cell_6t
Xbit_r88_c82 bl_82 br_82 wl_88 vdd gnd cell_6t
Xbit_r89_c82 bl_82 br_82 wl_89 vdd gnd cell_6t
Xbit_r90_c82 bl_82 br_82 wl_90 vdd gnd cell_6t
Xbit_r91_c82 bl_82 br_82 wl_91 vdd gnd cell_6t
Xbit_r92_c82 bl_82 br_82 wl_92 vdd gnd cell_6t
Xbit_r93_c82 bl_82 br_82 wl_93 vdd gnd cell_6t
Xbit_r94_c82 bl_82 br_82 wl_94 vdd gnd cell_6t
Xbit_r95_c82 bl_82 br_82 wl_95 vdd gnd cell_6t
Xbit_r96_c82 bl_82 br_82 wl_96 vdd gnd cell_6t
Xbit_r97_c82 bl_82 br_82 wl_97 vdd gnd cell_6t
Xbit_r98_c82 bl_82 br_82 wl_98 vdd gnd cell_6t
Xbit_r99_c82 bl_82 br_82 wl_99 vdd gnd cell_6t
Xbit_r100_c82 bl_82 br_82 wl_100 vdd gnd cell_6t
Xbit_r101_c82 bl_82 br_82 wl_101 vdd gnd cell_6t
Xbit_r102_c82 bl_82 br_82 wl_102 vdd gnd cell_6t
Xbit_r103_c82 bl_82 br_82 wl_103 vdd gnd cell_6t
Xbit_r104_c82 bl_82 br_82 wl_104 vdd gnd cell_6t
Xbit_r105_c82 bl_82 br_82 wl_105 vdd gnd cell_6t
Xbit_r106_c82 bl_82 br_82 wl_106 vdd gnd cell_6t
Xbit_r107_c82 bl_82 br_82 wl_107 vdd gnd cell_6t
Xbit_r108_c82 bl_82 br_82 wl_108 vdd gnd cell_6t
Xbit_r109_c82 bl_82 br_82 wl_109 vdd gnd cell_6t
Xbit_r110_c82 bl_82 br_82 wl_110 vdd gnd cell_6t
Xbit_r111_c82 bl_82 br_82 wl_111 vdd gnd cell_6t
Xbit_r112_c82 bl_82 br_82 wl_112 vdd gnd cell_6t
Xbit_r113_c82 bl_82 br_82 wl_113 vdd gnd cell_6t
Xbit_r114_c82 bl_82 br_82 wl_114 vdd gnd cell_6t
Xbit_r115_c82 bl_82 br_82 wl_115 vdd gnd cell_6t
Xbit_r116_c82 bl_82 br_82 wl_116 vdd gnd cell_6t
Xbit_r117_c82 bl_82 br_82 wl_117 vdd gnd cell_6t
Xbit_r118_c82 bl_82 br_82 wl_118 vdd gnd cell_6t
Xbit_r119_c82 bl_82 br_82 wl_119 vdd gnd cell_6t
Xbit_r120_c82 bl_82 br_82 wl_120 vdd gnd cell_6t
Xbit_r121_c82 bl_82 br_82 wl_121 vdd gnd cell_6t
Xbit_r122_c82 bl_82 br_82 wl_122 vdd gnd cell_6t
Xbit_r123_c82 bl_82 br_82 wl_123 vdd gnd cell_6t
Xbit_r124_c82 bl_82 br_82 wl_124 vdd gnd cell_6t
Xbit_r125_c82 bl_82 br_82 wl_125 vdd gnd cell_6t
Xbit_r126_c82 bl_82 br_82 wl_126 vdd gnd cell_6t
Xbit_r127_c82 bl_82 br_82 wl_127 vdd gnd cell_6t
Xbit_r128_c82 bl_82 br_82 wl_128 vdd gnd cell_6t
Xbit_r129_c82 bl_82 br_82 wl_129 vdd gnd cell_6t
Xbit_r130_c82 bl_82 br_82 wl_130 vdd gnd cell_6t
Xbit_r131_c82 bl_82 br_82 wl_131 vdd gnd cell_6t
Xbit_r132_c82 bl_82 br_82 wl_132 vdd gnd cell_6t
Xbit_r133_c82 bl_82 br_82 wl_133 vdd gnd cell_6t
Xbit_r134_c82 bl_82 br_82 wl_134 vdd gnd cell_6t
Xbit_r135_c82 bl_82 br_82 wl_135 vdd gnd cell_6t
Xbit_r136_c82 bl_82 br_82 wl_136 vdd gnd cell_6t
Xbit_r137_c82 bl_82 br_82 wl_137 vdd gnd cell_6t
Xbit_r138_c82 bl_82 br_82 wl_138 vdd gnd cell_6t
Xbit_r139_c82 bl_82 br_82 wl_139 vdd gnd cell_6t
Xbit_r140_c82 bl_82 br_82 wl_140 vdd gnd cell_6t
Xbit_r141_c82 bl_82 br_82 wl_141 vdd gnd cell_6t
Xbit_r142_c82 bl_82 br_82 wl_142 vdd gnd cell_6t
Xbit_r143_c82 bl_82 br_82 wl_143 vdd gnd cell_6t
Xbit_r144_c82 bl_82 br_82 wl_144 vdd gnd cell_6t
Xbit_r145_c82 bl_82 br_82 wl_145 vdd gnd cell_6t
Xbit_r146_c82 bl_82 br_82 wl_146 vdd gnd cell_6t
Xbit_r147_c82 bl_82 br_82 wl_147 vdd gnd cell_6t
Xbit_r148_c82 bl_82 br_82 wl_148 vdd gnd cell_6t
Xbit_r149_c82 bl_82 br_82 wl_149 vdd gnd cell_6t
Xbit_r150_c82 bl_82 br_82 wl_150 vdd gnd cell_6t
Xbit_r151_c82 bl_82 br_82 wl_151 vdd gnd cell_6t
Xbit_r152_c82 bl_82 br_82 wl_152 vdd gnd cell_6t
Xbit_r153_c82 bl_82 br_82 wl_153 vdd gnd cell_6t
Xbit_r154_c82 bl_82 br_82 wl_154 vdd gnd cell_6t
Xbit_r155_c82 bl_82 br_82 wl_155 vdd gnd cell_6t
Xbit_r156_c82 bl_82 br_82 wl_156 vdd gnd cell_6t
Xbit_r157_c82 bl_82 br_82 wl_157 vdd gnd cell_6t
Xbit_r158_c82 bl_82 br_82 wl_158 vdd gnd cell_6t
Xbit_r159_c82 bl_82 br_82 wl_159 vdd gnd cell_6t
Xbit_r160_c82 bl_82 br_82 wl_160 vdd gnd cell_6t
Xbit_r161_c82 bl_82 br_82 wl_161 vdd gnd cell_6t
Xbit_r162_c82 bl_82 br_82 wl_162 vdd gnd cell_6t
Xbit_r163_c82 bl_82 br_82 wl_163 vdd gnd cell_6t
Xbit_r164_c82 bl_82 br_82 wl_164 vdd gnd cell_6t
Xbit_r165_c82 bl_82 br_82 wl_165 vdd gnd cell_6t
Xbit_r166_c82 bl_82 br_82 wl_166 vdd gnd cell_6t
Xbit_r167_c82 bl_82 br_82 wl_167 vdd gnd cell_6t
Xbit_r168_c82 bl_82 br_82 wl_168 vdd gnd cell_6t
Xbit_r169_c82 bl_82 br_82 wl_169 vdd gnd cell_6t
Xbit_r170_c82 bl_82 br_82 wl_170 vdd gnd cell_6t
Xbit_r171_c82 bl_82 br_82 wl_171 vdd gnd cell_6t
Xbit_r172_c82 bl_82 br_82 wl_172 vdd gnd cell_6t
Xbit_r173_c82 bl_82 br_82 wl_173 vdd gnd cell_6t
Xbit_r174_c82 bl_82 br_82 wl_174 vdd gnd cell_6t
Xbit_r175_c82 bl_82 br_82 wl_175 vdd gnd cell_6t
Xbit_r176_c82 bl_82 br_82 wl_176 vdd gnd cell_6t
Xbit_r177_c82 bl_82 br_82 wl_177 vdd gnd cell_6t
Xbit_r178_c82 bl_82 br_82 wl_178 vdd gnd cell_6t
Xbit_r179_c82 bl_82 br_82 wl_179 vdd gnd cell_6t
Xbit_r180_c82 bl_82 br_82 wl_180 vdd gnd cell_6t
Xbit_r181_c82 bl_82 br_82 wl_181 vdd gnd cell_6t
Xbit_r182_c82 bl_82 br_82 wl_182 vdd gnd cell_6t
Xbit_r183_c82 bl_82 br_82 wl_183 vdd gnd cell_6t
Xbit_r184_c82 bl_82 br_82 wl_184 vdd gnd cell_6t
Xbit_r185_c82 bl_82 br_82 wl_185 vdd gnd cell_6t
Xbit_r186_c82 bl_82 br_82 wl_186 vdd gnd cell_6t
Xbit_r187_c82 bl_82 br_82 wl_187 vdd gnd cell_6t
Xbit_r188_c82 bl_82 br_82 wl_188 vdd gnd cell_6t
Xbit_r189_c82 bl_82 br_82 wl_189 vdd gnd cell_6t
Xbit_r190_c82 bl_82 br_82 wl_190 vdd gnd cell_6t
Xbit_r191_c82 bl_82 br_82 wl_191 vdd gnd cell_6t
Xbit_r192_c82 bl_82 br_82 wl_192 vdd gnd cell_6t
Xbit_r193_c82 bl_82 br_82 wl_193 vdd gnd cell_6t
Xbit_r194_c82 bl_82 br_82 wl_194 vdd gnd cell_6t
Xbit_r195_c82 bl_82 br_82 wl_195 vdd gnd cell_6t
Xbit_r196_c82 bl_82 br_82 wl_196 vdd gnd cell_6t
Xbit_r197_c82 bl_82 br_82 wl_197 vdd gnd cell_6t
Xbit_r198_c82 bl_82 br_82 wl_198 vdd gnd cell_6t
Xbit_r199_c82 bl_82 br_82 wl_199 vdd gnd cell_6t
Xbit_r200_c82 bl_82 br_82 wl_200 vdd gnd cell_6t
Xbit_r201_c82 bl_82 br_82 wl_201 vdd gnd cell_6t
Xbit_r202_c82 bl_82 br_82 wl_202 vdd gnd cell_6t
Xbit_r203_c82 bl_82 br_82 wl_203 vdd gnd cell_6t
Xbit_r204_c82 bl_82 br_82 wl_204 vdd gnd cell_6t
Xbit_r205_c82 bl_82 br_82 wl_205 vdd gnd cell_6t
Xbit_r206_c82 bl_82 br_82 wl_206 vdd gnd cell_6t
Xbit_r207_c82 bl_82 br_82 wl_207 vdd gnd cell_6t
Xbit_r208_c82 bl_82 br_82 wl_208 vdd gnd cell_6t
Xbit_r209_c82 bl_82 br_82 wl_209 vdd gnd cell_6t
Xbit_r210_c82 bl_82 br_82 wl_210 vdd gnd cell_6t
Xbit_r211_c82 bl_82 br_82 wl_211 vdd gnd cell_6t
Xbit_r212_c82 bl_82 br_82 wl_212 vdd gnd cell_6t
Xbit_r213_c82 bl_82 br_82 wl_213 vdd gnd cell_6t
Xbit_r214_c82 bl_82 br_82 wl_214 vdd gnd cell_6t
Xbit_r215_c82 bl_82 br_82 wl_215 vdd gnd cell_6t
Xbit_r216_c82 bl_82 br_82 wl_216 vdd gnd cell_6t
Xbit_r217_c82 bl_82 br_82 wl_217 vdd gnd cell_6t
Xbit_r218_c82 bl_82 br_82 wl_218 vdd gnd cell_6t
Xbit_r219_c82 bl_82 br_82 wl_219 vdd gnd cell_6t
Xbit_r220_c82 bl_82 br_82 wl_220 vdd gnd cell_6t
Xbit_r221_c82 bl_82 br_82 wl_221 vdd gnd cell_6t
Xbit_r222_c82 bl_82 br_82 wl_222 vdd gnd cell_6t
Xbit_r223_c82 bl_82 br_82 wl_223 vdd gnd cell_6t
Xbit_r224_c82 bl_82 br_82 wl_224 vdd gnd cell_6t
Xbit_r225_c82 bl_82 br_82 wl_225 vdd gnd cell_6t
Xbit_r226_c82 bl_82 br_82 wl_226 vdd gnd cell_6t
Xbit_r227_c82 bl_82 br_82 wl_227 vdd gnd cell_6t
Xbit_r228_c82 bl_82 br_82 wl_228 vdd gnd cell_6t
Xbit_r229_c82 bl_82 br_82 wl_229 vdd gnd cell_6t
Xbit_r230_c82 bl_82 br_82 wl_230 vdd gnd cell_6t
Xbit_r231_c82 bl_82 br_82 wl_231 vdd gnd cell_6t
Xbit_r232_c82 bl_82 br_82 wl_232 vdd gnd cell_6t
Xbit_r233_c82 bl_82 br_82 wl_233 vdd gnd cell_6t
Xbit_r234_c82 bl_82 br_82 wl_234 vdd gnd cell_6t
Xbit_r235_c82 bl_82 br_82 wl_235 vdd gnd cell_6t
Xbit_r236_c82 bl_82 br_82 wl_236 vdd gnd cell_6t
Xbit_r237_c82 bl_82 br_82 wl_237 vdd gnd cell_6t
Xbit_r238_c82 bl_82 br_82 wl_238 vdd gnd cell_6t
Xbit_r239_c82 bl_82 br_82 wl_239 vdd gnd cell_6t
Xbit_r240_c82 bl_82 br_82 wl_240 vdd gnd cell_6t
Xbit_r241_c82 bl_82 br_82 wl_241 vdd gnd cell_6t
Xbit_r242_c82 bl_82 br_82 wl_242 vdd gnd cell_6t
Xbit_r243_c82 bl_82 br_82 wl_243 vdd gnd cell_6t
Xbit_r244_c82 bl_82 br_82 wl_244 vdd gnd cell_6t
Xbit_r245_c82 bl_82 br_82 wl_245 vdd gnd cell_6t
Xbit_r246_c82 bl_82 br_82 wl_246 vdd gnd cell_6t
Xbit_r247_c82 bl_82 br_82 wl_247 vdd gnd cell_6t
Xbit_r248_c82 bl_82 br_82 wl_248 vdd gnd cell_6t
Xbit_r249_c82 bl_82 br_82 wl_249 vdd gnd cell_6t
Xbit_r250_c82 bl_82 br_82 wl_250 vdd gnd cell_6t
Xbit_r251_c82 bl_82 br_82 wl_251 vdd gnd cell_6t
Xbit_r252_c82 bl_82 br_82 wl_252 vdd gnd cell_6t
Xbit_r253_c82 bl_82 br_82 wl_253 vdd gnd cell_6t
Xbit_r254_c82 bl_82 br_82 wl_254 vdd gnd cell_6t
Xbit_r255_c82 bl_82 br_82 wl_255 vdd gnd cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd cell_6t
Xbit_r1_c83 bl_83 br_83 wl_1 vdd gnd cell_6t
Xbit_r2_c83 bl_83 br_83 wl_2 vdd gnd cell_6t
Xbit_r3_c83 bl_83 br_83 wl_3 vdd gnd cell_6t
Xbit_r4_c83 bl_83 br_83 wl_4 vdd gnd cell_6t
Xbit_r5_c83 bl_83 br_83 wl_5 vdd gnd cell_6t
Xbit_r6_c83 bl_83 br_83 wl_6 vdd gnd cell_6t
Xbit_r7_c83 bl_83 br_83 wl_7 vdd gnd cell_6t
Xbit_r8_c83 bl_83 br_83 wl_8 vdd gnd cell_6t
Xbit_r9_c83 bl_83 br_83 wl_9 vdd gnd cell_6t
Xbit_r10_c83 bl_83 br_83 wl_10 vdd gnd cell_6t
Xbit_r11_c83 bl_83 br_83 wl_11 vdd gnd cell_6t
Xbit_r12_c83 bl_83 br_83 wl_12 vdd gnd cell_6t
Xbit_r13_c83 bl_83 br_83 wl_13 vdd gnd cell_6t
Xbit_r14_c83 bl_83 br_83 wl_14 vdd gnd cell_6t
Xbit_r15_c83 bl_83 br_83 wl_15 vdd gnd cell_6t
Xbit_r16_c83 bl_83 br_83 wl_16 vdd gnd cell_6t
Xbit_r17_c83 bl_83 br_83 wl_17 vdd gnd cell_6t
Xbit_r18_c83 bl_83 br_83 wl_18 vdd gnd cell_6t
Xbit_r19_c83 bl_83 br_83 wl_19 vdd gnd cell_6t
Xbit_r20_c83 bl_83 br_83 wl_20 vdd gnd cell_6t
Xbit_r21_c83 bl_83 br_83 wl_21 vdd gnd cell_6t
Xbit_r22_c83 bl_83 br_83 wl_22 vdd gnd cell_6t
Xbit_r23_c83 bl_83 br_83 wl_23 vdd gnd cell_6t
Xbit_r24_c83 bl_83 br_83 wl_24 vdd gnd cell_6t
Xbit_r25_c83 bl_83 br_83 wl_25 vdd gnd cell_6t
Xbit_r26_c83 bl_83 br_83 wl_26 vdd gnd cell_6t
Xbit_r27_c83 bl_83 br_83 wl_27 vdd gnd cell_6t
Xbit_r28_c83 bl_83 br_83 wl_28 vdd gnd cell_6t
Xbit_r29_c83 bl_83 br_83 wl_29 vdd gnd cell_6t
Xbit_r30_c83 bl_83 br_83 wl_30 vdd gnd cell_6t
Xbit_r31_c83 bl_83 br_83 wl_31 vdd gnd cell_6t
Xbit_r32_c83 bl_83 br_83 wl_32 vdd gnd cell_6t
Xbit_r33_c83 bl_83 br_83 wl_33 vdd gnd cell_6t
Xbit_r34_c83 bl_83 br_83 wl_34 vdd gnd cell_6t
Xbit_r35_c83 bl_83 br_83 wl_35 vdd gnd cell_6t
Xbit_r36_c83 bl_83 br_83 wl_36 vdd gnd cell_6t
Xbit_r37_c83 bl_83 br_83 wl_37 vdd gnd cell_6t
Xbit_r38_c83 bl_83 br_83 wl_38 vdd gnd cell_6t
Xbit_r39_c83 bl_83 br_83 wl_39 vdd gnd cell_6t
Xbit_r40_c83 bl_83 br_83 wl_40 vdd gnd cell_6t
Xbit_r41_c83 bl_83 br_83 wl_41 vdd gnd cell_6t
Xbit_r42_c83 bl_83 br_83 wl_42 vdd gnd cell_6t
Xbit_r43_c83 bl_83 br_83 wl_43 vdd gnd cell_6t
Xbit_r44_c83 bl_83 br_83 wl_44 vdd gnd cell_6t
Xbit_r45_c83 bl_83 br_83 wl_45 vdd gnd cell_6t
Xbit_r46_c83 bl_83 br_83 wl_46 vdd gnd cell_6t
Xbit_r47_c83 bl_83 br_83 wl_47 vdd gnd cell_6t
Xbit_r48_c83 bl_83 br_83 wl_48 vdd gnd cell_6t
Xbit_r49_c83 bl_83 br_83 wl_49 vdd gnd cell_6t
Xbit_r50_c83 bl_83 br_83 wl_50 vdd gnd cell_6t
Xbit_r51_c83 bl_83 br_83 wl_51 vdd gnd cell_6t
Xbit_r52_c83 bl_83 br_83 wl_52 vdd gnd cell_6t
Xbit_r53_c83 bl_83 br_83 wl_53 vdd gnd cell_6t
Xbit_r54_c83 bl_83 br_83 wl_54 vdd gnd cell_6t
Xbit_r55_c83 bl_83 br_83 wl_55 vdd gnd cell_6t
Xbit_r56_c83 bl_83 br_83 wl_56 vdd gnd cell_6t
Xbit_r57_c83 bl_83 br_83 wl_57 vdd gnd cell_6t
Xbit_r58_c83 bl_83 br_83 wl_58 vdd gnd cell_6t
Xbit_r59_c83 bl_83 br_83 wl_59 vdd gnd cell_6t
Xbit_r60_c83 bl_83 br_83 wl_60 vdd gnd cell_6t
Xbit_r61_c83 bl_83 br_83 wl_61 vdd gnd cell_6t
Xbit_r62_c83 bl_83 br_83 wl_62 vdd gnd cell_6t
Xbit_r63_c83 bl_83 br_83 wl_63 vdd gnd cell_6t
Xbit_r64_c83 bl_83 br_83 wl_64 vdd gnd cell_6t
Xbit_r65_c83 bl_83 br_83 wl_65 vdd gnd cell_6t
Xbit_r66_c83 bl_83 br_83 wl_66 vdd gnd cell_6t
Xbit_r67_c83 bl_83 br_83 wl_67 vdd gnd cell_6t
Xbit_r68_c83 bl_83 br_83 wl_68 vdd gnd cell_6t
Xbit_r69_c83 bl_83 br_83 wl_69 vdd gnd cell_6t
Xbit_r70_c83 bl_83 br_83 wl_70 vdd gnd cell_6t
Xbit_r71_c83 bl_83 br_83 wl_71 vdd gnd cell_6t
Xbit_r72_c83 bl_83 br_83 wl_72 vdd gnd cell_6t
Xbit_r73_c83 bl_83 br_83 wl_73 vdd gnd cell_6t
Xbit_r74_c83 bl_83 br_83 wl_74 vdd gnd cell_6t
Xbit_r75_c83 bl_83 br_83 wl_75 vdd gnd cell_6t
Xbit_r76_c83 bl_83 br_83 wl_76 vdd gnd cell_6t
Xbit_r77_c83 bl_83 br_83 wl_77 vdd gnd cell_6t
Xbit_r78_c83 bl_83 br_83 wl_78 vdd gnd cell_6t
Xbit_r79_c83 bl_83 br_83 wl_79 vdd gnd cell_6t
Xbit_r80_c83 bl_83 br_83 wl_80 vdd gnd cell_6t
Xbit_r81_c83 bl_83 br_83 wl_81 vdd gnd cell_6t
Xbit_r82_c83 bl_83 br_83 wl_82 vdd gnd cell_6t
Xbit_r83_c83 bl_83 br_83 wl_83 vdd gnd cell_6t
Xbit_r84_c83 bl_83 br_83 wl_84 vdd gnd cell_6t
Xbit_r85_c83 bl_83 br_83 wl_85 vdd gnd cell_6t
Xbit_r86_c83 bl_83 br_83 wl_86 vdd gnd cell_6t
Xbit_r87_c83 bl_83 br_83 wl_87 vdd gnd cell_6t
Xbit_r88_c83 bl_83 br_83 wl_88 vdd gnd cell_6t
Xbit_r89_c83 bl_83 br_83 wl_89 vdd gnd cell_6t
Xbit_r90_c83 bl_83 br_83 wl_90 vdd gnd cell_6t
Xbit_r91_c83 bl_83 br_83 wl_91 vdd gnd cell_6t
Xbit_r92_c83 bl_83 br_83 wl_92 vdd gnd cell_6t
Xbit_r93_c83 bl_83 br_83 wl_93 vdd gnd cell_6t
Xbit_r94_c83 bl_83 br_83 wl_94 vdd gnd cell_6t
Xbit_r95_c83 bl_83 br_83 wl_95 vdd gnd cell_6t
Xbit_r96_c83 bl_83 br_83 wl_96 vdd gnd cell_6t
Xbit_r97_c83 bl_83 br_83 wl_97 vdd gnd cell_6t
Xbit_r98_c83 bl_83 br_83 wl_98 vdd gnd cell_6t
Xbit_r99_c83 bl_83 br_83 wl_99 vdd gnd cell_6t
Xbit_r100_c83 bl_83 br_83 wl_100 vdd gnd cell_6t
Xbit_r101_c83 bl_83 br_83 wl_101 vdd gnd cell_6t
Xbit_r102_c83 bl_83 br_83 wl_102 vdd gnd cell_6t
Xbit_r103_c83 bl_83 br_83 wl_103 vdd gnd cell_6t
Xbit_r104_c83 bl_83 br_83 wl_104 vdd gnd cell_6t
Xbit_r105_c83 bl_83 br_83 wl_105 vdd gnd cell_6t
Xbit_r106_c83 bl_83 br_83 wl_106 vdd gnd cell_6t
Xbit_r107_c83 bl_83 br_83 wl_107 vdd gnd cell_6t
Xbit_r108_c83 bl_83 br_83 wl_108 vdd gnd cell_6t
Xbit_r109_c83 bl_83 br_83 wl_109 vdd gnd cell_6t
Xbit_r110_c83 bl_83 br_83 wl_110 vdd gnd cell_6t
Xbit_r111_c83 bl_83 br_83 wl_111 vdd gnd cell_6t
Xbit_r112_c83 bl_83 br_83 wl_112 vdd gnd cell_6t
Xbit_r113_c83 bl_83 br_83 wl_113 vdd gnd cell_6t
Xbit_r114_c83 bl_83 br_83 wl_114 vdd gnd cell_6t
Xbit_r115_c83 bl_83 br_83 wl_115 vdd gnd cell_6t
Xbit_r116_c83 bl_83 br_83 wl_116 vdd gnd cell_6t
Xbit_r117_c83 bl_83 br_83 wl_117 vdd gnd cell_6t
Xbit_r118_c83 bl_83 br_83 wl_118 vdd gnd cell_6t
Xbit_r119_c83 bl_83 br_83 wl_119 vdd gnd cell_6t
Xbit_r120_c83 bl_83 br_83 wl_120 vdd gnd cell_6t
Xbit_r121_c83 bl_83 br_83 wl_121 vdd gnd cell_6t
Xbit_r122_c83 bl_83 br_83 wl_122 vdd gnd cell_6t
Xbit_r123_c83 bl_83 br_83 wl_123 vdd gnd cell_6t
Xbit_r124_c83 bl_83 br_83 wl_124 vdd gnd cell_6t
Xbit_r125_c83 bl_83 br_83 wl_125 vdd gnd cell_6t
Xbit_r126_c83 bl_83 br_83 wl_126 vdd gnd cell_6t
Xbit_r127_c83 bl_83 br_83 wl_127 vdd gnd cell_6t
Xbit_r128_c83 bl_83 br_83 wl_128 vdd gnd cell_6t
Xbit_r129_c83 bl_83 br_83 wl_129 vdd gnd cell_6t
Xbit_r130_c83 bl_83 br_83 wl_130 vdd gnd cell_6t
Xbit_r131_c83 bl_83 br_83 wl_131 vdd gnd cell_6t
Xbit_r132_c83 bl_83 br_83 wl_132 vdd gnd cell_6t
Xbit_r133_c83 bl_83 br_83 wl_133 vdd gnd cell_6t
Xbit_r134_c83 bl_83 br_83 wl_134 vdd gnd cell_6t
Xbit_r135_c83 bl_83 br_83 wl_135 vdd gnd cell_6t
Xbit_r136_c83 bl_83 br_83 wl_136 vdd gnd cell_6t
Xbit_r137_c83 bl_83 br_83 wl_137 vdd gnd cell_6t
Xbit_r138_c83 bl_83 br_83 wl_138 vdd gnd cell_6t
Xbit_r139_c83 bl_83 br_83 wl_139 vdd gnd cell_6t
Xbit_r140_c83 bl_83 br_83 wl_140 vdd gnd cell_6t
Xbit_r141_c83 bl_83 br_83 wl_141 vdd gnd cell_6t
Xbit_r142_c83 bl_83 br_83 wl_142 vdd gnd cell_6t
Xbit_r143_c83 bl_83 br_83 wl_143 vdd gnd cell_6t
Xbit_r144_c83 bl_83 br_83 wl_144 vdd gnd cell_6t
Xbit_r145_c83 bl_83 br_83 wl_145 vdd gnd cell_6t
Xbit_r146_c83 bl_83 br_83 wl_146 vdd gnd cell_6t
Xbit_r147_c83 bl_83 br_83 wl_147 vdd gnd cell_6t
Xbit_r148_c83 bl_83 br_83 wl_148 vdd gnd cell_6t
Xbit_r149_c83 bl_83 br_83 wl_149 vdd gnd cell_6t
Xbit_r150_c83 bl_83 br_83 wl_150 vdd gnd cell_6t
Xbit_r151_c83 bl_83 br_83 wl_151 vdd gnd cell_6t
Xbit_r152_c83 bl_83 br_83 wl_152 vdd gnd cell_6t
Xbit_r153_c83 bl_83 br_83 wl_153 vdd gnd cell_6t
Xbit_r154_c83 bl_83 br_83 wl_154 vdd gnd cell_6t
Xbit_r155_c83 bl_83 br_83 wl_155 vdd gnd cell_6t
Xbit_r156_c83 bl_83 br_83 wl_156 vdd gnd cell_6t
Xbit_r157_c83 bl_83 br_83 wl_157 vdd gnd cell_6t
Xbit_r158_c83 bl_83 br_83 wl_158 vdd gnd cell_6t
Xbit_r159_c83 bl_83 br_83 wl_159 vdd gnd cell_6t
Xbit_r160_c83 bl_83 br_83 wl_160 vdd gnd cell_6t
Xbit_r161_c83 bl_83 br_83 wl_161 vdd gnd cell_6t
Xbit_r162_c83 bl_83 br_83 wl_162 vdd gnd cell_6t
Xbit_r163_c83 bl_83 br_83 wl_163 vdd gnd cell_6t
Xbit_r164_c83 bl_83 br_83 wl_164 vdd gnd cell_6t
Xbit_r165_c83 bl_83 br_83 wl_165 vdd gnd cell_6t
Xbit_r166_c83 bl_83 br_83 wl_166 vdd gnd cell_6t
Xbit_r167_c83 bl_83 br_83 wl_167 vdd gnd cell_6t
Xbit_r168_c83 bl_83 br_83 wl_168 vdd gnd cell_6t
Xbit_r169_c83 bl_83 br_83 wl_169 vdd gnd cell_6t
Xbit_r170_c83 bl_83 br_83 wl_170 vdd gnd cell_6t
Xbit_r171_c83 bl_83 br_83 wl_171 vdd gnd cell_6t
Xbit_r172_c83 bl_83 br_83 wl_172 vdd gnd cell_6t
Xbit_r173_c83 bl_83 br_83 wl_173 vdd gnd cell_6t
Xbit_r174_c83 bl_83 br_83 wl_174 vdd gnd cell_6t
Xbit_r175_c83 bl_83 br_83 wl_175 vdd gnd cell_6t
Xbit_r176_c83 bl_83 br_83 wl_176 vdd gnd cell_6t
Xbit_r177_c83 bl_83 br_83 wl_177 vdd gnd cell_6t
Xbit_r178_c83 bl_83 br_83 wl_178 vdd gnd cell_6t
Xbit_r179_c83 bl_83 br_83 wl_179 vdd gnd cell_6t
Xbit_r180_c83 bl_83 br_83 wl_180 vdd gnd cell_6t
Xbit_r181_c83 bl_83 br_83 wl_181 vdd gnd cell_6t
Xbit_r182_c83 bl_83 br_83 wl_182 vdd gnd cell_6t
Xbit_r183_c83 bl_83 br_83 wl_183 vdd gnd cell_6t
Xbit_r184_c83 bl_83 br_83 wl_184 vdd gnd cell_6t
Xbit_r185_c83 bl_83 br_83 wl_185 vdd gnd cell_6t
Xbit_r186_c83 bl_83 br_83 wl_186 vdd gnd cell_6t
Xbit_r187_c83 bl_83 br_83 wl_187 vdd gnd cell_6t
Xbit_r188_c83 bl_83 br_83 wl_188 vdd gnd cell_6t
Xbit_r189_c83 bl_83 br_83 wl_189 vdd gnd cell_6t
Xbit_r190_c83 bl_83 br_83 wl_190 vdd gnd cell_6t
Xbit_r191_c83 bl_83 br_83 wl_191 vdd gnd cell_6t
Xbit_r192_c83 bl_83 br_83 wl_192 vdd gnd cell_6t
Xbit_r193_c83 bl_83 br_83 wl_193 vdd gnd cell_6t
Xbit_r194_c83 bl_83 br_83 wl_194 vdd gnd cell_6t
Xbit_r195_c83 bl_83 br_83 wl_195 vdd gnd cell_6t
Xbit_r196_c83 bl_83 br_83 wl_196 vdd gnd cell_6t
Xbit_r197_c83 bl_83 br_83 wl_197 vdd gnd cell_6t
Xbit_r198_c83 bl_83 br_83 wl_198 vdd gnd cell_6t
Xbit_r199_c83 bl_83 br_83 wl_199 vdd gnd cell_6t
Xbit_r200_c83 bl_83 br_83 wl_200 vdd gnd cell_6t
Xbit_r201_c83 bl_83 br_83 wl_201 vdd gnd cell_6t
Xbit_r202_c83 bl_83 br_83 wl_202 vdd gnd cell_6t
Xbit_r203_c83 bl_83 br_83 wl_203 vdd gnd cell_6t
Xbit_r204_c83 bl_83 br_83 wl_204 vdd gnd cell_6t
Xbit_r205_c83 bl_83 br_83 wl_205 vdd gnd cell_6t
Xbit_r206_c83 bl_83 br_83 wl_206 vdd gnd cell_6t
Xbit_r207_c83 bl_83 br_83 wl_207 vdd gnd cell_6t
Xbit_r208_c83 bl_83 br_83 wl_208 vdd gnd cell_6t
Xbit_r209_c83 bl_83 br_83 wl_209 vdd gnd cell_6t
Xbit_r210_c83 bl_83 br_83 wl_210 vdd gnd cell_6t
Xbit_r211_c83 bl_83 br_83 wl_211 vdd gnd cell_6t
Xbit_r212_c83 bl_83 br_83 wl_212 vdd gnd cell_6t
Xbit_r213_c83 bl_83 br_83 wl_213 vdd gnd cell_6t
Xbit_r214_c83 bl_83 br_83 wl_214 vdd gnd cell_6t
Xbit_r215_c83 bl_83 br_83 wl_215 vdd gnd cell_6t
Xbit_r216_c83 bl_83 br_83 wl_216 vdd gnd cell_6t
Xbit_r217_c83 bl_83 br_83 wl_217 vdd gnd cell_6t
Xbit_r218_c83 bl_83 br_83 wl_218 vdd gnd cell_6t
Xbit_r219_c83 bl_83 br_83 wl_219 vdd gnd cell_6t
Xbit_r220_c83 bl_83 br_83 wl_220 vdd gnd cell_6t
Xbit_r221_c83 bl_83 br_83 wl_221 vdd gnd cell_6t
Xbit_r222_c83 bl_83 br_83 wl_222 vdd gnd cell_6t
Xbit_r223_c83 bl_83 br_83 wl_223 vdd gnd cell_6t
Xbit_r224_c83 bl_83 br_83 wl_224 vdd gnd cell_6t
Xbit_r225_c83 bl_83 br_83 wl_225 vdd gnd cell_6t
Xbit_r226_c83 bl_83 br_83 wl_226 vdd gnd cell_6t
Xbit_r227_c83 bl_83 br_83 wl_227 vdd gnd cell_6t
Xbit_r228_c83 bl_83 br_83 wl_228 vdd gnd cell_6t
Xbit_r229_c83 bl_83 br_83 wl_229 vdd gnd cell_6t
Xbit_r230_c83 bl_83 br_83 wl_230 vdd gnd cell_6t
Xbit_r231_c83 bl_83 br_83 wl_231 vdd gnd cell_6t
Xbit_r232_c83 bl_83 br_83 wl_232 vdd gnd cell_6t
Xbit_r233_c83 bl_83 br_83 wl_233 vdd gnd cell_6t
Xbit_r234_c83 bl_83 br_83 wl_234 vdd gnd cell_6t
Xbit_r235_c83 bl_83 br_83 wl_235 vdd gnd cell_6t
Xbit_r236_c83 bl_83 br_83 wl_236 vdd gnd cell_6t
Xbit_r237_c83 bl_83 br_83 wl_237 vdd gnd cell_6t
Xbit_r238_c83 bl_83 br_83 wl_238 vdd gnd cell_6t
Xbit_r239_c83 bl_83 br_83 wl_239 vdd gnd cell_6t
Xbit_r240_c83 bl_83 br_83 wl_240 vdd gnd cell_6t
Xbit_r241_c83 bl_83 br_83 wl_241 vdd gnd cell_6t
Xbit_r242_c83 bl_83 br_83 wl_242 vdd gnd cell_6t
Xbit_r243_c83 bl_83 br_83 wl_243 vdd gnd cell_6t
Xbit_r244_c83 bl_83 br_83 wl_244 vdd gnd cell_6t
Xbit_r245_c83 bl_83 br_83 wl_245 vdd gnd cell_6t
Xbit_r246_c83 bl_83 br_83 wl_246 vdd gnd cell_6t
Xbit_r247_c83 bl_83 br_83 wl_247 vdd gnd cell_6t
Xbit_r248_c83 bl_83 br_83 wl_248 vdd gnd cell_6t
Xbit_r249_c83 bl_83 br_83 wl_249 vdd gnd cell_6t
Xbit_r250_c83 bl_83 br_83 wl_250 vdd gnd cell_6t
Xbit_r251_c83 bl_83 br_83 wl_251 vdd gnd cell_6t
Xbit_r252_c83 bl_83 br_83 wl_252 vdd gnd cell_6t
Xbit_r253_c83 bl_83 br_83 wl_253 vdd gnd cell_6t
Xbit_r254_c83 bl_83 br_83 wl_254 vdd gnd cell_6t
Xbit_r255_c83 bl_83 br_83 wl_255 vdd gnd cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd cell_6t
Xbit_r1_c84 bl_84 br_84 wl_1 vdd gnd cell_6t
Xbit_r2_c84 bl_84 br_84 wl_2 vdd gnd cell_6t
Xbit_r3_c84 bl_84 br_84 wl_3 vdd gnd cell_6t
Xbit_r4_c84 bl_84 br_84 wl_4 vdd gnd cell_6t
Xbit_r5_c84 bl_84 br_84 wl_5 vdd gnd cell_6t
Xbit_r6_c84 bl_84 br_84 wl_6 vdd gnd cell_6t
Xbit_r7_c84 bl_84 br_84 wl_7 vdd gnd cell_6t
Xbit_r8_c84 bl_84 br_84 wl_8 vdd gnd cell_6t
Xbit_r9_c84 bl_84 br_84 wl_9 vdd gnd cell_6t
Xbit_r10_c84 bl_84 br_84 wl_10 vdd gnd cell_6t
Xbit_r11_c84 bl_84 br_84 wl_11 vdd gnd cell_6t
Xbit_r12_c84 bl_84 br_84 wl_12 vdd gnd cell_6t
Xbit_r13_c84 bl_84 br_84 wl_13 vdd gnd cell_6t
Xbit_r14_c84 bl_84 br_84 wl_14 vdd gnd cell_6t
Xbit_r15_c84 bl_84 br_84 wl_15 vdd gnd cell_6t
Xbit_r16_c84 bl_84 br_84 wl_16 vdd gnd cell_6t
Xbit_r17_c84 bl_84 br_84 wl_17 vdd gnd cell_6t
Xbit_r18_c84 bl_84 br_84 wl_18 vdd gnd cell_6t
Xbit_r19_c84 bl_84 br_84 wl_19 vdd gnd cell_6t
Xbit_r20_c84 bl_84 br_84 wl_20 vdd gnd cell_6t
Xbit_r21_c84 bl_84 br_84 wl_21 vdd gnd cell_6t
Xbit_r22_c84 bl_84 br_84 wl_22 vdd gnd cell_6t
Xbit_r23_c84 bl_84 br_84 wl_23 vdd gnd cell_6t
Xbit_r24_c84 bl_84 br_84 wl_24 vdd gnd cell_6t
Xbit_r25_c84 bl_84 br_84 wl_25 vdd gnd cell_6t
Xbit_r26_c84 bl_84 br_84 wl_26 vdd gnd cell_6t
Xbit_r27_c84 bl_84 br_84 wl_27 vdd gnd cell_6t
Xbit_r28_c84 bl_84 br_84 wl_28 vdd gnd cell_6t
Xbit_r29_c84 bl_84 br_84 wl_29 vdd gnd cell_6t
Xbit_r30_c84 bl_84 br_84 wl_30 vdd gnd cell_6t
Xbit_r31_c84 bl_84 br_84 wl_31 vdd gnd cell_6t
Xbit_r32_c84 bl_84 br_84 wl_32 vdd gnd cell_6t
Xbit_r33_c84 bl_84 br_84 wl_33 vdd gnd cell_6t
Xbit_r34_c84 bl_84 br_84 wl_34 vdd gnd cell_6t
Xbit_r35_c84 bl_84 br_84 wl_35 vdd gnd cell_6t
Xbit_r36_c84 bl_84 br_84 wl_36 vdd gnd cell_6t
Xbit_r37_c84 bl_84 br_84 wl_37 vdd gnd cell_6t
Xbit_r38_c84 bl_84 br_84 wl_38 vdd gnd cell_6t
Xbit_r39_c84 bl_84 br_84 wl_39 vdd gnd cell_6t
Xbit_r40_c84 bl_84 br_84 wl_40 vdd gnd cell_6t
Xbit_r41_c84 bl_84 br_84 wl_41 vdd gnd cell_6t
Xbit_r42_c84 bl_84 br_84 wl_42 vdd gnd cell_6t
Xbit_r43_c84 bl_84 br_84 wl_43 vdd gnd cell_6t
Xbit_r44_c84 bl_84 br_84 wl_44 vdd gnd cell_6t
Xbit_r45_c84 bl_84 br_84 wl_45 vdd gnd cell_6t
Xbit_r46_c84 bl_84 br_84 wl_46 vdd gnd cell_6t
Xbit_r47_c84 bl_84 br_84 wl_47 vdd gnd cell_6t
Xbit_r48_c84 bl_84 br_84 wl_48 vdd gnd cell_6t
Xbit_r49_c84 bl_84 br_84 wl_49 vdd gnd cell_6t
Xbit_r50_c84 bl_84 br_84 wl_50 vdd gnd cell_6t
Xbit_r51_c84 bl_84 br_84 wl_51 vdd gnd cell_6t
Xbit_r52_c84 bl_84 br_84 wl_52 vdd gnd cell_6t
Xbit_r53_c84 bl_84 br_84 wl_53 vdd gnd cell_6t
Xbit_r54_c84 bl_84 br_84 wl_54 vdd gnd cell_6t
Xbit_r55_c84 bl_84 br_84 wl_55 vdd gnd cell_6t
Xbit_r56_c84 bl_84 br_84 wl_56 vdd gnd cell_6t
Xbit_r57_c84 bl_84 br_84 wl_57 vdd gnd cell_6t
Xbit_r58_c84 bl_84 br_84 wl_58 vdd gnd cell_6t
Xbit_r59_c84 bl_84 br_84 wl_59 vdd gnd cell_6t
Xbit_r60_c84 bl_84 br_84 wl_60 vdd gnd cell_6t
Xbit_r61_c84 bl_84 br_84 wl_61 vdd gnd cell_6t
Xbit_r62_c84 bl_84 br_84 wl_62 vdd gnd cell_6t
Xbit_r63_c84 bl_84 br_84 wl_63 vdd gnd cell_6t
Xbit_r64_c84 bl_84 br_84 wl_64 vdd gnd cell_6t
Xbit_r65_c84 bl_84 br_84 wl_65 vdd gnd cell_6t
Xbit_r66_c84 bl_84 br_84 wl_66 vdd gnd cell_6t
Xbit_r67_c84 bl_84 br_84 wl_67 vdd gnd cell_6t
Xbit_r68_c84 bl_84 br_84 wl_68 vdd gnd cell_6t
Xbit_r69_c84 bl_84 br_84 wl_69 vdd gnd cell_6t
Xbit_r70_c84 bl_84 br_84 wl_70 vdd gnd cell_6t
Xbit_r71_c84 bl_84 br_84 wl_71 vdd gnd cell_6t
Xbit_r72_c84 bl_84 br_84 wl_72 vdd gnd cell_6t
Xbit_r73_c84 bl_84 br_84 wl_73 vdd gnd cell_6t
Xbit_r74_c84 bl_84 br_84 wl_74 vdd gnd cell_6t
Xbit_r75_c84 bl_84 br_84 wl_75 vdd gnd cell_6t
Xbit_r76_c84 bl_84 br_84 wl_76 vdd gnd cell_6t
Xbit_r77_c84 bl_84 br_84 wl_77 vdd gnd cell_6t
Xbit_r78_c84 bl_84 br_84 wl_78 vdd gnd cell_6t
Xbit_r79_c84 bl_84 br_84 wl_79 vdd gnd cell_6t
Xbit_r80_c84 bl_84 br_84 wl_80 vdd gnd cell_6t
Xbit_r81_c84 bl_84 br_84 wl_81 vdd gnd cell_6t
Xbit_r82_c84 bl_84 br_84 wl_82 vdd gnd cell_6t
Xbit_r83_c84 bl_84 br_84 wl_83 vdd gnd cell_6t
Xbit_r84_c84 bl_84 br_84 wl_84 vdd gnd cell_6t
Xbit_r85_c84 bl_84 br_84 wl_85 vdd gnd cell_6t
Xbit_r86_c84 bl_84 br_84 wl_86 vdd gnd cell_6t
Xbit_r87_c84 bl_84 br_84 wl_87 vdd gnd cell_6t
Xbit_r88_c84 bl_84 br_84 wl_88 vdd gnd cell_6t
Xbit_r89_c84 bl_84 br_84 wl_89 vdd gnd cell_6t
Xbit_r90_c84 bl_84 br_84 wl_90 vdd gnd cell_6t
Xbit_r91_c84 bl_84 br_84 wl_91 vdd gnd cell_6t
Xbit_r92_c84 bl_84 br_84 wl_92 vdd gnd cell_6t
Xbit_r93_c84 bl_84 br_84 wl_93 vdd gnd cell_6t
Xbit_r94_c84 bl_84 br_84 wl_94 vdd gnd cell_6t
Xbit_r95_c84 bl_84 br_84 wl_95 vdd gnd cell_6t
Xbit_r96_c84 bl_84 br_84 wl_96 vdd gnd cell_6t
Xbit_r97_c84 bl_84 br_84 wl_97 vdd gnd cell_6t
Xbit_r98_c84 bl_84 br_84 wl_98 vdd gnd cell_6t
Xbit_r99_c84 bl_84 br_84 wl_99 vdd gnd cell_6t
Xbit_r100_c84 bl_84 br_84 wl_100 vdd gnd cell_6t
Xbit_r101_c84 bl_84 br_84 wl_101 vdd gnd cell_6t
Xbit_r102_c84 bl_84 br_84 wl_102 vdd gnd cell_6t
Xbit_r103_c84 bl_84 br_84 wl_103 vdd gnd cell_6t
Xbit_r104_c84 bl_84 br_84 wl_104 vdd gnd cell_6t
Xbit_r105_c84 bl_84 br_84 wl_105 vdd gnd cell_6t
Xbit_r106_c84 bl_84 br_84 wl_106 vdd gnd cell_6t
Xbit_r107_c84 bl_84 br_84 wl_107 vdd gnd cell_6t
Xbit_r108_c84 bl_84 br_84 wl_108 vdd gnd cell_6t
Xbit_r109_c84 bl_84 br_84 wl_109 vdd gnd cell_6t
Xbit_r110_c84 bl_84 br_84 wl_110 vdd gnd cell_6t
Xbit_r111_c84 bl_84 br_84 wl_111 vdd gnd cell_6t
Xbit_r112_c84 bl_84 br_84 wl_112 vdd gnd cell_6t
Xbit_r113_c84 bl_84 br_84 wl_113 vdd gnd cell_6t
Xbit_r114_c84 bl_84 br_84 wl_114 vdd gnd cell_6t
Xbit_r115_c84 bl_84 br_84 wl_115 vdd gnd cell_6t
Xbit_r116_c84 bl_84 br_84 wl_116 vdd gnd cell_6t
Xbit_r117_c84 bl_84 br_84 wl_117 vdd gnd cell_6t
Xbit_r118_c84 bl_84 br_84 wl_118 vdd gnd cell_6t
Xbit_r119_c84 bl_84 br_84 wl_119 vdd gnd cell_6t
Xbit_r120_c84 bl_84 br_84 wl_120 vdd gnd cell_6t
Xbit_r121_c84 bl_84 br_84 wl_121 vdd gnd cell_6t
Xbit_r122_c84 bl_84 br_84 wl_122 vdd gnd cell_6t
Xbit_r123_c84 bl_84 br_84 wl_123 vdd gnd cell_6t
Xbit_r124_c84 bl_84 br_84 wl_124 vdd gnd cell_6t
Xbit_r125_c84 bl_84 br_84 wl_125 vdd gnd cell_6t
Xbit_r126_c84 bl_84 br_84 wl_126 vdd gnd cell_6t
Xbit_r127_c84 bl_84 br_84 wl_127 vdd gnd cell_6t
Xbit_r128_c84 bl_84 br_84 wl_128 vdd gnd cell_6t
Xbit_r129_c84 bl_84 br_84 wl_129 vdd gnd cell_6t
Xbit_r130_c84 bl_84 br_84 wl_130 vdd gnd cell_6t
Xbit_r131_c84 bl_84 br_84 wl_131 vdd gnd cell_6t
Xbit_r132_c84 bl_84 br_84 wl_132 vdd gnd cell_6t
Xbit_r133_c84 bl_84 br_84 wl_133 vdd gnd cell_6t
Xbit_r134_c84 bl_84 br_84 wl_134 vdd gnd cell_6t
Xbit_r135_c84 bl_84 br_84 wl_135 vdd gnd cell_6t
Xbit_r136_c84 bl_84 br_84 wl_136 vdd gnd cell_6t
Xbit_r137_c84 bl_84 br_84 wl_137 vdd gnd cell_6t
Xbit_r138_c84 bl_84 br_84 wl_138 vdd gnd cell_6t
Xbit_r139_c84 bl_84 br_84 wl_139 vdd gnd cell_6t
Xbit_r140_c84 bl_84 br_84 wl_140 vdd gnd cell_6t
Xbit_r141_c84 bl_84 br_84 wl_141 vdd gnd cell_6t
Xbit_r142_c84 bl_84 br_84 wl_142 vdd gnd cell_6t
Xbit_r143_c84 bl_84 br_84 wl_143 vdd gnd cell_6t
Xbit_r144_c84 bl_84 br_84 wl_144 vdd gnd cell_6t
Xbit_r145_c84 bl_84 br_84 wl_145 vdd gnd cell_6t
Xbit_r146_c84 bl_84 br_84 wl_146 vdd gnd cell_6t
Xbit_r147_c84 bl_84 br_84 wl_147 vdd gnd cell_6t
Xbit_r148_c84 bl_84 br_84 wl_148 vdd gnd cell_6t
Xbit_r149_c84 bl_84 br_84 wl_149 vdd gnd cell_6t
Xbit_r150_c84 bl_84 br_84 wl_150 vdd gnd cell_6t
Xbit_r151_c84 bl_84 br_84 wl_151 vdd gnd cell_6t
Xbit_r152_c84 bl_84 br_84 wl_152 vdd gnd cell_6t
Xbit_r153_c84 bl_84 br_84 wl_153 vdd gnd cell_6t
Xbit_r154_c84 bl_84 br_84 wl_154 vdd gnd cell_6t
Xbit_r155_c84 bl_84 br_84 wl_155 vdd gnd cell_6t
Xbit_r156_c84 bl_84 br_84 wl_156 vdd gnd cell_6t
Xbit_r157_c84 bl_84 br_84 wl_157 vdd gnd cell_6t
Xbit_r158_c84 bl_84 br_84 wl_158 vdd gnd cell_6t
Xbit_r159_c84 bl_84 br_84 wl_159 vdd gnd cell_6t
Xbit_r160_c84 bl_84 br_84 wl_160 vdd gnd cell_6t
Xbit_r161_c84 bl_84 br_84 wl_161 vdd gnd cell_6t
Xbit_r162_c84 bl_84 br_84 wl_162 vdd gnd cell_6t
Xbit_r163_c84 bl_84 br_84 wl_163 vdd gnd cell_6t
Xbit_r164_c84 bl_84 br_84 wl_164 vdd gnd cell_6t
Xbit_r165_c84 bl_84 br_84 wl_165 vdd gnd cell_6t
Xbit_r166_c84 bl_84 br_84 wl_166 vdd gnd cell_6t
Xbit_r167_c84 bl_84 br_84 wl_167 vdd gnd cell_6t
Xbit_r168_c84 bl_84 br_84 wl_168 vdd gnd cell_6t
Xbit_r169_c84 bl_84 br_84 wl_169 vdd gnd cell_6t
Xbit_r170_c84 bl_84 br_84 wl_170 vdd gnd cell_6t
Xbit_r171_c84 bl_84 br_84 wl_171 vdd gnd cell_6t
Xbit_r172_c84 bl_84 br_84 wl_172 vdd gnd cell_6t
Xbit_r173_c84 bl_84 br_84 wl_173 vdd gnd cell_6t
Xbit_r174_c84 bl_84 br_84 wl_174 vdd gnd cell_6t
Xbit_r175_c84 bl_84 br_84 wl_175 vdd gnd cell_6t
Xbit_r176_c84 bl_84 br_84 wl_176 vdd gnd cell_6t
Xbit_r177_c84 bl_84 br_84 wl_177 vdd gnd cell_6t
Xbit_r178_c84 bl_84 br_84 wl_178 vdd gnd cell_6t
Xbit_r179_c84 bl_84 br_84 wl_179 vdd gnd cell_6t
Xbit_r180_c84 bl_84 br_84 wl_180 vdd gnd cell_6t
Xbit_r181_c84 bl_84 br_84 wl_181 vdd gnd cell_6t
Xbit_r182_c84 bl_84 br_84 wl_182 vdd gnd cell_6t
Xbit_r183_c84 bl_84 br_84 wl_183 vdd gnd cell_6t
Xbit_r184_c84 bl_84 br_84 wl_184 vdd gnd cell_6t
Xbit_r185_c84 bl_84 br_84 wl_185 vdd gnd cell_6t
Xbit_r186_c84 bl_84 br_84 wl_186 vdd gnd cell_6t
Xbit_r187_c84 bl_84 br_84 wl_187 vdd gnd cell_6t
Xbit_r188_c84 bl_84 br_84 wl_188 vdd gnd cell_6t
Xbit_r189_c84 bl_84 br_84 wl_189 vdd gnd cell_6t
Xbit_r190_c84 bl_84 br_84 wl_190 vdd gnd cell_6t
Xbit_r191_c84 bl_84 br_84 wl_191 vdd gnd cell_6t
Xbit_r192_c84 bl_84 br_84 wl_192 vdd gnd cell_6t
Xbit_r193_c84 bl_84 br_84 wl_193 vdd gnd cell_6t
Xbit_r194_c84 bl_84 br_84 wl_194 vdd gnd cell_6t
Xbit_r195_c84 bl_84 br_84 wl_195 vdd gnd cell_6t
Xbit_r196_c84 bl_84 br_84 wl_196 vdd gnd cell_6t
Xbit_r197_c84 bl_84 br_84 wl_197 vdd gnd cell_6t
Xbit_r198_c84 bl_84 br_84 wl_198 vdd gnd cell_6t
Xbit_r199_c84 bl_84 br_84 wl_199 vdd gnd cell_6t
Xbit_r200_c84 bl_84 br_84 wl_200 vdd gnd cell_6t
Xbit_r201_c84 bl_84 br_84 wl_201 vdd gnd cell_6t
Xbit_r202_c84 bl_84 br_84 wl_202 vdd gnd cell_6t
Xbit_r203_c84 bl_84 br_84 wl_203 vdd gnd cell_6t
Xbit_r204_c84 bl_84 br_84 wl_204 vdd gnd cell_6t
Xbit_r205_c84 bl_84 br_84 wl_205 vdd gnd cell_6t
Xbit_r206_c84 bl_84 br_84 wl_206 vdd gnd cell_6t
Xbit_r207_c84 bl_84 br_84 wl_207 vdd gnd cell_6t
Xbit_r208_c84 bl_84 br_84 wl_208 vdd gnd cell_6t
Xbit_r209_c84 bl_84 br_84 wl_209 vdd gnd cell_6t
Xbit_r210_c84 bl_84 br_84 wl_210 vdd gnd cell_6t
Xbit_r211_c84 bl_84 br_84 wl_211 vdd gnd cell_6t
Xbit_r212_c84 bl_84 br_84 wl_212 vdd gnd cell_6t
Xbit_r213_c84 bl_84 br_84 wl_213 vdd gnd cell_6t
Xbit_r214_c84 bl_84 br_84 wl_214 vdd gnd cell_6t
Xbit_r215_c84 bl_84 br_84 wl_215 vdd gnd cell_6t
Xbit_r216_c84 bl_84 br_84 wl_216 vdd gnd cell_6t
Xbit_r217_c84 bl_84 br_84 wl_217 vdd gnd cell_6t
Xbit_r218_c84 bl_84 br_84 wl_218 vdd gnd cell_6t
Xbit_r219_c84 bl_84 br_84 wl_219 vdd gnd cell_6t
Xbit_r220_c84 bl_84 br_84 wl_220 vdd gnd cell_6t
Xbit_r221_c84 bl_84 br_84 wl_221 vdd gnd cell_6t
Xbit_r222_c84 bl_84 br_84 wl_222 vdd gnd cell_6t
Xbit_r223_c84 bl_84 br_84 wl_223 vdd gnd cell_6t
Xbit_r224_c84 bl_84 br_84 wl_224 vdd gnd cell_6t
Xbit_r225_c84 bl_84 br_84 wl_225 vdd gnd cell_6t
Xbit_r226_c84 bl_84 br_84 wl_226 vdd gnd cell_6t
Xbit_r227_c84 bl_84 br_84 wl_227 vdd gnd cell_6t
Xbit_r228_c84 bl_84 br_84 wl_228 vdd gnd cell_6t
Xbit_r229_c84 bl_84 br_84 wl_229 vdd gnd cell_6t
Xbit_r230_c84 bl_84 br_84 wl_230 vdd gnd cell_6t
Xbit_r231_c84 bl_84 br_84 wl_231 vdd gnd cell_6t
Xbit_r232_c84 bl_84 br_84 wl_232 vdd gnd cell_6t
Xbit_r233_c84 bl_84 br_84 wl_233 vdd gnd cell_6t
Xbit_r234_c84 bl_84 br_84 wl_234 vdd gnd cell_6t
Xbit_r235_c84 bl_84 br_84 wl_235 vdd gnd cell_6t
Xbit_r236_c84 bl_84 br_84 wl_236 vdd gnd cell_6t
Xbit_r237_c84 bl_84 br_84 wl_237 vdd gnd cell_6t
Xbit_r238_c84 bl_84 br_84 wl_238 vdd gnd cell_6t
Xbit_r239_c84 bl_84 br_84 wl_239 vdd gnd cell_6t
Xbit_r240_c84 bl_84 br_84 wl_240 vdd gnd cell_6t
Xbit_r241_c84 bl_84 br_84 wl_241 vdd gnd cell_6t
Xbit_r242_c84 bl_84 br_84 wl_242 vdd gnd cell_6t
Xbit_r243_c84 bl_84 br_84 wl_243 vdd gnd cell_6t
Xbit_r244_c84 bl_84 br_84 wl_244 vdd gnd cell_6t
Xbit_r245_c84 bl_84 br_84 wl_245 vdd gnd cell_6t
Xbit_r246_c84 bl_84 br_84 wl_246 vdd gnd cell_6t
Xbit_r247_c84 bl_84 br_84 wl_247 vdd gnd cell_6t
Xbit_r248_c84 bl_84 br_84 wl_248 vdd gnd cell_6t
Xbit_r249_c84 bl_84 br_84 wl_249 vdd gnd cell_6t
Xbit_r250_c84 bl_84 br_84 wl_250 vdd gnd cell_6t
Xbit_r251_c84 bl_84 br_84 wl_251 vdd gnd cell_6t
Xbit_r252_c84 bl_84 br_84 wl_252 vdd gnd cell_6t
Xbit_r253_c84 bl_84 br_84 wl_253 vdd gnd cell_6t
Xbit_r254_c84 bl_84 br_84 wl_254 vdd gnd cell_6t
Xbit_r255_c84 bl_84 br_84 wl_255 vdd gnd cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd cell_6t
Xbit_r1_c85 bl_85 br_85 wl_1 vdd gnd cell_6t
Xbit_r2_c85 bl_85 br_85 wl_2 vdd gnd cell_6t
Xbit_r3_c85 bl_85 br_85 wl_3 vdd gnd cell_6t
Xbit_r4_c85 bl_85 br_85 wl_4 vdd gnd cell_6t
Xbit_r5_c85 bl_85 br_85 wl_5 vdd gnd cell_6t
Xbit_r6_c85 bl_85 br_85 wl_6 vdd gnd cell_6t
Xbit_r7_c85 bl_85 br_85 wl_7 vdd gnd cell_6t
Xbit_r8_c85 bl_85 br_85 wl_8 vdd gnd cell_6t
Xbit_r9_c85 bl_85 br_85 wl_9 vdd gnd cell_6t
Xbit_r10_c85 bl_85 br_85 wl_10 vdd gnd cell_6t
Xbit_r11_c85 bl_85 br_85 wl_11 vdd gnd cell_6t
Xbit_r12_c85 bl_85 br_85 wl_12 vdd gnd cell_6t
Xbit_r13_c85 bl_85 br_85 wl_13 vdd gnd cell_6t
Xbit_r14_c85 bl_85 br_85 wl_14 vdd gnd cell_6t
Xbit_r15_c85 bl_85 br_85 wl_15 vdd gnd cell_6t
Xbit_r16_c85 bl_85 br_85 wl_16 vdd gnd cell_6t
Xbit_r17_c85 bl_85 br_85 wl_17 vdd gnd cell_6t
Xbit_r18_c85 bl_85 br_85 wl_18 vdd gnd cell_6t
Xbit_r19_c85 bl_85 br_85 wl_19 vdd gnd cell_6t
Xbit_r20_c85 bl_85 br_85 wl_20 vdd gnd cell_6t
Xbit_r21_c85 bl_85 br_85 wl_21 vdd gnd cell_6t
Xbit_r22_c85 bl_85 br_85 wl_22 vdd gnd cell_6t
Xbit_r23_c85 bl_85 br_85 wl_23 vdd gnd cell_6t
Xbit_r24_c85 bl_85 br_85 wl_24 vdd gnd cell_6t
Xbit_r25_c85 bl_85 br_85 wl_25 vdd gnd cell_6t
Xbit_r26_c85 bl_85 br_85 wl_26 vdd gnd cell_6t
Xbit_r27_c85 bl_85 br_85 wl_27 vdd gnd cell_6t
Xbit_r28_c85 bl_85 br_85 wl_28 vdd gnd cell_6t
Xbit_r29_c85 bl_85 br_85 wl_29 vdd gnd cell_6t
Xbit_r30_c85 bl_85 br_85 wl_30 vdd gnd cell_6t
Xbit_r31_c85 bl_85 br_85 wl_31 vdd gnd cell_6t
Xbit_r32_c85 bl_85 br_85 wl_32 vdd gnd cell_6t
Xbit_r33_c85 bl_85 br_85 wl_33 vdd gnd cell_6t
Xbit_r34_c85 bl_85 br_85 wl_34 vdd gnd cell_6t
Xbit_r35_c85 bl_85 br_85 wl_35 vdd gnd cell_6t
Xbit_r36_c85 bl_85 br_85 wl_36 vdd gnd cell_6t
Xbit_r37_c85 bl_85 br_85 wl_37 vdd gnd cell_6t
Xbit_r38_c85 bl_85 br_85 wl_38 vdd gnd cell_6t
Xbit_r39_c85 bl_85 br_85 wl_39 vdd gnd cell_6t
Xbit_r40_c85 bl_85 br_85 wl_40 vdd gnd cell_6t
Xbit_r41_c85 bl_85 br_85 wl_41 vdd gnd cell_6t
Xbit_r42_c85 bl_85 br_85 wl_42 vdd gnd cell_6t
Xbit_r43_c85 bl_85 br_85 wl_43 vdd gnd cell_6t
Xbit_r44_c85 bl_85 br_85 wl_44 vdd gnd cell_6t
Xbit_r45_c85 bl_85 br_85 wl_45 vdd gnd cell_6t
Xbit_r46_c85 bl_85 br_85 wl_46 vdd gnd cell_6t
Xbit_r47_c85 bl_85 br_85 wl_47 vdd gnd cell_6t
Xbit_r48_c85 bl_85 br_85 wl_48 vdd gnd cell_6t
Xbit_r49_c85 bl_85 br_85 wl_49 vdd gnd cell_6t
Xbit_r50_c85 bl_85 br_85 wl_50 vdd gnd cell_6t
Xbit_r51_c85 bl_85 br_85 wl_51 vdd gnd cell_6t
Xbit_r52_c85 bl_85 br_85 wl_52 vdd gnd cell_6t
Xbit_r53_c85 bl_85 br_85 wl_53 vdd gnd cell_6t
Xbit_r54_c85 bl_85 br_85 wl_54 vdd gnd cell_6t
Xbit_r55_c85 bl_85 br_85 wl_55 vdd gnd cell_6t
Xbit_r56_c85 bl_85 br_85 wl_56 vdd gnd cell_6t
Xbit_r57_c85 bl_85 br_85 wl_57 vdd gnd cell_6t
Xbit_r58_c85 bl_85 br_85 wl_58 vdd gnd cell_6t
Xbit_r59_c85 bl_85 br_85 wl_59 vdd gnd cell_6t
Xbit_r60_c85 bl_85 br_85 wl_60 vdd gnd cell_6t
Xbit_r61_c85 bl_85 br_85 wl_61 vdd gnd cell_6t
Xbit_r62_c85 bl_85 br_85 wl_62 vdd gnd cell_6t
Xbit_r63_c85 bl_85 br_85 wl_63 vdd gnd cell_6t
Xbit_r64_c85 bl_85 br_85 wl_64 vdd gnd cell_6t
Xbit_r65_c85 bl_85 br_85 wl_65 vdd gnd cell_6t
Xbit_r66_c85 bl_85 br_85 wl_66 vdd gnd cell_6t
Xbit_r67_c85 bl_85 br_85 wl_67 vdd gnd cell_6t
Xbit_r68_c85 bl_85 br_85 wl_68 vdd gnd cell_6t
Xbit_r69_c85 bl_85 br_85 wl_69 vdd gnd cell_6t
Xbit_r70_c85 bl_85 br_85 wl_70 vdd gnd cell_6t
Xbit_r71_c85 bl_85 br_85 wl_71 vdd gnd cell_6t
Xbit_r72_c85 bl_85 br_85 wl_72 vdd gnd cell_6t
Xbit_r73_c85 bl_85 br_85 wl_73 vdd gnd cell_6t
Xbit_r74_c85 bl_85 br_85 wl_74 vdd gnd cell_6t
Xbit_r75_c85 bl_85 br_85 wl_75 vdd gnd cell_6t
Xbit_r76_c85 bl_85 br_85 wl_76 vdd gnd cell_6t
Xbit_r77_c85 bl_85 br_85 wl_77 vdd gnd cell_6t
Xbit_r78_c85 bl_85 br_85 wl_78 vdd gnd cell_6t
Xbit_r79_c85 bl_85 br_85 wl_79 vdd gnd cell_6t
Xbit_r80_c85 bl_85 br_85 wl_80 vdd gnd cell_6t
Xbit_r81_c85 bl_85 br_85 wl_81 vdd gnd cell_6t
Xbit_r82_c85 bl_85 br_85 wl_82 vdd gnd cell_6t
Xbit_r83_c85 bl_85 br_85 wl_83 vdd gnd cell_6t
Xbit_r84_c85 bl_85 br_85 wl_84 vdd gnd cell_6t
Xbit_r85_c85 bl_85 br_85 wl_85 vdd gnd cell_6t
Xbit_r86_c85 bl_85 br_85 wl_86 vdd gnd cell_6t
Xbit_r87_c85 bl_85 br_85 wl_87 vdd gnd cell_6t
Xbit_r88_c85 bl_85 br_85 wl_88 vdd gnd cell_6t
Xbit_r89_c85 bl_85 br_85 wl_89 vdd gnd cell_6t
Xbit_r90_c85 bl_85 br_85 wl_90 vdd gnd cell_6t
Xbit_r91_c85 bl_85 br_85 wl_91 vdd gnd cell_6t
Xbit_r92_c85 bl_85 br_85 wl_92 vdd gnd cell_6t
Xbit_r93_c85 bl_85 br_85 wl_93 vdd gnd cell_6t
Xbit_r94_c85 bl_85 br_85 wl_94 vdd gnd cell_6t
Xbit_r95_c85 bl_85 br_85 wl_95 vdd gnd cell_6t
Xbit_r96_c85 bl_85 br_85 wl_96 vdd gnd cell_6t
Xbit_r97_c85 bl_85 br_85 wl_97 vdd gnd cell_6t
Xbit_r98_c85 bl_85 br_85 wl_98 vdd gnd cell_6t
Xbit_r99_c85 bl_85 br_85 wl_99 vdd gnd cell_6t
Xbit_r100_c85 bl_85 br_85 wl_100 vdd gnd cell_6t
Xbit_r101_c85 bl_85 br_85 wl_101 vdd gnd cell_6t
Xbit_r102_c85 bl_85 br_85 wl_102 vdd gnd cell_6t
Xbit_r103_c85 bl_85 br_85 wl_103 vdd gnd cell_6t
Xbit_r104_c85 bl_85 br_85 wl_104 vdd gnd cell_6t
Xbit_r105_c85 bl_85 br_85 wl_105 vdd gnd cell_6t
Xbit_r106_c85 bl_85 br_85 wl_106 vdd gnd cell_6t
Xbit_r107_c85 bl_85 br_85 wl_107 vdd gnd cell_6t
Xbit_r108_c85 bl_85 br_85 wl_108 vdd gnd cell_6t
Xbit_r109_c85 bl_85 br_85 wl_109 vdd gnd cell_6t
Xbit_r110_c85 bl_85 br_85 wl_110 vdd gnd cell_6t
Xbit_r111_c85 bl_85 br_85 wl_111 vdd gnd cell_6t
Xbit_r112_c85 bl_85 br_85 wl_112 vdd gnd cell_6t
Xbit_r113_c85 bl_85 br_85 wl_113 vdd gnd cell_6t
Xbit_r114_c85 bl_85 br_85 wl_114 vdd gnd cell_6t
Xbit_r115_c85 bl_85 br_85 wl_115 vdd gnd cell_6t
Xbit_r116_c85 bl_85 br_85 wl_116 vdd gnd cell_6t
Xbit_r117_c85 bl_85 br_85 wl_117 vdd gnd cell_6t
Xbit_r118_c85 bl_85 br_85 wl_118 vdd gnd cell_6t
Xbit_r119_c85 bl_85 br_85 wl_119 vdd gnd cell_6t
Xbit_r120_c85 bl_85 br_85 wl_120 vdd gnd cell_6t
Xbit_r121_c85 bl_85 br_85 wl_121 vdd gnd cell_6t
Xbit_r122_c85 bl_85 br_85 wl_122 vdd gnd cell_6t
Xbit_r123_c85 bl_85 br_85 wl_123 vdd gnd cell_6t
Xbit_r124_c85 bl_85 br_85 wl_124 vdd gnd cell_6t
Xbit_r125_c85 bl_85 br_85 wl_125 vdd gnd cell_6t
Xbit_r126_c85 bl_85 br_85 wl_126 vdd gnd cell_6t
Xbit_r127_c85 bl_85 br_85 wl_127 vdd gnd cell_6t
Xbit_r128_c85 bl_85 br_85 wl_128 vdd gnd cell_6t
Xbit_r129_c85 bl_85 br_85 wl_129 vdd gnd cell_6t
Xbit_r130_c85 bl_85 br_85 wl_130 vdd gnd cell_6t
Xbit_r131_c85 bl_85 br_85 wl_131 vdd gnd cell_6t
Xbit_r132_c85 bl_85 br_85 wl_132 vdd gnd cell_6t
Xbit_r133_c85 bl_85 br_85 wl_133 vdd gnd cell_6t
Xbit_r134_c85 bl_85 br_85 wl_134 vdd gnd cell_6t
Xbit_r135_c85 bl_85 br_85 wl_135 vdd gnd cell_6t
Xbit_r136_c85 bl_85 br_85 wl_136 vdd gnd cell_6t
Xbit_r137_c85 bl_85 br_85 wl_137 vdd gnd cell_6t
Xbit_r138_c85 bl_85 br_85 wl_138 vdd gnd cell_6t
Xbit_r139_c85 bl_85 br_85 wl_139 vdd gnd cell_6t
Xbit_r140_c85 bl_85 br_85 wl_140 vdd gnd cell_6t
Xbit_r141_c85 bl_85 br_85 wl_141 vdd gnd cell_6t
Xbit_r142_c85 bl_85 br_85 wl_142 vdd gnd cell_6t
Xbit_r143_c85 bl_85 br_85 wl_143 vdd gnd cell_6t
Xbit_r144_c85 bl_85 br_85 wl_144 vdd gnd cell_6t
Xbit_r145_c85 bl_85 br_85 wl_145 vdd gnd cell_6t
Xbit_r146_c85 bl_85 br_85 wl_146 vdd gnd cell_6t
Xbit_r147_c85 bl_85 br_85 wl_147 vdd gnd cell_6t
Xbit_r148_c85 bl_85 br_85 wl_148 vdd gnd cell_6t
Xbit_r149_c85 bl_85 br_85 wl_149 vdd gnd cell_6t
Xbit_r150_c85 bl_85 br_85 wl_150 vdd gnd cell_6t
Xbit_r151_c85 bl_85 br_85 wl_151 vdd gnd cell_6t
Xbit_r152_c85 bl_85 br_85 wl_152 vdd gnd cell_6t
Xbit_r153_c85 bl_85 br_85 wl_153 vdd gnd cell_6t
Xbit_r154_c85 bl_85 br_85 wl_154 vdd gnd cell_6t
Xbit_r155_c85 bl_85 br_85 wl_155 vdd gnd cell_6t
Xbit_r156_c85 bl_85 br_85 wl_156 vdd gnd cell_6t
Xbit_r157_c85 bl_85 br_85 wl_157 vdd gnd cell_6t
Xbit_r158_c85 bl_85 br_85 wl_158 vdd gnd cell_6t
Xbit_r159_c85 bl_85 br_85 wl_159 vdd gnd cell_6t
Xbit_r160_c85 bl_85 br_85 wl_160 vdd gnd cell_6t
Xbit_r161_c85 bl_85 br_85 wl_161 vdd gnd cell_6t
Xbit_r162_c85 bl_85 br_85 wl_162 vdd gnd cell_6t
Xbit_r163_c85 bl_85 br_85 wl_163 vdd gnd cell_6t
Xbit_r164_c85 bl_85 br_85 wl_164 vdd gnd cell_6t
Xbit_r165_c85 bl_85 br_85 wl_165 vdd gnd cell_6t
Xbit_r166_c85 bl_85 br_85 wl_166 vdd gnd cell_6t
Xbit_r167_c85 bl_85 br_85 wl_167 vdd gnd cell_6t
Xbit_r168_c85 bl_85 br_85 wl_168 vdd gnd cell_6t
Xbit_r169_c85 bl_85 br_85 wl_169 vdd gnd cell_6t
Xbit_r170_c85 bl_85 br_85 wl_170 vdd gnd cell_6t
Xbit_r171_c85 bl_85 br_85 wl_171 vdd gnd cell_6t
Xbit_r172_c85 bl_85 br_85 wl_172 vdd gnd cell_6t
Xbit_r173_c85 bl_85 br_85 wl_173 vdd gnd cell_6t
Xbit_r174_c85 bl_85 br_85 wl_174 vdd gnd cell_6t
Xbit_r175_c85 bl_85 br_85 wl_175 vdd gnd cell_6t
Xbit_r176_c85 bl_85 br_85 wl_176 vdd gnd cell_6t
Xbit_r177_c85 bl_85 br_85 wl_177 vdd gnd cell_6t
Xbit_r178_c85 bl_85 br_85 wl_178 vdd gnd cell_6t
Xbit_r179_c85 bl_85 br_85 wl_179 vdd gnd cell_6t
Xbit_r180_c85 bl_85 br_85 wl_180 vdd gnd cell_6t
Xbit_r181_c85 bl_85 br_85 wl_181 vdd gnd cell_6t
Xbit_r182_c85 bl_85 br_85 wl_182 vdd gnd cell_6t
Xbit_r183_c85 bl_85 br_85 wl_183 vdd gnd cell_6t
Xbit_r184_c85 bl_85 br_85 wl_184 vdd gnd cell_6t
Xbit_r185_c85 bl_85 br_85 wl_185 vdd gnd cell_6t
Xbit_r186_c85 bl_85 br_85 wl_186 vdd gnd cell_6t
Xbit_r187_c85 bl_85 br_85 wl_187 vdd gnd cell_6t
Xbit_r188_c85 bl_85 br_85 wl_188 vdd gnd cell_6t
Xbit_r189_c85 bl_85 br_85 wl_189 vdd gnd cell_6t
Xbit_r190_c85 bl_85 br_85 wl_190 vdd gnd cell_6t
Xbit_r191_c85 bl_85 br_85 wl_191 vdd gnd cell_6t
Xbit_r192_c85 bl_85 br_85 wl_192 vdd gnd cell_6t
Xbit_r193_c85 bl_85 br_85 wl_193 vdd gnd cell_6t
Xbit_r194_c85 bl_85 br_85 wl_194 vdd gnd cell_6t
Xbit_r195_c85 bl_85 br_85 wl_195 vdd gnd cell_6t
Xbit_r196_c85 bl_85 br_85 wl_196 vdd gnd cell_6t
Xbit_r197_c85 bl_85 br_85 wl_197 vdd gnd cell_6t
Xbit_r198_c85 bl_85 br_85 wl_198 vdd gnd cell_6t
Xbit_r199_c85 bl_85 br_85 wl_199 vdd gnd cell_6t
Xbit_r200_c85 bl_85 br_85 wl_200 vdd gnd cell_6t
Xbit_r201_c85 bl_85 br_85 wl_201 vdd gnd cell_6t
Xbit_r202_c85 bl_85 br_85 wl_202 vdd gnd cell_6t
Xbit_r203_c85 bl_85 br_85 wl_203 vdd gnd cell_6t
Xbit_r204_c85 bl_85 br_85 wl_204 vdd gnd cell_6t
Xbit_r205_c85 bl_85 br_85 wl_205 vdd gnd cell_6t
Xbit_r206_c85 bl_85 br_85 wl_206 vdd gnd cell_6t
Xbit_r207_c85 bl_85 br_85 wl_207 vdd gnd cell_6t
Xbit_r208_c85 bl_85 br_85 wl_208 vdd gnd cell_6t
Xbit_r209_c85 bl_85 br_85 wl_209 vdd gnd cell_6t
Xbit_r210_c85 bl_85 br_85 wl_210 vdd gnd cell_6t
Xbit_r211_c85 bl_85 br_85 wl_211 vdd gnd cell_6t
Xbit_r212_c85 bl_85 br_85 wl_212 vdd gnd cell_6t
Xbit_r213_c85 bl_85 br_85 wl_213 vdd gnd cell_6t
Xbit_r214_c85 bl_85 br_85 wl_214 vdd gnd cell_6t
Xbit_r215_c85 bl_85 br_85 wl_215 vdd gnd cell_6t
Xbit_r216_c85 bl_85 br_85 wl_216 vdd gnd cell_6t
Xbit_r217_c85 bl_85 br_85 wl_217 vdd gnd cell_6t
Xbit_r218_c85 bl_85 br_85 wl_218 vdd gnd cell_6t
Xbit_r219_c85 bl_85 br_85 wl_219 vdd gnd cell_6t
Xbit_r220_c85 bl_85 br_85 wl_220 vdd gnd cell_6t
Xbit_r221_c85 bl_85 br_85 wl_221 vdd gnd cell_6t
Xbit_r222_c85 bl_85 br_85 wl_222 vdd gnd cell_6t
Xbit_r223_c85 bl_85 br_85 wl_223 vdd gnd cell_6t
Xbit_r224_c85 bl_85 br_85 wl_224 vdd gnd cell_6t
Xbit_r225_c85 bl_85 br_85 wl_225 vdd gnd cell_6t
Xbit_r226_c85 bl_85 br_85 wl_226 vdd gnd cell_6t
Xbit_r227_c85 bl_85 br_85 wl_227 vdd gnd cell_6t
Xbit_r228_c85 bl_85 br_85 wl_228 vdd gnd cell_6t
Xbit_r229_c85 bl_85 br_85 wl_229 vdd gnd cell_6t
Xbit_r230_c85 bl_85 br_85 wl_230 vdd gnd cell_6t
Xbit_r231_c85 bl_85 br_85 wl_231 vdd gnd cell_6t
Xbit_r232_c85 bl_85 br_85 wl_232 vdd gnd cell_6t
Xbit_r233_c85 bl_85 br_85 wl_233 vdd gnd cell_6t
Xbit_r234_c85 bl_85 br_85 wl_234 vdd gnd cell_6t
Xbit_r235_c85 bl_85 br_85 wl_235 vdd gnd cell_6t
Xbit_r236_c85 bl_85 br_85 wl_236 vdd gnd cell_6t
Xbit_r237_c85 bl_85 br_85 wl_237 vdd gnd cell_6t
Xbit_r238_c85 bl_85 br_85 wl_238 vdd gnd cell_6t
Xbit_r239_c85 bl_85 br_85 wl_239 vdd gnd cell_6t
Xbit_r240_c85 bl_85 br_85 wl_240 vdd gnd cell_6t
Xbit_r241_c85 bl_85 br_85 wl_241 vdd gnd cell_6t
Xbit_r242_c85 bl_85 br_85 wl_242 vdd gnd cell_6t
Xbit_r243_c85 bl_85 br_85 wl_243 vdd gnd cell_6t
Xbit_r244_c85 bl_85 br_85 wl_244 vdd gnd cell_6t
Xbit_r245_c85 bl_85 br_85 wl_245 vdd gnd cell_6t
Xbit_r246_c85 bl_85 br_85 wl_246 vdd gnd cell_6t
Xbit_r247_c85 bl_85 br_85 wl_247 vdd gnd cell_6t
Xbit_r248_c85 bl_85 br_85 wl_248 vdd gnd cell_6t
Xbit_r249_c85 bl_85 br_85 wl_249 vdd gnd cell_6t
Xbit_r250_c85 bl_85 br_85 wl_250 vdd gnd cell_6t
Xbit_r251_c85 bl_85 br_85 wl_251 vdd gnd cell_6t
Xbit_r252_c85 bl_85 br_85 wl_252 vdd gnd cell_6t
Xbit_r253_c85 bl_85 br_85 wl_253 vdd gnd cell_6t
Xbit_r254_c85 bl_85 br_85 wl_254 vdd gnd cell_6t
Xbit_r255_c85 bl_85 br_85 wl_255 vdd gnd cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd cell_6t
Xbit_r1_c86 bl_86 br_86 wl_1 vdd gnd cell_6t
Xbit_r2_c86 bl_86 br_86 wl_2 vdd gnd cell_6t
Xbit_r3_c86 bl_86 br_86 wl_3 vdd gnd cell_6t
Xbit_r4_c86 bl_86 br_86 wl_4 vdd gnd cell_6t
Xbit_r5_c86 bl_86 br_86 wl_5 vdd gnd cell_6t
Xbit_r6_c86 bl_86 br_86 wl_6 vdd gnd cell_6t
Xbit_r7_c86 bl_86 br_86 wl_7 vdd gnd cell_6t
Xbit_r8_c86 bl_86 br_86 wl_8 vdd gnd cell_6t
Xbit_r9_c86 bl_86 br_86 wl_9 vdd gnd cell_6t
Xbit_r10_c86 bl_86 br_86 wl_10 vdd gnd cell_6t
Xbit_r11_c86 bl_86 br_86 wl_11 vdd gnd cell_6t
Xbit_r12_c86 bl_86 br_86 wl_12 vdd gnd cell_6t
Xbit_r13_c86 bl_86 br_86 wl_13 vdd gnd cell_6t
Xbit_r14_c86 bl_86 br_86 wl_14 vdd gnd cell_6t
Xbit_r15_c86 bl_86 br_86 wl_15 vdd gnd cell_6t
Xbit_r16_c86 bl_86 br_86 wl_16 vdd gnd cell_6t
Xbit_r17_c86 bl_86 br_86 wl_17 vdd gnd cell_6t
Xbit_r18_c86 bl_86 br_86 wl_18 vdd gnd cell_6t
Xbit_r19_c86 bl_86 br_86 wl_19 vdd gnd cell_6t
Xbit_r20_c86 bl_86 br_86 wl_20 vdd gnd cell_6t
Xbit_r21_c86 bl_86 br_86 wl_21 vdd gnd cell_6t
Xbit_r22_c86 bl_86 br_86 wl_22 vdd gnd cell_6t
Xbit_r23_c86 bl_86 br_86 wl_23 vdd gnd cell_6t
Xbit_r24_c86 bl_86 br_86 wl_24 vdd gnd cell_6t
Xbit_r25_c86 bl_86 br_86 wl_25 vdd gnd cell_6t
Xbit_r26_c86 bl_86 br_86 wl_26 vdd gnd cell_6t
Xbit_r27_c86 bl_86 br_86 wl_27 vdd gnd cell_6t
Xbit_r28_c86 bl_86 br_86 wl_28 vdd gnd cell_6t
Xbit_r29_c86 bl_86 br_86 wl_29 vdd gnd cell_6t
Xbit_r30_c86 bl_86 br_86 wl_30 vdd gnd cell_6t
Xbit_r31_c86 bl_86 br_86 wl_31 vdd gnd cell_6t
Xbit_r32_c86 bl_86 br_86 wl_32 vdd gnd cell_6t
Xbit_r33_c86 bl_86 br_86 wl_33 vdd gnd cell_6t
Xbit_r34_c86 bl_86 br_86 wl_34 vdd gnd cell_6t
Xbit_r35_c86 bl_86 br_86 wl_35 vdd gnd cell_6t
Xbit_r36_c86 bl_86 br_86 wl_36 vdd gnd cell_6t
Xbit_r37_c86 bl_86 br_86 wl_37 vdd gnd cell_6t
Xbit_r38_c86 bl_86 br_86 wl_38 vdd gnd cell_6t
Xbit_r39_c86 bl_86 br_86 wl_39 vdd gnd cell_6t
Xbit_r40_c86 bl_86 br_86 wl_40 vdd gnd cell_6t
Xbit_r41_c86 bl_86 br_86 wl_41 vdd gnd cell_6t
Xbit_r42_c86 bl_86 br_86 wl_42 vdd gnd cell_6t
Xbit_r43_c86 bl_86 br_86 wl_43 vdd gnd cell_6t
Xbit_r44_c86 bl_86 br_86 wl_44 vdd gnd cell_6t
Xbit_r45_c86 bl_86 br_86 wl_45 vdd gnd cell_6t
Xbit_r46_c86 bl_86 br_86 wl_46 vdd gnd cell_6t
Xbit_r47_c86 bl_86 br_86 wl_47 vdd gnd cell_6t
Xbit_r48_c86 bl_86 br_86 wl_48 vdd gnd cell_6t
Xbit_r49_c86 bl_86 br_86 wl_49 vdd gnd cell_6t
Xbit_r50_c86 bl_86 br_86 wl_50 vdd gnd cell_6t
Xbit_r51_c86 bl_86 br_86 wl_51 vdd gnd cell_6t
Xbit_r52_c86 bl_86 br_86 wl_52 vdd gnd cell_6t
Xbit_r53_c86 bl_86 br_86 wl_53 vdd gnd cell_6t
Xbit_r54_c86 bl_86 br_86 wl_54 vdd gnd cell_6t
Xbit_r55_c86 bl_86 br_86 wl_55 vdd gnd cell_6t
Xbit_r56_c86 bl_86 br_86 wl_56 vdd gnd cell_6t
Xbit_r57_c86 bl_86 br_86 wl_57 vdd gnd cell_6t
Xbit_r58_c86 bl_86 br_86 wl_58 vdd gnd cell_6t
Xbit_r59_c86 bl_86 br_86 wl_59 vdd gnd cell_6t
Xbit_r60_c86 bl_86 br_86 wl_60 vdd gnd cell_6t
Xbit_r61_c86 bl_86 br_86 wl_61 vdd gnd cell_6t
Xbit_r62_c86 bl_86 br_86 wl_62 vdd gnd cell_6t
Xbit_r63_c86 bl_86 br_86 wl_63 vdd gnd cell_6t
Xbit_r64_c86 bl_86 br_86 wl_64 vdd gnd cell_6t
Xbit_r65_c86 bl_86 br_86 wl_65 vdd gnd cell_6t
Xbit_r66_c86 bl_86 br_86 wl_66 vdd gnd cell_6t
Xbit_r67_c86 bl_86 br_86 wl_67 vdd gnd cell_6t
Xbit_r68_c86 bl_86 br_86 wl_68 vdd gnd cell_6t
Xbit_r69_c86 bl_86 br_86 wl_69 vdd gnd cell_6t
Xbit_r70_c86 bl_86 br_86 wl_70 vdd gnd cell_6t
Xbit_r71_c86 bl_86 br_86 wl_71 vdd gnd cell_6t
Xbit_r72_c86 bl_86 br_86 wl_72 vdd gnd cell_6t
Xbit_r73_c86 bl_86 br_86 wl_73 vdd gnd cell_6t
Xbit_r74_c86 bl_86 br_86 wl_74 vdd gnd cell_6t
Xbit_r75_c86 bl_86 br_86 wl_75 vdd gnd cell_6t
Xbit_r76_c86 bl_86 br_86 wl_76 vdd gnd cell_6t
Xbit_r77_c86 bl_86 br_86 wl_77 vdd gnd cell_6t
Xbit_r78_c86 bl_86 br_86 wl_78 vdd gnd cell_6t
Xbit_r79_c86 bl_86 br_86 wl_79 vdd gnd cell_6t
Xbit_r80_c86 bl_86 br_86 wl_80 vdd gnd cell_6t
Xbit_r81_c86 bl_86 br_86 wl_81 vdd gnd cell_6t
Xbit_r82_c86 bl_86 br_86 wl_82 vdd gnd cell_6t
Xbit_r83_c86 bl_86 br_86 wl_83 vdd gnd cell_6t
Xbit_r84_c86 bl_86 br_86 wl_84 vdd gnd cell_6t
Xbit_r85_c86 bl_86 br_86 wl_85 vdd gnd cell_6t
Xbit_r86_c86 bl_86 br_86 wl_86 vdd gnd cell_6t
Xbit_r87_c86 bl_86 br_86 wl_87 vdd gnd cell_6t
Xbit_r88_c86 bl_86 br_86 wl_88 vdd gnd cell_6t
Xbit_r89_c86 bl_86 br_86 wl_89 vdd gnd cell_6t
Xbit_r90_c86 bl_86 br_86 wl_90 vdd gnd cell_6t
Xbit_r91_c86 bl_86 br_86 wl_91 vdd gnd cell_6t
Xbit_r92_c86 bl_86 br_86 wl_92 vdd gnd cell_6t
Xbit_r93_c86 bl_86 br_86 wl_93 vdd gnd cell_6t
Xbit_r94_c86 bl_86 br_86 wl_94 vdd gnd cell_6t
Xbit_r95_c86 bl_86 br_86 wl_95 vdd gnd cell_6t
Xbit_r96_c86 bl_86 br_86 wl_96 vdd gnd cell_6t
Xbit_r97_c86 bl_86 br_86 wl_97 vdd gnd cell_6t
Xbit_r98_c86 bl_86 br_86 wl_98 vdd gnd cell_6t
Xbit_r99_c86 bl_86 br_86 wl_99 vdd gnd cell_6t
Xbit_r100_c86 bl_86 br_86 wl_100 vdd gnd cell_6t
Xbit_r101_c86 bl_86 br_86 wl_101 vdd gnd cell_6t
Xbit_r102_c86 bl_86 br_86 wl_102 vdd gnd cell_6t
Xbit_r103_c86 bl_86 br_86 wl_103 vdd gnd cell_6t
Xbit_r104_c86 bl_86 br_86 wl_104 vdd gnd cell_6t
Xbit_r105_c86 bl_86 br_86 wl_105 vdd gnd cell_6t
Xbit_r106_c86 bl_86 br_86 wl_106 vdd gnd cell_6t
Xbit_r107_c86 bl_86 br_86 wl_107 vdd gnd cell_6t
Xbit_r108_c86 bl_86 br_86 wl_108 vdd gnd cell_6t
Xbit_r109_c86 bl_86 br_86 wl_109 vdd gnd cell_6t
Xbit_r110_c86 bl_86 br_86 wl_110 vdd gnd cell_6t
Xbit_r111_c86 bl_86 br_86 wl_111 vdd gnd cell_6t
Xbit_r112_c86 bl_86 br_86 wl_112 vdd gnd cell_6t
Xbit_r113_c86 bl_86 br_86 wl_113 vdd gnd cell_6t
Xbit_r114_c86 bl_86 br_86 wl_114 vdd gnd cell_6t
Xbit_r115_c86 bl_86 br_86 wl_115 vdd gnd cell_6t
Xbit_r116_c86 bl_86 br_86 wl_116 vdd gnd cell_6t
Xbit_r117_c86 bl_86 br_86 wl_117 vdd gnd cell_6t
Xbit_r118_c86 bl_86 br_86 wl_118 vdd gnd cell_6t
Xbit_r119_c86 bl_86 br_86 wl_119 vdd gnd cell_6t
Xbit_r120_c86 bl_86 br_86 wl_120 vdd gnd cell_6t
Xbit_r121_c86 bl_86 br_86 wl_121 vdd gnd cell_6t
Xbit_r122_c86 bl_86 br_86 wl_122 vdd gnd cell_6t
Xbit_r123_c86 bl_86 br_86 wl_123 vdd gnd cell_6t
Xbit_r124_c86 bl_86 br_86 wl_124 vdd gnd cell_6t
Xbit_r125_c86 bl_86 br_86 wl_125 vdd gnd cell_6t
Xbit_r126_c86 bl_86 br_86 wl_126 vdd gnd cell_6t
Xbit_r127_c86 bl_86 br_86 wl_127 vdd gnd cell_6t
Xbit_r128_c86 bl_86 br_86 wl_128 vdd gnd cell_6t
Xbit_r129_c86 bl_86 br_86 wl_129 vdd gnd cell_6t
Xbit_r130_c86 bl_86 br_86 wl_130 vdd gnd cell_6t
Xbit_r131_c86 bl_86 br_86 wl_131 vdd gnd cell_6t
Xbit_r132_c86 bl_86 br_86 wl_132 vdd gnd cell_6t
Xbit_r133_c86 bl_86 br_86 wl_133 vdd gnd cell_6t
Xbit_r134_c86 bl_86 br_86 wl_134 vdd gnd cell_6t
Xbit_r135_c86 bl_86 br_86 wl_135 vdd gnd cell_6t
Xbit_r136_c86 bl_86 br_86 wl_136 vdd gnd cell_6t
Xbit_r137_c86 bl_86 br_86 wl_137 vdd gnd cell_6t
Xbit_r138_c86 bl_86 br_86 wl_138 vdd gnd cell_6t
Xbit_r139_c86 bl_86 br_86 wl_139 vdd gnd cell_6t
Xbit_r140_c86 bl_86 br_86 wl_140 vdd gnd cell_6t
Xbit_r141_c86 bl_86 br_86 wl_141 vdd gnd cell_6t
Xbit_r142_c86 bl_86 br_86 wl_142 vdd gnd cell_6t
Xbit_r143_c86 bl_86 br_86 wl_143 vdd gnd cell_6t
Xbit_r144_c86 bl_86 br_86 wl_144 vdd gnd cell_6t
Xbit_r145_c86 bl_86 br_86 wl_145 vdd gnd cell_6t
Xbit_r146_c86 bl_86 br_86 wl_146 vdd gnd cell_6t
Xbit_r147_c86 bl_86 br_86 wl_147 vdd gnd cell_6t
Xbit_r148_c86 bl_86 br_86 wl_148 vdd gnd cell_6t
Xbit_r149_c86 bl_86 br_86 wl_149 vdd gnd cell_6t
Xbit_r150_c86 bl_86 br_86 wl_150 vdd gnd cell_6t
Xbit_r151_c86 bl_86 br_86 wl_151 vdd gnd cell_6t
Xbit_r152_c86 bl_86 br_86 wl_152 vdd gnd cell_6t
Xbit_r153_c86 bl_86 br_86 wl_153 vdd gnd cell_6t
Xbit_r154_c86 bl_86 br_86 wl_154 vdd gnd cell_6t
Xbit_r155_c86 bl_86 br_86 wl_155 vdd gnd cell_6t
Xbit_r156_c86 bl_86 br_86 wl_156 vdd gnd cell_6t
Xbit_r157_c86 bl_86 br_86 wl_157 vdd gnd cell_6t
Xbit_r158_c86 bl_86 br_86 wl_158 vdd gnd cell_6t
Xbit_r159_c86 bl_86 br_86 wl_159 vdd gnd cell_6t
Xbit_r160_c86 bl_86 br_86 wl_160 vdd gnd cell_6t
Xbit_r161_c86 bl_86 br_86 wl_161 vdd gnd cell_6t
Xbit_r162_c86 bl_86 br_86 wl_162 vdd gnd cell_6t
Xbit_r163_c86 bl_86 br_86 wl_163 vdd gnd cell_6t
Xbit_r164_c86 bl_86 br_86 wl_164 vdd gnd cell_6t
Xbit_r165_c86 bl_86 br_86 wl_165 vdd gnd cell_6t
Xbit_r166_c86 bl_86 br_86 wl_166 vdd gnd cell_6t
Xbit_r167_c86 bl_86 br_86 wl_167 vdd gnd cell_6t
Xbit_r168_c86 bl_86 br_86 wl_168 vdd gnd cell_6t
Xbit_r169_c86 bl_86 br_86 wl_169 vdd gnd cell_6t
Xbit_r170_c86 bl_86 br_86 wl_170 vdd gnd cell_6t
Xbit_r171_c86 bl_86 br_86 wl_171 vdd gnd cell_6t
Xbit_r172_c86 bl_86 br_86 wl_172 vdd gnd cell_6t
Xbit_r173_c86 bl_86 br_86 wl_173 vdd gnd cell_6t
Xbit_r174_c86 bl_86 br_86 wl_174 vdd gnd cell_6t
Xbit_r175_c86 bl_86 br_86 wl_175 vdd gnd cell_6t
Xbit_r176_c86 bl_86 br_86 wl_176 vdd gnd cell_6t
Xbit_r177_c86 bl_86 br_86 wl_177 vdd gnd cell_6t
Xbit_r178_c86 bl_86 br_86 wl_178 vdd gnd cell_6t
Xbit_r179_c86 bl_86 br_86 wl_179 vdd gnd cell_6t
Xbit_r180_c86 bl_86 br_86 wl_180 vdd gnd cell_6t
Xbit_r181_c86 bl_86 br_86 wl_181 vdd gnd cell_6t
Xbit_r182_c86 bl_86 br_86 wl_182 vdd gnd cell_6t
Xbit_r183_c86 bl_86 br_86 wl_183 vdd gnd cell_6t
Xbit_r184_c86 bl_86 br_86 wl_184 vdd gnd cell_6t
Xbit_r185_c86 bl_86 br_86 wl_185 vdd gnd cell_6t
Xbit_r186_c86 bl_86 br_86 wl_186 vdd gnd cell_6t
Xbit_r187_c86 bl_86 br_86 wl_187 vdd gnd cell_6t
Xbit_r188_c86 bl_86 br_86 wl_188 vdd gnd cell_6t
Xbit_r189_c86 bl_86 br_86 wl_189 vdd gnd cell_6t
Xbit_r190_c86 bl_86 br_86 wl_190 vdd gnd cell_6t
Xbit_r191_c86 bl_86 br_86 wl_191 vdd gnd cell_6t
Xbit_r192_c86 bl_86 br_86 wl_192 vdd gnd cell_6t
Xbit_r193_c86 bl_86 br_86 wl_193 vdd gnd cell_6t
Xbit_r194_c86 bl_86 br_86 wl_194 vdd gnd cell_6t
Xbit_r195_c86 bl_86 br_86 wl_195 vdd gnd cell_6t
Xbit_r196_c86 bl_86 br_86 wl_196 vdd gnd cell_6t
Xbit_r197_c86 bl_86 br_86 wl_197 vdd gnd cell_6t
Xbit_r198_c86 bl_86 br_86 wl_198 vdd gnd cell_6t
Xbit_r199_c86 bl_86 br_86 wl_199 vdd gnd cell_6t
Xbit_r200_c86 bl_86 br_86 wl_200 vdd gnd cell_6t
Xbit_r201_c86 bl_86 br_86 wl_201 vdd gnd cell_6t
Xbit_r202_c86 bl_86 br_86 wl_202 vdd gnd cell_6t
Xbit_r203_c86 bl_86 br_86 wl_203 vdd gnd cell_6t
Xbit_r204_c86 bl_86 br_86 wl_204 vdd gnd cell_6t
Xbit_r205_c86 bl_86 br_86 wl_205 vdd gnd cell_6t
Xbit_r206_c86 bl_86 br_86 wl_206 vdd gnd cell_6t
Xbit_r207_c86 bl_86 br_86 wl_207 vdd gnd cell_6t
Xbit_r208_c86 bl_86 br_86 wl_208 vdd gnd cell_6t
Xbit_r209_c86 bl_86 br_86 wl_209 vdd gnd cell_6t
Xbit_r210_c86 bl_86 br_86 wl_210 vdd gnd cell_6t
Xbit_r211_c86 bl_86 br_86 wl_211 vdd gnd cell_6t
Xbit_r212_c86 bl_86 br_86 wl_212 vdd gnd cell_6t
Xbit_r213_c86 bl_86 br_86 wl_213 vdd gnd cell_6t
Xbit_r214_c86 bl_86 br_86 wl_214 vdd gnd cell_6t
Xbit_r215_c86 bl_86 br_86 wl_215 vdd gnd cell_6t
Xbit_r216_c86 bl_86 br_86 wl_216 vdd gnd cell_6t
Xbit_r217_c86 bl_86 br_86 wl_217 vdd gnd cell_6t
Xbit_r218_c86 bl_86 br_86 wl_218 vdd gnd cell_6t
Xbit_r219_c86 bl_86 br_86 wl_219 vdd gnd cell_6t
Xbit_r220_c86 bl_86 br_86 wl_220 vdd gnd cell_6t
Xbit_r221_c86 bl_86 br_86 wl_221 vdd gnd cell_6t
Xbit_r222_c86 bl_86 br_86 wl_222 vdd gnd cell_6t
Xbit_r223_c86 bl_86 br_86 wl_223 vdd gnd cell_6t
Xbit_r224_c86 bl_86 br_86 wl_224 vdd gnd cell_6t
Xbit_r225_c86 bl_86 br_86 wl_225 vdd gnd cell_6t
Xbit_r226_c86 bl_86 br_86 wl_226 vdd gnd cell_6t
Xbit_r227_c86 bl_86 br_86 wl_227 vdd gnd cell_6t
Xbit_r228_c86 bl_86 br_86 wl_228 vdd gnd cell_6t
Xbit_r229_c86 bl_86 br_86 wl_229 vdd gnd cell_6t
Xbit_r230_c86 bl_86 br_86 wl_230 vdd gnd cell_6t
Xbit_r231_c86 bl_86 br_86 wl_231 vdd gnd cell_6t
Xbit_r232_c86 bl_86 br_86 wl_232 vdd gnd cell_6t
Xbit_r233_c86 bl_86 br_86 wl_233 vdd gnd cell_6t
Xbit_r234_c86 bl_86 br_86 wl_234 vdd gnd cell_6t
Xbit_r235_c86 bl_86 br_86 wl_235 vdd gnd cell_6t
Xbit_r236_c86 bl_86 br_86 wl_236 vdd gnd cell_6t
Xbit_r237_c86 bl_86 br_86 wl_237 vdd gnd cell_6t
Xbit_r238_c86 bl_86 br_86 wl_238 vdd gnd cell_6t
Xbit_r239_c86 bl_86 br_86 wl_239 vdd gnd cell_6t
Xbit_r240_c86 bl_86 br_86 wl_240 vdd gnd cell_6t
Xbit_r241_c86 bl_86 br_86 wl_241 vdd gnd cell_6t
Xbit_r242_c86 bl_86 br_86 wl_242 vdd gnd cell_6t
Xbit_r243_c86 bl_86 br_86 wl_243 vdd gnd cell_6t
Xbit_r244_c86 bl_86 br_86 wl_244 vdd gnd cell_6t
Xbit_r245_c86 bl_86 br_86 wl_245 vdd gnd cell_6t
Xbit_r246_c86 bl_86 br_86 wl_246 vdd gnd cell_6t
Xbit_r247_c86 bl_86 br_86 wl_247 vdd gnd cell_6t
Xbit_r248_c86 bl_86 br_86 wl_248 vdd gnd cell_6t
Xbit_r249_c86 bl_86 br_86 wl_249 vdd gnd cell_6t
Xbit_r250_c86 bl_86 br_86 wl_250 vdd gnd cell_6t
Xbit_r251_c86 bl_86 br_86 wl_251 vdd gnd cell_6t
Xbit_r252_c86 bl_86 br_86 wl_252 vdd gnd cell_6t
Xbit_r253_c86 bl_86 br_86 wl_253 vdd gnd cell_6t
Xbit_r254_c86 bl_86 br_86 wl_254 vdd gnd cell_6t
Xbit_r255_c86 bl_86 br_86 wl_255 vdd gnd cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd cell_6t
Xbit_r1_c87 bl_87 br_87 wl_1 vdd gnd cell_6t
Xbit_r2_c87 bl_87 br_87 wl_2 vdd gnd cell_6t
Xbit_r3_c87 bl_87 br_87 wl_3 vdd gnd cell_6t
Xbit_r4_c87 bl_87 br_87 wl_4 vdd gnd cell_6t
Xbit_r5_c87 bl_87 br_87 wl_5 vdd gnd cell_6t
Xbit_r6_c87 bl_87 br_87 wl_6 vdd gnd cell_6t
Xbit_r7_c87 bl_87 br_87 wl_7 vdd gnd cell_6t
Xbit_r8_c87 bl_87 br_87 wl_8 vdd gnd cell_6t
Xbit_r9_c87 bl_87 br_87 wl_9 vdd gnd cell_6t
Xbit_r10_c87 bl_87 br_87 wl_10 vdd gnd cell_6t
Xbit_r11_c87 bl_87 br_87 wl_11 vdd gnd cell_6t
Xbit_r12_c87 bl_87 br_87 wl_12 vdd gnd cell_6t
Xbit_r13_c87 bl_87 br_87 wl_13 vdd gnd cell_6t
Xbit_r14_c87 bl_87 br_87 wl_14 vdd gnd cell_6t
Xbit_r15_c87 bl_87 br_87 wl_15 vdd gnd cell_6t
Xbit_r16_c87 bl_87 br_87 wl_16 vdd gnd cell_6t
Xbit_r17_c87 bl_87 br_87 wl_17 vdd gnd cell_6t
Xbit_r18_c87 bl_87 br_87 wl_18 vdd gnd cell_6t
Xbit_r19_c87 bl_87 br_87 wl_19 vdd gnd cell_6t
Xbit_r20_c87 bl_87 br_87 wl_20 vdd gnd cell_6t
Xbit_r21_c87 bl_87 br_87 wl_21 vdd gnd cell_6t
Xbit_r22_c87 bl_87 br_87 wl_22 vdd gnd cell_6t
Xbit_r23_c87 bl_87 br_87 wl_23 vdd gnd cell_6t
Xbit_r24_c87 bl_87 br_87 wl_24 vdd gnd cell_6t
Xbit_r25_c87 bl_87 br_87 wl_25 vdd gnd cell_6t
Xbit_r26_c87 bl_87 br_87 wl_26 vdd gnd cell_6t
Xbit_r27_c87 bl_87 br_87 wl_27 vdd gnd cell_6t
Xbit_r28_c87 bl_87 br_87 wl_28 vdd gnd cell_6t
Xbit_r29_c87 bl_87 br_87 wl_29 vdd gnd cell_6t
Xbit_r30_c87 bl_87 br_87 wl_30 vdd gnd cell_6t
Xbit_r31_c87 bl_87 br_87 wl_31 vdd gnd cell_6t
Xbit_r32_c87 bl_87 br_87 wl_32 vdd gnd cell_6t
Xbit_r33_c87 bl_87 br_87 wl_33 vdd gnd cell_6t
Xbit_r34_c87 bl_87 br_87 wl_34 vdd gnd cell_6t
Xbit_r35_c87 bl_87 br_87 wl_35 vdd gnd cell_6t
Xbit_r36_c87 bl_87 br_87 wl_36 vdd gnd cell_6t
Xbit_r37_c87 bl_87 br_87 wl_37 vdd gnd cell_6t
Xbit_r38_c87 bl_87 br_87 wl_38 vdd gnd cell_6t
Xbit_r39_c87 bl_87 br_87 wl_39 vdd gnd cell_6t
Xbit_r40_c87 bl_87 br_87 wl_40 vdd gnd cell_6t
Xbit_r41_c87 bl_87 br_87 wl_41 vdd gnd cell_6t
Xbit_r42_c87 bl_87 br_87 wl_42 vdd gnd cell_6t
Xbit_r43_c87 bl_87 br_87 wl_43 vdd gnd cell_6t
Xbit_r44_c87 bl_87 br_87 wl_44 vdd gnd cell_6t
Xbit_r45_c87 bl_87 br_87 wl_45 vdd gnd cell_6t
Xbit_r46_c87 bl_87 br_87 wl_46 vdd gnd cell_6t
Xbit_r47_c87 bl_87 br_87 wl_47 vdd gnd cell_6t
Xbit_r48_c87 bl_87 br_87 wl_48 vdd gnd cell_6t
Xbit_r49_c87 bl_87 br_87 wl_49 vdd gnd cell_6t
Xbit_r50_c87 bl_87 br_87 wl_50 vdd gnd cell_6t
Xbit_r51_c87 bl_87 br_87 wl_51 vdd gnd cell_6t
Xbit_r52_c87 bl_87 br_87 wl_52 vdd gnd cell_6t
Xbit_r53_c87 bl_87 br_87 wl_53 vdd gnd cell_6t
Xbit_r54_c87 bl_87 br_87 wl_54 vdd gnd cell_6t
Xbit_r55_c87 bl_87 br_87 wl_55 vdd gnd cell_6t
Xbit_r56_c87 bl_87 br_87 wl_56 vdd gnd cell_6t
Xbit_r57_c87 bl_87 br_87 wl_57 vdd gnd cell_6t
Xbit_r58_c87 bl_87 br_87 wl_58 vdd gnd cell_6t
Xbit_r59_c87 bl_87 br_87 wl_59 vdd gnd cell_6t
Xbit_r60_c87 bl_87 br_87 wl_60 vdd gnd cell_6t
Xbit_r61_c87 bl_87 br_87 wl_61 vdd gnd cell_6t
Xbit_r62_c87 bl_87 br_87 wl_62 vdd gnd cell_6t
Xbit_r63_c87 bl_87 br_87 wl_63 vdd gnd cell_6t
Xbit_r64_c87 bl_87 br_87 wl_64 vdd gnd cell_6t
Xbit_r65_c87 bl_87 br_87 wl_65 vdd gnd cell_6t
Xbit_r66_c87 bl_87 br_87 wl_66 vdd gnd cell_6t
Xbit_r67_c87 bl_87 br_87 wl_67 vdd gnd cell_6t
Xbit_r68_c87 bl_87 br_87 wl_68 vdd gnd cell_6t
Xbit_r69_c87 bl_87 br_87 wl_69 vdd gnd cell_6t
Xbit_r70_c87 bl_87 br_87 wl_70 vdd gnd cell_6t
Xbit_r71_c87 bl_87 br_87 wl_71 vdd gnd cell_6t
Xbit_r72_c87 bl_87 br_87 wl_72 vdd gnd cell_6t
Xbit_r73_c87 bl_87 br_87 wl_73 vdd gnd cell_6t
Xbit_r74_c87 bl_87 br_87 wl_74 vdd gnd cell_6t
Xbit_r75_c87 bl_87 br_87 wl_75 vdd gnd cell_6t
Xbit_r76_c87 bl_87 br_87 wl_76 vdd gnd cell_6t
Xbit_r77_c87 bl_87 br_87 wl_77 vdd gnd cell_6t
Xbit_r78_c87 bl_87 br_87 wl_78 vdd gnd cell_6t
Xbit_r79_c87 bl_87 br_87 wl_79 vdd gnd cell_6t
Xbit_r80_c87 bl_87 br_87 wl_80 vdd gnd cell_6t
Xbit_r81_c87 bl_87 br_87 wl_81 vdd gnd cell_6t
Xbit_r82_c87 bl_87 br_87 wl_82 vdd gnd cell_6t
Xbit_r83_c87 bl_87 br_87 wl_83 vdd gnd cell_6t
Xbit_r84_c87 bl_87 br_87 wl_84 vdd gnd cell_6t
Xbit_r85_c87 bl_87 br_87 wl_85 vdd gnd cell_6t
Xbit_r86_c87 bl_87 br_87 wl_86 vdd gnd cell_6t
Xbit_r87_c87 bl_87 br_87 wl_87 vdd gnd cell_6t
Xbit_r88_c87 bl_87 br_87 wl_88 vdd gnd cell_6t
Xbit_r89_c87 bl_87 br_87 wl_89 vdd gnd cell_6t
Xbit_r90_c87 bl_87 br_87 wl_90 vdd gnd cell_6t
Xbit_r91_c87 bl_87 br_87 wl_91 vdd gnd cell_6t
Xbit_r92_c87 bl_87 br_87 wl_92 vdd gnd cell_6t
Xbit_r93_c87 bl_87 br_87 wl_93 vdd gnd cell_6t
Xbit_r94_c87 bl_87 br_87 wl_94 vdd gnd cell_6t
Xbit_r95_c87 bl_87 br_87 wl_95 vdd gnd cell_6t
Xbit_r96_c87 bl_87 br_87 wl_96 vdd gnd cell_6t
Xbit_r97_c87 bl_87 br_87 wl_97 vdd gnd cell_6t
Xbit_r98_c87 bl_87 br_87 wl_98 vdd gnd cell_6t
Xbit_r99_c87 bl_87 br_87 wl_99 vdd gnd cell_6t
Xbit_r100_c87 bl_87 br_87 wl_100 vdd gnd cell_6t
Xbit_r101_c87 bl_87 br_87 wl_101 vdd gnd cell_6t
Xbit_r102_c87 bl_87 br_87 wl_102 vdd gnd cell_6t
Xbit_r103_c87 bl_87 br_87 wl_103 vdd gnd cell_6t
Xbit_r104_c87 bl_87 br_87 wl_104 vdd gnd cell_6t
Xbit_r105_c87 bl_87 br_87 wl_105 vdd gnd cell_6t
Xbit_r106_c87 bl_87 br_87 wl_106 vdd gnd cell_6t
Xbit_r107_c87 bl_87 br_87 wl_107 vdd gnd cell_6t
Xbit_r108_c87 bl_87 br_87 wl_108 vdd gnd cell_6t
Xbit_r109_c87 bl_87 br_87 wl_109 vdd gnd cell_6t
Xbit_r110_c87 bl_87 br_87 wl_110 vdd gnd cell_6t
Xbit_r111_c87 bl_87 br_87 wl_111 vdd gnd cell_6t
Xbit_r112_c87 bl_87 br_87 wl_112 vdd gnd cell_6t
Xbit_r113_c87 bl_87 br_87 wl_113 vdd gnd cell_6t
Xbit_r114_c87 bl_87 br_87 wl_114 vdd gnd cell_6t
Xbit_r115_c87 bl_87 br_87 wl_115 vdd gnd cell_6t
Xbit_r116_c87 bl_87 br_87 wl_116 vdd gnd cell_6t
Xbit_r117_c87 bl_87 br_87 wl_117 vdd gnd cell_6t
Xbit_r118_c87 bl_87 br_87 wl_118 vdd gnd cell_6t
Xbit_r119_c87 bl_87 br_87 wl_119 vdd gnd cell_6t
Xbit_r120_c87 bl_87 br_87 wl_120 vdd gnd cell_6t
Xbit_r121_c87 bl_87 br_87 wl_121 vdd gnd cell_6t
Xbit_r122_c87 bl_87 br_87 wl_122 vdd gnd cell_6t
Xbit_r123_c87 bl_87 br_87 wl_123 vdd gnd cell_6t
Xbit_r124_c87 bl_87 br_87 wl_124 vdd gnd cell_6t
Xbit_r125_c87 bl_87 br_87 wl_125 vdd gnd cell_6t
Xbit_r126_c87 bl_87 br_87 wl_126 vdd gnd cell_6t
Xbit_r127_c87 bl_87 br_87 wl_127 vdd gnd cell_6t
Xbit_r128_c87 bl_87 br_87 wl_128 vdd gnd cell_6t
Xbit_r129_c87 bl_87 br_87 wl_129 vdd gnd cell_6t
Xbit_r130_c87 bl_87 br_87 wl_130 vdd gnd cell_6t
Xbit_r131_c87 bl_87 br_87 wl_131 vdd gnd cell_6t
Xbit_r132_c87 bl_87 br_87 wl_132 vdd gnd cell_6t
Xbit_r133_c87 bl_87 br_87 wl_133 vdd gnd cell_6t
Xbit_r134_c87 bl_87 br_87 wl_134 vdd gnd cell_6t
Xbit_r135_c87 bl_87 br_87 wl_135 vdd gnd cell_6t
Xbit_r136_c87 bl_87 br_87 wl_136 vdd gnd cell_6t
Xbit_r137_c87 bl_87 br_87 wl_137 vdd gnd cell_6t
Xbit_r138_c87 bl_87 br_87 wl_138 vdd gnd cell_6t
Xbit_r139_c87 bl_87 br_87 wl_139 vdd gnd cell_6t
Xbit_r140_c87 bl_87 br_87 wl_140 vdd gnd cell_6t
Xbit_r141_c87 bl_87 br_87 wl_141 vdd gnd cell_6t
Xbit_r142_c87 bl_87 br_87 wl_142 vdd gnd cell_6t
Xbit_r143_c87 bl_87 br_87 wl_143 vdd gnd cell_6t
Xbit_r144_c87 bl_87 br_87 wl_144 vdd gnd cell_6t
Xbit_r145_c87 bl_87 br_87 wl_145 vdd gnd cell_6t
Xbit_r146_c87 bl_87 br_87 wl_146 vdd gnd cell_6t
Xbit_r147_c87 bl_87 br_87 wl_147 vdd gnd cell_6t
Xbit_r148_c87 bl_87 br_87 wl_148 vdd gnd cell_6t
Xbit_r149_c87 bl_87 br_87 wl_149 vdd gnd cell_6t
Xbit_r150_c87 bl_87 br_87 wl_150 vdd gnd cell_6t
Xbit_r151_c87 bl_87 br_87 wl_151 vdd gnd cell_6t
Xbit_r152_c87 bl_87 br_87 wl_152 vdd gnd cell_6t
Xbit_r153_c87 bl_87 br_87 wl_153 vdd gnd cell_6t
Xbit_r154_c87 bl_87 br_87 wl_154 vdd gnd cell_6t
Xbit_r155_c87 bl_87 br_87 wl_155 vdd gnd cell_6t
Xbit_r156_c87 bl_87 br_87 wl_156 vdd gnd cell_6t
Xbit_r157_c87 bl_87 br_87 wl_157 vdd gnd cell_6t
Xbit_r158_c87 bl_87 br_87 wl_158 vdd gnd cell_6t
Xbit_r159_c87 bl_87 br_87 wl_159 vdd gnd cell_6t
Xbit_r160_c87 bl_87 br_87 wl_160 vdd gnd cell_6t
Xbit_r161_c87 bl_87 br_87 wl_161 vdd gnd cell_6t
Xbit_r162_c87 bl_87 br_87 wl_162 vdd gnd cell_6t
Xbit_r163_c87 bl_87 br_87 wl_163 vdd gnd cell_6t
Xbit_r164_c87 bl_87 br_87 wl_164 vdd gnd cell_6t
Xbit_r165_c87 bl_87 br_87 wl_165 vdd gnd cell_6t
Xbit_r166_c87 bl_87 br_87 wl_166 vdd gnd cell_6t
Xbit_r167_c87 bl_87 br_87 wl_167 vdd gnd cell_6t
Xbit_r168_c87 bl_87 br_87 wl_168 vdd gnd cell_6t
Xbit_r169_c87 bl_87 br_87 wl_169 vdd gnd cell_6t
Xbit_r170_c87 bl_87 br_87 wl_170 vdd gnd cell_6t
Xbit_r171_c87 bl_87 br_87 wl_171 vdd gnd cell_6t
Xbit_r172_c87 bl_87 br_87 wl_172 vdd gnd cell_6t
Xbit_r173_c87 bl_87 br_87 wl_173 vdd gnd cell_6t
Xbit_r174_c87 bl_87 br_87 wl_174 vdd gnd cell_6t
Xbit_r175_c87 bl_87 br_87 wl_175 vdd gnd cell_6t
Xbit_r176_c87 bl_87 br_87 wl_176 vdd gnd cell_6t
Xbit_r177_c87 bl_87 br_87 wl_177 vdd gnd cell_6t
Xbit_r178_c87 bl_87 br_87 wl_178 vdd gnd cell_6t
Xbit_r179_c87 bl_87 br_87 wl_179 vdd gnd cell_6t
Xbit_r180_c87 bl_87 br_87 wl_180 vdd gnd cell_6t
Xbit_r181_c87 bl_87 br_87 wl_181 vdd gnd cell_6t
Xbit_r182_c87 bl_87 br_87 wl_182 vdd gnd cell_6t
Xbit_r183_c87 bl_87 br_87 wl_183 vdd gnd cell_6t
Xbit_r184_c87 bl_87 br_87 wl_184 vdd gnd cell_6t
Xbit_r185_c87 bl_87 br_87 wl_185 vdd gnd cell_6t
Xbit_r186_c87 bl_87 br_87 wl_186 vdd gnd cell_6t
Xbit_r187_c87 bl_87 br_87 wl_187 vdd gnd cell_6t
Xbit_r188_c87 bl_87 br_87 wl_188 vdd gnd cell_6t
Xbit_r189_c87 bl_87 br_87 wl_189 vdd gnd cell_6t
Xbit_r190_c87 bl_87 br_87 wl_190 vdd gnd cell_6t
Xbit_r191_c87 bl_87 br_87 wl_191 vdd gnd cell_6t
Xbit_r192_c87 bl_87 br_87 wl_192 vdd gnd cell_6t
Xbit_r193_c87 bl_87 br_87 wl_193 vdd gnd cell_6t
Xbit_r194_c87 bl_87 br_87 wl_194 vdd gnd cell_6t
Xbit_r195_c87 bl_87 br_87 wl_195 vdd gnd cell_6t
Xbit_r196_c87 bl_87 br_87 wl_196 vdd gnd cell_6t
Xbit_r197_c87 bl_87 br_87 wl_197 vdd gnd cell_6t
Xbit_r198_c87 bl_87 br_87 wl_198 vdd gnd cell_6t
Xbit_r199_c87 bl_87 br_87 wl_199 vdd gnd cell_6t
Xbit_r200_c87 bl_87 br_87 wl_200 vdd gnd cell_6t
Xbit_r201_c87 bl_87 br_87 wl_201 vdd gnd cell_6t
Xbit_r202_c87 bl_87 br_87 wl_202 vdd gnd cell_6t
Xbit_r203_c87 bl_87 br_87 wl_203 vdd gnd cell_6t
Xbit_r204_c87 bl_87 br_87 wl_204 vdd gnd cell_6t
Xbit_r205_c87 bl_87 br_87 wl_205 vdd gnd cell_6t
Xbit_r206_c87 bl_87 br_87 wl_206 vdd gnd cell_6t
Xbit_r207_c87 bl_87 br_87 wl_207 vdd gnd cell_6t
Xbit_r208_c87 bl_87 br_87 wl_208 vdd gnd cell_6t
Xbit_r209_c87 bl_87 br_87 wl_209 vdd gnd cell_6t
Xbit_r210_c87 bl_87 br_87 wl_210 vdd gnd cell_6t
Xbit_r211_c87 bl_87 br_87 wl_211 vdd gnd cell_6t
Xbit_r212_c87 bl_87 br_87 wl_212 vdd gnd cell_6t
Xbit_r213_c87 bl_87 br_87 wl_213 vdd gnd cell_6t
Xbit_r214_c87 bl_87 br_87 wl_214 vdd gnd cell_6t
Xbit_r215_c87 bl_87 br_87 wl_215 vdd gnd cell_6t
Xbit_r216_c87 bl_87 br_87 wl_216 vdd gnd cell_6t
Xbit_r217_c87 bl_87 br_87 wl_217 vdd gnd cell_6t
Xbit_r218_c87 bl_87 br_87 wl_218 vdd gnd cell_6t
Xbit_r219_c87 bl_87 br_87 wl_219 vdd gnd cell_6t
Xbit_r220_c87 bl_87 br_87 wl_220 vdd gnd cell_6t
Xbit_r221_c87 bl_87 br_87 wl_221 vdd gnd cell_6t
Xbit_r222_c87 bl_87 br_87 wl_222 vdd gnd cell_6t
Xbit_r223_c87 bl_87 br_87 wl_223 vdd gnd cell_6t
Xbit_r224_c87 bl_87 br_87 wl_224 vdd gnd cell_6t
Xbit_r225_c87 bl_87 br_87 wl_225 vdd gnd cell_6t
Xbit_r226_c87 bl_87 br_87 wl_226 vdd gnd cell_6t
Xbit_r227_c87 bl_87 br_87 wl_227 vdd gnd cell_6t
Xbit_r228_c87 bl_87 br_87 wl_228 vdd gnd cell_6t
Xbit_r229_c87 bl_87 br_87 wl_229 vdd gnd cell_6t
Xbit_r230_c87 bl_87 br_87 wl_230 vdd gnd cell_6t
Xbit_r231_c87 bl_87 br_87 wl_231 vdd gnd cell_6t
Xbit_r232_c87 bl_87 br_87 wl_232 vdd gnd cell_6t
Xbit_r233_c87 bl_87 br_87 wl_233 vdd gnd cell_6t
Xbit_r234_c87 bl_87 br_87 wl_234 vdd gnd cell_6t
Xbit_r235_c87 bl_87 br_87 wl_235 vdd gnd cell_6t
Xbit_r236_c87 bl_87 br_87 wl_236 vdd gnd cell_6t
Xbit_r237_c87 bl_87 br_87 wl_237 vdd gnd cell_6t
Xbit_r238_c87 bl_87 br_87 wl_238 vdd gnd cell_6t
Xbit_r239_c87 bl_87 br_87 wl_239 vdd gnd cell_6t
Xbit_r240_c87 bl_87 br_87 wl_240 vdd gnd cell_6t
Xbit_r241_c87 bl_87 br_87 wl_241 vdd gnd cell_6t
Xbit_r242_c87 bl_87 br_87 wl_242 vdd gnd cell_6t
Xbit_r243_c87 bl_87 br_87 wl_243 vdd gnd cell_6t
Xbit_r244_c87 bl_87 br_87 wl_244 vdd gnd cell_6t
Xbit_r245_c87 bl_87 br_87 wl_245 vdd gnd cell_6t
Xbit_r246_c87 bl_87 br_87 wl_246 vdd gnd cell_6t
Xbit_r247_c87 bl_87 br_87 wl_247 vdd gnd cell_6t
Xbit_r248_c87 bl_87 br_87 wl_248 vdd gnd cell_6t
Xbit_r249_c87 bl_87 br_87 wl_249 vdd gnd cell_6t
Xbit_r250_c87 bl_87 br_87 wl_250 vdd gnd cell_6t
Xbit_r251_c87 bl_87 br_87 wl_251 vdd gnd cell_6t
Xbit_r252_c87 bl_87 br_87 wl_252 vdd gnd cell_6t
Xbit_r253_c87 bl_87 br_87 wl_253 vdd gnd cell_6t
Xbit_r254_c87 bl_87 br_87 wl_254 vdd gnd cell_6t
Xbit_r255_c87 bl_87 br_87 wl_255 vdd gnd cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd cell_6t
Xbit_r1_c88 bl_88 br_88 wl_1 vdd gnd cell_6t
Xbit_r2_c88 bl_88 br_88 wl_2 vdd gnd cell_6t
Xbit_r3_c88 bl_88 br_88 wl_3 vdd gnd cell_6t
Xbit_r4_c88 bl_88 br_88 wl_4 vdd gnd cell_6t
Xbit_r5_c88 bl_88 br_88 wl_5 vdd gnd cell_6t
Xbit_r6_c88 bl_88 br_88 wl_6 vdd gnd cell_6t
Xbit_r7_c88 bl_88 br_88 wl_7 vdd gnd cell_6t
Xbit_r8_c88 bl_88 br_88 wl_8 vdd gnd cell_6t
Xbit_r9_c88 bl_88 br_88 wl_9 vdd gnd cell_6t
Xbit_r10_c88 bl_88 br_88 wl_10 vdd gnd cell_6t
Xbit_r11_c88 bl_88 br_88 wl_11 vdd gnd cell_6t
Xbit_r12_c88 bl_88 br_88 wl_12 vdd gnd cell_6t
Xbit_r13_c88 bl_88 br_88 wl_13 vdd gnd cell_6t
Xbit_r14_c88 bl_88 br_88 wl_14 vdd gnd cell_6t
Xbit_r15_c88 bl_88 br_88 wl_15 vdd gnd cell_6t
Xbit_r16_c88 bl_88 br_88 wl_16 vdd gnd cell_6t
Xbit_r17_c88 bl_88 br_88 wl_17 vdd gnd cell_6t
Xbit_r18_c88 bl_88 br_88 wl_18 vdd gnd cell_6t
Xbit_r19_c88 bl_88 br_88 wl_19 vdd gnd cell_6t
Xbit_r20_c88 bl_88 br_88 wl_20 vdd gnd cell_6t
Xbit_r21_c88 bl_88 br_88 wl_21 vdd gnd cell_6t
Xbit_r22_c88 bl_88 br_88 wl_22 vdd gnd cell_6t
Xbit_r23_c88 bl_88 br_88 wl_23 vdd gnd cell_6t
Xbit_r24_c88 bl_88 br_88 wl_24 vdd gnd cell_6t
Xbit_r25_c88 bl_88 br_88 wl_25 vdd gnd cell_6t
Xbit_r26_c88 bl_88 br_88 wl_26 vdd gnd cell_6t
Xbit_r27_c88 bl_88 br_88 wl_27 vdd gnd cell_6t
Xbit_r28_c88 bl_88 br_88 wl_28 vdd gnd cell_6t
Xbit_r29_c88 bl_88 br_88 wl_29 vdd gnd cell_6t
Xbit_r30_c88 bl_88 br_88 wl_30 vdd gnd cell_6t
Xbit_r31_c88 bl_88 br_88 wl_31 vdd gnd cell_6t
Xbit_r32_c88 bl_88 br_88 wl_32 vdd gnd cell_6t
Xbit_r33_c88 bl_88 br_88 wl_33 vdd gnd cell_6t
Xbit_r34_c88 bl_88 br_88 wl_34 vdd gnd cell_6t
Xbit_r35_c88 bl_88 br_88 wl_35 vdd gnd cell_6t
Xbit_r36_c88 bl_88 br_88 wl_36 vdd gnd cell_6t
Xbit_r37_c88 bl_88 br_88 wl_37 vdd gnd cell_6t
Xbit_r38_c88 bl_88 br_88 wl_38 vdd gnd cell_6t
Xbit_r39_c88 bl_88 br_88 wl_39 vdd gnd cell_6t
Xbit_r40_c88 bl_88 br_88 wl_40 vdd gnd cell_6t
Xbit_r41_c88 bl_88 br_88 wl_41 vdd gnd cell_6t
Xbit_r42_c88 bl_88 br_88 wl_42 vdd gnd cell_6t
Xbit_r43_c88 bl_88 br_88 wl_43 vdd gnd cell_6t
Xbit_r44_c88 bl_88 br_88 wl_44 vdd gnd cell_6t
Xbit_r45_c88 bl_88 br_88 wl_45 vdd gnd cell_6t
Xbit_r46_c88 bl_88 br_88 wl_46 vdd gnd cell_6t
Xbit_r47_c88 bl_88 br_88 wl_47 vdd gnd cell_6t
Xbit_r48_c88 bl_88 br_88 wl_48 vdd gnd cell_6t
Xbit_r49_c88 bl_88 br_88 wl_49 vdd gnd cell_6t
Xbit_r50_c88 bl_88 br_88 wl_50 vdd gnd cell_6t
Xbit_r51_c88 bl_88 br_88 wl_51 vdd gnd cell_6t
Xbit_r52_c88 bl_88 br_88 wl_52 vdd gnd cell_6t
Xbit_r53_c88 bl_88 br_88 wl_53 vdd gnd cell_6t
Xbit_r54_c88 bl_88 br_88 wl_54 vdd gnd cell_6t
Xbit_r55_c88 bl_88 br_88 wl_55 vdd gnd cell_6t
Xbit_r56_c88 bl_88 br_88 wl_56 vdd gnd cell_6t
Xbit_r57_c88 bl_88 br_88 wl_57 vdd gnd cell_6t
Xbit_r58_c88 bl_88 br_88 wl_58 vdd gnd cell_6t
Xbit_r59_c88 bl_88 br_88 wl_59 vdd gnd cell_6t
Xbit_r60_c88 bl_88 br_88 wl_60 vdd gnd cell_6t
Xbit_r61_c88 bl_88 br_88 wl_61 vdd gnd cell_6t
Xbit_r62_c88 bl_88 br_88 wl_62 vdd gnd cell_6t
Xbit_r63_c88 bl_88 br_88 wl_63 vdd gnd cell_6t
Xbit_r64_c88 bl_88 br_88 wl_64 vdd gnd cell_6t
Xbit_r65_c88 bl_88 br_88 wl_65 vdd gnd cell_6t
Xbit_r66_c88 bl_88 br_88 wl_66 vdd gnd cell_6t
Xbit_r67_c88 bl_88 br_88 wl_67 vdd gnd cell_6t
Xbit_r68_c88 bl_88 br_88 wl_68 vdd gnd cell_6t
Xbit_r69_c88 bl_88 br_88 wl_69 vdd gnd cell_6t
Xbit_r70_c88 bl_88 br_88 wl_70 vdd gnd cell_6t
Xbit_r71_c88 bl_88 br_88 wl_71 vdd gnd cell_6t
Xbit_r72_c88 bl_88 br_88 wl_72 vdd gnd cell_6t
Xbit_r73_c88 bl_88 br_88 wl_73 vdd gnd cell_6t
Xbit_r74_c88 bl_88 br_88 wl_74 vdd gnd cell_6t
Xbit_r75_c88 bl_88 br_88 wl_75 vdd gnd cell_6t
Xbit_r76_c88 bl_88 br_88 wl_76 vdd gnd cell_6t
Xbit_r77_c88 bl_88 br_88 wl_77 vdd gnd cell_6t
Xbit_r78_c88 bl_88 br_88 wl_78 vdd gnd cell_6t
Xbit_r79_c88 bl_88 br_88 wl_79 vdd gnd cell_6t
Xbit_r80_c88 bl_88 br_88 wl_80 vdd gnd cell_6t
Xbit_r81_c88 bl_88 br_88 wl_81 vdd gnd cell_6t
Xbit_r82_c88 bl_88 br_88 wl_82 vdd gnd cell_6t
Xbit_r83_c88 bl_88 br_88 wl_83 vdd gnd cell_6t
Xbit_r84_c88 bl_88 br_88 wl_84 vdd gnd cell_6t
Xbit_r85_c88 bl_88 br_88 wl_85 vdd gnd cell_6t
Xbit_r86_c88 bl_88 br_88 wl_86 vdd gnd cell_6t
Xbit_r87_c88 bl_88 br_88 wl_87 vdd gnd cell_6t
Xbit_r88_c88 bl_88 br_88 wl_88 vdd gnd cell_6t
Xbit_r89_c88 bl_88 br_88 wl_89 vdd gnd cell_6t
Xbit_r90_c88 bl_88 br_88 wl_90 vdd gnd cell_6t
Xbit_r91_c88 bl_88 br_88 wl_91 vdd gnd cell_6t
Xbit_r92_c88 bl_88 br_88 wl_92 vdd gnd cell_6t
Xbit_r93_c88 bl_88 br_88 wl_93 vdd gnd cell_6t
Xbit_r94_c88 bl_88 br_88 wl_94 vdd gnd cell_6t
Xbit_r95_c88 bl_88 br_88 wl_95 vdd gnd cell_6t
Xbit_r96_c88 bl_88 br_88 wl_96 vdd gnd cell_6t
Xbit_r97_c88 bl_88 br_88 wl_97 vdd gnd cell_6t
Xbit_r98_c88 bl_88 br_88 wl_98 vdd gnd cell_6t
Xbit_r99_c88 bl_88 br_88 wl_99 vdd gnd cell_6t
Xbit_r100_c88 bl_88 br_88 wl_100 vdd gnd cell_6t
Xbit_r101_c88 bl_88 br_88 wl_101 vdd gnd cell_6t
Xbit_r102_c88 bl_88 br_88 wl_102 vdd gnd cell_6t
Xbit_r103_c88 bl_88 br_88 wl_103 vdd gnd cell_6t
Xbit_r104_c88 bl_88 br_88 wl_104 vdd gnd cell_6t
Xbit_r105_c88 bl_88 br_88 wl_105 vdd gnd cell_6t
Xbit_r106_c88 bl_88 br_88 wl_106 vdd gnd cell_6t
Xbit_r107_c88 bl_88 br_88 wl_107 vdd gnd cell_6t
Xbit_r108_c88 bl_88 br_88 wl_108 vdd gnd cell_6t
Xbit_r109_c88 bl_88 br_88 wl_109 vdd gnd cell_6t
Xbit_r110_c88 bl_88 br_88 wl_110 vdd gnd cell_6t
Xbit_r111_c88 bl_88 br_88 wl_111 vdd gnd cell_6t
Xbit_r112_c88 bl_88 br_88 wl_112 vdd gnd cell_6t
Xbit_r113_c88 bl_88 br_88 wl_113 vdd gnd cell_6t
Xbit_r114_c88 bl_88 br_88 wl_114 vdd gnd cell_6t
Xbit_r115_c88 bl_88 br_88 wl_115 vdd gnd cell_6t
Xbit_r116_c88 bl_88 br_88 wl_116 vdd gnd cell_6t
Xbit_r117_c88 bl_88 br_88 wl_117 vdd gnd cell_6t
Xbit_r118_c88 bl_88 br_88 wl_118 vdd gnd cell_6t
Xbit_r119_c88 bl_88 br_88 wl_119 vdd gnd cell_6t
Xbit_r120_c88 bl_88 br_88 wl_120 vdd gnd cell_6t
Xbit_r121_c88 bl_88 br_88 wl_121 vdd gnd cell_6t
Xbit_r122_c88 bl_88 br_88 wl_122 vdd gnd cell_6t
Xbit_r123_c88 bl_88 br_88 wl_123 vdd gnd cell_6t
Xbit_r124_c88 bl_88 br_88 wl_124 vdd gnd cell_6t
Xbit_r125_c88 bl_88 br_88 wl_125 vdd gnd cell_6t
Xbit_r126_c88 bl_88 br_88 wl_126 vdd gnd cell_6t
Xbit_r127_c88 bl_88 br_88 wl_127 vdd gnd cell_6t
Xbit_r128_c88 bl_88 br_88 wl_128 vdd gnd cell_6t
Xbit_r129_c88 bl_88 br_88 wl_129 vdd gnd cell_6t
Xbit_r130_c88 bl_88 br_88 wl_130 vdd gnd cell_6t
Xbit_r131_c88 bl_88 br_88 wl_131 vdd gnd cell_6t
Xbit_r132_c88 bl_88 br_88 wl_132 vdd gnd cell_6t
Xbit_r133_c88 bl_88 br_88 wl_133 vdd gnd cell_6t
Xbit_r134_c88 bl_88 br_88 wl_134 vdd gnd cell_6t
Xbit_r135_c88 bl_88 br_88 wl_135 vdd gnd cell_6t
Xbit_r136_c88 bl_88 br_88 wl_136 vdd gnd cell_6t
Xbit_r137_c88 bl_88 br_88 wl_137 vdd gnd cell_6t
Xbit_r138_c88 bl_88 br_88 wl_138 vdd gnd cell_6t
Xbit_r139_c88 bl_88 br_88 wl_139 vdd gnd cell_6t
Xbit_r140_c88 bl_88 br_88 wl_140 vdd gnd cell_6t
Xbit_r141_c88 bl_88 br_88 wl_141 vdd gnd cell_6t
Xbit_r142_c88 bl_88 br_88 wl_142 vdd gnd cell_6t
Xbit_r143_c88 bl_88 br_88 wl_143 vdd gnd cell_6t
Xbit_r144_c88 bl_88 br_88 wl_144 vdd gnd cell_6t
Xbit_r145_c88 bl_88 br_88 wl_145 vdd gnd cell_6t
Xbit_r146_c88 bl_88 br_88 wl_146 vdd gnd cell_6t
Xbit_r147_c88 bl_88 br_88 wl_147 vdd gnd cell_6t
Xbit_r148_c88 bl_88 br_88 wl_148 vdd gnd cell_6t
Xbit_r149_c88 bl_88 br_88 wl_149 vdd gnd cell_6t
Xbit_r150_c88 bl_88 br_88 wl_150 vdd gnd cell_6t
Xbit_r151_c88 bl_88 br_88 wl_151 vdd gnd cell_6t
Xbit_r152_c88 bl_88 br_88 wl_152 vdd gnd cell_6t
Xbit_r153_c88 bl_88 br_88 wl_153 vdd gnd cell_6t
Xbit_r154_c88 bl_88 br_88 wl_154 vdd gnd cell_6t
Xbit_r155_c88 bl_88 br_88 wl_155 vdd gnd cell_6t
Xbit_r156_c88 bl_88 br_88 wl_156 vdd gnd cell_6t
Xbit_r157_c88 bl_88 br_88 wl_157 vdd gnd cell_6t
Xbit_r158_c88 bl_88 br_88 wl_158 vdd gnd cell_6t
Xbit_r159_c88 bl_88 br_88 wl_159 vdd gnd cell_6t
Xbit_r160_c88 bl_88 br_88 wl_160 vdd gnd cell_6t
Xbit_r161_c88 bl_88 br_88 wl_161 vdd gnd cell_6t
Xbit_r162_c88 bl_88 br_88 wl_162 vdd gnd cell_6t
Xbit_r163_c88 bl_88 br_88 wl_163 vdd gnd cell_6t
Xbit_r164_c88 bl_88 br_88 wl_164 vdd gnd cell_6t
Xbit_r165_c88 bl_88 br_88 wl_165 vdd gnd cell_6t
Xbit_r166_c88 bl_88 br_88 wl_166 vdd gnd cell_6t
Xbit_r167_c88 bl_88 br_88 wl_167 vdd gnd cell_6t
Xbit_r168_c88 bl_88 br_88 wl_168 vdd gnd cell_6t
Xbit_r169_c88 bl_88 br_88 wl_169 vdd gnd cell_6t
Xbit_r170_c88 bl_88 br_88 wl_170 vdd gnd cell_6t
Xbit_r171_c88 bl_88 br_88 wl_171 vdd gnd cell_6t
Xbit_r172_c88 bl_88 br_88 wl_172 vdd gnd cell_6t
Xbit_r173_c88 bl_88 br_88 wl_173 vdd gnd cell_6t
Xbit_r174_c88 bl_88 br_88 wl_174 vdd gnd cell_6t
Xbit_r175_c88 bl_88 br_88 wl_175 vdd gnd cell_6t
Xbit_r176_c88 bl_88 br_88 wl_176 vdd gnd cell_6t
Xbit_r177_c88 bl_88 br_88 wl_177 vdd gnd cell_6t
Xbit_r178_c88 bl_88 br_88 wl_178 vdd gnd cell_6t
Xbit_r179_c88 bl_88 br_88 wl_179 vdd gnd cell_6t
Xbit_r180_c88 bl_88 br_88 wl_180 vdd gnd cell_6t
Xbit_r181_c88 bl_88 br_88 wl_181 vdd gnd cell_6t
Xbit_r182_c88 bl_88 br_88 wl_182 vdd gnd cell_6t
Xbit_r183_c88 bl_88 br_88 wl_183 vdd gnd cell_6t
Xbit_r184_c88 bl_88 br_88 wl_184 vdd gnd cell_6t
Xbit_r185_c88 bl_88 br_88 wl_185 vdd gnd cell_6t
Xbit_r186_c88 bl_88 br_88 wl_186 vdd gnd cell_6t
Xbit_r187_c88 bl_88 br_88 wl_187 vdd gnd cell_6t
Xbit_r188_c88 bl_88 br_88 wl_188 vdd gnd cell_6t
Xbit_r189_c88 bl_88 br_88 wl_189 vdd gnd cell_6t
Xbit_r190_c88 bl_88 br_88 wl_190 vdd gnd cell_6t
Xbit_r191_c88 bl_88 br_88 wl_191 vdd gnd cell_6t
Xbit_r192_c88 bl_88 br_88 wl_192 vdd gnd cell_6t
Xbit_r193_c88 bl_88 br_88 wl_193 vdd gnd cell_6t
Xbit_r194_c88 bl_88 br_88 wl_194 vdd gnd cell_6t
Xbit_r195_c88 bl_88 br_88 wl_195 vdd gnd cell_6t
Xbit_r196_c88 bl_88 br_88 wl_196 vdd gnd cell_6t
Xbit_r197_c88 bl_88 br_88 wl_197 vdd gnd cell_6t
Xbit_r198_c88 bl_88 br_88 wl_198 vdd gnd cell_6t
Xbit_r199_c88 bl_88 br_88 wl_199 vdd gnd cell_6t
Xbit_r200_c88 bl_88 br_88 wl_200 vdd gnd cell_6t
Xbit_r201_c88 bl_88 br_88 wl_201 vdd gnd cell_6t
Xbit_r202_c88 bl_88 br_88 wl_202 vdd gnd cell_6t
Xbit_r203_c88 bl_88 br_88 wl_203 vdd gnd cell_6t
Xbit_r204_c88 bl_88 br_88 wl_204 vdd gnd cell_6t
Xbit_r205_c88 bl_88 br_88 wl_205 vdd gnd cell_6t
Xbit_r206_c88 bl_88 br_88 wl_206 vdd gnd cell_6t
Xbit_r207_c88 bl_88 br_88 wl_207 vdd gnd cell_6t
Xbit_r208_c88 bl_88 br_88 wl_208 vdd gnd cell_6t
Xbit_r209_c88 bl_88 br_88 wl_209 vdd gnd cell_6t
Xbit_r210_c88 bl_88 br_88 wl_210 vdd gnd cell_6t
Xbit_r211_c88 bl_88 br_88 wl_211 vdd gnd cell_6t
Xbit_r212_c88 bl_88 br_88 wl_212 vdd gnd cell_6t
Xbit_r213_c88 bl_88 br_88 wl_213 vdd gnd cell_6t
Xbit_r214_c88 bl_88 br_88 wl_214 vdd gnd cell_6t
Xbit_r215_c88 bl_88 br_88 wl_215 vdd gnd cell_6t
Xbit_r216_c88 bl_88 br_88 wl_216 vdd gnd cell_6t
Xbit_r217_c88 bl_88 br_88 wl_217 vdd gnd cell_6t
Xbit_r218_c88 bl_88 br_88 wl_218 vdd gnd cell_6t
Xbit_r219_c88 bl_88 br_88 wl_219 vdd gnd cell_6t
Xbit_r220_c88 bl_88 br_88 wl_220 vdd gnd cell_6t
Xbit_r221_c88 bl_88 br_88 wl_221 vdd gnd cell_6t
Xbit_r222_c88 bl_88 br_88 wl_222 vdd gnd cell_6t
Xbit_r223_c88 bl_88 br_88 wl_223 vdd gnd cell_6t
Xbit_r224_c88 bl_88 br_88 wl_224 vdd gnd cell_6t
Xbit_r225_c88 bl_88 br_88 wl_225 vdd gnd cell_6t
Xbit_r226_c88 bl_88 br_88 wl_226 vdd gnd cell_6t
Xbit_r227_c88 bl_88 br_88 wl_227 vdd gnd cell_6t
Xbit_r228_c88 bl_88 br_88 wl_228 vdd gnd cell_6t
Xbit_r229_c88 bl_88 br_88 wl_229 vdd gnd cell_6t
Xbit_r230_c88 bl_88 br_88 wl_230 vdd gnd cell_6t
Xbit_r231_c88 bl_88 br_88 wl_231 vdd gnd cell_6t
Xbit_r232_c88 bl_88 br_88 wl_232 vdd gnd cell_6t
Xbit_r233_c88 bl_88 br_88 wl_233 vdd gnd cell_6t
Xbit_r234_c88 bl_88 br_88 wl_234 vdd gnd cell_6t
Xbit_r235_c88 bl_88 br_88 wl_235 vdd gnd cell_6t
Xbit_r236_c88 bl_88 br_88 wl_236 vdd gnd cell_6t
Xbit_r237_c88 bl_88 br_88 wl_237 vdd gnd cell_6t
Xbit_r238_c88 bl_88 br_88 wl_238 vdd gnd cell_6t
Xbit_r239_c88 bl_88 br_88 wl_239 vdd gnd cell_6t
Xbit_r240_c88 bl_88 br_88 wl_240 vdd gnd cell_6t
Xbit_r241_c88 bl_88 br_88 wl_241 vdd gnd cell_6t
Xbit_r242_c88 bl_88 br_88 wl_242 vdd gnd cell_6t
Xbit_r243_c88 bl_88 br_88 wl_243 vdd gnd cell_6t
Xbit_r244_c88 bl_88 br_88 wl_244 vdd gnd cell_6t
Xbit_r245_c88 bl_88 br_88 wl_245 vdd gnd cell_6t
Xbit_r246_c88 bl_88 br_88 wl_246 vdd gnd cell_6t
Xbit_r247_c88 bl_88 br_88 wl_247 vdd gnd cell_6t
Xbit_r248_c88 bl_88 br_88 wl_248 vdd gnd cell_6t
Xbit_r249_c88 bl_88 br_88 wl_249 vdd gnd cell_6t
Xbit_r250_c88 bl_88 br_88 wl_250 vdd gnd cell_6t
Xbit_r251_c88 bl_88 br_88 wl_251 vdd gnd cell_6t
Xbit_r252_c88 bl_88 br_88 wl_252 vdd gnd cell_6t
Xbit_r253_c88 bl_88 br_88 wl_253 vdd gnd cell_6t
Xbit_r254_c88 bl_88 br_88 wl_254 vdd gnd cell_6t
Xbit_r255_c88 bl_88 br_88 wl_255 vdd gnd cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd cell_6t
Xbit_r1_c89 bl_89 br_89 wl_1 vdd gnd cell_6t
Xbit_r2_c89 bl_89 br_89 wl_2 vdd gnd cell_6t
Xbit_r3_c89 bl_89 br_89 wl_3 vdd gnd cell_6t
Xbit_r4_c89 bl_89 br_89 wl_4 vdd gnd cell_6t
Xbit_r5_c89 bl_89 br_89 wl_5 vdd gnd cell_6t
Xbit_r6_c89 bl_89 br_89 wl_6 vdd gnd cell_6t
Xbit_r7_c89 bl_89 br_89 wl_7 vdd gnd cell_6t
Xbit_r8_c89 bl_89 br_89 wl_8 vdd gnd cell_6t
Xbit_r9_c89 bl_89 br_89 wl_9 vdd gnd cell_6t
Xbit_r10_c89 bl_89 br_89 wl_10 vdd gnd cell_6t
Xbit_r11_c89 bl_89 br_89 wl_11 vdd gnd cell_6t
Xbit_r12_c89 bl_89 br_89 wl_12 vdd gnd cell_6t
Xbit_r13_c89 bl_89 br_89 wl_13 vdd gnd cell_6t
Xbit_r14_c89 bl_89 br_89 wl_14 vdd gnd cell_6t
Xbit_r15_c89 bl_89 br_89 wl_15 vdd gnd cell_6t
Xbit_r16_c89 bl_89 br_89 wl_16 vdd gnd cell_6t
Xbit_r17_c89 bl_89 br_89 wl_17 vdd gnd cell_6t
Xbit_r18_c89 bl_89 br_89 wl_18 vdd gnd cell_6t
Xbit_r19_c89 bl_89 br_89 wl_19 vdd gnd cell_6t
Xbit_r20_c89 bl_89 br_89 wl_20 vdd gnd cell_6t
Xbit_r21_c89 bl_89 br_89 wl_21 vdd gnd cell_6t
Xbit_r22_c89 bl_89 br_89 wl_22 vdd gnd cell_6t
Xbit_r23_c89 bl_89 br_89 wl_23 vdd gnd cell_6t
Xbit_r24_c89 bl_89 br_89 wl_24 vdd gnd cell_6t
Xbit_r25_c89 bl_89 br_89 wl_25 vdd gnd cell_6t
Xbit_r26_c89 bl_89 br_89 wl_26 vdd gnd cell_6t
Xbit_r27_c89 bl_89 br_89 wl_27 vdd gnd cell_6t
Xbit_r28_c89 bl_89 br_89 wl_28 vdd gnd cell_6t
Xbit_r29_c89 bl_89 br_89 wl_29 vdd gnd cell_6t
Xbit_r30_c89 bl_89 br_89 wl_30 vdd gnd cell_6t
Xbit_r31_c89 bl_89 br_89 wl_31 vdd gnd cell_6t
Xbit_r32_c89 bl_89 br_89 wl_32 vdd gnd cell_6t
Xbit_r33_c89 bl_89 br_89 wl_33 vdd gnd cell_6t
Xbit_r34_c89 bl_89 br_89 wl_34 vdd gnd cell_6t
Xbit_r35_c89 bl_89 br_89 wl_35 vdd gnd cell_6t
Xbit_r36_c89 bl_89 br_89 wl_36 vdd gnd cell_6t
Xbit_r37_c89 bl_89 br_89 wl_37 vdd gnd cell_6t
Xbit_r38_c89 bl_89 br_89 wl_38 vdd gnd cell_6t
Xbit_r39_c89 bl_89 br_89 wl_39 vdd gnd cell_6t
Xbit_r40_c89 bl_89 br_89 wl_40 vdd gnd cell_6t
Xbit_r41_c89 bl_89 br_89 wl_41 vdd gnd cell_6t
Xbit_r42_c89 bl_89 br_89 wl_42 vdd gnd cell_6t
Xbit_r43_c89 bl_89 br_89 wl_43 vdd gnd cell_6t
Xbit_r44_c89 bl_89 br_89 wl_44 vdd gnd cell_6t
Xbit_r45_c89 bl_89 br_89 wl_45 vdd gnd cell_6t
Xbit_r46_c89 bl_89 br_89 wl_46 vdd gnd cell_6t
Xbit_r47_c89 bl_89 br_89 wl_47 vdd gnd cell_6t
Xbit_r48_c89 bl_89 br_89 wl_48 vdd gnd cell_6t
Xbit_r49_c89 bl_89 br_89 wl_49 vdd gnd cell_6t
Xbit_r50_c89 bl_89 br_89 wl_50 vdd gnd cell_6t
Xbit_r51_c89 bl_89 br_89 wl_51 vdd gnd cell_6t
Xbit_r52_c89 bl_89 br_89 wl_52 vdd gnd cell_6t
Xbit_r53_c89 bl_89 br_89 wl_53 vdd gnd cell_6t
Xbit_r54_c89 bl_89 br_89 wl_54 vdd gnd cell_6t
Xbit_r55_c89 bl_89 br_89 wl_55 vdd gnd cell_6t
Xbit_r56_c89 bl_89 br_89 wl_56 vdd gnd cell_6t
Xbit_r57_c89 bl_89 br_89 wl_57 vdd gnd cell_6t
Xbit_r58_c89 bl_89 br_89 wl_58 vdd gnd cell_6t
Xbit_r59_c89 bl_89 br_89 wl_59 vdd gnd cell_6t
Xbit_r60_c89 bl_89 br_89 wl_60 vdd gnd cell_6t
Xbit_r61_c89 bl_89 br_89 wl_61 vdd gnd cell_6t
Xbit_r62_c89 bl_89 br_89 wl_62 vdd gnd cell_6t
Xbit_r63_c89 bl_89 br_89 wl_63 vdd gnd cell_6t
Xbit_r64_c89 bl_89 br_89 wl_64 vdd gnd cell_6t
Xbit_r65_c89 bl_89 br_89 wl_65 vdd gnd cell_6t
Xbit_r66_c89 bl_89 br_89 wl_66 vdd gnd cell_6t
Xbit_r67_c89 bl_89 br_89 wl_67 vdd gnd cell_6t
Xbit_r68_c89 bl_89 br_89 wl_68 vdd gnd cell_6t
Xbit_r69_c89 bl_89 br_89 wl_69 vdd gnd cell_6t
Xbit_r70_c89 bl_89 br_89 wl_70 vdd gnd cell_6t
Xbit_r71_c89 bl_89 br_89 wl_71 vdd gnd cell_6t
Xbit_r72_c89 bl_89 br_89 wl_72 vdd gnd cell_6t
Xbit_r73_c89 bl_89 br_89 wl_73 vdd gnd cell_6t
Xbit_r74_c89 bl_89 br_89 wl_74 vdd gnd cell_6t
Xbit_r75_c89 bl_89 br_89 wl_75 vdd gnd cell_6t
Xbit_r76_c89 bl_89 br_89 wl_76 vdd gnd cell_6t
Xbit_r77_c89 bl_89 br_89 wl_77 vdd gnd cell_6t
Xbit_r78_c89 bl_89 br_89 wl_78 vdd gnd cell_6t
Xbit_r79_c89 bl_89 br_89 wl_79 vdd gnd cell_6t
Xbit_r80_c89 bl_89 br_89 wl_80 vdd gnd cell_6t
Xbit_r81_c89 bl_89 br_89 wl_81 vdd gnd cell_6t
Xbit_r82_c89 bl_89 br_89 wl_82 vdd gnd cell_6t
Xbit_r83_c89 bl_89 br_89 wl_83 vdd gnd cell_6t
Xbit_r84_c89 bl_89 br_89 wl_84 vdd gnd cell_6t
Xbit_r85_c89 bl_89 br_89 wl_85 vdd gnd cell_6t
Xbit_r86_c89 bl_89 br_89 wl_86 vdd gnd cell_6t
Xbit_r87_c89 bl_89 br_89 wl_87 vdd gnd cell_6t
Xbit_r88_c89 bl_89 br_89 wl_88 vdd gnd cell_6t
Xbit_r89_c89 bl_89 br_89 wl_89 vdd gnd cell_6t
Xbit_r90_c89 bl_89 br_89 wl_90 vdd gnd cell_6t
Xbit_r91_c89 bl_89 br_89 wl_91 vdd gnd cell_6t
Xbit_r92_c89 bl_89 br_89 wl_92 vdd gnd cell_6t
Xbit_r93_c89 bl_89 br_89 wl_93 vdd gnd cell_6t
Xbit_r94_c89 bl_89 br_89 wl_94 vdd gnd cell_6t
Xbit_r95_c89 bl_89 br_89 wl_95 vdd gnd cell_6t
Xbit_r96_c89 bl_89 br_89 wl_96 vdd gnd cell_6t
Xbit_r97_c89 bl_89 br_89 wl_97 vdd gnd cell_6t
Xbit_r98_c89 bl_89 br_89 wl_98 vdd gnd cell_6t
Xbit_r99_c89 bl_89 br_89 wl_99 vdd gnd cell_6t
Xbit_r100_c89 bl_89 br_89 wl_100 vdd gnd cell_6t
Xbit_r101_c89 bl_89 br_89 wl_101 vdd gnd cell_6t
Xbit_r102_c89 bl_89 br_89 wl_102 vdd gnd cell_6t
Xbit_r103_c89 bl_89 br_89 wl_103 vdd gnd cell_6t
Xbit_r104_c89 bl_89 br_89 wl_104 vdd gnd cell_6t
Xbit_r105_c89 bl_89 br_89 wl_105 vdd gnd cell_6t
Xbit_r106_c89 bl_89 br_89 wl_106 vdd gnd cell_6t
Xbit_r107_c89 bl_89 br_89 wl_107 vdd gnd cell_6t
Xbit_r108_c89 bl_89 br_89 wl_108 vdd gnd cell_6t
Xbit_r109_c89 bl_89 br_89 wl_109 vdd gnd cell_6t
Xbit_r110_c89 bl_89 br_89 wl_110 vdd gnd cell_6t
Xbit_r111_c89 bl_89 br_89 wl_111 vdd gnd cell_6t
Xbit_r112_c89 bl_89 br_89 wl_112 vdd gnd cell_6t
Xbit_r113_c89 bl_89 br_89 wl_113 vdd gnd cell_6t
Xbit_r114_c89 bl_89 br_89 wl_114 vdd gnd cell_6t
Xbit_r115_c89 bl_89 br_89 wl_115 vdd gnd cell_6t
Xbit_r116_c89 bl_89 br_89 wl_116 vdd gnd cell_6t
Xbit_r117_c89 bl_89 br_89 wl_117 vdd gnd cell_6t
Xbit_r118_c89 bl_89 br_89 wl_118 vdd gnd cell_6t
Xbit_r119_c89 bl_89 br_89 wl_119 vdd gnd cell_6t
Xbit_r120_c89 bl_89 br_89 wl_120 vdd gnd cell_6t
Xbit_r121_c89 bl_89 br_89 wl_121 vdd gnd cell_6t
Xbit_r122_c89 bl_89 br_89 wl_122 vdd gnd cell_6t
Xbit_r123_c89 bl_89 br_89 wl_123 vdd gnd cell_6t
Xbit_r124_c89 bl_89 br_89 wl_124 vdd gnd cell_6t
Xbit_r125_c89 bl_89 br_89 wl_125 vdd gnd cell_6t
Xbit_r126_c89 bl_89 br_89 wl_126 vdd gnd cell_6t
Xbit_r127_c89 bl_89 br_89 wl_127 vdd gnd cell_6t
Xbit_r128_c89 bl_89 br_89 wl_128 vdd gnd cell_6t
Xbit_r129_c89 bl_89 br_89 wl_129 vdd gnd cell_6t
Xbit_r130_c89 bl_89 br_89 wl_130 vdd gnd cell_6t
Xbit_r131_c89 bl_89 br_89 wl_131 vdd gnd cell_6t
Xbit_r132_c89 bl_89 br_89 wl_132 vdd gnd cell_6t
Xbit_r133_c89 bl_89 br_89 wl_133 vdd gnd cell_6t
Xbit_r134_c89 bl_89 br_89 wl_134 vdd gnd cell_6t
Xbit_r135_c89 bl_89 br_89 wl_135 vdd gnd cell_6t
Xbit_r136_c89 bl_89 br_89 wl_136 vdd gnd cell_6t
Xbit_r137_c89 bl_89 br_89 wl_137 vdd gnd cell_6t
Xbit_r138_c89 bl_89 br_89 wl_138 vdd gnd cell_6t
Xbit_r139_c89 bl_89 br_89 wl_139 vdd gnd cell_6t
Xbit_r140_c89 bl_89 br_89 wl_140 vdd gnd cell_6t
Xbit_r141_c89 bl_89 br_89 wl_141 vdd gnd cell_6t
Xbit_r142_c89 bl_89 br_89 wl_142 vdd gnd cell_6t
Xbit_r143_c89 bl_89 br_89 wl_143 vdd gnd cell_6t
Xbit_r144_c89 bl_89 br_89 wl_144 vdd gnd cell_6t
Xbit_r145_c89 bl_89 br_89 wl_145 vdd gnd cell_6t
Xbit_r146_c89 bl_89 br_89 wl_146 vdd gnd cell_6t
Xbit_r147_c89 bl_89 br_89 wl_147 vdd gnd cell_6t
Xbit_r148_c89 bl_89 br_89 wl_148 vdd gnd cell_6t
Xbit_r149_c89 bl_89 br_89 wl_149 vdd gnd cell_6t
Xbit_r150_c89 bl_89 br_89 wl_150 vdd gnd cell_6t
Xbit_r151_c89 bl_89 br_89 wl_151 vdd gnd cell_6t
Xbit_r152_c89 bl_89 br_89 wl_152 vdd gnd cell_6t
Xbit_r153_c89 bl_89 br_89 wl_153 vdd gnd cell_6t
Xbit_r154_c89 bl_89 br_89 wl_154 vdd gnd cell_6t
Xbit_r155_c89 bl_89 br_89 wl_155 vdd gnd cell_6t
Xbit_r156_c89 bl_89 br_89 wl_156 vdd gnd cell_6t
Xbit_r157_c89 bl_89 br_89 wl_157 vdd gnd cell_6t
Xbit_r158_c89 bl_89 br_89 wl_158 vdd gnd cell_6t
Xbit_r159_c89 bl_89 br_89 wl_159 vdd gnd cell_6t
Xbit_r160_c89 bl_89 br_89 wl_160 vdd gnd cell_6t
Xbit_r161_c89 bl_89 br_89 wl_161 vdd gnd cell_6t
Xbit_r162_c89 bl_89 br_89 wl_162 vdd gnd cell_6t
Xbit_r163_c89 bl_89 br_89 wl_163 vdd gnd cell_6t
Xbit_r164_c89 bl_89 br_89 wl_164 vdd gnd cell_6t
Xbit_r165_c89 bl_89 br_89 wl_165 vdd gnd cell_6t
Xbit_r166_c89 bl_89 br_89 wl_166 vdd gnd cell_6t
Xbit_r167_c89 bl_89 br_89 wl_167 vdd gnd cell_6t
Xbit_r168_c89 bl_89 br_89 wl_168 vdd gnd cell_6t
Xbit_r169_c89 bl_89 br_89 wl_169 vdd gnd cell_6t
Xbit_r170_c89 bl_89 br_89 wl_170 vdd gnd cell_6t
Xbit_r171_c89 bl_89 br_89 wl_171 vdd gnd cell_6t
Xbit_r172_c89 bl_89 br_89 wl_172 vdd gnd cell_6t
Xbit_r173_c89 bl_89 br_89 wl_173 vdd gnd cell_6t
Xbit_r174_c89 bl_89 br_89 wl_174 vdd gnd cell_6t
Xbit_r175_c89 bl_89 br_89 wl_175 vdd gnd cell_6t
Xbit_r176_c89 bl_89 br_89 wl_176 vdd gnd cell_6t
Xbit_r177_c89 bl_89 br_89 wl_177 vdd gnd cell_6t
Xbit_r178_c89 bl_89 br_89 wl_178 vdd gnd cell_6t
Xbit_r179_c89 bl_89 br_89 wl_179 vdd gnd cell_6t
Xbit_r180_c89 bl_89 br_89 wl_180 vdd gnd cell_6t
Xbit_r181_c89 bl_89 br_89 wl_181 vdd gnd cell_6t
Xbit_r182_c89 bl_89 br_89 wl_182 vdd gnd cell_6t
Xbit_r183_c89 bl_89 br_89 wl_183 vdd gnd cell_6t
Xbit_r184_c89 bl_89 br_89 wl_184 vdd gnd cell_6t
Xbit_r185_c89 bl_89 br_89 wl_185 vdd gnd cell_6t
Xbit_r186_c89 bl_89 br_89 wl_186 vdd gnd cell_6t
Xbit_r187_c89 bl_89 br_89 wl_187 vdd gnd cell_6t
Xbit_r188_c89 bl_89 br_89 wl_188 vdd gnd cell_6t
Xbit_r189_c89 bl_89 br_89 wl_189 vdd gnd cell_6t
Xbit_r190_c89 bl_89 br_89 wl_190 vdd gnd cell_6t
Xbit_r191_c89 bl_89 br_89 wl_191 vdd gnd cell_6t
Xbit_r192_c89 bl_89 br_89 wl_192 vdd gnd cell_6t
Xbit_r193_c89 bl_89 br_89 wl_193 vdd gnd cell_6t
Xbit_r194_c89 bl_89 br_89 wl_194 vdd gnd cell_6t
Xbit_r195_c89 bl_89 br_89 wl_195 vdd gnd cell_6t
Xbit_r196_c89 bl_89 br_89 wl_196 vdd gnd cell_6t
Xbit_r197_c89 bl_89 br_89 wl_197 vdd gnd cell_6t
Xbit_r198_c89 bl_89 br_89 wl_198 vdd gnd cell_6t
Xbit_r199_c89 bl_89 br_89 wl_199 vdd gnd cell_6t
Xbit_r200_c89 bl_89 br_89 wl_200 vdd gnd cell_6t
Xbit_r201_c89 bl_89 br_89 wl_201 vdd gnd cell_6t
Xbit_r202_c89 bl_89 br_89 wl_202 vdd gnd cell_6t
Xbit_r203_c89 bl_89 br_89 wl_203 vdd gnd cell_6t
Xbit_r204_c89 bl_89 br_89 wl_204 vdd gnd cell_6t
Xbit_r205_c89 bl_89 br_89 wl_205 vdd gnd cell_6t
Xbit_r206_c89 bl_89 br_89 wl_206 vdd gnd cell_6t
Xbit_r207_c89 bl_89 br_89 wl_207 vdd gnd cell_6t
Xbit_r208_c89 bl_89 br_89 wl_208 vdd gnd cell_6t
Xbit_r209_c89 bl_89 br_89 wl_209 vdd gnd cell_6t
Xbit_r210_c89 bl_89 br_89 wl_210 vdd gnd cell_6t
Xbit_r211_c89 bl_89 br_89 wl_211 vdd gnd cell_6t
Xbit_r212_c89 bl_89 br_89 wl_212 vdd gnd cell_6t
Xbit_r213_c89 bl_89 br_89 wl_213 vdd gnd cell_6t
Xbit_r214_c89 bl_89 br_89 wl_214 vdd gnd cell_6t
Xbit_r215_c89 bl_89 br_89 wl_215 vdd gnd cell_6t
Xbit_r216_c89 bl_89 br_89 wl_216 vdd gnd cell_6t
Xbit_r217_c89 bl_89 br_89 wl_217 vdd gnd cell_6t
Xbit_r218_c89 bl_89 br_89 wl_218 vdd gnd cell_6t
Xbit_r219_c89 bl_89 br_89 wl_219 vdd gnd cell_6t
Xbit_r220_c89 bl_89 br_89 wl_220 vdd gnd cell_6t
Xbit_r221_c89 bl_89 br_89 wl_221 vdd gnd cell_6t
Xbit_r222_c89 bl_89 br_89 wl_222 vdd gnd cell_6t
Xbit_r223_c89 bl_89 br_89 wl_223 vdd gnd cell_6t
Xbit_r224_c89 bl_89 br_89 wl_224 vdd gnd cell_6t
Xbit_r225_c89 bl_89 br_89 wl_225 vdd gnd cell_6t
Xbit_r226_c89 bl_89 br_89 wl_226 vdd gnd cell_6t
Xbit_r227_c89 bl_89 br_89 wl_227 vdd gnd cell_6t
Xbit_r228_c89 bl_89 br_89 wl_228 vdd gnd cell_6t
Xbit_r229_c89 bl_89 br_89 wl_229 vdd gnd cell_6t
Xbit_r230_c89 bl_89 br_89 wl_230 vdd gnd cell_6t
Xbit_r231_c89 bl_89 br_89 wl_231 vdd gnd cell_6t
Xbit_r232_c89 bl_89 br_89 wl_232 vdd gnd cell_6t
Xbit_r233_c89 bl_89 br_89 wl_233 vdd gnd cell_6t
Xbit_r234_c89 bl_89 br_89 wl_234 vdd gnd cell_6t
Xbit_r235_c89 bl_89 br_89 wl_235 vdd gnd cell_6t
Xbit_r236_c89 bl_89 br_89 wl_236 vdd gnd cell_6t
Xbit_r237_c89 bl_89 br_89 wl_237 vdd gnd cell_6t
Xbit_r238_c89 bl_89 br_89 wl_238 vdd gnd cell_6t
Xbit_r239_c89 bl_89 br_89 wl_239 vdd gnd cell_6t
Xbit_r240_c89 bl_89 br_89 wl_240 vdd gnd cell_6t
Xbit_r241_c89 bl_89 br_89 wl_241 vdd gnd cell_6t
Xbit_r242_c89 bl_89 br_89 wl_242 vdd gnd cell_6t
Xbit_r243_c89 bl_89 br_89 wl_243 vdd gnd cell_6t
Xbit_r244_c89 bl_89 br_89 wl_244 vdd gnd cell_6t
Xbit_r245_c89 bl_89 br_89 wl_245 vdd gnd cell_6t
Xbit_r246_c89 bl_89 br_89 wl_246 vdd gnd cell_6t
Xbit_r247_c89 bl_89 br_89 wl_247 vdd gnd cell_6t
Xbit_r248_c89 bl_89 br_89 wl_248 vdd gnd cell_6t
Xbit_r249_c89 bl_89 br_89 wl_249 vdd gnd cell_6t
Xbit_r250_c89 bl_89 br_89 wl_250 vdd gnd cell_6t
Xbit_r251_c89 bl_89 br_89 wl_251 vdd gnd cell_6t
Xbit_r252_c89 bl_89 br_89 wl_252 vdd gnd cell_6t
Xbit_r253_c89 bl_89 br_89 wl_253 vdd gnd cell_6t
Xbit_r254_c89 bl_89 br_89 wl_254 vdd gnd cell_6t
Xbit_r255_c89 bl_89 br_89 wl_255 vdd gnd cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd cell_6t
Xbit_r1_c90 bl_90 br_90 wl_1 vdd gnd cell_6t
Xbit_r2_c90 bl_90 br_90 wl_2 vdd gnd cell_6t
Xbit_r3_c90 bl_90 br_90 wl_3 vdd gnd cell_6t
Xbit_r4_c90 bl_90 br_90 wl_4 vdd gnd cell_6t
Xbit_r5_c90 bl_90 br_90 wl_5 vdd gnd cell_6t
Xbit_r6_c90 bl_90 br_90 wl_6 vdd gnd cell_6t
Xbit_r7_c90 bl_90 br_90 wl_7 vdd gnd cell_6t
Xbit_r8_c90 bl_90 br_90 wl_8 vdd gnd cell_6t
Xbit_r9_c90 bl_90 br_90 wl_9 vdd gnd cell_6t
Xbit_r10_c90 bl_90 br_90 wl_10 vdd gnd cell_6t
Xbit_r11_c90 bl_90 br_90 wl_11 vdd gnd cell_6t
Xbit_r12_c90 bl_90 br_90 wl_12 vdd gnd cell_6t
Xbit_r13_c90 bl_90 br_90 wl_13 vdd gnd cell_6t
Xbit_r14_c90 bl_90 br_90 wl_14 vdd gnd cell_6t
Xbit_r15_c90 bl_90 br_90 wl_15 vdd gnd cell_6t
Xbit_r16_c90 bl_90 br_90 wl_16 vdd gnd cell_6t
Xbit_r17_c90 bl_90 br_90 wl_17 vdd gnd cell_6t
Xbit_r18_c90 bl_90 br_90 wl_18 vdd gnd cell_6t
Xbit_r19_c90 bl_90 br_90 wl_19 vdd gnd cell_6t
Xbit_r20_c90 bl_90 br_90 wl_20 vdd gnd cell_6t
Xbit_r21_c90 bl_90 br_90 wl_21 vdd gnd cell_6t
Xbit_r22_c90 bl_90 br_90 wl_22 vdd gnd cell_6t
Xbit_r23_c90 bl_90 br_90 wl_23 vdd gnd cell_6t
Xbit_r24_c90 bl_90 br_90 wl_24 vdd gnd cell_6t
Xbit_r25_c90 bl_90 br_90 wl_25 vdd gnd cell_6t
Xbit_r26_c90 bl_90 br_90 wl_26 vdd gnd cell_6t
Xbit_r27_c90 bl_90 br_90 wl_27 vdd gnd cell_6t
Xbit_r28_c90 bl_90 br_90 wl_28 vdd gnd cell_6t
Xbit_r29_c90 bl_90 br_90 wl_29 vdd gnd cell_6t
Xbit_r30_c90 bl_90 br_90 wl_30 vdd gnd cell_6t
Xbit_r31_c90 bl_90 br_90 wl_31 vdd gnd cell_6t
Xbit_r32_c90 bl_90 br_90 wl_32 vdd gnd cell_6t
Xbit_r33_c90 bl_90 br_90 wl_33 vdd gnd cell_6t
Xbit_r34_c90 bl_90 br_90 wl_34 vdd gnd cell_6t
Xbit_r35_c90 bl_90 br_90 wl_35 vdd gnd cell_6t
Xbit_r36_c90 bl_90 br_90 wl_36 vdd gnd cell_6t
Xbit_r37_c90 bl_90 br_90 wl_37 vdd gnd cell_6t
Xbit_r38_c90 bl_90 br_90 wl_38 vdd gnd cell_6t
Xbit_r39_c90 bl_90 br_90 wl_39 vdd gnd cell_6t
Xbit_r40_c90 bl_90 br_90 wl_40 vdd gnd cell_6t
Xbit_r41_c90 bl_90 br_90 wl_41 vdd gnd cell_6t
Xbit_r42_c90 bl_90 br_90 wl_42 vdd gnd cell_6t
Xbit_r43_c90 bl_90 br_90 wl_43 vdd gnd cell_6t
Xbit_r44_c90 bl_90 br_90 wl_44 vdd gnd cell_6t
Xbit_r45_c90 bl_90 br_90 wl_45 vdd gnd cell_6t
Xbit_r46_c90 bl_90 br_90 wl_46 vdd gnd cell_6t
Xbit_r47_c90 bl_90 br_90 wl_47 vdd gnd cell_6t
Xbit_r48_c90 bl_90 br_90 wl_48 vdd gnd cell_6t
Xbit_r49_c90 bl_90 br_90 wl_49 vdd gnd cell_6t
Xbit_r50_c90 bl_90 br_90 wl_50 vdd gnd cell_6t
Xbit_r51_c90 bl_90 br_90 wl_51 vdd gnd cell_6t
Xbit_r52_c90 bl_90 br_90 wl_52 vdd gnd cell_6t
Xbit_r53_c90 bl_90 br_90 wl_53 vdd gnd cell_6t
Xbit_r54_c90 bl_90 br_90 wl_54 vdd gnd cell_6t
Xbit_r55_c90 bl_90 br_90 wl_55 vdd gnd cell_6t
Xbit_r56_c90 bl_90 br_90 wl_56 vdd gnd cell_6t
Xbit_r57_c90 bl_90 br_90 wl_57 vdd gnd cell_6t
Xbit_r58_c90 bl_90 br_90 wl_58 vdd gnd cell_6t
Xbit_r59_c90 bl_90 br_90 wl_59 vdd gnd cell_6t
Xbit_r60_c90 bl_90 br_90 wl_60 vdd gnd cell_6t
Xbit_r61_c90 bl_90 br_90 wl_61 vdd gnd cell_6t
Xbit_r62_c90 bl_90 br_90 wl_62 vdd gnd cell_6t
Xbit_r63_c90 bl_90 br_90 wl_63 vdd gnd cell_6t
Xbit_r64_c90 bl_90 br_90 wl_64 vdd gnd cell_6t
Xbit_r65_c90 bl_90 br_90 wl_65 vdd gnd cell_6t
Xbit_r66_c90 bl_90 br_90 wl_66 vdd gnd cell_6t
Xbit_r67_c90 bl_90 br_90 wl_67 vdd gnd cell_6t
Xbit_r68_c90 bl_90 br_90 wl_68 vdd gnd cell_6t
Xbit_r69_c90 bl_90 br_90 wl_69 vdd gnd cell_6t
Xbit_r70_c90 bl_90 br_90 wl_70 vdd gnd cell_6t
Xbit_r71_c90 bl_90 br_90 wl_71 vdd gnd cell_6t
Xbit_r72_c90 bl_90 br_90 wl_72 vdd gnd cell_6t
Xbit_r73_c90 bl_90 br_90 wl_73 vdd gnd cell_6t
Xbit_r74_c90 bl_90 br_90 wl_74 vdd gnd cell_6t
Xbit_r75_c90 bl_90 br_90 wl_75 vdd gnd cell_6t
Xbit_r76_c90 bl_90 br_90 wl_76 vdd gnd cell_6t
Xbit_r77_c90 bl_90 br_90 wl_77 vdd gnd cell_6t
Xbit_r78_c90 bl_90 br_90 wl_78 vdd gnd cell_6t
Xbit_r79_c90 bl_90 br_90 wl_79 vdd gnd cell_6t
Xbit_r80_c90 bl_90 br_90 wl_80 vdd gnd cell_6t
Xbit_r81_c90 bl_90 br_90 wl_81 vdd gnd cell_6t
Xbit_r82_c90 bl_90 br_90 wl_82 vdd gnd cell_6t
Xbit_r83_c90 bl_90 br_90 wl_83 vdd gnd cell_6t
Xbit_r84_c90 bl_90 br_90 wl_84 vdd gnd cell_6t
Xbit_r85_c90 bl_90 br_90 wl_85 vdd gnd cell_6t
Xbit_r86_c90 bl_90 br_90 wl_86 vdd gnd cell_6t
Xbit_r87_c90 bl_90 br_90 wl_87 vdd gnd cell_6t
Xbit_r88_c90 bl_90 br_90 wl_88 vdd gnd cell_6t
Xbit_r89_c90 bl_90 br_90 wl_89 vdd gnd cell_6t
Xbit_r90_c90 bl_90 br_90 wl_90 vdd gnd cell_6t
Xbit_r91_c90 bl_90 br_90 wl_91 vdd gnd cell_6t
Xbit_r92_c90 bl_90 br_90 wl_92 vdd gnd cell_6t
Xbit_r93_c90 bl_90 br_90 wl_93 vdd gnd cell_6t
Xbit_r94_c90 bl_90 br_90 wl_94 vdd gnd cell_6t
Xbit_r95_c90 bl_90 br_90 wl_95 vdd gnd cell_6t
Xbit_r96_c90 bl_90 br_90 wl_96 vdd gnd cell_6t
Xbit_r97_c90 bl_90 br_90 wl_97 vdd gnd cell_6t
Xbit_r98_c90 bl_90 br_90 wl_98 vdd gnd cell_6t
Xbit_r99_c90 bl_90 br_90 wl_99 vdd gnd cell_6t
Xbit_r100_c90 bl_90 br_90 wl_100 vdd gnd cell_6t
Xbit_r101_c90 bl_90 br_90 wl_101 vdd gnd cell_6t
Xbit_r102_c90 bl_90 br_90 wl_102 vdd gnd cell_6t
Xbit_r103_c90 bl_90 br_90 wl_103 vdd gnd cell_6t
Xbit_r104_c90 bl_90 br_90 wl_104 vdd gnd cell_6t
Xbit_r105_c90 bl_90 br_90 wl_105 vdd gnd cell_6t
Xbit_r106_c90 bl_90 br_90 wl_106 vdd gnd cell_6t
Xbit_r107_c90 bl_90 br_90 wl_107 vdd gnd cell_6t
Xbit_r108_c90 bl_90 br_90 wl_108 vdd gnd cell_6t
Xbit_r109_c90 bl_90 br_90 wl_109 vdd gnd cell_6t
Xbit_r110_c90 bl_90 br_90 wl_110 vdd gnd cell_6t
Xbit_r111_c90 bl_90 br_90 wl_111 vdd gnd cell_6t
Xbit_r112_c90 bl_90 br_90 wl_112 vdd gnd cell_6t
Xbit_r113_c90 bl_90 br_90 wl_113 vdd gnd cell_6t
Xbit_r114_c90 bl_90 br_90 wl_114 vdd gnd cell_6t
Xbit_r115_c90 bl_90 br_90 wl_115 vdd gnd cell_6t
Xbit_r116_c90 bl_90 br_90 wl_116 vdd gnd cell_6t
Xbit_r117_c90 bl_90 br_90 wl_117 vdd gnd cell_6t
Xbit_r118_c90 bl_90 br_90 wl_118 vdd gnd cell_6t
Xbit_r119_c90 bl_90 br_90 wl_119 vdd gnd cell_6t
Xbit_r120_c90 bl_90 br_90 wl_120 vdd gnd cell_6t
Xbit_r121_c90 bl_90 br_90 wl_121 vdd gnd cell_6t
Xbit_r122_c90 bl_90 br_90 wl_122 vdd gnd cell_6t
Xbit_r123_c90 bl_90 br_90 wl_123 vdd gnd cell_6t
Xbit_r124_c90 bl_90 br_90 wl_124 vdd gnd cell_6t
Xbit_r125_c90 bl_90 br_90 wl_125 vdd gnd cell_6t
Xbit_r126_c90 bl_90 br_90 wl_126 vdd gnd cell_6t
Xbit_r127_c90 bl_90 br_90 wl_127 vdd gnd cell_6t
Xbit_r128_c90 bl_90 br_90 wl_128 vdd gnd cell_6t
Xbit_r129_c90 bl_90 br_90 wl_129 vdd gnd cell_6t
Xbit_r130_c90 bl_90 br_90 wl_130 vdd gnd cell_6t
Xbit_r131_c90 bl_90 br_90 wl_131 vdd gnd cell_6t
Xbit_r132_c90 bl_90 br_90 wl_132 vdd gnd cell_6t
Xbit_r133_c90 bl_90 br_90 wl_133 vdd gnd cell_6t
Xbit_r134_c90 bl_90 br_90 wl_134 vdd gnd cell_6t
Xbit_r135_c90 bl_90 br_90 wl_135 vdd gnd cell_6t
Xbit_r136_c90 bl_90 br_90 wl_136 vdd gnd cell_6t
Xbit_r137_c90 bl_90 br_90 wl_137 vdd gnd cell_6t
Xbit_r138_c90 bl_90 br_90 wl_138 vdd gnd cell_6t
Xbit_r139_c90 bl_90 br_90 wl_139 vdd gnd cell_6t
Xbit_r140_c90 bl_90 br_90 wl_140 vdd gnd cell_6t
Xbit_r141_c90 bl_90 br_90 wl_141 vdd gnd cell_6t
Xbit_r142_c90 bl_90 br_90 wl_142 vdd gnd cell_6t
Xbit_r143_c90 bl_90 br_90 wl_143 vdd gnd cell_6t
Xbit_r144_c90 bl_90 br_90 wl_144 vdd gnd cell_6t
Xbit_r145_c90 bl_90 br_90 wl_145 vdd gnd cell_6t
Xbit_r146_c90 bl_90 br_90 wl_146 vdd gnd cell_6t
Xbit_r147_c90 bl_90 br_90 wl_147 vdd gnd cell_6t
Xbit_r148_c90 bl_90 br_90 wl_148 vdd gnd cell_6t
Xbit_r149_c90 bl_90 br_90 wl_149 vdd gnd cell_6t
Xbit_r150_c90 bl_90 br_90 wl_150 vdd gnd cell_6t
Xbit_r151_c90 bl_90 br_90 wl_151 vdd gnd cell_6t
Xbit_r152_c90 bl_90 br_90 wl_152 vdd gnd cell_6t
Xbit_r153_c90 bl_90 br_90 wl_153 vdd gnd cell_6t
Xbit_r154_c90 bl_90 br_90 wl_154 vdd gnd cell_6t
Xbit_r155_c90 bl_90 br_90 wl_155 vdd gnd cell_6t
Xbit_r156_c90 bl_90 br_90 wl_156 vdd gnd cell_6t
Xbit_r157_c90 bl_90 br_90 wl_157 vdd gnd cell_6t
Xbit_r158_c90 bl_90 br_90 wl_158 vdd gnd cell_6t
Xbit_r159_c90 bl_90 br_90 wl_159 vdd gnd cell_6t
Xbit_r160_c90 bl_90 br_90 wl_160 vdd gnd cell_6t
Xbit_r161_c90 bl_90 br_90 wl_161 vdd gnd cell_6t
Xbit_r162_c90 bl_90 br_90 wl_162 vdd gnd cell_6t
Xbit_r163_c90 bl_90 br_90 wl_163 vdd gnd cell_6t
Xbit_r164_c90 bl_90 br_90 wl_164 vdd gnd cell_6t
Xbit_r165_c90 bl_90 br_90 wl_165 vdd gnd cell_6t
Xbit_r166_c90 bl_90 br_90 wl_166 vdd gnd cell_6t
Xbit_r167_c90 bl_90 br_90 wl_167 vdd gnd cell_6t
Xbit_r168_c90 bl_90 br_90 wl_168 vdd gnd cell_6t
Xbit_r169_c90 bl_90 br_90 wl_169 vdd gnd cell_6t
Xbit_r170_c90 bl_90 br_90 wl_170 vdd gnd cell_6t
Xbit_r171_c90 bl_90 br_90 wl_171 vdd gnd cell_6t
Xbit_r172_c90 bl_90 br_90 wl_172 vdd gnd cell_6t
Xbit_r173_c90 bl_90 br_90 wl_173 vdd gnd cell_6t
Xbit_r174_c90 bl_90 br_90 wl_174 vdd gnd cell_6t
Xbit_r175_c90 bl_90 br_90 wl_175 vdd gnd cell_6t
Xbit_r176_c90 bl_90 br_90 wl_176 vdd gnd cell_6t
Xbit_r177_c90 bl_90 br_90 wl_177 vdd gnd cell_6t
Xbit_r178_c90 bl_90 br_90 wl_178 vdd gnd cell_6t
Xbit_r179_c90 bl_90 br_90 wl_179 vdd gnd cell_6t
Xbit_r180_c90 bl_90 br_90 wl_180 vdd gnd cell_6t
Xbit_r181_c90 bl_90 br_90 wl_181 vdd gnd cell_6t
Xbit_r182_c90 bl_90 br_90 wl_182 vdd gnd cell_6t
Xbit_r183_c90 bl_90 br_90 wl_183 vdd gnd cell_6t
Xbit_r184_c90 bl_90 br_90 wl_184 vdd gnd cell_6t
Xbit_r185_c90 bl_90 br_90 wl_185 vdd gnd cell_6t
Xbit_r186_c90 bl_90 br_90 wl_186 vdd gnd cell_6t
Xbit_r187_c90 bl_90 br_90 wl_187 vdd gnd cell_6t
Xbit_r188_c90 bl_90 br_90 wl_188 vdd gnd cell_6t
Xbit_r189_c90 bl_90 br_90 wl_189 vdd gnd cell_6t
Xbit_r190_c90 bl_90 br_90 wl_190 vdd gnd cell_6t
Xbit_r191_c90 bl_90 br_90 wl_191 vdd gnd cell_6t
Xbit_r192_c90 bl_90 br_90 wl_192 vdd gnd cell_6t
Xbit_r193_c90 bl_90 br_90 wl_193 vdd gnd cell_6t
Xbit_r194_c90 bl_90 br_90 wl_194 vdd gnd cell_6t
Xbit_r195_c90 bl_90 br_90 wl_195 vdd gnd cell_6t
Xbit_r196_c90 bl_90 br_90 wl_196 vdd gnd cell_6t
Xbit_r197_c90 bl_90 br_90 wl_197 vdd gnd cell_6t
Xbit_r198_c90 bl_90 br_90 wl_198 vdd gnd cell_6t
Xbit_r199_c90 bl_90 br_90 wl_199 vdd gnd cell_6t
Xbit_r200_c90 bl_90 br_90 wl_200 vdd gnd cell_6t
Xbit_r201_c90 bl_90 br_90 wl_201 vdd gnd cell_6t
Xbit_r202_c90 bl_90 br_90 wl_202 vdd gnd cell_6t
Xbit_r203_c90 bl_90 br_90 wl_203 vdd gnd cell_6t
Xbit_r204_c90 bl_90 br_90 wl_204 vdd gnd cell_6t
Xbit_r205_c90 bl_90 br_90 wl_205 vdd gnd cell_6t
Xbit_r206_c90 bl_90 br_90 wl_206 vdd gnd cell_6t
Xbit_r207_c90 bl_90 br_90 wl_207 vdd gnd cell_6t
Xbit_r208_c90 bl_90 br_90 wl_208 vdd gnd cell_6t
Xbit_r209_c90 bl_90 br_90 wl_209 vdd gnd cell_6t
Xbit_r210_c90 bl_90 br_90 wl_210 vdd gnd cell_6t
Xbit_r211_c90 bl_90 br_90 wl_211 vdd gnd cell_6t
Xbit_r212_c90 bl_90 br_90 wl_212 vdd gnd cell_6t
Xbit_r213_c90 bl_90 br_90 wl_213 vdd gnd cell_6t
Xbit_r214_c90 bl_90 br_90 wl_214 vdd gnd cell_6t
Xbit_r215_c90 bl_90 br_90 wl_215 vdd gnd cell_6t
Xbit_r216_c90 bl_90 br_90 wl_216 vdd gnd cell_6t
Xbit_r217_c90 bl_90 br_90 wl_217 vdd gnd cell_6t
Xbit_r218_c90 bl_90 br_90 wl_218 vdd gnd cell_6t
Xbit_r219_c90 bl_90 br_90 wl_219 vdd gnd cell_6t
Xbit_r220_c90 bl_90 br_90 wl_220 vdd gnd cell_6t
Xbit_r221_c90 bl_90 br_90 wl_221 vdd gnd cell_6t
Xbit_r222_c90 bl_90 br_90 wl_222 vdd gnd cell_6t
Xbit_r223_c90 bl_90 br_90 wl_223 vdd gnd cell_6t
Xbit_r224_c90 bl_90 br_90 wl_224 vdd gnd cell_6t
Xbit_r225_c90 bl_90 br_90 wl_225 vdd gnd cell_6t
Xbit_r226_c90 bl_90 br_90 wl_226 vdd gnd cell_6t
Xbit_r227_c90 bl_90 br_90 wl_227 vdd gnd cell_6t
Xbit_r228_c90 bl_90 br_90 wl_228 vdd gnd cell_6t
Xbit_r229_c90 bl_90 br_90 wl_229 vdd gnd cell_6t
Xbit_r230_c90 bl_90 br_90 wl_230 vdd gnd cell_6t
Xbit_r231_c90 bl_90 br_90 wl_231 vdd gnd cell_6t
Xbit_r232_c90 bl_90 br_90 wl_232 vdd gnd cell_6t
Xbit_r233_c90 bl_90 br_90 wl_233 vdd gnd cell_6t
Xbit_r234_c90 bl_90 br_90 wl_234 vdd gnd cell_6t
Xbit_r235_c90 bl_90 br_90 wl_235 vdd gnd cell_6t
Xbit_r236_c90 bl_90 br_90 wl_236 vdd gnd cell_6t
Xbit_r237_c90 bl_90 br_90 wl_237 vdd gnd cell_6t
Xbit_r238_c90 bl_90 br_90 wl_238 vdd gnd cell_6t
Xbit_r239_c90 bl_90 br_90 wl_239 vdd gnd cell_6t
Xbit_r240_c90 bl_90 br_90 wl_240 vdd gnd cell_6t
Xbit_r241_c90 bl_90 br_90 wl_241 vdd gnd cell_6t
Xbit_r242_c90 bl_90 br_90 wl_242 vdd gnd cell_6t
Xbit_r243_c90 bl_90 br_90 wl_243 vdd gnd cell_6t
Xbit_r244_c90 bl_90 br_90 wl_244 vdd gnd cell_6t
Xbit_r245_c90 bl_90 br_90 wl_245 vdd gnd cell_6t
Xbit_r246_c90 bl_90 br_90 wl_246 vdd gnd cell_6t
Xbit_r247_c90 bl_90 br_90 wl_247 vdd gnd cell_6t
Xbit_r248_c90 bl_90 br_90 wl_248 vdd gnd cell_6t
Xbit_r249_c90 bl_90 br_90 wl_249 vdd gnd cell_6t
Xbit_r250_c90 bl_90 br_90 wl_250 vdd gnd cell_6t
Xbit_r251_c90 bl_90 br_90 wl_251 vdd gnd cell_6t
Xbit_r252_c90 bl_90 br_90 wl_252 vdd gnd cell_6t
Xbit_r253_c90 bl_90 br_90 wl_253 vdd gnd cell_6t
Xbit_r254_c90 bl_90 br_90 wl_254 vdd gnd cell_6t
Xbit_r255_c90 bl_90 br_90 wl_255 vdd gnd cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd cell_6t
Xbit_r1_c91 bl_91 br_91 wl_1 vdd gnd cell_6t
Xbit_r2_c91 bl_91 br_91 wl_2 vdd gnd cell_6t
Xbit_r3_c91 bl_91 br_91 wl_3 vdd gnd cell_6t
Xbit_r4_c91 bl_91 br_91 wl_4 vdd gnd cell_6t
Xbit_r5_c91 bl_91 br_91 wl_5 vdd gnd cell_6t
Xbit_r6_c91 bl_91 br_91 wl_6 vdd gnd cell_6t
Xbit_r7_c91 bl_91 br_91 wl_7 vdd gnd cell_6t
Xbit_r8_c91 bl_91 br_91 wl_8 vdd gnd cell_6t
Xbit_r9_c91 bl_91 br_91 wl_9 vdd gnd cell_6t
Xbit_r10_c91 bl_91 br_91 wl_10 vdd gnd cell_6t
Xbit_r11_c91 bl_91 br_91 wl_11 vdd gnd cell_6t
Xbit_r12_c91 bl_91 br_91 wl_12 vdd gnd cell_6t
Xbit_r13_c91 bl_91 br_91 wl_13 vdd gnd cell_6t
Xbit_r14_c91 bl_91 br_91 wl_14 vdd gnd cell_6t
Xbit_r15_c91 bl_91 br_91 wl_15 vdd gnd cell_6t
Xbit_r16_c91 bl_91 br_91 wl_16 vdd gnd cell_6t
Xbit_r17_c91 bl_91 br_91 wl_17 vdd gnd cell_6t
Xbit_r18_c91 bl_91 br_91 wl_18 vdd gnd cell_6t
Xbit_r19_c91 bl_91 br_91 wl_19 vdd gnd cell_6t
Xbit_r20_c91 bl_91 br_91 wl_20 vdd gnd cell_6t
Xbit_r21_c91 bl_91 br_91 wl_21 vdd gnd cell_6t
Xbit_r22_c91 bl_91 br_91 wl_22 vdd gnd cell_6t
Xbit_r23_c91 bl_91 br_91 wl_23 vdd gnd cell_6t
Xbit_r24_c91 bl_91 br_91 wl_24 vdd gnd cell_6t
Xbit_r25_c91 bl_91 br_91 wl_25 vdd gnd cell_6t
Xbit_r26_c91 bl_91 br_91 wl_26 vdd gnd cell_6t
Xbit_r27_c91 bl_91 br_91 wl_27 vdd gnd cell_6t
Xbit_r28_c91 bl_91 br_91 wl_28 vdd gnd cell_6t
Xbit_r29_c91 bl_91 br_91 wl_29 vdd gnd cell_6t
Xbit_r30_c91 bl_91 br_91 wl_30 vdd gnd cell_6t
Xbit_r31_c91 bl_91 br_91 wl_31 vdd gnd cell_6t
Xbit_r32_c91 bl_91 br_91 wl_32 vdd gnd cell_6t
Xbit_r33_c91 bl_91 br_91 wl_33 vdd gnd cell_6t
Xbit_r34_c91 bl_91 br_91 wl_34 vdd gnd cell_6t
Xbit_r35_c91 bl_91 br_91 wl_35 vdd gnd cell_6t
Xbit_r36_c91 bl_91 br_91 wl_36 vdd gnd cell_6t
Xbit_r37_c91 bl_91 br_91 wl_37 vdd gnd cell_6t
Xbit_r38_c91 bl_91 br_91 wl_38 vdd gnd cell_6t
Xbit_r39_c91 bl_91 br_91 wl_39 vdd gnd cell_6t
Xbit_r40_c91 bl_91 br_91 wl_40 vdd gnd cell_6t
Xbit_r41_c91 bl_91 br_91 wl_41 vdd gnd cell_6t
Xbit_r42_c91 bl_91 br_91 wl_42 vdd gnd cell_6t
Xbit_r43_c91 bl_91 br_91 wl_43 vdd gnd cell_6t
Xbit_r44_c91 bl_91 br_91 wl_44 vdd gnd cell_6t
Xbit_r45_c91 bl_91 br_91 wl_45 vdd gnd cell_6t
Xbit_r46_c91 bl_91 br_91 wl_46 vdd gnd cell_6t
Xbit_r47_c91 bl_91 br_91 wl_47 vdd gnd cell_6t
Xbit_r48_c91 bl_91 br_91 wl_48 vdd gnd cell_6t
Xbit_r49_c91 bl_91 br_91 wl_49 vdd gnd cell_6t
Xbit_r50_c91 bl_91 br_91 wl_50 vdd gnd cell_6t
Xbit_r51_c91 bl_91 br_91 wl_51 vdd gnd cell_6t
Xbit_r52_c91 bl_91 br_91 wl_52 vdd gnd cell_6t
Xbit_r53_c91 bl_91 br_91 wl_53 vdd gnd cell_6t
Xbit_r54_c91 bl_91 br_91 wl_54 vdd gnd cell_6t
Xbit_r55_c91 bl_91 br_91 wl_55 vdd gnd cell_6t
Xbit_r56_c91 bl_91 br_91 wl_56 vdd gnd cell_6t
Xbit_r57_c91 bl_91 br_91 wl_57 vdd gnd cell_6t
Xbit_r58_c91 bl_91 br_91 wl_58 vdd gnd cell_6t
Xbit_r59_c91 bl_91 br_91 wl_59 vdd gnd cell_6t
Xbit_r60_c91 bl_91 br_91 wl_60 vdd gnd cell_6t
Xbit_r61_c91 bl_91 br_91 wl_61 vdd gnd cell_6t
Xbit_r62_c91 bl_91 br_91 wl_62 vdd gnd cell_6t
Xbit_r63_c91 bl_91 br_91 wl_63 vdd gnd cell_6t
Xbit_r64_c91 bl_91 br_91 wl_64 vdd gnd cell_6t
Xbit_r65_c91 bl_91 br_91 wl_65 vdd gnd cell_6t
Xbit_r66_c91 bl_91 br_91 wl_66 vdd gnd cell_6t
Xbit_r67_c91 bl_91 br_91 wl_67 vdd gnd cell_6t
Xbit_r68_c91 bl_91 br_91 wl_68 vdd gnd cell_6t
Xbit_r69_c91 bl_91 br_91 wl_69 vdd gnd cell_6t
Xbit_r70_c91 bl_91 br_91 wl_70 vdd gnd cell_6t
Xbit_r71_c91 bl_91 br_91 wl_71 vdd gnd cell_6t
Xbit_r72_c91 bl_91 br_91 wl_72 vdd gnd cell_6t
Xbit_r73_c91 bl_91 br_91 wl_73 vdd gnd cell_6t
Xbit_r74_c91 bl_91 br_91 wl_74 vdd gnd cell_6t
Xbit_r75_c91 bl_91 br_91 wl_75 vdd gnd cell_6t
Xbit_r76_c91 bl_91 br_91 wl_76 vdd gnd cell_6t
Xbit_r77_c91 bl_91 br_91 wl_77 vdd gnd cell_6t
Xbit_r78_c91 bl_91 br_91 wl_78 vdd gnd cell_6t
Xbit_r79_c91 bl_91 br_91 wl_79 vdd gnd cell_6t
Xbit_r80_c91 bl_91 br_91 wl_80 vdd gnd cell_6t
Xbit_r81_c91 bl_91 br_91 wl_81 vdd gnd cell_6t
Xbit_r82_c91 bl_91 br_91 wl_82 vdd gnd cell_6t
Xbit_r83_c91 bl_91 br_91 wl_83 vdd gnd cell_6t
Xbit_r84_c91 bl_91 br_91 wl_84 vdd gnd cell_6t
Xbit_r85_c91 bl_91 br_91 wl_85 vdd gnd cell_6t
Xbit_r86_c91 bl_91 br_91 wl_86 vdd gnd cell_6t
Xbit_r87_c91 bl_91 br_91 wl_87 vdd gnd cell_6t
Xbit_r88_c91 bl_91 br_91 wl_88 vdd gnd cell_6t
Xbit_r89_c91 bl_91 br_91 wl_89 vdd gnd cell_6t
Xbit_r90_c91 bl_91 br_91 wl_90 vdd gnd cell_6t
Xbit_r91_c91 bl_91 br_91 wl_91 vdd gnd cell_6t
Xbit_r92_c91 bl_91 br_91 wl_92 vdd gnd cell_6t
Xbit_r93_c91 bl_91 br_91 wl_93 vdd gnd cell_6t
Xbit_r94_c91 bl_91 br_91 wl_94 vdd gnd cell_6t
Xbit_r95_c91 bl_91 br_91 wl_95 vdd gnd cell_6t
Xbit_r96_c91 bl_91 br_91 wl_96 vdd gnd cell_6t
Xbit_r97_c91 bl_91 br_91 wl_97 vdd gnd cell_6t
Xbit_r98_c91 bl_91 br_91 wl_98 vdd gnd cell_6t
Xbit_r99_c91 bl_91 br_91 wl_99 vdd gnd cell_6t
Xbit_r100_c91 bl_91 br_91 wl_100 vdd gnd cell_6t
Xbit_r101_c91 bl_91 br_91 wl_101 vdd gnd cell_6t
Xbit_r102_c91 bl_91 br_91 wl_102 vdd gnd cell_6t
Xbit_r103_c91 bl_91 br_91 wl_103 vdd gnd cell_6t
Xbit_r104_c91 bl_91 br_91 wl_104 vdd gnd cell_6t
Xbit_r105_c91 bl_91 br_91 wl_105 vdd gnd cell_6t
Xbit_r106_c91 bl_91 br_91 wl_106 vdd gnd cell_6t
Xbit_r107_c91 bl_91 br_91 wl_107 vdd gnd cell_6t
Xbit_r108_c91 bl_91 br_91 wl_108 vdd gnd cell_6t
Xbit_r109_c91 bl_91 br_91 wl_109 vdd gnd cell_6t
Xbit_r110_c91 bl_91 br_91 wl_110 vdd gnd cell_6t
Xbit_r111_c91 bl_91 br_91 wl_111 vdd gnd cell_6t
Xbit_r112_c91 bl_91 br_91 wl_112 vdd gnd cell_6t
Xbit_r113_c91 bl_91 br_91 wl_113 vdd gnd cell_6t
Xbit_r114_c91 bl_91 br_91 wl_114 vdd gnd cell_6t
Xbit_r115_c91 bl_91 br_91 wl_115 vdd gnd cell_6t
Xbit_r116_c91 bl_91 br_91 wl_116 vdd gnd cell_6t
Xbit_r117_c91 bl_91 br_91 wl_117 vdd gnd cell_6t
Xbit_r118_c91 bl_91 br_91 wl_118 vdd gnd cell_6t
Xbit_r119_c91 bl_91 br_91 wl_119 vdd gnd cell_6t
Xbit_r120_c91 bl_91 br_91 wl_120 vdd gnd cell_6t
Xbit_r121_c91 bl_91 br_91 wl_121 vdd gnd cell_6t
Xbit_r122_c91 bl_91 br_91 wl_122 vdd gnd cell_6t
Xbit_r123_c91 bl_91 br_91 wl_123 vdd gnd cell_6t
Xbit_r124_c91 bl_91 br_91 wl_124 vdd gnd cell_6t
Xbit_r125_c91 bl_91 br_91 wl_125 vdd gnd cell_6t
Xbit_r126_c91 bl_91 br_91 wl_126 vdd gnd cell_6t
Xbit_r127_c91 bl_91 br_91 wl_127 vdd gnd cell_6t
Xbit_r128_c91 bl_91 br_91 wl_128 vdd gnd cell_6t
Xbit_r129_c91 bl_91 br_91 wl_129 vdd gnd cell_6t
Xbit_r130_c91 bl_91 br_91 wl_130 vdd gnd cell_6t
Xbit_r131_c91 bl_91 br_91 wl_131 vdd gnd cell_6t
Xbit_r132_c91 bl_91 br_91 wl_132 vdd gnd cell_6t
Xbit_r133_c91 bl_91 br_91 wl_133 vdd gnd cell_6t
Xbit_r134_c91 bl_91 br_91 wl_134 vdd gnd cell_6t
Xbit_r135_c91 bl_91 br_91 wl_135 vdd gnd cell_6t
Xbit_r136_c91 bl_91 br_91 wl_136 vdd gnd cell_6t
Xbit_r137_c91 bl_91 br_91 wl_137 vdd gnd cell_6t
Xbit_r138_c91 bl_91 br_91 wl_138 vdd gnd cell_6t
Xbit_r139_c91 bl_91 br_91 wl_139 vdd gnd cell_6t
Xbit_r140_c91 bl_91 br_91 wl_140 vdd gnd cell_6t
Xbit_r141_c91 bl_91 br_91 wl_141 vdd gnd cell_6t
Xbit_r142_c91 bl_91 br_91 wl_142 vdd gnd cell_6t
Xbit_r143_c91 bl_91 br_91 wl_143 vdd gnd cell_6t
Xbit_r144_c91 bl_91 br_91 wl_144 vdd gnd cell_6t
Xbit_r145_c91 bl_91 br_91 wl_145 vdd gnd cell_6t
Xbit_r146_c91 bl_91 br_91 wl_146 vdd gnd cell_6t
Xbit_r147_c91 bl_91 br_91 wl_147 vdd gnd cell_6t
Xbit_r148_c91 bl_91 br_91 wl_148 vdd gnd cell_6t
Xbit_r149_c91 bl_91 br_91 wl_149 vdd gnd cell_6t
Xbit_r150_c91 bl_91 br_91 wl_150 vdd gnd cell_6t
Xbit_r151_c91 bl_91 br_91 wl_151 vdd gnd cell_6t
Xbit_r152_c91 bl_91 br_91 wl_152 vdd gnd cell_6t
Xbit_r153_c91 bl_91 br_91 wl_153 vdd gnd cell_6t
Xbit_r154_c91 bl_91 br_91 wl_154 vdd gnd cell_6t
Xbit_r155_c91 bl_91 br_91 wl_155 vdd gnd cell_6t
Xbit_r156_c91 bl_91 br_91 wl_156 vdd gnd cell_6t
Xbit_r157_c91 bl_91 br_91 wl_157 vdd gnd cell_6t
Xbit_r158_c91 bl_91 br_91 wl_158 vdd gnd cell_6t
Xbit_r159_c91 bl_91 br_91 wl_159 vdd gnd cell_6t
Xbit_r160_c91 bl_91 br_91 wl_160 vdd gnd cell_6t
Xbit_r161_c91 bl_91 br_91 wl_161 vdd gnd cell_6t
Xbit_r162_c91 bl_91 br_91 wl_162 vdd gnd cell_6t
Xbit_r163_c91 bl_91 br_91 wl_163 vdd gnd cell_6t
Xbit_r164_c91 bl_91 br_91 wl_164 vdd gnd cell_6t
Xbit_r165_c91 bl_91 br_91 wl_165 vdd gnd cell_6t
Xbit_r166_c91 bl_91 br_91 wl_166 vdd gnd cell_6t
Xbit_r167_c91 bl_91 br_91 wl_167 vdd gnd cell_6t
Xbit_r168_c91 bl_91 br_91 wl_168 vdd gnd cell_6t
Xbit_r169_c91 bl_91 br_91 wl_169 vdd gnd cell_6t
Xbit_r170_c91 bl_91 br_91 wl_170 vdd gnd cell_6t
Xbit_r171_c91 bl_91 br_91 wl_171 vdd gnd cell_6t
Xbit_r172_c91 bl_91 br_91 wl_172 vdd gnd cell_6t
Xbit_r173_c91 bl_91 br_91 wl_173 vdd gnd cell_6t
Xbit_r174_c91 bl_91 br_91 wl_174 vdd gnd cell_6t
Xbit_r175_c91 bl_91 br_91 wl_175 vdd gnd cell_6t
Xbit_r176_c91 bl_91 br_91 wl_176 vdd gnd cell_6t
Xbit_r177_c91 bl_91 br_91 wl_177 vdd gnd cell_6t
Xbit_r178_c91 bl_91 br_91 wl_178 vdd gnd cell_6t
Xbit_r179_c91 bl_91 br_91 wl_179 vdd gnd cell_6t
Xbit_r180_c91 bl_91 br_91 wl_180 vdd gnd cell_6t
Xbit_r181_c91 bl_91 br_91 wl_181 vdd gnd cell_6t
Xbit_r182_c91 bl_91 br_91 wl_182 vdd gnd cell_6t
Xbit_r183_c91 bl_91 br_91 wl_183 vdd gnd cell_6t
Xbit_r184_c91 bl_91 br_91 wl_184 vdd gnd cell_6t
Xbit_r185_c91 bl_91 br_91 wl_185 vdd gnd cell_6t
Xbit_r186_c91 bl_91 br_91 wl_186 vdd gnd cell_6t
Xbit_r187_c91 bl_91 br_91 wl_187 vdd gnd cell_6t
Xbit_r188_c91 bl_91 br_91 wl_188 vdd gnd cell_6t
Xbit_r189_c91 bl_91 br_91 wl_189 vdd gnd cell_6t
Xbit_r190_c91 bl_91 br_91 wl_190 vdd gnd cell_6t
Xbit_r191_c91 bl_91 br_91 wl_191 vdd gnd cell_6t
Xbit_r192_c91 bl_91 br_91 wl_192 vdd gnd cell_6t
Xbit_r193_c91 bl_91 br_91 wl_193 vdd gnd cell_6t
Xbit_r194_c91 bl_91 br_91 wl_194 vdd gnd cell_6t
Xbit_r195_c91 bl_91 br_91 wl_195 vdd gnd cell_6t
Xbit_r196_c91 bl_91 br_91 wl_196 vdd gnd cell_6t
Xbit_r197_c91 bl_91 br_91 wl_197 vdd gnd cell_6t
Xbit_r198_c91 bl_91 br_91 wl_198 vdd gnd cell_6t
Xbit_r199_c91 bl_91 br_91 wl_199 vdd gnd cell_6t
Xbit_r200_c91 bl_91 br_91 wl_200 vdd gnd cell_6t
Xbit_r201_c91 bl_91 br_91 wl_201 vdd gnd cell_6t
Xbit_r202_c91 bl_91 br_91 wl_202 vdd gnd cell_6t
Xbit_r203_c91 bl_91 br_91 wl_203 vdd gnd cell_6t
Xbit_r204_c91 bl_91 br_91 wl_204 vdd gnd cell_6t
Xbit_r205_c91 bl_91 br_91 wl_205 vdd gnd cell_6t
Xbit_r206_c91 bl_91 br_91 wl_206 vdd gnd cell_6t
Xbit_r207_c91 bl_91 br_91 wl_207 vdd gnd cell_6t
Xbit_r208_c91 bl_91 br_91 wl_208 vdd gnd cell_6t
Xbit_r209_c91 bl_91 br_91 wl_209 vdd gnd cell_6t
Xbit_r210_c91 bl_91 br_91 wl_210 vdd gnd cell_6t
Xbit_r211_c91 bl_91 br_91 wl_211 vdd gnd cell_6t
Xbit_r212_c91 bl_91 br_91 wl_212 vdd gnd cell_6t
Xbit_r213_c91 bl_91 br_91 wl_213 vdd gnd cell_6t
Xbit_r214_c91 bl_91 br_91 wl_214 vdd gnd cell_6t
Xbit_r215_c91 bl_91 br_91 wl_215 vdd gnd cell_6t
Xbit_r216_c91 bl_91 br_91 wl_216 vdd gnd cell_6t
Xbit_r217_c91 bl_91 br_91 wl_217 vdd gnd cell_6t
Xbit_r218_c91 bl_91 br_91 wl_218 vdd gnd cell_6t
Xbit_r219_c91 bl_91 br_91 wl_219 vdd gnd cell_6t
Xbit_r220_c91 bl_91 br_91 wl_220 vdd gnd cell_6t
Xbit_r221_c91 bl_91 br_91 wl_221 vdd gnd cell_6t
Xbit_r222_c91 bl_91 br_91 wl_222 vdd gnd cell_6t
Xbit_r223_c91 bl_91 br_91 wl_223 vdd gnd cell_6t
Xbit_r224_c91 bl_91 br_91 wl_224 vdd gnd cell_6t
Xbit_r225_c91 bl_91 br_91 wl_225 vdd gnd cell_6t
Xbit_r226_c91 bl_91 br_91 wl_226 vdd gnd cell_6t
Xbit_r227_c91 bl_91 br_91 wl_227 vdd gnd cell_6t
Xbit_r228_c91 bl_91 br_91 wl_228 vdd gnd cell_6t
Xbit_r229_c91 bl_91 br_91 wl_229 vdd gnd cell_6t
Xbit_r230_c91 bl_91 br_91 wl_230 vdd gnd cell_6t
Xbit_r231_c91 bl_91 br_91 wl_231 vdd gnd cell_6t
Xbit_r232_c91 bl_91 br_91 wl_232 vdd gnd cell_6t
Xbit_r233_c91 bl_91 br_91 wl_233 vdd gnd cell_6t
Xbit_r234_c91 bl_91 br_91 wl_234 vdd gnd cell_6t
Xbit_r235_c91 bl_91 br_91 wl_235 vdd gnd cell_6t
Xbit_r236_c91 bl_91 br_91 wl_236 vdd gnd cell_6t
Xbit_r237_c91 bl_91 br_91 wl_237 vdd gnd cell_6t
Xbit_r238_c91 bl_91 br_91 wl_238 vdd gnd cell_6t
Xbit_r239_c91 bl_91 br_91 wl_239 vdd gnd cell_6t
Xbit_r240_c91 bl_91 br_91 wl_240 vdd gnd cell_6t
Xbit_r241_c91 bl_91 br_91 wl_241 vdd gnd cell_6t
Xbit_r242_c91 bl_91 br_91 wl_242 vdd gnd cell_6t
Xbit_r243_c91 bl_91 br_91 wl_243 vdd gnd cell_6t
Xbit_r244_c91 bl_91 br_91 wl_244 vdd gnd cell_6t
Xbit_r245_c91 bl_91 br_91 wl_245 vdd gnd cell_6t
Xbit_r246_c91 bl_91 br_91 wl_246 vdd gnd cell_6t
Xbit_r247_c91 bl_91 br_91 wl_247 vdd gnd cell_6t
Xbit_r248_c91 bl_91 br_91 wl_248 vdd gnd cell_6t
Xbit_r249_c91 bl_91 br_91 wl_249 vdd gnd cell_6t
Xbit_r250_c91 bl_91 br_91 wl_250 vdd gnd cell_6t
Xbit_r251_c91 bl_91 br_91 wl_251 vdd gnd cell_6t
Xbit_r252_c91 bl_91 br_91 wl_252 vdd gnd cell_6t
Xbit_r253_c91 bl_91 br_91 wl_253 vdd gnd cell_6t
Xbit_r254_c91 bl_91 br_91 wl_254 vdd gnd cell_6t
Xbit_r255_c91 bl_91 br_91 wl_255 vdd gnd cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd cell_6t
Xbit_r1_c92 bl_92 br_92 wl_1 vdd gnd cell_6t
Xbit_r2_c92 bl_92 br_92 wl_2 vdd gnd cell_6t
Xbit_r3_c92 bl_92 br_92 wl_3 vdd gnd cell_6t
Xbit_r4_c92 bl_92 br_92 wl_4 vdd gnd cell_6t
Xbit_r5_c92 bl_92 br_92 wl_5 vdd gnd cell_6t
Xbit_r6_c92 bl_92 br_92 wl_6 vdd gnd cell_6t
Xbit_r7_c92 bl_92 br_92 wl_7 vdd gnd cell_6t
Xbit_r8_c92 bl_92 br_92 wl_8 vdd gnd cell_6t
Xbit_r9_c92 bl_92 br_92 wl_9 vdd gnd cell_6t
Xbit_r10_c92 bl_92 br_92 wl_10 vdd gnd cell_6t
Xbit_r11_c92 bl_92 br_92 wl_11 vdd gnd cell_6t
Xbit_r12_c92 bl_92 br_92 wl_12 vdd gnd cell_6t
Xbit_r13_c92 bl_92 br_92 wl_13 vdd gnd cell_6t
Xbit_r14_c92 bl_92 br_92 wl_14 vdd gnd cell_6t
Xbit_r15_c92 bl_92 br_92 wl_15 vdd gnd cell_6t
Xbit_r16_c92 bl_92 br_92 wl_16 vdd gnd cell_6t
Xbit_r17_c92 bl_92 br_92 wl_17 vdd gnd cell_6t
Xbit_r18_c92 bl_92 br_92 wl_18 vdd gnd cell_6t
Xbit_r19_c92 bl_92 br_92 wl_19 vdd gnd cell_6t
Xbit_r20_c92 bl_92 br_92 wl_20 vdd gnd cell_6t
Xbit_r21_c92 bl_92 br_92 wl_21 vdd gnd cell_6t
Xbit_r22_c92 bl_92 br_92 wl_22 vdd gnd cell_6t
Xbit_r23_c92 bl_92 br_92 wl_23 vdd gnd cell_6t
Xbit_r24_c92 bl_92 br_92 wl_24 vdd gnd cell_6t
Xbit_r25_c92 bl_92 br_92 wl_25 vdd gnd cell_6t
Xbit_r26_c92 bl_92 br_92 wl_26 vdd gnd cell_6t
Xbit_r27_c92 bl_92 br_92 wl_27 vdd gnd cell_6t
Xbit_r28_c92 bl_92 br_92 wl_28 vdd gnd cell_6t
Xbit_r29_c92 bl_92 br_92 wl_29 vdd gnd cell_6t
Xbit_r30_c92 bl_92 br_92 wl_30 vdd gnd cell_6t
Xbit_r31_c92 bl_92 br_92 wl_31 vdd gnd cell_6t
Xbit_r32_c92 bl_92 br_92 wl_32 vdd gnd cell_6t
Xbit_r33_c92 bl_92 br_92 wl_33 vdd gnd cell_6t
Xbit_r34_c92 bl_92 br_92 wl_34 vdd gnd cell_6t
Xbit_r35_c92 bl_92 br_92 wl_35 vdd gnd cell_6t
Xbit_r36_c92 bl_92 br_92 wl_36 vdd gnd cell_6t
Xbit_r37_c92 bl_92 br_92 wl_37 vdd gnd cell_6t
Xbit_r38_c92 bl_92 br_92 wl_38 vdd gnd cell_6t
Xbit_r39_c92 bl_92 br_92 wl_39 vdd gnd cell_6t
Xbit_r40_c92 bl_92 br_92 wl_40 vdd gnd cell_6t
Xbit_r41_c92 bl_92 br_92 wl_41 vdd gnd cell_6t
Xbit_r42_c92 bl_92 br_92 wl_42 vdd gnd cell_6t
Xbit_r43_c92 bl_92 br_92 wl_43 vdd gnd cell_6t
Xbit_r44_c92 bl_92 br_92 wl_44 vdd gnd cell_6t
Xbit_r45_c92 bl_92 br_92 wl_45 vdd gnd cell_6t
Xbit_r46_c92 bl_92 br_92 wl_46 vdd gnd cell_6t
Xbit_r47_c92 bl_92 br_92 wl_47 vdd gnd cell_6t
Xbit_r48_c92 bl_92 br_92 wl_48 vdd gnd cell_6t
Xbit_r49_c92 bl_92 br_92 wl_49 vdd gnd cell_6t
Xbit_r50_c92 bl_92 br_92 wl_50 vdd gnd cell_6t
Xbit_r51_c92 bl_92 br_92 wl_51 vdd gnd cell_6t
Xbit_r52_c92 bl_92 br_92 wl_52 vdd gnd cell_6t
Xbit_r53_c92 bl_92 br_92 wl_53 vdd gnd cell_6t
Xbit_r54_c92 bl_92 br_92 wl_54 vdd gnd cell_6t
Xbit_r55_c92 bl_92 br_92 wl_55 vdd gnd cell_6t
Xbit_r56_c92 bl_92 br_92 wl_56 vdd gnd cell_6t
Xbit_r57_c92 bl_92 br_92 wl_57 vdd gnd cell_6t
Xbit_r58_c92 bl_92 br_92 wl_58 vdd gnd cell_6t
Xbit_r59_c92 bl_92 br_92 wl_59 vdd gnd cell_6t
Xbit_r60_c92 bl_92 br_92 wl_60 vdd gnd cell_6t
Xbit_r61_c92 bl_92 br_92 wl_61 vdd gnd cell_6t
Xbit_r62_c92 bl_92 br_92 wl_62 vdd gnd cell_6t
Xbit_r63_c92 bl_92 br_92 wl_63 vdd gnd cell_6t
Xbit_r64_c92 bl_92 br_92 wl_64 vdd gnd cell_6t
Xbit_r65_c92 bl_92 br_92 wl_65 vdd gnd cell_6t
Xbit_r66_c92 bl_92 br_92 wl_66 vdd gnd cell_6t
Xbit_r67_c92 bl_92 br_92 wl_67 vdd gnd cell_6t
Xbit_r68_c92 bl_92 br_92 wl_68 vdd gnd cell_6t
Xbit_r69_c92 bl_92 br_92 wl_69 vdd gnd cell_6t
Xbit_r70_c92 bl_92 br_92 wl_70 vdd gnd cell_6t
Xbit_r71_c92 bl_92 br_92 wl_71 vdd gnd cell_6t
Xbit_r72_c92 bl_92 br_92 wl_72 vdd gnd cell_6t
Xbit_r73_c92 bl_92 br_92 wl_73 vdd gnd cell_6t
Xbit_r74_c92 bl_92 br_92 wl_74 vdd gnd cell_6t
Xbit_r75_c92 bl_92 br_92 wl_75 vdd gnd cell_6t
Xbit_r76_c92 bl_92 br_92 wl_76 vdd gnd cell_6t
Xbit_r77_c92 bl_92 br_92 wl_77 vdd gnd cell_6t
Xbit_r78_c92 bl_92 br_92 wl_78 vdd gnd cell_6t
Xbit_r79_c92 bl_92 br_92 wl_79 vdd gnd cell_6t
Xbit_r80_c92 bl_92 br_92 wl_80 vdd gnd cell_6t
Xbit_r81_c92 bl_92 br_92 wl_81 vdd gnd cell_6t
Xbit_r82_c92 bl_92 br_92 wl_82 vdd gnd cell_6t
Xbit_r83_c92 bl_92 br_92 wl_83 vdd gnd cell_6t
Xbit_r84_c92 bl_92 br_92 wl_84 vdd gnd cell_6t
Xbit_r85_c92 bl_92 br_92 wl_85 vdd gnd cell_6t
Xbit_r86_c92 bl_92 br_92 wl_86 vdd gnd cell_6t
Xbit_r87_c92 bl_92 br_92 wl_87 vdd gnd cell_6t
Xbit_r88_c92 bl_92 br_92 wl_88 vdd gnd cell_6t
Xbit_r89_c92 bl_92 br_92 wl_89 vdd gnd cell_6t
Xbit_r90_c92 bl_92 br_92 wl_90 vdd gnd cell_6t
Xbit_r91_c92 bl_92 br_92 wl_91 vdd gnd cell_6t
Xbit_r92_c92 bl_92 br_92 wl_92 vdd gnd cell_6t
Xbit_r93_c92 bl_92 br_92 wl_93 vdd gnd cell_6t
Xbit_r94_c92 bl_92 br_92 wl_94 vdd gnd cell_6t
Xbit_r95_c92 bl_92 br_92 wl_95 vdd gnd cell_6t
Xbit_r96_c92 bl_92 br_92 wl_96 vdd gnd cell_6t
Xbit_r97_c92 bl_92 br_92 wl_97 vdd gnd cell_6t
Xbit_r98_c92 bl_92 br_92 wl_98 vdd gnd cell_6t
Xbit_r99_c92 bl_92 br_92 wl_99 vdd gnd cell_6t
Xbit_r100_c92 bl_92 br_92 wl_100 vdd gnd cell_6t
Xbit_r101_c92 bl_92 br_92 wl_101 vdd gnd cell_6t
Xbit_r102_c92 bl_92 br_92 wl_102 vdd gnd cell_6t
Xbit_r103_c92 bl_92 br_92 wl_103 vdd gnd cell_6t
Xbit_r104_c92 bl_92 br_92 wl_104 vdd gnd cell_6t
Xbit_r105_c92 bl_92 br_92 wl_105 vdd gnd cell_6t
Xbit_r106_c92 bl_92 br_92 wl_106 vdd gnd cell_6t
Xbit_r107_c92 bl_92 br_92 wl_107 vdd gnd cell_6t
Xbit_r108_c92 bl_92 br_92 wl_108 vdd gnd cell_6t
Xbit_r109_c92 bl_92 br_92 wl_109 vdd gnd cell_6t
Xbit_r110_c92 bl_92 br_92 wl_110 vdd gnd cell_6t
Xbit_r111_c92 bl_92 br_92 wl_111 vdd gnd cell_6t
Xbit_r112_c92 bl_92 br_92 wl_112 vdd gnd cell_6t
Xbit_r113_c92 bl_92 br_92 wl_113 vdd gnd cell_6t
Xbit_r114_c92 bl_92 br_92 wl_114 vdd gnd cell_6t
Xbit_r115_c92 bl_92 br_92 wl_115 vdd gnd cell_6t
Xbit_r116_c92 bl_92 br_92 wl_116 vdd gnd cell_6t
Xbit_r117_c92 bl_92 br_92 wl_117 vdd gnd cell_6t
Xbit_r118_c92 bl_92 br_92 wl_118 vdd gnd cell_6t
Xbit_r119_c92 bl_92 br_92 wl_119 vdd gnd cell_6t
Xbit_r120_c92 bl_92 br_92 wl_120 vdd gnd cell_6t
Xbit_r121_c92 bl_92 br_92 wl_121 vdd gnd cell_6t
Xbit_r122_c92 bl_92 br_92 wl_122 vdd gnd cell_6t
Xbit_r123_c92 bl_92 br_92 wl_123 vdd gnd cell_6t
Xbit_r124_c92 bl_92 br_92 wl_124 vdd gnd cell_6t
Xbit_r125_c92 bl_92 br_92 wl_125 vdd gnd cell_6t
Xbit_r126_c92 bl_92 br_92 wl_126 vdd gnd cell_6t
Xbit_r127_c92 bl_92 br_92 wl_127 vdd gnd cell_6t
Xbit_r128_c92 bl_92 br_92 wl_128 vdd gnd cell_6t
Xbit_r129_c92 bl_92 br_92 wl_129 vdd gnd cell_6t
Xbit_r130_c92 bl_92 br_92 wl_130 vdd gnd cell_6t
Xbit_r131_c92 bl_92 br_92 wl_131 vdd gnd cell_6t
Xbit_r132_c92 bl_92 br_92 wl_132 vdd gnd cell_6t
Xbit_r133_c92 bl_92 br_92 wl_133 vdd gnd cell_6t
Xbit_r134_c92 bl_92 br_92 wl_134 vdd gnd cell_6t
Xbit_r135_c92 bl_92 br_92 wl_135 vdd gnd cell_6t
Xbit_r136_c92 bl_92 br_92 wl_136 vdd gnd cell_6t
Xbit_r137_c92 bl_92 br_92 wl_137 vdd gnd cell_6t
Xbit_r138_c92 bl_92 br_92 wl_138 vdd gnd cell_6t
Xbit_r139_c92 bl_92 br_92 wl_139 vdd gnd cell_6t
Xbit_r140_c92 bl_92 br_92 wl_140 vdd gnd cell_6t
Xbit_r141_c92 bl_92 br_92 wl_141 vdd gnd cell_6t
Xbit_r142_c92 bl_92 br_92 wl_142 vdd gnd cell_6t
Xbit_r143_c92 bl_92 br_92 wl_143 vdd gnd cell_6t
Xbit_r144_c92 bl_92 br_92 wl_144 vdd gnd cell_6t
Xbit_r145_c92 bl_92 br_92 wl_145 vdd gnd cell_6t
Xbit_r146_c92 bl_92 br_92 wl_146 vdd gnd cell_6t
Xbit_r147_c92 bl_92 br_92 wl_147 vdd gnd cell_6t
Xbit_r148_c92 bl_92 br_92 wl_148 vdd gnd cell_6t
Xbit_r149_c92 bl_92 br_92 wl_149 vdd gnd cell_6t
Xbit_r150_c92 bl_92 br_92 wl_150 vdd gnd cell_6t
Xbit_r151_c92 bl_92 br_92 wl_151 vdd gnd cell_6t
Xbit_r152_c92 bl_92 br_92 wl_152 vdd gnd cell_6t
Xbit_r153_c92 bl_92 br_92 wl_153 vdd gnd cell_6t
Xbit_r154_c92 bl_92 br_92 wl_154 vdd gnd cell_6t
Xbit_r155_c92 bl_92 br_92 wl_155 vdd gnd cell_6t
Xbit_r156_c92 bl_92 br_92 wl_156 vdd gnd cell_6t
Xbit_r157_c92 bl_92 br_92 wl_157 vdd gnd cell_6t
Xbit_r158_c92 bl_92 br_92 wl_158 vdd gnd cell_6t
Xbit_r159_c92 bl_92 br_92 wl_159 vdd gnd cell_6t
Xbit_r160_c92 bl_92 br_92 wl_160 vdd gnd cell_6t
Xbit_r161_c92 bl_92 br_92 wl_161 vdd gnd cell_6t
Xbit_r162_c92 bl_92 br_92 wl_162 vdd gnd cell_6t
Xbit_r163_c92 bl_92 br_92 wl_163 vdd gnd cell_6t
Xbit_r164_c92 bl_92 br_92 wl_164 vdd gnd cell_6t
Xbit_r165_c92 bl_92 br_92 wl_165 vdd gnd cell_6t
Xbit_r166_c92 bl_92 br_92 wl_166 vdd gnd cell_6t
Xbit_r167_c92 bl_92 br_92 wl_167 vdd gnd cell_6t
Xbit_r168_c92 bl_92 br_92 wl_168 vdd gnd cell_6t
Xbit_r169_c92 bl_92 br_92 wl_169 vdd gnd cell_6t
Xbit_r170_c92 bl_92 br_92 wl_170 vdd gnd cell_6t
Xbit_r171_c92 bl_92 br_92 wl_171 vdd gnd cell_6t
Xbit_r172_c92 bl_92 br_92 wl_172 vdd gnd cell_6t
Xbit_r173_c92 bl_92 br_92 wl_173 vdd gnd cell_6t
Xbit_r174_c92 bl_92 br_92 wl_174 vdd gnd cell_6t
Xbit_r175_c92 bl_92 br_92 wl_175 vdd gnd cell_6t
Xbit_r176_c92 bl_92 br_92 wl_176 vdd gnd cell_6t
Xbit_r177_c92 bl_92 br_92 wl_177 vdd gnd cell_6t
Xbit_r178_c92 bl_92 br_92 wl_178 vdd gnd cell_6t
Xbit_r179_c92 bl_92 br_92 wl_179 vdd gnd cell_6t
Xbit_r180_c92 bl_92 br_92 wl_180 vdd gnd cell_6t
Xbit_r181_c92 bl_92 br_92 wl_181 vdd gnd cell_6t
Xbit_r182_c92 bl_92 br_92 wl_182 vdd gnd cell_6t
Xbit_r183_c92 bl_92 br_92 wl_183 vdd gnd cell_6t
Xbit_r184_c92 bl_92 br_92 wl_184 vdd gnd cell_6t
Xbit_r185_c92 bl_92 br_92 wl_185 vdd gnd cell_6t
Xbit_r186_c92 bl_92 br_92 wl_186 vdd gnd cell_6t
Xbit_r187_c92 bl_92 br_92 wl_187 vdd gnd cell_6t
Xbit_r188_c92 bl_92 br_92 wl_188 vdd gnd cell_6t
Xbit_r189_c92 bl_92 br_92 wl_189 vdd gnd cell_6t
Xbit_r190_c92 bl_92 br_92 wl_190 vdd gnd cell_6t
Xbit_r191_c92 bl_92 br_92 wl_191 vdd gnd cell_6t
Xbit_r192_c92 bl_92 br_92 wl_192 vdd gnd cell_6t
Xbit_r193_c92 bl_92 br_92 wl_193 vdd gnd cell_6t
Xbit_r194_c92 bl_92 br_92 wl_194 vdd gnd cell_6t
Xbit_r195_c92 bl_92 br_92 wl_195 vdd gnd cell_6t
Xbit_r196_c92 bl_92 br_92 wl_196 vdd gnd cell_6t
Xbit_r197_c92 bl_92 br_92 wl_197 vdd gnd cell_6t
Xbit_r198_c92 bl_92 br_92 wl_198 vdd gnd cell_6t
Xbit_r199_c92 bl_92 br_92 wl_199 vdd gnd cell_6t
Xbit_r200_c92 bl_92 br_92 wl_200 vdd gnd cell_6t
Xbit_r201_c92 bl_92 br_92 wl_201 vdd gnd cell_6t
Xbit_r202_c92 bl_92 br_92 wl_202 vdd gnd cell_6t
Xbit_r203_c92 bl_92 br_92 wl_203 vdd gnd cell_6t
Xbit_r204_c92 bl_92 br_92 wl_204 vdd gnd cell_6t
Xbit_r205_c92 bl_92 br_92 wl_205 vdd gnd cell_6t
Xbit_r206_c92 bl_92 br_92 wl_206 vdd gnd cell_6t
Xbit_r207_c92 bl_92 br_92 wl_207 vdd gnd cell_6t
Xbit_r208_c92 bl_92 br_92 wl_208 vdd gnd cell_6t
Xbit_r209_c92 bl_92 br_92 wl_209 vdd gnd cell_6t
Xbit_r210_c92 bl_92 br_92 wl_210 vdd gnd cell_6t
Xbit_r211_c92 bl_92 br_92 wl_211 vdd gnd cell_6t
Xbit_r212_c92 bl_92 br_92 wl_212 vdd gnd cell_6t
Xbit_r213_c92 bl_92 br_92 wl_213 vdd gnd cell_6t
Xbit_r214_c92 bl_92 br_92 wl_214 vdd gnd cell_6t
Xbit_r215_c92 bl_92 br_92 wl_215 vdd gnd cell_6t
Xbit_r216_c92 bl_92 br_92 wl_216 vdd gnd cell_6t
Xbit_r217_c92 bl_92 br_92 wl_217 vdd gnd cell_6t
Xbit_r218_c92 bl_92 br_92 wl_218 vdd gnd cell_6t
Xbit_r219_c92 bl_92 br_92 wl_219 vdd gnd cell_6t
Xbit_r220_c92 bl_92 br_92 wl_220 vdd gnd cell_6t
Xbit_r221_c92 bl_92 br_92 wl_221 vdd gnd cell_6t
Xbit_r222_c92 bl_92 br_92 wl_222 vdd gnd cell_6t
Xbit_r223_c92 bl_92 br_92 wl_223 vdd gnd cell_6t
Xbit_r224_c92 bl_92 br_92 wl_224 vdd gnd cell_6t
Xbit_r225_c92 bl_92 br_92 wl_225 vdd gnd cell_6t
Xbit_r226_c92 bl_92 br_92 wl_226 vdd gnd cell_6t
Xbit_r227_c92 bl_92 br_92 wl_227 vdd gnd cell_6t
Xbit_r228_c92 bl_92 br_92 wl_228 vdd gnd cell_6t
Xbit_r229_c92 bl_92 br_92 wl_229 vdd gnd cell_6t
Xbit_r230_c92 bl_92 br_92 wl_230 vdd gnd cell_6t
Xbit_r231_c92 bl_92 br_92 wl_231 vdd gnd cell_6t
Xbit_r232_c92 bl_92 br_92 wl_232 vdd gnd cell_6t
Xbit_r233_c92 bl_92 br_92 wl_233 vdd gnd cell_6t
Xbit_r234_c92 bl_92 br_92 wl_234 vdd gnd cell_6t
Xbit_r235_c92 bl_92 br_92 wl_235 vdd gnd cell_6t
Xbit_r236_c92 bl_92 br_92 wl_236 vdd gnd cell_6t
Xbit_r237_c92 bl_92 br_92 wl_237 vdd gnd cell_6t
Xbit_r238_c92 bl_92 br_92 wl_238 vdd gnd cell_6t
Xbit_r239_c92 bl_92 br_92 wl_239 vdd gnd cell_6t
Xbit_r240_c92 bl_92 br_92 wl_240 vdd gnd cell_6t
Xbit_r241_c92 bl_92 br_92 wl_241 vdd gnd cell_6t
Xbit_r242_c92 bl_92 br_92 wl_242 vdd gnd cell_6t
Xbit_r243_c92 bl_92 br_92 wl_243 vdd gnd cell_6t
Xbit_r244_c92 bl_92 br_92 wl_244 vdd gnd cell_6t
Xbit_r245_c92 bl_92 br_92 wl_245 vdd gnd cell_6t
Xbit_r246_c92 bl_92 br_92 wl_246 vdd gnd cell_6t
Xbit_r247_c92 bl_92 br_92 wl_247 vdd gnd cell_6t
Xbit_r248_c92 bl_92 br_92 wl_248 vdd gnd cell_6t
Xbit_r249_c92 bl_92 br_92 wl_249 vdd gnd cell_6t
Xbit_r250_c92 bl_92 br_92 wl_250 vdd gnd cell_6t
Xbit_r251_c92 bl_92 br_92 wl_251 vdd gnd cell_6t
Xbit_r252_c92 bl_92 br_92 wl_252 vdd gnd cell_6t
Xbit_r253_c92 bl_92 br_92 wl_253 vdd gnd cell_6t
Xbit_r254_c92 bl_92 br_92 wl_254 vdd gnd cell_6t
Xbit_r255_c92 bl_92 br_92 wl_255 vdd gnd cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd cell_6t
Xbit_r1_c93 bl_93 br_93 wl_1 vdd gnd cell_6t
Xbit_r2_c93 bl_93 br_93 wl_2 vdd gnd cell_6t
Xbit_r3_c93 bl_93 br_93 wl_3 vdd gnd cell_6t
Xbit_r4_c93 bl_93 br_93 wl_4 vdd gnd cell_6t
Xbit_r5_c93 bl_93 br_93 wl_5 vdd gnd cell_6t
Xbit_r6_c93 bl_93 br_93 wl_6 vdd gnd cell_6t
Xbit_r7_c93 bl_93 br_93 wl_7 vdd gnd cell_6t
Xbit_r8_c93 bl_93 br_93 wl_8 vdd gnd cell_6t
Xbit_r9_c93 bl_93 br_93 wl_9 vdd gnd cell_6t
Xbit_r10_c93 bl_93 br_93 wl_10 vdd gnd cell_6t
Xbit_r11_c93 bl_93 br_93 wl_11 vdd gnd cell_6t
Xbit_r12_c93 bl_93 br_93 wl_12 vdd gnd cell_6t
Xbit_r13_c93 bl_93 br_93 wl_13 vdd gnd cell_6t
Xbit_r14_c93 bl_93 br_93 wl_14 vdd gnd cell_6t
Xbit_r15_c93 bl_93 br_93 wl_15 vdd gnd cell_6t
Xbit_r16_c93 bl_93 br_93 wl_16 vdd gnd cell_6t
Xbit_r17_c93 bl_93 br_93 wl_17 vdd gnd cell_6t
Xbit_r18_c93 bl_93 br_93 wl_18 vdd gnd cell_6t
Xbit_r19_c93 bl_93 br_93 wl_19 vdd gnd cell_6t
Xbit_r20_c93 bl_93 br_93 wl_20 vdd gnd cell_6t
Xbit_r21_c93 bl_93 br_93 wl_21 vdd gnd cell_6t
Xbit_r22_c93 bl_93 br_93 wl_22 vdd gnd cell_6t
Xbit_r23_c93 bl_93 br_93 wl_23 vdd gnd cell_6t
Xbit_r24_c93 bl_93 br_93 wl_24 vdd gnd cell_6t
Xbit_r25_c93 bl_93 br_93 wl_25 vdd gnd cell_6t
Xbit_r26_c93 bl_93 br_93 wl_26 vdd gnd cell_6t
Xbit_r27_c93 bl_93 br_93 wl_27 vdd gnd cell_6t
Xbit_r28_c93 bl_93 br_93 wl_28 vdd gnd cell_6t
Xbit_r29_c93 bl_93 br_93 wl_29 vdd gnd cell_6t
Xbit_r30_c93 bl_93 br_93 wl_30 vdd gnd cell_6t
Xbit_r31_c93 bl_93 br_93 wl_31 vdd gnd cell_6t
Xbit_r32_c93 bl_93 br_93 wl_32 vdd gnd cell_6t
Xbit_r33_c93 bl_93 br_93 wl_33 vdd gnd cell_6t
Xbit_r34_c93 bl_93 br_93 wl_34 vdd gnd cell_6t
Xbit_r35_c93 bl_93 br_93 wl_35 vdd gnd cell_6t
Xbit_r36_c93 bl_93 br_93 wl_36 vdd gnd cell_6t
Xbit_r37_c93 bl_93 br_93 wl_37 vdd gnd cell_6t
Xbit_r38_c93 bl_93 br_93 wl_38 vdd gnd cell_6t
Xbit_r39_c93 bl_93 br_93 wl_39 vdd gnd cell_6t
Xbit_r40_c93 bl_93 br_93 wl_40 vdd gnd cell_6t
Xbit_r41_c93 bl_93 br_93 wl_41 vdd gnd cell_6t
Xbit_r42_c93 bl_93 br_93 wl_42 vdd gnd cell_6t
Xbit_r43_c93 bl_93 br_93 wl_43 vdd gnd cell_6t
Xbit_r44_c93 bl_93 br_93 wl_44 vdd gnd cell_6t
Xbit_r45_c93 bl_93 br_93 wl_45 vdd gnd cell_6t
Xbit_r46_c93 bl_93 br_93 wl_46 vdd gnd cell_6t
Xbit_r47_c93 bl_93 br_93 wl_47 vdd gnd cell_6t
Xbit_r48_c93 bl_93 br_93 wl_48 vdd gnd cell_6t
Xbit_r49_c93 bl_93 br_93 wl_49 vdd gnd cell_6t
Xbit_r50_c93 bl_93 br_93 wl_50 vdd gnd cell_6t
Xbit_r51_c93 bl_93 br_93 wl_51 vdd gnd cell_6t
Xbit_r52_c93 bl_93 br_93 wl_52 vdd gnd cell_6t
Xbit_r53_c93 bl_93 br_93 wl_53 vdd gnd cell_6t
Xbit_r54_c93 bl_93 br_93 wl_54 vdd gnd cell_6t
Xbit_r55_c93 bl_93 br_93 wl_55 vdd gnd cell_6t
Xbit_r56_c93 bl_93 br_93 wl_56 vdd gnd cell_6t
Xbit_r57_c93 bl_93 br_93 wl_57 vdd gnd cell_6t
Xbit_r58_c93 bl_93 br_93 wl_58 vdd gnd cell_6t
Xbit_r59_c93 bl_93 br_93 wl_59 vdd gnd cell_6t
Xbit_r60_c93 bl_93 br_93 wl_60 vdd gnd cell_6t
Xbit_r61_c93 bl_93 br_93 wl_61 vdd gnd cell_6t
Xbit_r62_c93 bl_93 br_93 wl_62 vdd gnd cell_6t
Xbit_r63_c93 bl_93 br_93 wl_63 vdd gnd cell_6t
Xbit_r64_c93 bl_93 br_93 wl_64 vdd gnd cell_6t
Xbit_r65_c93 bl_93 br_93 wl_65 vdd gnd cell_6t
Xbit_r66_c93 bl_93 br_93 wl_66 vdd gnd cell_6t
Xbit_r67_c93 bl_93 br_93 wl_67 vdd gnd cell_6t
Xbit_r68_c93 bl_93 br_93 wl_68 vdd gnd cell_6t
Xbit_r69_c93 bl_93 br_93 wl_69 vdd gnd cell_6t
Xbit_r70_c93 bl_93 br_93 wl_70 vdd gnd cell_6t
Xbit_r71_c93 bl_93 br_93 wl_71 vdd gnd cell_6t
Xbit_r72_c93 bl_93 br_93 wl_72 vdd gnd cell_6t
Xbit_r73_c93 bl_93 br_93 wl_73 vdd gnd cell_6t
Xbit_r74_c93 bl_93 br_93 wl_74 vdd gnd cell_6t
Xbit_r75_c93 bl_93 br_93 wl_75 vdd gnd cell_6t
Xbit_r76_c93 bl_93 br_93 wl_76 vdd gnd cell_6t
Xbit_r77_c93 bl_93 br_93 wl_77 vdd gnd cell_6t
Xbit_r78_c93 bl_93 br_93 wl_78 vdd gnd cell_6t
Xbit_r79_c93 bl_93 br_93 wl_79 vdd gnd cell_6t
Xbit_r80_c93 bl_93 br_93 wl_80 vdd gnd cell_6t
Xbit_r81_c93 bl_93 br_93 wl_81 vdd gnd cell_6t
Xbit_r82_c93 bl_93 br_93 wl_82 vdd gnd cell_6t
Xbit_r83_c93 bl_93 br_93 wl_83 vdd gnd cell_6t
Xbit_r84_c93 bl_93 br_93 wl_84 vdd gnd cell_6t
Xbit_r85_c93 bl_93 br_93 wl_85 vdd gnd cell_6t
Xbit_r86_c93 bl_93 br_93 wl_86 vdd gnd cell_6t
Xbit_r87_c93 bl_93 br_93 wl_87 vdd gnd cell_6t
Xbit_r88_c93 bl_93 br_93 wl_88 vdd gnd cell_6t
Xbit_r89_c93 bl_93 br_93 wl_89 vdd gnd cell_6t
Xbit_r90_c93 bl_93 br_93 wl_90 vdd gnd cell_6t
Xbit_r91_c93 bl_93 br_93 wl_91 vdd gnd cell_6t
Xbit_r92_c93 bl_93 br_93 wl_92 vdd gnd cell_6t
Xbit_r93_c93 bl_93 br_93 wl_93 vdd gnd cell_6t
Xbit_r94_c93 bl_93 br_93 wl_94 vdd gnd cell_6t
Xbit_r95_c93 bl_93 br_93 wl_95 vdd gnd cell_6t
Xbit_r96_c93 bl_93 br_93 wl_96 vdd gnd cell_6t
Xbit_r97_c93 bl_93 br_93 wl_97 vdd gnd cell_6t
Xbit_r98_c93 bl_93 br_93 wl_98 vdd gnd cell_6t
Xbit_r99_c93 bl_93 br_93 wl_99 vdd gnd cell_6t
Xbit_r100_c93 bl_93 br_93 wl_100 vdd gnd cell_6t
Xbit_r101_c93 bl_93 br_93 wl_101 vdd gnd cell_6t
Xbit_r102_c93 bl_93 br_93 wl_102 vdd gnd cell_6t
Xbit_r103_c93 bl_93 br_93 wl_103 vdd gnd cell_6t
Xbit_r104_c93 bl_93 br_93 wl_104 vdd gnd cell_6t
Xbit_r105_c93 bl_93 br_93 wl_105 vdd gnd cell_6t
Xbit_r106_c93 bl_93 br_93 wl_106 vdd gnd cell_6t
Xbit_r107_c93 bl_93 br_93 wl_107 vdd gnd cell_6t
Xbit_r108_c93 bl_93 br_93 wl_108 vdd gnd cell_6t
Xbit_r109_c93 bl_93 br_93 wl_109 vdd gnd cell_6t
Xbit_r110_c93 bl_93 br_93 wl_110 vdd gnd cell_6t
Xbit_r111_c93 bl_93 br_93 wl_111 vdd gnd cell_6t
Xbit_r112_c93 bl_93 br_93 wl_112 vdd gnd cell_6t
Xbit_r113_c93 bl_93 br_93 wl_113 vdd gnd cell_6t
Xbit_r114_c93 bl_93 br_93 wl_114 vdd gnd cell_6t
Xbit_r115_c93 bl_93 br_93 wl_115 vdd gnd cell_6t
Xbit_r116_c93 bl_93 br_93 wl_116 vdd gnd cell_6t
Xbit_r117_c93 bl_93 br_93 wl_117 vdd gnd cell_6t
Xbit_r118_c93 bl_93 br_93 wl_118 vdd gnd cell_6t
Xbit_r119_c93 bl_93 br_93 wl_119 vdd gnd cell_6t
Xbit_r120_c93 bl_93 br_93 wl_120 vdd gnd cell_6t
Xbit_r121_c93 bl_93 br_93 wl_121 vdd gnd cell_6t
Xbit_r122_c93 bl_93 br_93 wl_122 vdd gnd cell_6t
Xbit_r123_c93 bl_93 br_93 wl_123 vdd gnd cell_6t
Xbit_r124_c93 bl_93 br_93 wl_124 vdd gnd cell_6t
Xbit_r125_c93 bl_93 br_93 wl_125 vdd gnd cell_6t
Xbit_r126_c93 bl_93 br_93 wl_126 vdd gnd cell_6t
Xbit_r127_c93 bl_93 br_93 wl_127 vdd gnd cell_6t
Xbit_r128_c93 bl_93 br_93 wl_128 vdd gnd cell_6t
Xbit_r129_c93 bl_93 br_93 wl_129 vdd gnd cell_6t
Xbit_r130_c93 bl_93 br_93 wl_130 vdd gnd cell_6t
Xbit_r131_c93 bl_93 br_93 wl_131 vdd gnd cell_6t
Xbit_r132_c93 bl_93 br_93 wl_132 vdd gnd cell_6t
Xbit_r133_c93 bl_93 br_93 wl_133 vdd gnd cell_6t
Xbit_r134_c93 bl_93 br_93 wl_134 vdd gnd cell_6t
Xbit_r135_c93 bl_93 br_93 wl_135 vdd gnd cell_6t
Xbit_r136_c93 bl_93 br_93 wl_136 vdd gnd cell_6t
Xbit_r137_c93 bl_93 br_93 wl_137 vdd gnd cell_6t
Xbit_r138_c93 bl_93 br_93 wl_138 vdd gnd cell_6t
Xbit_r139_c93 bl_93 br_93 wl_139 vdd gnd cell_6t
Xbit_r140_c93 bl_93 br_93 wl_140 vdd gnd cell_6t
Xbit_r141_c93 bl_93 br_93 wl_141 vdd gnd cell_6t
Xbit_r142_c93 bl_93 br_93 wl_142 vdd gnd cell_6t
Xbit_r143_c93 bl_93 br_93 wl_143 vdd gnd cell_6t
Xbit_r144_c93 bl_93 br_93 wl_144 vdd gnd cell_6t
Xbit_r145_c93 bl_93 br_93 wl_145 vdd gnd cell_6t
Xbit_r146_c93 bl_93 br_93 wl_146 vdd gnd cell_6t
Xbit_r147_c93 bl_93 br_93 wl_147 vdd gnd cell_6t
Xbit_r148_c93 bl_93 br_93 wl_148 vdd gnd cell_6t
Xbit_r149_c93 bl_93 br_93 wl_149 vdd gnd cell_6t
Xbit_r150_c93 bl_93 br_93 wl_150 vdd gnd cell_6t
Xbit_r151_c93 bl_93 br_93 wl_151 vdd gnd cell_6t
Xbit_r152_c93 bl_93 br_93 wl_152 vdd gnd cell_6t
Xbit_r153_c93 bl_93 br_93 wl_153 vdd gnd cell_6t
Xbit_r154_c93 bl_93 br_93 wl_154 vdd gnd cell_6t
Xbit_r155_c93 bl_93 br_93 wl_155 vdd gnd cell_6t
Xbit_r156_c93 bl_93 br_93 wl_156 vdd gnd cell_6t
Xbit_r157_c93 bl_93 br_93 wl_157 vdd gnd cell_6t
Xbit_r158_c93 bl_93 br_93 wl_158 vdd gnd cell_6t
Xbit_r159_c93 bl_93 br_93 wl_159 vdd gnd cell_6t
Xbit_r160_c93 bl_93 br_93 wl_160 vdd gnd cell_6t
Xbit_r161_c93 bl_93 br_93 wl_161 vdd gnd cell_6t
Xbit_r162_c93 bl_93 br_93 wl_162 vdd gnd cell_6t
Xbit_r163_c93 bl_93 br_93 wl_163 vdd gnd cell_6t
Xbit_r164_c93 bl_93 br_93 wl_164 vdd gnd cell_6t
Xbit_r165_c93 bl_93 br_93 wl_165 vdd gnd cell_6t
Xbit_r166_c93 bl_93 br_93 wl_166 vdd gnd cell_6t
Xbit_r167_c93 bl_93 br_93 wl_167 vdd gnd cell_6t
Xbit_r168_c93 bl_93 br_93 wl_168 vdd gnd cell_6t
Xbit_r169_c93 bl_93 br_93 wl_169 vdd gnd cell_6t
Xbit_r170_c93 bl_93 br_93 wl_170 vdd gnd cell_6t
Xbit_r171_c93 bl_93 br_93 wl_171 vdd gnd cell_6t
Xbit_r172_c93 bl_93 br_93 wl_172 vdd gnd cell_6t
Xbit_r173_c93 bl_93 br_93 wl_173 vdd gnd cell_6t
Xbit_r174_c93 bl_93 br_93 wl_174 vdd gnd cell_6t
Xbit_r175_c93 bl_93 br_93 wl_175 vdd gnd cell_6t
Xbit_r176_c93 bl_93 br_93 wl_176 vdd gnd cell_6t
Xbit_r177_c93 bl_93 br_93 wl_177 vdd gnd cell_6t
Xbit_r178_c93 bl_93 br_93 wl_178 vdd gnd cell_6t
Xbit_r179_c93 bl_93 br_93 wl_179 vdd gnd cell_6t
Xbit_r180_c93 bl_93 br_93 wl_180 vdd gnd cell_6t
Xbit_r181_c93 bl_93 br_93 wl_181 vdd gnd cell_6t
Xbit_r182_c93 bl_93 br_93 wl_182 vdd gnd cell_6t
Xbit_r183_c93 bl_93 br_93 wl_183 vdd gnd cell_6t
Xbit_r184_c93 bl_93 br_93 wl_184 vdd gnd cell_6t
Xbit_r185_c93 bl_93 br_93 wl_185 vdd gnd cell_6t
Xbit_r186_c93 bl_93 br_93 wl_186 vdd gnd cell_6t
Xbit_r187_c93 bl_93 br_93 wl_187 vdd gnd cell_6t
Xbit_r188_c93 bl_93 br_93 wl_188 vdd gnd cell_6t
Xbit_r189_c93 bl_93 br_93 wl_189 vdd gnd cell_6t
Xbit_r190_c93 bl_93 br_93 wl_190 vdd gnd cell_6t
Xbit_r191_c93 bl_93 br_93 wl_191 vdd gnd cell_6t
Xbit_r192_c93 bl_93 br_93 wl_192 vdd gnd cell_6t
Xbit_r193_c93 bl_93 br_93 wl_193 vdd gnd cell_6t
Xbit_r194_c93 bl_93 br_93 wl_194 vdd gnd cell_6t
Xbit_r195_c93 bl_93 br_93 wl_195 vdd gnd cell_6t
Xbit_r196_c93 bl_93 br_93 wl_196 vdd gnd cell_6t
Xbit_r197_c93 bl_93 br_93 wl_197 vdd gnd cell_6t
Xbit_r198_c93 bl_93 br_93 wl_198 vdd gnd cell_6t
Xbit_r199_c93 bl_93 br_93 wl_199 vdd gnd cell_6t
Xbit_r200_c93 bl_93 br_93 wl_200 vdd gnd cell_6t
Xbit_r201_c93 bl_93 br_93 wl_201 vdd gnd cell_6t
Xbit_r202_c93 bl_93 br_93 wl_202 vdd gnd cell_6t
Xbit_r203_c93 bl_93 br_93 wl_203 vdd gnd cell_6t
Xbit_r204_c93 bl_93 br_93 wl_204 vdd gnd cell_6t
Xbit_r205_c93 bl_93 br_93 wl_205 vdd gnd cell_6t
Xbit_r206_c93 bl_93 br_93 wl_206 vdd gnd cell_6t
Xbit_r207_c93 bl_93 br_93 wl_207 vdd gnd cell_6t
Xbit_r208_c93 bl_93 br_93 wl_208 vdd gnd cell_6t
Xbit_r209_c93 bl_93 br_93 wl_209 vdd gnd cell_6t
Xbit_r210_c93 bl_93 br_93 wl_210 vdd gnd cell_6t
Xbit_r211_c93 bl_93 br_93 wl_211 vdd gnd cell_6t
Xbit_r212_c93 bl_93 br_93 wl_212 vdd gnd cell_6t
Xbit_r213_c93 bl_93 br_93 wl_213 vdd gnd cell_6t
Xbit_r214_c93 bl_93 br_93 wl_214 vdd gnd cell_6t
Xbit_r215_c93 bl_93 br_93 wl_215 vdd gnd cell_6t
Xbit_r216_c93 bl_93 br_93 wl_216 vdd gnd cell_6t
Xbit_r217_c93 bl_93 br_93 wl_217 vdd gnd cell_6t
Xbit_r218_c93 bl_93 br_93 wl_218 vdd gnd cell_6t
Xbit_r219_c93 bl_93 br_93 wl_219 vdd gnd cell_6t
Xbit_r220_c93 bl_93 br_93 wl_220 vdd gnd cell_6t
Xbit_r221_c93 bl_93 br_93 wl_221 vdd gnd cell_6t
Xbit_r222_c93 bl_93 br_93 wl_222 vdd gnd cell_6t
Xbit_r223_c93 bl_93 br_93 wl_223 vdd gnd cell_6t
Xbit_r224_c93 bl_93 br_93 wl_224 vdd gnd cell_6t
Xbit_r225_c93 bl_93 br_93 wl_225 vdd gnd cell_6t
Xbit_r226_c93 bl_93 br_93 wl_226 vdd gnd cell_6t
Xbit_r227_c93 bl_93 br_93 wl_227 vdd gnd cell_6t
Xbit_r228_c93 bl_93 br_93 wl_228 vdd gnd cell_6t
Xbit_r229_c93 bl_93 br_93 wl_229 vdd gnd cell_6t
Xbit_r230_c93 bl_93 br_93 wl_230 vdd gnd cell_6t
Xbit_r231_c93 bl_93 br_93 wl_231 vdd gnd cell_6t
Xbit_r232_c93 bl_93 br_93 wl_232 vdd gnd cell_6t
Xbit_r233_c93 bl_93 br_93 wl_233 vdd gnd cell_6t
Xbit_r234_c93 bl_93 br_93 wl_234 vdd gnd cell_6t
Xbit_r235_c93 bl_93 br_93 wl_235 vdd gnd cell_6t
Xbit_r236_c93 bl_93 br_93 wl_236 vdd gnd cell_6t
Xbit_r237_c93 bl_93 br_93 wl_237 vdd gnd cell_6t
Xbit_r238_c93 bl_93 br_93 wl_238 vdd gnd cell_6t
Xbit_r239_c93 bl_93 br_93 wl_239 vdd gnd cell_6t
Xbit_r240_c93 bl_93 br_93 wl_240 vdd gnd cell_6t
Xbit_r241_c93 bl_93 br_93 wl_241 vdd gnd cell_6t
Xbit_r242_c93 bl_93 br_93 wl_242 vdd gnd cell_6t
Xbit_r243_c93 bl_93 br_93 wl_243 vdd gnd cell_6t
Xbit_r244_c93 bl_93 br_93 wl_244 vdd gnd cell_6t
Xbit_r245_c93 bl_93 br_93 wl_245 vdd gnd cell_6t
Xbit_r246_c93 bl_93 br_93 wl_246 vdd gnd cell_6t
Xbit_r247_c93 bl_93 br_93 wl_247 vdd gnd cell_6t
Xbit_r248_c93 bl_93 br_93 wl_248 vdd gnd cell_6t
Xbit_r249_c93 bl_93 br_93 wl_249 vdd gnd cell_6t
Xbit_r250_c93 bl_93 br_93 wl_250 vdd gnd cell_6t
Xbit_r251_c93 bl_93 br_93 wl_251 vdd gnd cell_6t
Xbit_r252_c93 bl_93 br_93 wl_252 vdd gnd cell_6t
Xbit_r253_c93 bl_93 br_93 wl_253 vdd gnd cell_6t
Xbit_r254_c93 bl_93 br_93 wl_254 vdd gnd cell_6t
Xbit_r255_c93 bl_93 br_93 wl_255 vdd gnd cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd cell_6t
Xbit_r1_c94 bl_94 br_94 wl_1 vdd gnd cell_6t
Xbit_r2_c94 bl_94 br_94 wl_2 vdd gnd cell_6t
Xbit_r3_c94 bl_94 br_94 wl_3 vdd gnd cell_6t
Xbit_r4_c94 bl_94 br_94 wl_4 vdd gnd cell_6t
Xbit_r5_c94 bl_94 br_94 wl_5 vdd gnd cell_6t
Xbit_r6_c94 bl_94 br_94 wl_6 vdd gnd cell_6t
Xbit_r7_c94 bl_94 br_94 wl_7 vdd gnd cell_6t
Xbit_r8_c94 bl_94 br_94 wl_8 vdd gnd cell_6t
Xbit_r9_c94 bl_94 br_94 wl_9 vdd gnd cell_6t
Xbit_r10_c94 bl_94 br_94 wl_10 vdd gnd cell_6t
Xbit_r11_c94 bl_94 br_94 wl_11 vdd gnd cell_6t
Xbit_r12_c94 bl_94 br_94 wl_12 vdd gnd cell_6t
Xbit_r13_c94 bl_94 br_94 wl_13 vdd gnd cell_6t
Xbit_r14_c94 bl_94 br_94 wl_14 vdd gnd cell_6t
Xbit_r15_c94 bl_94 br_94 wl_15 vdd gnd cell_6t
Xbit_r16_c94 bl_94 br_94 wl_16 vdd gnd cell_6t
Xbit_r17_c94 bl_94 br_94 wl_17 vdd gnd cell_6t
Xbit_r18_c94 bl_94 br_94 wl_18 vdd gnd cell_6t
Xbit_r19_c94 bl_94 br_94 wl_19 vdd gnd cell_6t
Xbit_r20_c94 bl_94 br_94 wl_20 vdd gnd cell_6t
Xbit_r21_c94 bl_94 br_94 wl_21 vdd gnd cell_6t
Xbit_r22_c94 bl_94 br_94 wl_22 vdd gnd cell_6t
Xbit_r23_c94 bl_94 br_94 wl_23 vdd gnd cell_6t
Xbit_r24_c94 bl_94 br_94 wl_24 vdd gnd cell_6t
Xbit_r25_c94 bl_94 br_94 wl_25 vdd gnd cell_6t
Xbit_r26_c94 bl_94 br_94 wl_26 vdd gnd cell_6t
Xbit_r27_c94 bl_94 br_94 wl_27 vdd gnd cell_6t
Xbit_r28_c94 bl_94 br_94 wl_28 vdd gnd cell_6t
Xbit_r29_c94 bl_94 br_94 wl_29 vdd gnd cell_6t
Xbit_r30_c94 bl_94 br_94 wl_30 vdd gnd cell_6t
Xbit_r31_c94 bl_94 br_94 wl_31 vdd gnd cell_6t
Xbit_r32_c94 bl_94 br_94 wl_32 vdd gnd cell_6t
Xbit_r33_c94 bl_94 br_94 wl_33 vdd gnd cell_6t
Xbit_r34_c94 bl_94 br_94 wl_34 vdd gnd cell_6t
Xbit_r35_c94 bl_94 br_94 wl_35 vdd gnd cell_6t
Xbit_r36_c94 bl_94 br_94 wl_36 vdd gnd cell_6t
Xbit_r37_c94 bl_94 br_94 wl_37 vdd gnd cell_6t
Xbit_r38_c94 bl_94 br_94 wl_38 vdd gnd cell_6t
Xbit_r39_c94 bl_94 br_94 wl_39 vdd gnd cell_6t
Xbit_r40_c94 bl_94 br_94 wl_40 vdd gnd cell_6t
Xbit_r41_c94 bl_94 br_94 wl_41 vdd gnd cell_6t
Xbit_r42_c94 bl_94 br_94 wl_42 vdd gnd cell_6t
Xbit_r43_c94 bl_94 br_94 wl_43 vdd gnd cell_6t
Xbit_r44_c94 bl_94 br_94 wl_44 vdd gnd cell_6t
Xbit_r45_c94 bl_94 br_94 wl_45 vdd gnd cell_6t
Xbit_r46_c94 bl_94 br_94 wl_46 vdd gnd cell_6t
Xbit_r47_c94 bl_94 br_94 wl_47 vdd gnd cell_6t
Xbit_r48_c94 bl_94 br_94 wl_48 vdd gnd cell_6t
Xbit_r49_c94 bl_94 br_94 wl_49 vdd gnd cell_6t
Xbit_r50_c94 bl_94 br_94 wl_50 vdd gnd cell_6t
Xbit_r51_c94 bl_94 br_94 wl_51 vdd gnd cell_6t
Xbit_r52_c94 bl_94 br_94 wl_52 vdd gnd cell_6t
Xbit_r53_c94 bl_94 br_94 wl_53 vdd gnd cell_6t
Xbit_r54_c94 bl_94 br_94 wl_54 vdd gnd cell_6t
Xbit_r55_c94 bl_94 br_94 wl_55 vdd gnd cell_6t
Xbit_r56_c94 bl_94 br_94 wl_56 vdd gnd cell_6t
Xbit_r57_c94 bl_94 br_94 wl_57 vdd gnd cell_6t
Xbit_r58_c94 bl_94 br_94 wl_58 vdd gnd cell_6t
Xbit_r59_c94 bl_94 br_94 wl_59 vdd gnd cell_6t
Xbit_r60_c94 bl_94 br_94 wl_60 vdd gnd cell_6t
Xbit_r61_c94 bl_94 br_94 wl_61 vdd gnd cell_6t
Xbit_r62_c94 bl_94 br_94 wl_62 vdd gnd cell_6t
Xbit_r63_c94 bl_94 br_94 wl_63 vdd gnd cell_6t
Xbit_r64_c94 bl_94 br_94 wl_64 vdd gnd cell_6t
Xbit_r65_c94 bl_94 br_94 wl_65 vdd gnd cell_6t
Xbit_r66_c94 bl_94 br_94 wl_66 vdd gnd cell_6t
Xbit_r67_c94 bl_94 br_94 wl_67 vdd gnd cell_6t
Xbit_r68_c94 bl_94 br_94 wl_68 vdd gnd cell_6t
Xbit_r69_c94 bl_94 br_94 wl_69 vdd gnd cell_6t
Xbit_r70_c94 bl_94 br_94 wl_70 vdd gnd cell_6t
Xbit_r71_c94 bl_94 br_94 wl_71 vdd gnd cell_6t
Xbit_r72_c94 bl_94 br_94 wl_72 vdd gnd cell_6t
Xbit_r73_c94 bl_94 br_94 wl_73 vdd gnd cell_6t
Xbit_r74_c94 bl_94 br_94 wl_74 vdd gnd cell_6t
Xbit_r75_c94 bl_94 br_94 wl_75 vdd gnd cell_6t
Xbit_r76_c94 bl_94 br_94 wl_76 vdd gnd cell_6t
Xbit_r77_c94 bl_94 br_94 wl_77 vdd gnd cell_6t
Xbit_r78_c94 bl_94 br_94 wl_78 vdd gnd cell_6t
Xbit_r79_c94 bl_94 br_94 wl_79 vdd gnd cell_6t
Xbit_r80_c94 bl_94 br_94 wl_80 vdd gnd cell_6t
Xbit_r81_c94 bl_94 br_94 wl_81 vdd gnd cell_6t
Xbit_r82_c94 bl_94 br_94 wl_82 vdd gnd cell_6t
Xbit_r83_c94 bl_94 br_94 wl_83 vdd gnd cell_6t
Xbit_r84_c94 bl_94 br_94 wl_84 vdd gnd cell_6t
Xbit_r85_c94 bl_94 br_94 wl_85 vdd gnd cell_6t
Xbit_r86_c94 bl_94 br_94 wl_86 vdd gnd cell_6t
Xbit_r87_c94 bl_94 br_94 wl_87 vdd gnd cell_6t
Xbit_r88_c94 bl_94 br_94 wl_88 vdd gnd cell_6t
Xbit_r89_c94 bl_94 br_94 wl_89 vdd gnd cell_6t
Xbit_r90_c94 bl_94 br_94 wl_90 vdd gnd cell_6t
Xbit_r91_c94 bl_94 br_94 wl_91 vdd gnd cell_6t
Xbit_r92_c94 bl_94 br_94 wl_92 vdd gnd cell_6t
Xbit_r93_c94 bl_94 br_94 wl_93 vdd gnd cell_6t
Xbit_r94_c94 bl_94 br_94 wl_94 vdd gnd cell_6t
Xbit_r95_c94 bl_94 br_94 wl_95 vdd gnd cell_6t
Xbit_r96_c94 bl_94 br_94 wl_96 vdd gnd cell_6t
Xbit_r97_c94 bl_94 br_94 wl_97 vdd gnd cell_6t
Xbit_r98_c94 bl_94 br_94 wl_98 vdd gnd cell_6t
Xbit_r99_c94 bl_94 br_94 wl_99 vdd gnd cell_6t
Xbit_r100_c94 bl_94 br_94 wl_100 vdd gnd cell_6t
Xbit_r101_c94 bl_94 br_94 wl_101 vdd gnd cell_6t
Xbit_r102_c94 bl_94 br_94 wl_102 vdd gnd cell_6t
Xbit_r103_c94 bl_94 br_94 wl_103 vdd gnd cell_6t
Xbit_r104_c94 bl_94 br_94 wl_104 vdd gnd cell_6t
Xbit_r105_c94 bl_94 br_94 wl_105 vdd gnd cell_6t
Xbit_r106_c94 bl_94 br_94 wl_106 vdd gnd cell_6t
Xbit_r107_c94 bl_94 br_94 wl_107 vdd gnd cell_6t
Xbit_r108_c94 bl_94 br_94 wl_108 vdd gnd cell_6t
Xbit_r109_c94 bl_94 br_94 wl_109 vdd gnd cell_6t
Xbit_r110_c94 bl_94 br_94 wl_110 vdd gnd cell_6t
Xbit_r111_c94 bl_94 br_94 wl_111 vdd gnd cell_6t
Xbit_r112_c94 bl_94 br_94 wl_112 vdd gnd cell_6t
Xbit_r113_c94 bl_94 br_94 wl_113 vdd gnd cell_6t
Xbit_r114_c94 bl_94 br_94 wl_114 vdd gnd cell_6t
Xbit_r115_c94 bl_94 br_94 wl_115 vdd gnd cell_6t
Xbit_r116_c94 bl_94 br_94 wl_116 vdd gnd cell_6t
Xbit_r117_c94 bl_94 br_94 wl_117 vdd gnd cell_6t
Xbit_r118_c94 bl_94 br_94 wl_118 vdd gnd cell_6t
Xbit_r119_c94 bl_94 br_94 wl_119 vdd gnd cell_6t
Xbit_r120_c94 bl_94 br_94 wl_120 vdd gnd cell_6t
Xbit_r121_c94 bl_94 br_94 wl_121 vdd gnd cell_6t
Xbit_r122_c94 bl_94 br_94 wl_122 vdd gnd cell_6t
Xbit_r123_c94 bl_94 br_94 wl_123 vdd gnd cell_6t
Xbit_r124_c94 bl_94 br_94 wl_124 vdd gnd cell_6t
Xbit_r125_c94 bl_94 br_94 wl_125 vdd gnd cell_6t
Xbit_r126_c94 bl_94 br_94 wl_126 vdd gnd cell_6t
Xbit_r127_c94 bl_94 br_94 wl_127 vdd gnd cell_6t
Xbit_r128_c94 bl_94 br_94 wl_128 vdd gnd cell_6t
Xbit_r129_c94 bl_94 br_94 wl_129 vdd gnd cell_6t
Xbit_r130_c94 bl_94 br_94 wl_130 vdd gnd cell_6t
Xbit_r131_c94 bl_94 br_94 wl_131 vdd gnd cell_6t
Xbit_r132_c94 bl_94 br_94 wl_132 vdd gnd cell_6t
Xbit_r133_c94 bl_94 br_94 wl_133 vdd gnd cell_6t
Xbit_r134_c94 bl_94 br_94 wl_134 vdd gnd cell_6t
Xbit_r135_c94 bl_94 br_94 wl_135 vdd gnd cell_6t
Xbit_r136_c94 bl_94 br_94 wl_136 vdd gnd cell_6t
Xbit_r137_c94 bl_94 br_94 wl_137 vdd gnd cell_6t
Xbit_r138_c94 bl_94 br_94 wl_138 vdd gnd cell_6t
Xbit_r139_c94 bl_94 br_94 wl_139 vdd gnd cell_6t
Xbit_r140_c94 bl_94 br_94 wl_140 vdd gnd cell_6t
Xbit_r141_c94 bl_94 br_94 wl_141 vdd gnd cell_6t
Xbit_r142_c94 bl_94 br_94 wl_142 vdd gnd cell_6t
Xbit_r143_c94 bl_94 br_94 wl_143 vdd gnd cell_6t
Xbit_r144_c94 bl_94 br_94 wl_144 vdd gnd cell_6t
Xbit_r145_c94 bl_94 br_94 wl_145 vdd gnd cell_6t
Xbit_r146_c94 bl_94 br_94 wl_146 vdd gnd cell_6t
Xbit_r147_c94 bl_94 br_94 wl_147 vdd gnd cell_6t
Xbit_r148_c94 bl_94 br_94 wl_148 vdd gnd cell_6t
Xbit_r149_c94 bl_94 br_94 wl_149 vdd gnd cell_6t
Xbit_r150_c94 bl_94 br_94 wl_150 vdd gnd cell_6t
Xbit_r151_c94 bl_94 br_94 wl_151 vdd gnd cell_6t
Xbit_r152_c94 bl_94 br_94 wl_152 vdd gnd cell_6t
Xbit_r153_c94 bl_94 br_94 wl_153 vdd gnd cell_6t
Xbit_r154_c94 bl_94 br_94 wl_154 vdd gnd cell_6t
Xbit_r155_c94 bl_94 br_94 wl_155 vdd gnd cell_6t
Xbit_r156_c94 bl_94 br_94 wl_156 vdd gnd cell_6t
Xbit_r157_c94 bl_94 br_94 wl_157 vdd gnd cell_6t
Xbit_r158_c94 bl_94 br_94 wl_158 vdd gnd cell_6t
Xbit_r159_c94 bl_94 br_94 wl_159 vdd gnd cell_6t
Xbit_r160_c94 bl_94 br_94 wl_160 vdd gnd cell_6t
Xbit_r161_c94 bl_94 br_94 wl_161 vdd gnd cell_6t
Xbit_r162_c94 bl_94 br_94 wl_162 vdd gnd cell_6t
Xbit_r163_c94 bl_94 br_94 wl_163 vdd gnd cell_6t
Xbit_r164_c94 bl_94 br_94 wl_164 vdd gnd cell_6t
Xbit_r165_c94 bl_94 br_94 wl_165 vdd gnd cell_6t
Xbit_r166_c94 bl_94 br_94 wl_166 vdd gnd cell_6t
Xbit_r167_c94 bl_94 br_94 wl_167 vdd gnd cell_6t
Xbit_r168_c94 bl_94 br_94 wl_168 vdd gnd cell_6t
Xbit_r169_c94 bl_94 br_94 wl_169 vdd gnd cell_6t
Xbit_r170_c94 bl_94 br_94 wl_170 vdd gnd cell_6t
Xbit_r171_c94 bl_94 br_94 wl_171 vdd gnd cell_6t
Xbit_r172_c94 bl_94 br_94 wl_172 vdd gnd cell_6t
Xbit_r173_c94 bl_94 br_94 wl_173 vdd gnd cell_6t
Xbit_r174_c94 bl_94 br_94 wl_174 vdd gnd cell_6t
Xbit_r175_c94 bl_94 br_94 wl_175 vdd gnd cell_6t
Xbit_r176_c94 bl_94 br_94 wl_176 vdd gnd cell_6t
Xbit_r177_c94 bl_94 br_94 wl_177 vdd gnd cell_6t
Xbit_r178_c94 bl_94 br_94 wl_178 vdd gnd cell_6t
Xbit_r179_c94 bl_94 br_94 wl_179 vdd gnd cell_6t
Xbit_r180_c94 bl_94 br_94 wl_180 vdd gnd cell_6t
Xbit_r181_c94 bl_94 br_94 wl_181 vdd gnd cell_6t
Xbit_r182_c94 bl_94 br_94 wl_182 vdd gnd cell_6t
Xbit_r183_c94 bl_94 br_94 wl_183 vdd gnd cell_6t
Xbit_r184_c94 bl_94 br_94 wl_184 vdd gnd cell_6t
Xbit_r185_c94 bl_94 br_94 wl_185 vdd gnd cell_6t
Xbit_r186_c94 bl_94 br_94 wl_186 vdd gnd cell_6t
Xbit_r187_c94 bl_94 br_94 wl_187 vdd gnd cell_6t
Xbit_r188_c94 bl_94 br_94 wl_188 vdd gnd cell_6t
Xbit_r189_c94 bl_94 br_94 wl_189 vdd gnd cell_6t
Xbit_r190_c94 bl_94 br_94 wl_190 vdd gnd cell_6t
Xbit_r191_c94 bl_94 br_94 wl_191 vdd gnd cell_6t
Xbit_r192_c94 bl_94 br_94 wl_192 vdd gnd cell_6t
Xbit_r193_c94 bl_94 br_94 wl_193 vdd gnd cell_6t
Xbit_r194_c94 bl_94 br_94 wl_194 vdd gnd cell_6t
Xbit_r195_c94 bl_94 br_94 wl_195 vdd gnd cell_6t
Xbit_r196_c94 bl_94 br_94 wl_196 vdd gnd cell_6t
Xbit_r197_c94 bl_94 br_94 wl_197 vdd gnd cell_6t
Xbit_r198_c94 bl_94 br_94 wl_198 vdd gnd cell_6t
Xbit_r199_c94 bl_94 br_94 wl_199 vdd gnd cell_6t
Xbit_r200_c94 bl_94 br_94 wl_200 vdd gnd cell_6t
Xbit_r201_c94 bl_94 br_94 wl_201 vdd gnd cell_6t
Xbit_r202_c94 bl_94 br_94 wl_202 vdd gnd cell_6t
Xbit_r203_c94 bl_94 br_94 wl_203 vdd gnd cell_6t
Xbit_r204_c94 bl_94 br_94 wl_204 vdd gnd cell_6t
Xbit_r205_c94 bl_94 br_94 wl_205 vdd gnd cell_6t
Xbit_r206_c94 bl_94 br_94 wl_206 vdd gnd cell_6t
Xbit_r207_c94 bl_94 br_94 wl_207 vdd gnd cell_6t
Xbit_r208_c94 bl_94 br_94 wl_208 vdd gnd cell_6t
Xbit_r209_c94 bl_94 br_94 wl_209 vdd gnd cell_6t
Xbit_r210_c94 bl_94 br_94 wl_210 vdd gnd cell_6t
Xbit_r211_c94 bl_94 br_94 wl_211 vdd gnd cell_6t
Xbit_r212_c94 bl_94 br_94 wl_212 vdd gnd cell_6t
Xbit_r213_c94 bl_94 br_94 wl_213 vdd gnd cell_6t
Xbit_r214_c94 bl_94 br_94 wl_214 vdd gnd cell_6t
Xbit_r215_c94 bl_94 br_94 wl_215 vdd gnd cell_6t
Xbit_r216_c94 bl_94 br_94 wl_216 vdd gnd cell_6t
Xbit_r217_c94 bl_94 br_94 wl_217 vdd gnd cell_6t
Xbit_r218_c94 bl_94 br_94 wl_218 vdd gnd cell_6t
Xbit_r219_c94 bl_94 br_94 wl_219 vdd gnd cell_6t
Xbit_r220_c94 bl_94 br_94 wl_220 vdd gnd cell_6t
Xbit_r221_c94 bl_94 br_94 wl_221 vdd gnd cell_6t
Xbit_r222_c94 bl_94 br_94 wl_222 vdd gnd cell_6t
Xbit_r223_c94 bl_94 br_94 wl_223 vdd gnd cell_6t
Xbit_r224_c94 bl_94 br_94 wl_224 vdd gnd cell_6t
Xbit_r225_c94 bl_94 br_94 wl_225 vdd gnd cell_6t
Xbit_r226_c94 bl_94 br_94 wl_226 vdd gnd cell_6t
Xbit_r227_c94 bl_94 br_94 wl_227 vdd gnd cell_6t
Xbit_r228_c94 bl_94 br_94 wl_228 vdd gnd cell_6t
Xbit_r229_c94 bl_94 br_94 wl_229 vdd gnd cell_6t
Xbit_r230_c94 bl_94 br_94 wl_230 vdd gnd cell_6t
Xbit_r231_c94 bl_94 br_94 wl_231 vdd gnd cell_6t
Xbit_r232_c94 bl_94 br_94 wl_232 vdd gnd cell_6t
Xbit_r233_c94 bl_94 br_94 wl_233 vdd gnd cell_6t
Xbit_r234_c94 bl_94 br_94 wl_234 vdd gnd cell_6t
Xbit_r235_c94 bl_94 br_94 wl_235 vdd gnd cell_6t
Xbit_r236_c94 bl_94 br_94 wl_236 vdd gnd cell_6t
Xbit_r237_c94 bl_94 br_94 wl_237 vdd gnd cell_6t
Xbit_r238_c94 bl_94 br_94 wl_238 vdd gnd cell_6t
Xbit_r239_c94 bl_94 br_94 wl_239 vdd gnd cell_6t
Xbit_r240_c94 bl_94 br_94 wl_240 vdd gnd cell_6t
Xbit_r241_c94 bl_94 br_94 wl_241 vdd gnd cell_6t
Xbit_r242_c94 bl_94 br_94 wl_242 vdd gnd cell_6t
Xbit_r243_c94 bl_94 br_94 wl_243 vdd gnd cell_6t
Xbit_r244_c94 bl_94 br_94 wl_244 vdd gnd cell_6t
Xbit_r245_c94 bl_94 br_94 wl_245 vdd gnd cell_6t
Xbit_r246_c94 bl_94 br_94 wl_246 vdd gnd cell_6t
Xbit_r247_c94 bl_94 br_94 wl_247 vdd gnd cell_6t
Xbit_r248_c94 bl_94 br_94 wl_248 vdd gnd cell_6t
Xbit_r249_c94 bl_94 br_94 wl_249 vdd gnd cell_6t
Xbit_r250_c94 bl_94 br_94 wl_250 vdd gnd cell_6t
Xbit_r251_c94 bl_94 br_94 wl_251 vdd gnd cell_6t
Xbit_r252_c94 bl_94 br_94 wl_252 vdd gnd cell_6t
Xbit_r253_c94 bl_94 br_94 wl_253 vdd gnd cell_6t
Xbit_r254_c94 bl_94 br_94 wl_254 vdd gnd cell_6t
Xbit_r255_c94 bl_94 br_94 wl_255 vdd gnd cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd cell_6t
Xbit_r1_c95 bl_95 br_95 wl_1 vdd gnd cell_6t
Xbit_r2_c95 bl_95 br_95 wl_2 vdd gnd cell_6t
Xbit_r3_c95 bl_95 br_95 wl_3 vdd gnd cell_6t
Xbit_r4_c95 bl_95 br_95 wl_4 vdd gnd cell_6t
Xbit_r5_c95 bl_95 br_95 wl_5 vdd gnd cell_6t
Xbit_r6_c95 bl_95 br_95 wl_6 vdd gnd cell_6t
Xbit_r7_c95 bl_95 br_95 wl_7 vdd gnd cell_6t
Xbit_r8_c95 bl_95 br_95 wl_8 vdd gnd cell_6t
Xbit_r9_c95 bl_95 br_95 wl_9 vdd gnd cell_6t
Xbit_r10_c95 bl_95 br_95 wl_10 vdd gnd cell_6t
Xbit_r11_c95 bl_95 br_95 wl_11 vdd gnd cell_6t
Xbit_r12_c95 bl_95 br_95 wl_12 vdd gnd cell_6t
Xbit_r13_c95 bl_95 br_95 wl_13 vdd gnd cell_6t
Xbit_r14_c95 bl_95 br_95 wl_14 vdd gnd cell_6t
Xbit_r15_c95 bl_95 br_95 wl_15 vdd gnd cell_6t
Xbit_r16_c95 bl_95 br_95 wl_16 vdd gnd cell_6t
Xbit_r17_c95 bl_95 br_95 wl_17 vdd gnd cell_6t
Xbit_r18_c95 bl_95 br_95 wl_18 vdd gnd cell_6t
Xbit_r19_c95 bl_95 br_95 wl_19 vdd gnd cell_6t
Xbit_r20_c95 bl_95 br_95 wl_20 vdd gnd cell_6t
Xbit_r21_c95 bl_95 br_95 wl_21 vdd gnd cell_6t
Xbit_r22_c95 bl_95 br_95 wl_22 vdd gnd cell_6t
Xbit_r23_c95 bl_95 br_95 wl_23 vdd gnd cell_6t
Xbit_r24_c95 bl_95 br_95 wl_24 vdd gnd cell_6t
Xbit_r25_c95 bl_95 br_95 wl_25 vdd gnd cell_6t
Xbit_r26_c95 bl_95 br_95 wl_26 vdd gnd cell_6t
Xbit_r27_c95 bl_95 br_95 wl_27 vdd gnd cell_6t
Xbit_r28_c95 bl_95 br_95 wl_28 vdd gnd cell_6t
Xbit_r29_c95 bl_95 br_95 wl_29 vdd gnd cell_6t
Xbit_r30_c95 bl_95 br_95 wl_30 vdd gnd cell_6t
Xbit_r31_c95 bl_95 br_95 wl_31 vdd gnd cell_6t
Xbit_r32_c95 bl_95 br_95 wl_32 vdd gnd cell_6t
Xbit_r33_c95 bl_95 br_95 wl_33 vdd gnd cell_6t
Xbit_r34_c95 bl_95 br_95 wl_34 vdd gnd cell_6t
Xbit_r35_c95 bl_95 br_95 wl_35 vdd gnd cell_6t
Xbit_r36_c95 bl_95 br_95 wl_36 vdd gnd cell_6t
Xbit_r37_c95 bl_95 br_95 wl_37 vdd gnd cell_6t
Xbit_r38_c95 bl_95 br_95 wl_38 vdd gnd cell_6t
Xbit_r39_c95 bl_95 br_95 wl_39 vdd gnd cell_6t
Xbit_r40_c95 bl_95 br_95 wl_40 vdd gnd cell_6t
Xbit_r41_c95 bl_95 br_95 wl_41 vdd gnd cell_6t
Xbit_r42_c95 bl_95 br_95 wl_42 vdd gnd cell_6t
Xbit_r43_c95 bl_95 br_95 wl_43 vdd gnd cell_6t
Xbit_r44_c95 bl_95 br_95 wl_44 vdd gnd cell_6t
Xbit_r45_c95 bl_95 br_95 wl_45 vdd gnd cell_6t
Xbit_r46_c95 bl_95 br_95 wl_46 vdd gnd cell_6t
Xbit_r47_c95 bl_95 br_95 wl_47 vdd gnd cell_6t
Xbit_r48_c95 bl_95 br_95 wl_48 vdd gnd cell_6t
Xbit_r49_c95 bl_95 br_95 wl_49 vdd gnd cell_6t
Xbit_r50_c95 bl_95 br_95 wl_50 vdd gnd cell_6t
Xbit_r51_c95 bl_95 br_95 wl_51 vdd gnd cell_6t
Xbit_r52_c95 bl_95 br_95 wl_52 vdd gnd cell_6t
Xbit_r53_c95 bl_95 br_95 wl_53 vdd gnd cell_6t
Xbit_r54_c95 bl_95 br_95 wl_54 vdd gnd cell_6t
Xbit_r55_c95 bl_95 br_95 wl_55 vdd gnd cell_6t
Xbit_r56_c95 bl_95 br_95 wl_56 vdd gnd cell_6t
Xbit_r57_c95 bl_95 br_95 wl_57 vdd gnd cell_6t
Xbit_r58_c95 bl_95 br_95 wl_58 vdd gnd cell_6t
Xbit_r59_c95 bl_95 br_95 wl_59 vdd gnd cell_6t
Xbit_r60_c95 bl_95 br_95 wl_60 vdd gnd cell_6t
Xbit_r61_c95 bl_95 br_95 wl_61 vdd gnd cell_6t
Xbit_r62_c95 bl_95 br_95 wl_62 vdd gnd cell_6t
Xbit_r63_c95 bl_95 br_95 wl_63 vdd gnd cell_6t
Xbit_r64_c95 bl_95 br_95 wl_64 vdd gnd cell_6t
Xbit_r65_c95 bl_95 br_95 wl_65 vdd gnd cell_6t
Xbit_r66_c95 bl_95 br_95 wl_66 vdd gnd cell_6t
Xbit_r67_c95 bl_95 br_95 wl_67 vdd gnd cell_6t
Xbit_r68_c95 bl_95 br_95 wl_68 vdd gnd cell_6t
Xbit_r69_c95 bl_95 br_95 wl_69 vdd gnd cell_6t
Xbit_r70_c95 bl_95 br_95 wl_70 vdd gnd cell_6t
Xbit_r71_c95 bl_95 br_95 wl_71 vdd gnd cell_6t
Xbit_r72_c95 bl_95 br_95 wl_72 vdd gnd cell_6t
Xbit_r73_c95 bl_95 br_95 wl_73 vdd gnd cell_6t
Xbit_r74_c95 bl_95 br_95 wl_74 vdd gnd cell_6t
Xbit_r75_c95 bl_95 br_95 wl_75 vdd gnd cell_6t
Xbit_r76_c95 bl_95 br_95 wl_76 vdd gnd cell_6t
Xbit_r77_c95 bl_95 br_95 wl_77 vdd gnd cell_6t
Xbit_r78_c95 bl_95 br_95 wl_78 vdd gnd cell_6t
Xbit_r79_c95 bl_95 br_95 wl_79 vdd gnd cell_6t
Xbit_r80_c95 bl_95 br_95 wl_80 vdd gnd cell_6t
Xbit_r81_c95 bl_95 br_95 wl_81 vdd gnd cell_6t
Xbit_r82_c95 bl_95 br_95 wl_82 vdd gnd cell_6t
Xbit_r83_c95 bl_95 br_95 wl_83 vdd gnd cell_6t
Xbit_r84_c95 bl_95 br_95 wl_84 vdd gnd cell_6t
Xbit_r85_c95 bl_95 br_95 wl_85 vdd gnd cell_6t
Xbit_r86_c95 bl_95 br_95 wl_86 vdd gnd cell_6t
Xbit_r87_c95 bl_95 br_95 wl_87 vdd gnd cell_6t
Xbit_r88_c95 bl_95 br_95 wl_88 vdd gnd cell_6t
Xbit_r89_c95 bl_95 br_95 wl_89 vdd gnd cell_6t
Xbit_r90_c95 bl_95 br_95 wl_90 vdd gnd cell_6t
Xbit_r91_c95 bl_95 br_95 wl_91 vdd gnd cell_6t
Xbit_r92_c95 bl_95 br_95 wl_92 vdd gnd cell_6t
Xbit_r93_c95 bl_95 br_95 wl_93 vdd gnd cell_6t
Xbit_r94_c95 bl_95 br_95 wl_94 vdd gnd cell_6t
Xbit_r95_c95 bl_95 br_95 wl_95 vdd gnd cell_6t
Xbit_r96_c95 bl_95 br_95 wl_96 vdd gnd cell_6t
Xbit_r97_c95 bl_95 br_95 wl_97 vdd gnd cell_6t
Xbit_r98_c95 bl_95 br_95 wl_98 vdd gnd cell_6t
Xbit_r99_c95 bl_95 br_95 wl_99 vdd gnd cell_6t
Xbit_r100_c95 bl_95 br_95 wl_100 vdd gnd cell_6t
Xbit_r101_c95 bl_95 br_95 wl_101 vdd gnd cell_6t
Xbit_r102_c95 bl_95 br_95 wl_102 vdd gnd cell_6t
Xbit_r103_c95 bl_95 br_95 wl_103 vdd gnd cell_6t
Xbit_r104_c95 bl_95 br_95 wl_104 vdd gnd cell_6t
Xbit_r105_c95 bl_95 br_95 wl_105 vdd gnd cell_6t
Xbit_r106_c95 bl_95 br_95 wl_106 vdd gnd cell_6t
Xbit_r107_c95 bl_95 br_95 wl_107 vdd gnd cell_6t
Xbit_r108_c95 bl_95 br_95 wl_108 vdd gnd cell_6t
Xbit_r109_c95 bl_95 br_95 wl_109 vdd gnd cell_6t
Xbit_r110_c95 bl_95 br_95 wl_110 vdd gnd cell_6t
Xbit_r111_c95 bl_95 br_95 wl_111 vdd gnd cell_6t
Xbit_r112_c95 bl_95 br_95 wl_112 vdd gnd cell_6t
Xbit_r113_c95 bl_95 br_95 wl_113 vdd gnd cell_6t
Xbit_r114_c95 bl_95 br_95 wl_114 vdd gnd cell_6t
Xbit_r115_c95 bl_95 br_95 wl_115 vdd gnd cell_6t
Xbit_r116_c95 bl_95 br_95 wl_116 vdd gnd cell_6t
Xbit_r117_c95 bl_95 br_95 wl_117 vdd gnd cell_6t
Xbit_r118_c95 bl_95 br_95 wl_118 vdd gnd cell_6t
Xbit_r119_c95 bl_95 br_95 wl_119 vdd gnd cell_6t
Xbit_r120_c95 bl_95 br_95 wl_120 vdd gnd cell_6t
Xbit_r121_c95 bl_95 br_95 wl_121 vdd gnd cell_6t
Xbit_r122_c95 bl_95 br_95 wl_122 vdd gnd cell_6t
Xbit_r123_c95 bl_95 br_95 wl_123 vdd gnd cell_6t
Xbit_r124_c95 bl_95 br_95 wl_124 vdd gnd cell_6t
Xbit_r125_c95 bl_95 br_95 wl_125 vdd gnd cell_6t
Xbit_r126_c95 bl_95 br_95 wl_126 vdd gnd cell_6t
Xbit_r127_c95 bl_95 br_95 wl_127 vdd gnd cell_6t
Xbit_r128_c95 bl_95 br_95 wl_128 vdd gnd cell_6t
Xbit_r129_c95 bl_95 br_95 wl_129 vdd gnd cell_6t
Xbit_r130_c95 bl_95 br_95 wl_130 vdd gnd cell_6t
Xbit_r131_c95 bl_95 br_95 wl_131 vdd gnd cell_6t
Xbit_r132_c95 bl_95 br_95 wl_132 vdd gnd cell_6t
Xbit_r133_c95 bl_95 br_95 wl_133 vdd gnd cell_6t
Xbit_r134_c95 bl_95 br_95 wl_134 vdd gnd cell_6t
Xbit_r135_c95 bl_95 br_95 wl_135 vdd gnd cell_6t
Xbit_r136_c95 bl_95 br_95 wl_136 vdd gnd cell_6t
Xbit_r137_c95 bl_95 br_95 wl_137 vdd gnd cell_6t
Xbit_r138_c95 bl_95 br_95 wl_138 vdd gnd cell_6t
Xbit_r139_c95 bl_95 br_95 wl_139 vdd gnd cell_6t
Xbit_r140_c95 bl_95 br_95 wl_140 vdd gnd cell_6t
Xbit_r141_c95 bl_95 br_95 wl_141 vdd gnd cell_6t
Xbit_r142_c95 bl_95 br_95 wl_142 vdd gnd cell_6t
Xbit_r143_c95 bl_95 br_95 wl_143 vdd gnd cell_6t
Xbit_r144_c95 bl_95 br_95 wl_144 vdd gnd cell_6t
Xbit_r145_c95 bl_95 br_95 wl_145 vdd gnd cell_6t
Xbit_r146_c95 bl_95 br_95 wl_146 vdd gnd cell_6t
Xbit_r147_c95 bl_95 br_95 wl_147 vdd gnd cell_6t
Xbit_r148_c95 bl_95 br_95 wl_148 vdd gnd cell_6t
Xbit_r149_c95 bl_95 br_95 wl_149 vdd gnd cell_6t
Xbit_r150_c95 bl_95 br_95 wl_150 vdd gnd cell_6t
Xbit_r151_c95 bl_95 br_95 wl_151 vdd gnd cell_6t
Xbit_r152_c95 bl_95 br_95 wl_152 vdd gnd cell_6t
Xbit_r153_c95 bl_95 br_95 wl_153 vdd gnd cell_6t
Xbit_r154_c95 bl_95 br_95 wl_154 vdd gnd cell_6t
Xbit_r155_c95 bl_95 br_95 wl_155 vdd gnd cell_6t
Xbit_r156_c95 bl_95 br_95 wl_156 vdd gnd cell_6t
Xbit_r157_c95 bl_95 br_95 wl_157 vdd gnd cell_6t
Xbit_r158_c95 bl_95 br_95 wl_158 vdd gnd cell_6t
Xbit_r159_c95 bl_95 br_95 wl_159 vdd gnd cell_6t
Xbit_r160_c95 bl_95 br_95 wl_160 vdd gnd cell_6t
Xbit_r161_c95 bl_95 br_95 wl_161 vdd gnd cell_6t
Xbit_r162_c95 bl_95 br_95 wl_162 vdd gnd cell_6t
Xbit_r163_c95 bl_95 br_95 wl_163 vdd gnd cell_6t
Xbit_r164_c95 bl_95 br_95 wl_164 vdd gnd cell_6t
Xbit_r165_c95 bl_95 br_95 wl_165 vdd gnd cell_6t
Xbit_r166_c95 bl_95 br_95 wl_166 vdd gnd cell_6t
Xbit_r167_c95 bl_95 br_95 wl_167 vdd gnd cell_6t
Xbit_r168_c95 bl_95 br_95 wl_168 vdd gnd cell_6t
Xbit_r169_c95 bl_95 br_95 wl_169 vdd gnd cell_6t
Xbit_r170_c95 bl_95 br_95 wl_170 vdd gnd cell_6t
Xbit_r171_c95 bl_95 br_95 wl_171 vdd gnd cell_6t
Xbit_r172_c95 bl_95 br_95 wl_172 vdd gnd cell_6t
Xbit_r173_c95 bl_95 br_95 wl_173 vdd gnd cell_6t
Xbit_r174_c95 bl_95 br_95 wl_174 vdd gnd cell_6t
Xbit_r175_c95 bl_95 br_95 wl_175 vdd gnd cell_6t
Xbit_r176_c95 bl_95 br_95 wl_176 vdd gnd cell_6t
Xbit_r177_c95 bl_95 br_95 wl_177 vdd gnd cell_6t
Xbit_r178_c95 bl_95 br_95 wl_178 vdd gnd cell_6t
Xbit_r179_c95 bl_95 br_95 wl_179 vdd gnd cell_6t
Xbit_r180_c95 bl_95 br_95 wl_180 vdd gnd cell_6t
Xbit_r181_c95 bl_95 br_95 wl_181 vdd gnd cell_6t
Xbit_r182_c95 bl_95 br_95 wl_182 vdd gnd cell_6t
Xbit_r183_c95 bl_95 br_95 wl_183 vdd gnd cell_6t
Xbit_r184_c95 bl_95 br_95 wl_184 vdd gnd cell_6t
Xbit_r185_c95 bl_95 br_95 wl_185 vdd gnd cell_6t
Xbit_r186_c95 bl_95 br_95 wl_186 vdd gnd cell_6t
Xbit_r187_c95 bl_95 br_95 wl_187 vdd gnd cell_6t
Xbit_r188_c95 bl_95 br_95 wl_188 vdd gnd cell_6t
Xbit_r189_c95 bl_95 br_95 wl_189 vdd gnd cell_6t
Xbit_r190_c95 bl_95 br_95 wl_190 vdd gnd cell_6t
Xbit_r191_c95 bl_95 br_95 wl_191 vdd gnd cell_6t
Xbit_r192_c95 bl_95 br_95 wl_192 vdd gnd cell_6t
Xbit_r193_c95 bl_95 br_95 wl_193 vdd gnd cell_6t
Xbit_r194_c95 bl_95 br_95 wl_194 vdd gnd cell_6t
Xbit_r195_c95 bl_95 br_95 wl_195 vdd gnd cell_6t
Xbit_r196_c95 bl_95 br_95 wl_196 vdd gnd cell_6t
Xbit_r197_c95 bl_95 br_95 wl_197 vdd gnd cell_6t
Xbit_r198_c95 bl_95 br_95 wl_198 vdd gnd cell_6t
Xbit_r199_c95 bl_95 br_95 wl_199 vdd gnd cell_6t
Xbit_r200_c95 bl_95 br_95 wl_200 vdd gnd cell_6t
Xbit_r201_c95 bl_95 br_95 wl_201 vdd gnd cell_6t
Xbit_r202_c95 bl_95 br_95 wl_202 vdd gnd cell_6t
Xbit_r203_c95 bl_95 br_95 wl_203 vdd gnd cell_6t
Xbit_r204_c95 bl_95 br_95 wl_204 vdd gnd cell_6t
Xbit_r205_c95 bl_95 br_95 wl_205 vdd gnd cell_6t
Xbit_r206_c95 bl_95 br_95 wl_206 vdd gnd cell_6t
Xbit_r207_c95 bl_95 br_95 wl_207 vdd gnd cell_6t
Xbit_r208_c95 bl_95 br_95 wl_208 vdd gnd cell_6t
Xbit_r209_c95 bl_95 br_95 wl_209 vdd gnd cell_6t
Xbit_r210_c95 bl_95 br_95 wl_210 vdd gnd cell_6t
Xbit_r211_c95 bl_95 br_95 wl_211 vdd gnd cell_6t
Xbit_r212_c95 bl_95 br_95 wl_212 vdd gnd cell_6t
Xbit_r213_c95 bl_95 br_95 wl_213 vdd gnd cell_6t
Xbit_r214_c95 bl_95 br_95 wl_214 vdd gnd cell_6t
Xbit_r215_c95 bl_95 br_95 wl_215 vdd gnd cell_6t
Xbit_r216_c95 bl_95 br_95 wl_216 vdd gnd cell_6t
Xbit_r217_c95 bl_95 br_95 wl_217 vdd gnd cell_6t
Xbit_r218_c95 bl_95 br_95 wl_218 vdd gnd cell_6t
Xbit_r219_c95 bl_95 br_95 wl_219 vdd gnd cell_6t
Xbit_r220_c95 bl_95 br_95 wl_220 vdd gnd cell_6t
Xbit_r221_c95 bl_95 br_95 wl_221 vdd gnd cell_6t
Xbit_r222_c95 bl_95 br_95 wl_222 vdd gnd cell_6t
Xbit_r223_c95 bl_95 br_95 wl_223 vdd gnd cell_6t
Xbit_r224_c95 bl_95 br_95 wl_224 vdd gnd cell_6t
Xbit_r225_c95 bl_95 br_95 wl_225 vdd gnd cell_6t
Xbit_r226_c95 bl_95 br_95 wl_226 vdd gnd cell_6t
Xbit_r227_c95 bl_95 br_95 wl_227 vdd gnd cell_6t
Xbit_r228_c95 bl_95 br_95 wl_228 vdd gnd cell_6t
Xbit_r229_c95 bl_95 br_95 wl_229 vdd gnd cell_6t
Xbit_r230_c95 bl_95 br_95 wl_230 vdd gnd cell_6t
Xbit_r231_c95 bl_95 br_95 wl_231 vdd gnd cell_6t
Xbit_r232_c95 bl_95 br_95 wl_232 vdd gnd cell_6t
Xbit_r233_c95 bl_95 br_95 wl_233 vdd gnd cell_6t
Xbit_r234_c95 bl_95 br_95 wl_234 vdd gnd cell_6t
Xbit_r235_c95 bl_95 br_95 wl_235 vdd gnd cell_6t
Xbit_r236_c95 bl_95 br_95 wl_236 vdd gnd cell_6t
Xbit_r237_c95 bl_95 br_95 wl_237 vdd gnd cell_6t
Xbit_r238_c95 bl_95 br_95 wl_238 vdd gnd cell_6t
Xbit_r239_c95 bl_95 br_95 wl_239 vdd gnd cell_6t
Xbit_r240_c95 bl_95 br_95 wl_240 vdd gnd cell_6t
Xbit_r241_c95 bl_95 br_95 wl_241 vdd gnd cell_6t
Xbit_r242_c95 bl_95 br_95 wl_242 vdd gnd cell_6t
Xbit_r243_c95 bl_95 br_95 wl_243 vdd gnd cell_6t
Xbit_r244_c95 bl_95 br_95 wl_244 vdd gnd cell_6t
Xbit_r245_c95 bl_95 br_95 wl_245 vdd gnd cell_6t
Xbit_r246_c95 bl_95 br_95 wl_246 vdd gnd cell_6t
Xbit_r247_c95 bl_95 br_95 wl_247 vdd gnd cell_6t
Xbit_r248_c95 bl_95 br_95 wl_248 vdd gnd cell_6t
Xbit_r249_c95 bl_95 br_95 wl_249 vdd gnd cell_6t
Xbit_r250_c95 bl_95 br_95 wl_250 vdd gnd cell_6t
Xbit_r251_c95 bl_95 br_95 wl_251 vdd gnd cell_6t
Xbit_r252_c95 bl_95 br_95 wl_252 vdd gnd cell_6t
Xbit_r253_c95 bl_95 br_95 wl_253 vdd gnd cell_6t
Xbit_r254_c95 bl_95 br_95 wl_254 vdd gnd cell_6t
Xbit_r255_c95 bl_95 br_95 wl_255 vdd gnd cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd cell_6t
Xbit_r1_c96 bl_96 br_96 wl_1 vdd gnd cell_6t
Xbit_r2_c96 bl_96 br_96 wl_2 vdd gnd cell_6t
Xbit_r3_c96 bl_96 br_96 wl_3 vdd gnd cell_6t
Xbit_r4_c96 bl_96 br_96 wl_4 vdd gnd cell_6t
Xbit_r5_c96 bl_96 br_96 wl_5 vdd gnd cell_6t
Xbit_r6_c96 bl_96 br_96 wl_6 vdd gnd cell_6t
Xbit_r7_c96 bl_96 br_96 wl_7 vdd gnd cell_6t
Xbit_r8_c96 bl_96 br_96 wl_8 vdd gnd cell_6t
Xbit_r9_c96 bl_96 br_96 wl_9 vdd gnd cell_6t
Xbit_r10_c96 bl_96 br_96 wl_10 vdd gnd cell_6t
Xbit_r11_c96 bl_96 br_96 wl_11 vdd gnd cell_6t
Xbit_r12_c96 bl_96 br_96 wl_12 vdd gnd cell_6t
Xbit_r13_c96 bl_96 br_96 wl_13 vdd gnd cell_6t
Xbit_r14_c96 bl_96 br_96 wl_14 vdd gnd cell_6t
Xbit_r15_c96 bl_96 br_96 wl_15 vdd gnd cell_6t
Xbit_r16_c96 bl_96 br_96 wl_16 vdd gnd cell_6t
Xbit_r17_c96 bl_96 br_96 wl_17 vdd gnd cell_6t
Xbit_r18_c96 bl_96 br_96 wl_18 vdd gnd cell_6t
Xbit_r19_c96 bl_96 br_96 wl_19 vdd gnd cell_6t
Xbit_r20_c96 bl_96 br_96 wl_20 vdd gnd cell_6t
Xbit_r21_c96 bl_96 br_96 wl_21 vdd gnd cell_6t
Xbit_r22_c96 bl_96 br_96 wl_22 vdd gnd cell_6t
Xbit_r23_c96 bl_96 br_96 wl_23 vdd gnd cell_6t
Xbit_r24_c96 bl_96 br_96 wl_24 vdd gnd cell_6t
Xbit_r25_c96 bl_96 br_96 wl_25 vdd gnd cell_6t
Xbit_r26_c96 bl_96 br_96 wl_26 vdd gnd cell_6t
Xbit_r27_c96 bl_96 br_96 wl_27 vdd gnd cell_6t
Xbit_r28_c96 bl_96 br_96 wl_28 vdd gnd cell_6t
Xbit_r29_c96 bl_96 br_96 wl_29 vdd gnd cell_6t
Xbit_r30_c96 bl_96 br_96 wl_30 vdd gnd cell_6t
Xbit_r31_c96 bl_96 br_96 wl_31 vdd gnd cell_6t
Xbit_r32_c96 bl_96 br_96 wl_32 vdd gnd cell_6t
Xbit_r33_c96 bl_96 br_96 wl_33 vdd gnd cell_6t
Xbit_r34_c96 bl_96 br_96 wl_34 vdd gnd cell_6t
Xbit_r35_c96 bl_96 br_96 wl_35 vdd gnd cell_6t
Xbit_r36_c96 bl_96 br_96 wl_36 vdd gnd cell_6t
Xbit_r37_c96 bl_96 br_96 wl_37 vdd gnd cell_6t
Xbit_r38_c96 bl_96 br_96 wl_38 vdd gnd cell_6t
Xbit_r39_c96 bl_96 br_96 wl_39 vdd gnd cell_6t
Xbit_r40_c96 bl_96 br_96 wl_40 vdd gnd cell_6t
Xbit_r41_c96 bl_96 br_96 wl_41 vdd gnd cell_6t
Xbit_r42_c96 bl_96 br_96 wl_42 vdd gnd cell_6t
Xbit_r43_c96 bl_96 br_96 wl_43 vdd gnd cell_6t
Xbit_r44_c96 bl_96 br_96 wl_44 vdd gnd cell_6t
Xbit_r45_c96 bl_96 br_96 wl_45 vdd gnd cell_6t
Xbit_r46_c96 bl_96 br_96 wl_46 vdd gnd cell_6t
Xbit_r47_c96 bl_96 br_96 wl_47 vdd gnd cell_6t
Xbit_r48_c96 bl_96 br_96 wl_48 vdd gnd cell_6t
Xbit_r49_c96 bl_96 br_96 wl_49 vdd gnd cell_6t
Xbit_r50_c96 bl_96 br_96 wl_50 vdd gnd cell_6t
Xbit_r51_c96 bl_96 br_96 wl_51 vdd gnd cell_6t
Xbit_r52_c96 bl_96 br_96 wl_52 vdd gnd cell_6t
Xbit_r53_c96 bl_96 br_96 wl_53 vdd gnd cell_6t
Xbit_r54_c96 bl_96 br_96 wl_54 vdd gnd cell_6t
Xbit_r55_c96 bl_96 br_96 wl_55 vdd gnd cell_6t
Xbit_r56_c96 bl_96 br_96 wl_56 vdd gnd cell_6t
Xbit_r57_c96 bl_96 br_96 wl_57 vdd gnd cell_6t
Xbit_r58_c96 bl_96 br_96 wl_58 vdd gnd cell_6t
Xbit_r59_c96 bl_96 br_96 wl_59 vdd gnd cell_6t
Xbit_r60_c96 bl_96 br_96 wl_60 vdd gnd cell_6t
Xbit_r61_c96 bl_96 br_96 wl_61 vdd gnd cell_6t
Xbit_r62_c96 bl_96 br_96 wl_62 vdd gnd cell_6t
Xbit_r63_c96 bl_96 br_96 wl_63 vdd gnd cell_6t
Xbit_r64_c96 bl_96 br_96 wl_64 vdd gnd cell_6t
Xbit_r65_c96 bl_96 br_96 wl_65 vdd gnd cell_6t
Xbit_r66_c96 bl_96 br_96 wl_66 vdd gnd cell_6t
Xbit_r67_c96 bl_96 br_96 wl_67 vdd gnd cell_6t
Xbit_r68_c96 bl_96 br_96 wl_68 vdd gnd cell_6t
Xbit_r69_c96 bl_96 br_96 wl_69 vdd gnd cell_6t
Xbit_r70_c96 bl_96 br_96 wl_70 vdd gnd cell_6t
Xbit_r71_c96 bl_96 br_96 wl_71 vdd gnd cell_6t
Xbit_r72_c96 bl_96 br_96 wl_72 vdd gnd cell_6t
Xbit_r73_c96 bl_96 br_96 wl_73 vdd gnd cell_6t
Xbit_r74_c96 bl_96 br_96 wl_74 vdd gnd cell_6t
Xbit_r75_c96 bl_96 br_96 wl_75 vdd gnd cell_6t
Xbit_r76_c96 bl_96 br_96 wl_76 vdd gnd cell_6t
Xbit_r77_c96 bl_96 br_96 wl_77 vdd gnd cell_6t
Xbit_r78_c96 bl_96 br_96 wl_78 vdd gnd cell_6t
Xbit_r79_c96 bl_96 br_96 wl_79 vdd gnd cell_6t
Xbit_r80_c96 bl_96 br_96 wl_80 vdd gnd cell_6t
Xbit_r81_c96 bl_96 br_96 wl_81 vdd gnd cell_6t
Xbit_r82_c96 bl_96 br_96 wl_82 vdd gnd cell_6t
Xbit_r83_c96 bl_96 br_96 wl_83 vdd gnd cell_6t
Xbit_r84_c96 bl_96 br_96 wl_84 vdd gnd cell_6t
Xbit_r85_c96 bl_96 br_96 wl_85 vdd gnd cell_6t
Xbit_r86_c96 bl_96 br_96 wl_86 vdd gnd cell_6t
Xbit_r87_c96 bl_96 br_96 wl_87 vdd gnd cell_6t
Xbit_r88_c96 bl_96 br_96 wl_88 vdd gnd cell_6t
Xbit_r89_c96 bl_96 br_96 wl_89 vdd gnd cell_6t
Xbit_r90_c96 bl_96 br_96 wl_90 vdd gnd cell_6t
Xbit_r91_c96 bl_96 br_96 wl_91 vdd gnd cell_6t
Xbit_r92_c96 bl_96 br_96 wl_92 vdd gnd cell_6t
Xbit_r93_c96 bl_96 br_96 wl_93 vdd gnd cell_6t
Xbit_r94_c96 bl_96 br_96 wl_94 vdd gnd cell_6t
Xbit_r95_c96 bl_96 br_96 wl_95 vdd gnd cell_6t
Xbit_r96_c96 bl_96 br_96 wl_96 vdd gnd cell_6t
Xbit_r97_c96 bl_96 br_96 wl_97 vdd gnd cell_6t
Xbit_r98_c96 bl_96 br_96 wl_98 vdd gnd cell_6t
Xbit_r99_c96 bl_96 br_96 wl_99 vdd gnd cell_6t
Xbit_r100_c96 bl_96 br_96 wl_100 vdd gnd cell_6t
Xbit_r101_c96 bl_96 br_96 wl_101 vdd gnd cell_6t
Xbit_r102_c96 bl_96 br_96 wl_102 vdd gnd cell_6t
Xbit_r103_c96 bl_96 br_96 wl_103 vdd gnd cell_6t
Xbit_r104_c96 bl_96 br_96 wl_104 vdd gnd cell_6t
Xbit_r105_c96 bl_96 br_96 wl_105 vdd gnd cell_6t
Xbit_r106_c96 bl_96 br_96 wl_106 vdd gnd cell_6t
Xbit_r107_c96 bl_96 br_96 wl_107 vdd gnd cell_6t
Xbit_r108_c96 bl_96 br_96 wl_108 vdd gnd cell_6t
Xbit_r109_c96 bl_96 br_96 wl_109 vdd gnd cell_6t
Xbit_r110_c96 bl_96 br_96 wl_110 vdd gnd cell_6t
Xbit_r111_c96 bl_96 br_96 wl_111 vdd gnd cell_6t
Xbit_r112_c96 bl_96 br_96 wl_112 vdd gnd cell_6t
Xbit_r113_c96 bl_96 br_96 wl_113 vdd gnd cell_6t
Xbit_r114_c96 bl_96 br_96 wl_114 vdd gnd cell_6t
Xbit_r115_c96 bl_96 br_96 wl_115 vdd gnd cell_6t
Xbit_r116_c96 bl_96 br_96 wl_116 vdd gnd cell_6t
Xbit_r117_c96 bl_96 br_96 wl_117 vdd gnd cell_6t
Xbit_r118_c96 bl_96 br_96 wl_118 vdd gnd cell_6t
Xbit_r119_c96 bl_96 br_96 wl_119 vdd gnd cell_6t
Xbit_r120_c96 bl_96 br_96 wl_120 vdd gnd cell_6t
Xbit_r121_c96 bl_96 br_96 wl_121 vdd gnd cell_6t
Xbit_r122_c96 bl_96 br_96 wl_122 vdd gnd cell_6t
Xbit_r123_c96 bl_96 br_96 wl_123 vdd gnd cell_6t
Xbit_r124_c96 bl_96 br_96 wl_124 vdd gnd cell_6t
Xbit_r125_c96 bl_96 br_96 wl_125 vdd gnd cell_6t
Xbit_r126_c96 bl_96 br_96 wl_126 vdd gnd cell_6t
Xbit_r127_c96 bl_96 br_96 wl_127 vdd gnd cell_6t
Xbit_r128_c96 bl_96 br_96 wl_128 vdd gnd cell_6t
Xbit_r129_c96 bl_96 br_96 wl_129 vdd gnd cell_6t
Xbit_r130_c96 bl_96 br_96 wl_130 vdd gnd cell_6t
Xbit_r131_c96 bl_96 br_96 wl_131 vdd gnd cell_6t
Xbit_r132_c96 bl_96 br_96 wl_132 vdd gnd cell_6t
Xbit_r133_c96 bl_96 br_96 wl_133 vdd gnd cell_6t
Xbit_r134_c96 bl_96 br_96 wl_134 vdd gnd cell_6t
Xbit_r135_c96 bl_96 br_96 wl_135 vdd gnd cell_6t
Xbit_r136_c96 bl_96 br_96 wl_136 vdd gnd cell_6t
Xbit_r137_c96 bl_96 br_96 wl_137 vdd gnd cell_6t
Xbit_r138_c96 bl_96 br_96 wl_138 vdd gnd cell_6t
Xbit_r139_c96 bl_96 br_96 wl_139 vdd gnd cell_6t
Xbit_r140_c96 bl_96 br_96 wl_140 vdd gnd cell_6t
Xbit_r141_c96 bl_96 br_96 wl_141 vdd gnd cell_6t
Xbit_r142_c96 bl_96 br_96 wl_142 vdd gnd cell_6t
Xbit_r143_c96 bl_96 br_96 wl_143 vdd gnd cell_6t
Xbit_r144_c96 bl_96 br_96 wl_144 vdd gnd cell_6t
Xbit_r145_c96 bl_96 br_96 wl_145 vdd gnd cell_6t
Xbit_r146_c96 bl_96 br_96 wl_146 vdd gnd cell_6t
Xbit_r147_c96 bl_96 br_96 wl_147 vdd gnd cell_6t
Xbit_r148_c96 bl_96 br_96 wl_148 vdd gnd cell_6t
Xbit_r149_c96 bl_96 br_96 wl_149 vdd gnd cell_6t
Xbit_r150_c96 bl_96 br_96 wl_150 vdd gnd cell_6t
Xbit_r151_c96 bl_96 br_96 wl_151 vdd gnd cell_6t
Xbit_r152_c96 bl_96 br_96 wl_152 vdd gnd cell_6t
Xbit_r153_c96 bl_96 br_96 wl_153 vdd gnd cell_6t
Xbit_r154_c96 bl_96 br_96 wl_154 vdd gnd cell_6t
Xbit_r155_c96 bl_96 br_96 wl_155 vdd gnd cell_6t
Xbit_r156_c96 bl_96 br_96 wl_156 vdd gnd cell_6t
Xbit_r157_c96 bl_96 br_96 wl_157 vdd gnd cell_6t
Xbit_r158_c96 bl_96 br_96 wl_158 vdd gnd cell_6t
Xbit_r159_c96 bl_96 br_96 wl_159 vdd gnd cell_6t
Xbit_r160_c96 bl_96 br_96 wl_160 vdd gnd cell_6t
Xbit_r161_c96 bl_96 br_96 wl_161 vdd gnd cell_6t
Xbit_r162_c96 bl_96 br_96 wl_162 vdd gnd cell_6t
Xbit_r163_c96 bl_96 br_96 wl_163 vdd gnd cell_6t
Xbit_r164_c96 bl_96 br_96 wl_164 vdd gnd cell_6t
Xbit_r165_c96 bl_96 br_96 wl_165 vdd gnd cell_6t
Xbit_r166_c96 bl_96 br_96 wl_166 vdd gnd cell_6t
Xbit_r167_c96 bl_96 br_96 wl_167 vdd gnd cell_6t
Xbit_r168_c96 bl_96 br_96 wl_168 vdd gnd cell_6t
Xbit_r169_c96 bl_96 br_96 wl_169 vdd gnd cell_6t
Xbit_r170_c96 bl_96 br_96 wl_170 vdd gnd cell_6t
Xbit_r171_c96 bl_96 br_96 wl_171 vdd gnd cell_6t
Xbit_r172_c96 bl_96 br_96 wl_172 vdd gnd cell_6t
Xbit_r173_c96 bl_96 br_96 wl_173 vdd gnd cell_6t
Xbit_r174_c96 bl_96 br_96 wl_174 vdd gnd cell_6t
Xbit_r175_c96 bl_96 br_96 wl_175 vdd gnd cell_6t
Xbit_r176_c96 bl_96 br_96 wl_176 vdd gnd cell_6t
Xbit_r177_c96 bl_96 br_96 wl_177 vdd gnd cell_6t
Xbit_r178_c96 bl_96 br_96 wl_178 vdd gnd cell_6t
Xbit_r179_c96 bl_96 br_96 wl_179 vdd gnd cell_6t
Xbit_r180_c96 bl_96 br_96 wl_180 vdd gnd cell_6t
Xbit_r181_c96 bl_96 br_96 wl_181 vdd gnd cell_6t
Xbit_r182_c96 bl_96 br_96 wl_182 vdd gnd cell_6t
Xbit_r183_c96 bl_96 br_96 wl_183 vdd gnd cell_6t
Xbit_r184_c96 bl_96 br_96 wl_184 vdd gnd cell_6t
Xbit_r185_c96 bl_96 br_96 wl_185 vdd gnd cell_6t
Xbit_r186_c96 bl_96 br_96 wl_186 vdd gnd cell_6t
Xbit_r187_c96 bl_96 br_96 wl_187 vdd gnd cell_6t
Xbit_r188_c96 bl_96 br_96 wl_188 vdd gnd cell_6t
Xbit_r189_c96 bl_96 br_96 wl_189 vdd gnd cell_6t
Xbit_r190_c96 bl_96 br_96 wl_190 vdd gnd cell_6t
Xbit_r191_c96 bl_96 br_96 wl_191 vdd gnd cell_6t
Xbit_r192_c96 bl_96 br_96 wl_192 vdd gnd cell_6t
Xbit_r193_c96 bl_96 br_96 wl_193 vdd gnd cell_6t
Xbit_r194_c96 bl_96 br_96 wl_194 vdd gnd cell_6t
Xbit_r195_c96 bl_96 br_96 wl_195 vdd gnd cell_6t
Xbit_r196_c96 bl_96 br_96 wl_196 vdd gnd cell_6t
Xbit_r197_c96 bl_96 br_96 wl_197 vdd gnd cell_6t
Xbit_r198_c96 bl_96 br_96 wl_198 vdd gnd cell_6t
Xbit_r199_c96 bl_96 br_96 wl_199 vdd gnd cell_6t
Xbit_r200_c96 bl_96 br_96 wl_200 vdd gnd cell_6t
Xbit_r201_c96 bl_96 br_96 wl_201 vdd gnd cell_6t
Xbit_r202_c96 bl_96 br_96 wl_202 vdd gnd cell_6t
Xbit_r203_c96 bl_96 br_96 wl_203 vdd gnd cell_6t
Xbit_r204_c96 bl_96 br_96 wl_204 vdd gnd cell_6t
Xbit_r205_c96 bl_96 br_96 wl_205 vdd gnd cell_6t
Xbit_r206_c96 bl_96 br_96 wl_206 vdd gnd cell_6t
Xbit_r207_c96 bl_96 br_96 wl_207 vdd gnd cell_6t
Xbit_r208_c96 bl_96 br_96 wl_208 vdd gnd cell_6t
Xbit_r209_c96 bl_96 br_96 wl_209 vdd gnd cell_6t
Xbit_r210_c96 bl_96 br_96 wl_210 vdd gnd cell_6t
Xbit_r211_c96 bl_96 br_96 wl_211 vdd gnd cell_6t
Xbit_r212_c96 bl_96 br_96 wl_212 vdd gnd cell_6t
Xbit_r213_c96 bl_96 br_96 wl_213 vdd gnd cell_6t
Xbit_r214_c96 bl_96 br_96 wl_214 vdd gnd cell_6t
Xbit_r215_c96 bl_96 br_96 wl_215 vdd gnd cell_6t
Xbit_r216_c96 bl_96 br_96 wl_216 vdd gnd cell_6t
Xbit_r217_c96 bl_96 br_96 wl_217 vdd gnd cell_6t
Xbit_r218_c96 bl_96 br_96 wl_218 vdd gnd cell_6t
Xbit_r219_c96 bl_96 br_96 wl_219 vdd gnd cell_6t
Xbit_r220_c96 bl_96 br_96 wl_220 vdd gnd cell_6t
Xbit_r221_c96 bl_96 br_96 wl_221 vdd gnd cell_6t
Xbit_r222_c96 bl_96 br_96 wl_222 vdd gnd cell_6t
Xbit_r223_c96 bl_96 br_96 wl_223 vdd gnd cell_6t
Xbit_r224_c96 bl_96 br_96 wl_224 vdd gnd cell_6t
Xbit_r225_c96 bl_96 br_96 wl_225 vdd gnd cell_6t
Xbit_r226_c96 bl_96 br_96 wl_226 vdd gnd cell_6t
Xbit_r227_c96 bl_96 br_96 wl_227 vdd gnd cell_6t
Xbit_r228_c96 bl_96 br_96 wl_228 vdd gnd cell_6t
Xbit_r229_c96 bl_96 br_96 wl_229 vdd gnd cell_6t
Xbit_r230_c96 bl_96 br_96 wl_230 vdd gnd cell_6t
Xbit_r231_c96 bl_96 br_96 wl_231 vdd gnd cell_6t
Xbit_r232_c96 bl_96 br_96 wl_232 vdd gnd cell_6t
Xbit_r233_c96 bl_96 br_96 wl_233 vdd gnd cell_6t
Xbit_r234_c96 bl_96 br_96 wl_234 vdd gnd cell_6t
Xbit_r235_c96 bl_96 br_96 wl_235 vdd gnd cell_6t
Xbit_r236_c96 bl_96 br_96 wl_236 vdd gnd cell_6t
Xbit_r237_c96 bl_96 br_96 wl_237 vdd gnd cell_6t
Xbit_r238_c96 bl_96 br_96 wl_238 vdd gnd cell_6t
Xbit_r239_c96 bl_96 br_96 wl_239 vdd gnd cell_6t
Xbit_r240_c96 bl_96 br_96 wl_240 vdd gnd cell_6t
Xbit_r241_c96 bl_96 br_96 wl_241 vdd gnd cell_6t
Xbit_r242_c96 bl_96 br_96 wl_242 vdd gnd cell_6t
Xbit_r243_c96 bl_96 br_96 wl_243 vdd gnd cell_6t
Xbit_r244_c96 bl_96 br_96 wl_244 vdd gnd cell_6t
Xbit_r245_c96 bl_96 br_96 wl_245 vdd gnd cell_6t
Xbit_r246_c96 bl_96 br_96 wl_246 vdd gnd cell_6t
Xbit_r247_c96 bl_96 br_96 wl_247 vdd gnd cell_6t
Xbit_r248_c96 bl_96 br_96 wl_248 vdd gnd cell_6t
Xbit_r249_c96 bl_96 br_96 wl_249 vdd gnd cell_6t
Xbit_r250_c96 bl_96 br_96 wl_250 vdd gnd cell_6t
Xbit_r251_c96 bl_96 br_96 wl_251 vdd gnd cell_6t
Xbit_r252_c96 bl_96 br_96 wl_252 vdd gnd cell_6t
Xbit_r253_c96 bl_96 br_96 wl_253 vdd gnd cell_6t
Xbit_r254_c96 bl_96 br_96 wl_254 vdd gnd cell_6t
Xbit_r255_c96 bl_96 br_96 wl_255 vdd gnd cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd cell_6t
Xbit_r1_c97 bl_97 br_97 wl_1 vdd gnd cell_6t
Xbit_r2_c97 bl_97 br_97 wl_2 vdd gnd cell_6t
Xbit_r3_c97 bl_97 br_97 wl_3 vdd gnd cell_6t
Xbit_r4_c97 bl_97 br_97 wl_4 vdd gnd cell_6t
Xbit_r5_c97 bl_97 br_97 wl_5 vdd gnd cell_6t
Xbit_r6_c97 bl_97 br_97 wl_6 vdd gnd cell_6t
Xbit_r7_c97 bl_97 br_97 wl_7 vdd gnd cell_6t
Xbit_r8_c97 bl_97 br_97 wl_8 vdd gnd cell_6t
Xbit_r9_c97 bl_97 br_97 wl_9 vdd gnd cell_6t
Xbit_r10_c97 bl_97 br_97 wl_10 vdd gnd cell_6t
Xbit_r11_c97 bl_97 br_97 wl_11 vdd gnd cell_6t
Xbit_r12_c97 bl_97 br_97 wl_12 vdd gnd cell_6t
Xbit_r13_c97 bl_97 br_97 wl_13 vdd gnd cell_6t
Xbit_r14_c97 bl_97 br_97 wl_14 vdd gnd cell_6t
Xbit_r15_c97 bl_97 br_97 wl_15 vdd gnd cell_6t
Xbit_r16_c97 bl_97 br_97 wl_16 vdd gnd cell_6t
Xbit_r17_c97 bl_97 br_97 wl_17 vdd gnd cell_6t
Xbit_r18_c97 bl_97 br_97 wl_18 vdd gnd cell_6t
Xbit_r19_c97 bl_97 br_97 wl_19 vdd gnd cell_6t
Xbit_r20_c97 bl_97 br_97 wl_20 vdd gnd cell_6t
Xbit_r21_c97 bl_97 br_97 wl_21 vdd gnd cell_6t
Xbit_r22_c97 bl_97 br_97 wl_22 vdd gnd cell_6t
Xbit_r23_c97 bl_97 br_97 wl_23 vdd gnd cell_6t
Xbit_r24_c97 bl_97 br_97 wl_24 vdd gnd cell_6t
Xbit_r25_c97 bl_97 br_97 wl_25 vdd gnd cell_6t
Xbit_r26_c97 bl_97 br_97 wl_26 vdd gnd cell_6t
Xbit_r27_c97 bl_97 br_97 wl_27 vdd gnd cell_6t
Xbit_r28_c97 bl_97 br_97 wl_28 vdd gnd cell_6t
Xbit_r29_c97 bl_97 br_97 wl_29 vdd gnd cell_6t
Xbit_r30_c97 bl_97 br_97 wl_30 vdd gnd cell_6t
Xbit_r31_c97 bl_97 br_97 wl_31 vdd gnd cell_6t
Xbit_r32_c97 bl_97 br_97 wl_32 vdd gnd cell_6t
Xbit_r33_c97 bl_97 br_97 wl_33 vdd gnd cell_6t
Xbit_r34_c97 bl_97 br_97 wl_34 vdd gnd cell_6t
Xbit_r35_c97 bl_97 br_97 wl_35 vdd gnd cell_6t
Xbit_r36_c97 bl_97 br_97 wl_36 vdd gnd cell_6t
Xbit_r37_c97 bl_97 br_97 wl_37 vdd gnd cell_6t
Xbit_r38_c97 bl_97 br_97 wl_38 vdd gnd cell_6t
Xbit_r39_c97 bl_97 br_97 wl_39 vdd gnd cell_6t
Xbit_r40_c97 bl_97 br_97 wl_40 vdd gnd cell_6t
Xbit_r41_c97 bl_97 br_97 wl_41 vdd gnd cell_6t
Xbit_r42_c97 bl_97 br_97 wl_42 vdd gnd cell_6t
Xbit_r43_c97 bl_97 br_97 wl_43 vdd gnd cell_6t
Xbit_r44_c97 bl_97 br_97 wl_44 vdd gnd cell_6t
Xbit_r45_c97 bl_97 br_97 wl_45 vdd gnd cell_6t
Xbit_r46_c97 bl_97 br_97 wl_46 vdd gnd cell_6t
Xbit_r47_c97 bl_97 br_97 wl_47 vdd gnd cell_6t
Xbit_r48_c97 bl_97 br_97 wl_48 vdd gnd cell_6t
Xbit_r49_c97 bl_97 br_97 wl_49 vdd gnd cell_6t
Xbit_r50_c97 bl_97 br_97 wl_50 vdd gnd cell_6t
Xbit_r51_c97 bl_97 br_97 wl_51 vdd gnd cell_6t
Xbit_r52_c97 bl_97 br_97 wl_52 vdd gnd cell_6t
Xbit_r53_c97 bl_97 br_97 wl_53 vdd gnd cell_6t
Xbit_r54_c97 bl_97 br_97 wl_54 vdd gnd cell_6t
Xbit_r55_c97 bl_97 br_97 wl_55 vdd gnd cell_6t
Xbit_r56_c97 bl_97 br_97 wl_56 vdd gnd cell_6t
Xbit_r57_c97 bl_97 br_97 wl_57 vdd gnd cell_6t
Xbit_r58_c97 bl_97 br_97 wl_58 vdd gnd cell_6t
Xbit_r59_c97 bl_97 br_97 wl_59 vdd gnd cell_6t
Xbit_r60_c97 bl_97 br_97 wl_60 vdd gnd cell_6t
Xbit_r61_c97 bl_97 br_97 wl_61 vdd gnd cell_6t
Xbit_r62_c97 bl_97 br_97 wl_62 vdd gnd cell_6t
Xbit_r63_c97 bl_97 br_97 wl_63 vdd gnd cell_6t
Xbit_r64_c97 bl_97 br_97 wl_64 vdd gnd cell_6t
Xbit_r65_c97 bl_97 br_97 wl_65 vdd gnd cell_6t
Xbit_r66_c97 bl_97 br_97 wl_66 vdd gnd cell_6t
Xbit_r67_c97 bl_97 br_97 wl_67 vdd gnd cell_6t
Xbit_r68_c97 bl_97 br_97 wl_68 vdd gnd cell_6t
Xbit_r69_c97 bl_97 br_97 wl_69 vdd gnd cell_6t
Xbit_r70_c97 bl_97 br_97 wl_70 vdd gnd cell_6t
Xbit_r71_c97 bl_97 br_97 wl_71 vdd gnd cell_6t
Xbit_r72_c97 bl_97 br_97 wl_72 vdd gnd cell_6t
Xbit_r73_c97 bl_97 br_97 wl_73 vdd gnd cell_6t
Xbit_r74_c97 bl_97 br_97 wl_74 vdd gnd cell_6t
Xbit_r75_c97 bl_97 br_97 wl_75 vdd gnd cell_6t
Xbit_r76_c97 bl_97 br_97 wl_76 vdd gnd cell_6t
Xbit_r77_c97 bl_97 br_97 wl_77 vdd gnd cell_6t
Xbit_r78_c97 bl_97 br_97 wl_78 vdd gnd cell_6t
Xbit_r79_c97 bl_97 br_97 wl_79 vdd gnd cell_6t
Xbit_r80_c97 bl_97 br_97 wl_80 vdd gnd cell_6t
Xbit_r81_c97 bl_97 br_97 wl_81 vdd gnd cell_6t
Xbit_r82_c97 bl_97 br_97 wl_82 vdd gnd cell_6t
Xbit_r83_c97 bl_97 br_97 wl_83 vdd gnd cell_6t
Xbit_r84_c97 bl_97 br_97 wl_84 vdd gnd cell_6t
Xbit_r85_c97 bl_97 br_97 wl_85 vdd gnd cell_6t
Xbit_r86_c97 bl_97 br_97 wl_86 vdd gnd cell_6t
Xbit_r87_c97 bl_97 br_97 wl_87 vdd gnd cell_6t
Xbit_r88_c97 bl_97 br_97 wl_88 vdd gnd cell_6t
Xbit_r89_c97 bl_97 br_97 wl_89 vdd gnd cell_6t
Xbit_r90_c97 bl_97 br_97 wl_90 vdd gnd cell_6t
Xbit_r91_c97 bl_97 br_97 wl_91 vdd gnd cell_6t
Xbit_r92_c97 bl_97 br_97 wl_92 vdd gnd cell_6t
Xbit_r93_c97 bl_97 br_97 wl_93 vdd gnd cell_6t
Xbit_r94_c97 bl_97 br_97 wl_94 vdd gnd cell_6t
Xbit_r95_c97 bl_97 br_97 wl_95 vdd gnd cell_6t
Xbit_r96_c97 bl_97 br_97 wl_96 vdd gnd cell_6t
Xbit_r97_c97 bl_97 br_97 wl_97 vdd gnd cell_6t
Xbit_r98_c97 bl_97 br_97 wl_98 vdd gnd cell_6t
Xbit_r99_c97 bl_97 br_97 wl_99 vdd gnd cell_6t
Xbit_r100_c97 bl_97 br_97 wl_100 vdd gnd cell_6t
Xbit_r101_c97 bl_97 br_97 wl_101 vdd gnd cell_6t
Xbit_r102_c97 bl_97 br_97 wl_102 vdd gnd cell_6t
Xbit_r103_c97 bl_97 br_97 wl_103 vdd gnd cell_6t
Xbit_r104_c97 bl_97 br_97 wl_104 vdd gnd cell_6t
Xbit_r105_c97 bl_97 br_97 wl_105 vdd gnd cell_6t
Xbit_r106_c97 bl_97 br_97 wl_106 vdd gnd cell_6t
Xbit_r107_c97 bl_97 br_97 wl_107 vdd gnd cell_6t
Xbit_r108_c97 bl_97 br_97 wl_108 vdd gnd cell_6t
Xbit_r109_c97 bl_97 br_97 wl_109 vdd gnd cell_6t
Xbit_r110_c97 bl_97 br_97 wl_110 vdd gnd cell_6t
Xbit_r111_c97 bl_97 br_97 wl_111 vdd gnd cell_6t
Xbit_r112_c97 bl_97 br_97 wl_112 vdd gnd cell_6t
Xbit_r113_c97 bl_97 br_97 wl_113 vdd gnd cell_6t
Xbit_r114_c97 bl_97 br_97 wl_114 vdd gnd cell_6t
Xbit_r115_c97 bl_97 br_97 wl_115 vdd gnd cell_6t
Xbit_r116_c97 bl_97 br_97 wl_116 vdd gnd cell_6t
Xbit_r117_c97 bl_97 br_97 wl_117 vdd gnd cell_6t
Xbit_r118_c97 bl_97 br_97 wl_118 vdd gnd cell_6t
Xbit_r119_c97 bl_97 br_97 wl_119 vdd gnd cell_6t
Xbit_r120_c97 bl_97 br_97 wl_120 vdd gnd cell_6t
Xbit_r121_c97 bl_97 br_97 wl_121 vdd gnd cell_6t
Xbit_r122_c97 bl_97 br_97 wl_122 vdd gnd cell_6t
Xbit_r123_c97 bl_97 br_97 wl_123 vdd gnd cell_6t
Xbit_r124_c97 bl_97 br_97 wl_124 vdd gnd cell_6t
Xbit_r125_c97 bl_97 br_97 wl_125 vdd gnd cell_6t
Xbit_r126_c97 bl_97 br_97 wl_126 vdd gnd cell_6t
Xbit_r127_c97 bl_97 br_97 wl_127 vdd gnd cell_6t
Xbit_r128_c97 bl_97 br_97 wl_128 vdd gnd cell_6t
Xbit_r129_c97 bl_97 br_97 wl_129 vdd gnd cell_6t
Xbit_r130_c97 bl_97 br_97 wl_130 vdd gnd cell_6t
Xbit_r131_c97 bl_97 br_97 wl_131 vdd gnd cell_6t
Xbit_r132_c97 bl_97 br_97 wl_132 vdd gnd cell_6t
Xbit_r133_c97 bl_97 br_97 wl_133 vdd gnd cell_6t
Xbit_r134_c97 bl_97 br_97 wl_134 vdd gnd cell_6t
Xbit_r135_c97 bl_97 br_97 wl_135 vdd gnd cell_6t
Xbit_r136_c97 bl_97 br_97 wl_136 vdd gnd cell_6t
Xbit_r137_c97 bl_97 br_97 wl_137 vdd gnd cell_6t
Xbit_r138_c97 bl_97 br_97 wl_138 vdd gnd cell_6t
Xbit_r139_c97 bl_97 br_97 wl_139 vdd gnd cell_6t
Xbit_r140_c97 bl_97 br_97 wl_140 vdd gnd cell_6t
Xbit_r141_c97 bl_97 br_97 wl_141 vdd gnd cell_6t
Xbit_r142_c97 bl_97 br_97 wl_142 vdd gnd cell_6t
Xbit_r143_c97 bl_97 br_97 wl_143 vdd gnd cell_6t
Xbit_r144_c97 bl_97 br_97 wl_144 vdd gnd cell_6t
Xbit_r145_c97 bl_97 br_97 wl_145 vdd gnd cell_6t
Xbit_r146_c97 bl_97 br_97 wl_146 vdd gnd cell_6t
Xbit_r147_c97 bl_97 br_97 wl_147 vdd gnd cell_6t
Xbit_r148_c97 bl_97 br_97 wl_148 vdd gnd cell_6t
Xbit_r149_c97 bl_97 br_97 wl_149 vdd gnd cell_6t
Xbit_r150_c97 bl_97 br_97 wl_150 vdd gnd cell_6t
Xbit_r151_c97 bl_97 br_97 wl_151 vdd gnd cell_6t
Xbit_r152_c97 bl_97 br_97 wl_152 vdd gnd cell_6t
Xbit_r153_c97 bl_97 br_97 wl_153 vdd gnd cell_6t
Xbit_r154_c97 bl_97 br_97 wl_154 vdd gnd cell_6t
Xbit_r155_c97 bl_97 br_97 wl_155 vdd gnd cell_6t
Xbit_r156_c97 bl_97 br_97 wl_156 vdd gnd cell_6t
Xbit_r157_c97 bl_97 br_97 wl_157 vdd gnd cell_6t
Xbit_r158_c97 bl_97 br_97 wl_158 vdd gnd cell_6t
Xbit_r159_c97 bl_97 br_97 wl_159 vdd gnd cell_6t
Xbit_r160_c97 bl_97 br_97 wl_160 vdd gnd cell_6t
Xbit_r161_c97 bl_97 br_97 wl_161 vdd gnd cell_6t
Xbit_r162_c97 bl_97 br_97 wl_162 vdd gnd cell_6t
Xbit_r163_c97 bl_97 br_97 wl_163 vdd gnd cell_6t
Xbit_r164_c97 bl_97 br_97 wl_164 vdd gnd cell_6t
Xbit_r165_c97 bl_97 br_97 wl_165 vdd gnd cell_6t
Xbit_r166_c97 bl_97 br_97 wl_166 vdd gnd cell_6t
Xbit_r167_c97 bl_97 br_97 wl_167 vdd gnd cell_6t
Xbit_r168_c97 bl_97 br_97 wl_168 vdd gnd cell_6t
Xbit_r169_c97 bl_97 br_97 wl_169 vdd gnd cell_6t
Xbit_r170_c97 bl_97 br_97 wl_170 vdd gnd cell_6t
Xbit_r171_c97 bl_97 br_97 wl_171 vdd gnd cell_6t
Xbit_r172_c97 bl_97 br_97 wl_172 vdd gnd cell_6t
Xbit_r173_c97 bl_97 br_97 wl_173 vdd gnd cell_6t
Xbit_r174_c97 bl_97 br_97 wl_174 vdd gnd cell_6t
Xbit_r175_c97 bl_97 br_97 wl_175 vdd gnd cell_6t
Xbit_r176_c97 bl_97 br_97 wl_176 vdd gnd cell_6t
Xbit_r177_c97 bl_97 br_97 wl_177 vdd gnd cell_6t
Xbit_r178_c97 bl_97 br_97 wl_178 vdd gnd cell_6t
Xbit_r179_c97 bl_97 br_97 wl_179 vdd gnd cell_6t
Xbit_r180_c97 bl_97 br_97 wl_180 vdd gnd cell_6t
Xbit_r181_c97 bl_97 br_97 wl_181 vdd gnd cell_6t
Xbit_r182_c97 bl_97 br_97 wl_182 vdd gnd cell_6t
Xbit_r183_c97 bl_97 br_97 wl_183 vdd gnd cell_6t
Xbit_r184_c97 bl_97 br_97 wl_184 vdd gnd cell_6t
Xbit_r185_c97 bl_97 br_97 wl_185 vdd gnd cell_6t
Xbit_r186_c97 bl_97 br_97 wl_186 vdd gnd cell_6t
Xbit_r187_c97 bl_97 br_97 wl_187 vdd gnd cell_6t
Xbit_r188_c97 bl_97 br_97 wl_188 vdd gnd cell_6t
Xbit_r189_c97 bl_97 br_97 wl_189 vdd gnd cell_6t
Xbit_r190_c97 bl_97 br_97 wl_190 vdd gnd cell_6t
Xbit_r191_c97 bl_97 br_97 wl_191 vdd gnd cell_6t
Xbit_r192_c97 bl_97 br_97 wl_192 vdd gnd cell_6t
Xbit_r193_c97 bl_97 br_97 wl_193 vdd gnd cell_6t
Xbit_r194_c97 bl_97 br_97 wl_194 vdd gnd cell_6t
Xbit_r195_c97 bl_97 br_97 wl_195 vdd gnd cell_6t
Xbit_r196_c97 bl_97 br_97 wl_196 vdd gnd cell_6t
Xbit_r197_c97 bl_97 br_97 wl_197 vdd gnd cell_6t
Xbit_r198_c97 bl_97 br_97 wl_198 vdd gnd cell_6t
Xbit_r199_c97 bl_97 br_97 wl_199 vdd gnd cell_6t
Xbit_r200_c97 bl_97 br_97 wl_200 vdd gnd cell_6t
Xbit_r201_c97 bl_97 br_97 wl_201 vdd gnd cell_6t
Xbit_r202_c97 bl_97 br_97 wl_202 vdd gnd cell_6t
Xbit_r203_c97 bl_97 br_97 wl_203 vdd gnd cell_6t
Xbit_r204_c97 bl_97 br_97 wl_204 vdd gnd cell_6t
Xbit_r205_c97 bl_97 br_97 wl_205 vdd gnd cell_6t
Xbit_r206_c97 bl_97 br_97 wl_206 vdd gnd cell_6t
Xbit_r207_c97 bl_97 br_97 wl_207 vdd gnd cell_6t
Xbit_r208_c97 bl_97 br_97 wl_208 vdd gnd cell_6t
Xbit_r209_c97 bl_97 br_97 wl_209 vdd gnd cell_6t
Xbit_r210_c97 bl_97 br_97 wl_210 vdd gnd cell_6t
Xbit_r211_c97 bl_97 br_97 wl_211 vdd gnd cell_6t
Xbit_r212_c97 bl_97 br_97 wl_212 vdd gnd cell_6t
Xbit_r213_c97 bl_97 br_97 wl_213 vdd gnd cell_6t
Xbit_r214_c97 bl_97 br_97 wl_214 vdd gnd cell_6t
Xbit_r215_c97 bl_97 br_97 wl_215 vdd gnd cell_6t
Xbit_r216_c97 bl_97 br_97 wl_216 vdd gnd cell_6t
Xbit_r217_c97 bl_97 br_97 wl_217 vdd gnd cell_6t
Xbit_r218_c97 bl_97 br_97 wl_218 vdd gnd cell_6t
Xbit_r219_c97 bl_97 br_97 wl_219 vdd gnd cell_6t
Xbit_r220_c97 bl_97 br_97 wl_220 vdd gnd cell_6t
Xbit_r221_c97 bl_97 br_97 wl_221 vdd gnd cell_6t
Xbit_r222_c97 bl_97 br_97 wl_222 vdd gnd cell_6t
Xbit_r223_c97 bl_97 br_97 wl_223 vdd gnd cell_6t
Xbit_r224_c97 bl_97 br_97 wl_224 vdd gnd cell_6t
Xbit_r225_c97 bl_97 br_97 wl_225 vdd gnd cell_6t
Xbit_r226_c97 bl_97 br_97 wl_226 vdd gnd cell_6t
Xbit_r227_c97 bl_97 br_97 wl_227 vdd gnd cell_6t
Xbit_r228_c97 bl_97 br_97 wl_228 vdd gnd cell_6t
Xbit_r229_c97 bl_97 br_97 wl_229 vdd gnd cell_6t
Xbit_r230_c97 bl_97 br_97 wl_230 vdd gnd cell_6t
Xbit_r231_c97 bl_97 br_97 wl_231 vdd gnd cell_6t
Xbit_r232_c97 bl_97 br_97 wl_232 vdd gnd cell_6t
Xbit_r233_c97 bl_97 br_97 wl_233 vdd gnd cell_6t
Xbit_r234_c97 bl_97 br_97 wl_234 vdd gnd cell_6t
Xbit_r235_c97 bl_97 br_97 wl_235 vdd gnd cell_6t
Xbit_r236_c97 bl_97 br_97 wl_236 vdd gnd cell_6t
Xbit_r237_c97 bl_97 br_97 wl_237 vdd gnd cell_6t
Xbit_r238_c97 bl_97 br_97 wl_238 vdd gnd cell_6t
Xbit_r239_c97 bl_97 br_97 wl_239 vdd gnd cell_6t
Xbit_r240_c97 bl_97 br_97 wl_240 vdd gnd cell_6t
Xbit_r241_c97 bl_97 br_97 wl_241 vdd gnd cell_6t
Xbit_r242_c97 bl_97 br_97 wl_242 vdd gnd cell_6t
Xbit_r243_c97 bl_97 br_97 wl_243 vdd gnd cell_6t
Xbit_r244_c97 bl_97 br_97 wl_244 vdd gnd cell_6t
Xbit_r245_c97 bl_97 br_97 wl_245 vdd gnd cell_6t
Xbit_r246_c97 bl_97 br_97 wl_246 vdd gnd cell_6t
Xbit_r247_c97 bl_97 br_97 wl_247 vdd gnd cell_6t
Xbit_r248_c97 bl_97 br_97 wl_248 vdd gnd cell_6t
Xbit_r249_c97 bl_97 br_97 wl_249 vdd gnd cell_6t
Xbit_r250_c97 bl_97 br_97 wl_250 vdd gnd cell_6t
Xbit_r251_c97 bl_97 br_97 wl_251 vdd gnd cell_6t
Xbit_r252_c97 bl_97 br_97 wl_252 vdd gnd cell_6t
Xbit_r253_c97 bl_97 br_97 wl_253 vdd gnd cell_6t
Xbit_r254_c97 bl_97 br_97 wl_254 vdd gnd cell_6t
Xbit_r255_c97 bl_97 br_97 wl_255 vdd gnd cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd cell_6t
Xbit_r1_c98 bl_98 br_98 wl_1 vdd gnd cell_6t
Xbit_r2_c98 bl_98 br_98 wl_2 vdd gnd cell_6t
Xbit_r3_c98 bl_98 br_98 wl_3 vdd gnd cell_6t
Xbit_r4_c98 bl_98 br_98 wl_4 vdd gnd cell_6t
Xbit_r5_c98 bl_98 br_98 wl_5 vdd gnd cell_6t
Xbit_r6_c98 bl_98 br_98 wl_6 vdd gnd cell_6t
Xbit_r7_c98 bl_98 br_98 wl_7 vdd gnd cell_6t
Xbit_r8_c98 bl_98 br_98 wl_8 vdd gnd cell_6t
Xbit_r9_c98 bl_98 br_98 wl_9 vdd gnd cell_6t
Xbit_r10_c98 bl_98 br_98 wl_10 vdd gnd cell_6t
Xbit_r11_c98 bl_98 br_98 wl_11 vdd gnd cell_6t
Xbit_r12_c98 bl_98 br_98 wl_12 vdd gnd cell_6t
Xbit_r13_c98 bl_98 br_98 wl_13 vdd gnd cell_6t
Xbit_r14_c98 bl_98 br_98 wl_14 vdd gnd cell_6t
Xbit_r15_c98 bl_98 br_98 wl_15 vdd gnd cell_6t
Xbit_r16_c98 bl_98 br_98 wl_16 vdd gnd cell_6t
Xbit_r17_c98 bl_98 br_98 wl_17 vdd gnd cell_6t
Xbit_r18_c98 bl_98 br_98 wl_18 vdd gnd cell_6t
Xbit_r19_c98 bl_98 br_98 wl_19 vdd gnd cell_6t
Xbit_r20_c98 bl_98 br_98 wl_20 vdd gnd cell_6t
Xbit_r21_c98 bl_98 br_98 wl_21 vdd gnd cell_6t
Xbit_r22_c98 bl_98 br_98 wl_22 vdd gnd cell_6t
Xbit_r23_c98 bl_98 br_98 wl_23 vdd gnd cell_6t
Xbit_r24_c98 bl_98 br_98 wl_24 vdd gnd cell_6t
Xbit_r25_c98 bl_98 br_98 wl_25 vdd gnd cell_6t
Xbit_r26_c98 bl_98 br_98 wl_26 vdd gnd cell_6t
Xbit_r27_c98 bl_98 br_98 wl_27 vdd gnd cell_6t
Xbit_r28_c98 bl_98 br_98 wl_28 vdd gnd cell_6t
Xbit_r29_c98 bl_98 br_98 wl_29 vdd gnd cell_6t
Xbit_r30_c98 bl_98 br_98 wl_30 vdd gnd cell_6t
Xbit_r31_c98 bl_98 br_98 wl_31 vdd gnd cell_6t
Xbit_r32_c98 bl_98 br_98 wl_32 vdd gnd cell_6t
Xbit_r33_c98 bl_98 br_98 wl_33 vdd gnd cell_6t
Xbit_r34_c98 bl_98 br_98 wl_34 vdd gnd cell_6t
Xbit_r35_c98 bl_98 br_98 wl_35 vdd gnd cell_6t
Xbit_r36_c98 bl_98 br_98 wl_36 vdd gnd cell_6t
Xbit_r37_c98 bl_98 br_98 wl_37 vdd gnd cell_6t
Xbit_r38_c98 bl_98 br_98 wl_38 vdd gnd cell_6t
Xbit_r39_c98 bl_98 br_98 wl_39 vdd gnd cell_6t
Xbit_r40_c98 bl_98 br_98 wl_40 vdd gnd cell_6t
Xbit_r41_c98 bl_98 br_98 wl_41 vdd gnd cell_6t
Xbit_r42_c98 bl_98 br_98 wl_42 vdd gnd cell_6t
Xbit_r43_c98 bl_98 br_98 wl_43 vdd gnd cell_6t
Xbit_r44_c98 bl_98 br_98 wl_44 vdd gnd cell_6t
Xbit_r45_c98 bl_98 br_98 wl_45 vdd gnd cell_6t
Xbit_r46_c98 bl_98 br_98 wl_46 vdd gnd cell_6t
Xbit_r47_c98 bl_98 br_98 wl_47 vdd gnd cell_6t
Xbit_r48_c98 bl_98 br_98 wl_48 vdd gnd cell_6t
Xbit_r49_c98 bl_98 br_98 wl_49 vdd gnd cell_6t
Xbit_r50_c98 bl_98 br_98 wl_50 vdd gnd cell_6t
Xbit_r51_c98 bl_98 br_98 wl_51 vdd gnd cell_6t
Xbit_r52_c98 bl_98 br_98 wl_52 vdd gnd cell_6t
Xbit_r53_c98 bl_98 br_98 wl_53 vdd gnd cell_6t
Xbit_r54_c98 bl_98 br_98 wl_54 vdd gnd cell_6t
Xbit_r55_c98 bl_98 br_98 wl_55 vdd gnd cell_6t
Xbit_r56_c98 bl_98 br_98 wl_56 vdd gnd cell_6t
Xbit_r57_c98 bl_98 br_98 wl_57 vdd gnd cell_6t
Xbit_r58_c98 bl_98 br_98 wl_58 vdd gnd cell_6t
Xbit_r59_c98 bl_98 br_98 wl_59 vdd gnd cell_6t
Xbit_r60_c98 bl_98 br_98 wl_60 vdd gnd cell_6t
Xbit_r61_c98 bl_98 br_98 wl_61 vdd gnd cell_6t
Xbit_r62_c98 bl_98 br_98 wl_62 vdd gnd cell_6t
Xbit_r63_c98 bl_98 br_98 wl_63 vdd gnd cell_6t
Xbit_r64_c98 bl_98 br_98 wl_64 vdd gnd cell_6t
Xbit_r65_c98 bl_98 br_98 wl_65 vdd gnd cell_6t
Xbit_r66_c98 bl_98 br_98 wl_66 vdd gnd cell_6t
Xbit_r67_c98 bl_98 br_98 wl_67 vdd gnd cell_6t
Xbit_r68_c98 bl_98 br_98 wl_68 vdd gnd cell_6t
Xbit_r69_c98 bl_98 br_98 wl_69 vdd gnd cell_6t
Xbit_r70_c98 bl_98 br_98 wl_70 vdd gnd cell_6t
Xbit_r71_c98 bl_98 br_98 wl_71 vdd gnd cell_6t
Xbit_r72_c98 bl_98 br_98 wl_72 vdd gnd cell_6t
Xbit_r73_c98 bl_98 br_98 wl_73 vdd gnd cell_6t
Xbit_r74_c98 bl_98 br_98 wl_74 vdd gnd cell_6t
Xbit_r75_c98 bl_98 br_98 wl_75 vdd gnd cell_6t
Xbit_r76_c98 bl_98 br_98 wl_76 vdd gnd cell_6t
Xbit_r77_c98 bl_98 br_98 wl_77 vdd gnd cell_6t
Xbit_r78_c98 bl_98 br_98 wl_78 vdd gnd cell_6t
Xbit_r79_c98 bl_98 br_98 wl_79 vdd gnd cell_6t
Xbit_r80_c98 bl_98 br_98 wl_80 vdd gnd cell_6t
Xbit_r81_c98 bl_98 br_98 wl_81 vdd gnd cell_6t
Xbit_r82_c98 bl_98 br_98 wl_82 vdd gnd cell_6t
Xbit_r83_c98 bl_98 br_98 wl_83 vdd gnd cell_6t
Xbit_r84_c98 bl_98 br_98 wl_84 vdd gnd cell_6t
Xbit_r85_c98 bl_98 br_98 wl_85 vdd gnd cell_6t
Xbit_r86_c98 bl_98 br_98 wl_86 vdd gnd cell_6t
Xbit_r87_c98 bl_98 br_98 wl_87 vdd gnd cell_6t
Xbit_r88_c98 bl_98 br_98 wl_88 vdd gnd cell_6t
Xbit_r89_c98 bl_98 br_98 wl_89 vdd gnd cell_6t
Xbit_r90_c98 bl_98 br_98 wl_90 vdd gnd cell_6t
Xbit_r91_c98 bl_98 br_98 wl_91 vdd gnd cell_6t
Xbit_r92_c98 bl_98 br_98 wl_92 vdd gnd cell_6t
Xbit_r93_c98 bl_98 br_98 wl_93 vdd gnd cell_6t
Xbit_r94_c98 bl_98 br_98 wl_94 vdd gnd cell_6t
Xbit_r95_c98 bl_98 br_98 wl_95 vdd gnd cell_6t
Xbit_r96_c98 bl_98 br_98 wl_96 vdd gnd cell_6t
Xbit_r97_c98 bl_98 br_98 wl_97 vdd gnd cell_6t
Xbit_r98_c98 bl_98 br_98 wl_98 vdd gnd cell_6t
Xbit_r99_c98 bl_98 br_98 wl_99 vdd gnd cell_6t
Xbit_r100_c98 bl_98 br_98 wl_100 vdd gnd cell_6t
Xbit_r101_c98 bl_98 br_98 wl_101 vdd gnd cell_6t
Xbit_r102_c98 bl_98 br_98 wl_102 vdd gnd cell_6t
Xbit_r103_c98 bl_98 br_98 wl_103 vdd gnd cell_6t
Xbit_r104_c98 bl_98 br_98 wl_104 vdd gnd cell_6t
Xbit_r105_c98 bl_98 br_98 wl_105 vdd gnd cell_6t
Xbit_r106_c98 bl_98 br_98 wl_106 vdd gnd cell_6t
Xbit_r107_c98 bl_98 br_98 wl_107 vdd gnd cell_6t
Xbit_r108_c98 bl_98 br_98 wl_108 vdd gnd cell_6t
Xbit_r109_c98 bl_98 br_98 wl_109 vdd gnd cell_6t
Xbit_r110_c98 bl_98 br_98 wl_110 vdd gnd cell_6t
Xbit_r111_c98 bl_98 br_98 wl_111 vdd gnd cell_6t
Xbit_r112_c98 bl_98 br_98 wl_112 vdd gnd cell_6t
Xbit_r113_c98 bl_98 br_98 wl_113 vdd gnd cell_6t
Xbit_r114_c98 bl_98 br_98 wl_114 vdd gnd cell_6t
Xbit_r115_c98 bl_98 br_98 wl_115 vdd gnd cell_6t
Xbit_r116_c98 bl_98 br_98 wl_116 vdd gnd cell_6t
Xbit_r117_c98 bl_98 br_98 wl_117 vdd gnd cell_6t
Xbit_r118_c98 bl_98 br_98 wl_118 vdd gnd cell_6t
Xbit_r119_c98 bl_98 br_98 wl_119 vdd gnd cell_6t
Xbit_r120_c98 bl_98 br_98 wl_120 vdd gnd cell_6t
Xbit_r121_c98 bl_98 br_98 wl_121 vdd gnd cell_6t
Xbit_r122_c98 bl_98 br_98 wl_122 vdd gnd cell_6t
Xbit_r123_c98 bl_98 br_98 wl_123 vdd gnd cell_6t
Xbit_r124_c98 bl_98 br_98 wl_124 vdd gnd cell_6t
Xbit_r125_c98 bl_98 br_98 wl_125 vdd gnd cell_6t
Xbit_r126_c98 bl_98 br_98 wl_126 vdd gnd cell_6t
Xbit_r127_c98 bl_98 br_98 wl_127 vdd gnd cell_6t
Xbit_r128_c98 bl_98 br_98 wl_128 vdd gnd cell_6t
Xbit_r129_c98 bl_98 br_98 wl_129 vdd gnd cell_6t
Xbit_r130_c98 bl_98 br_98 wl_130 vdd gnd cell_6t
Xbit_r131_c98 bl_98 br_98 wl_131 vdd gnd cell_6t
Xbit_r132_c98 bl_98 br_98 wl_132 vdd gnd cell_6t
Xbit_r133_c98 bl_98 br_98 wl_133 vdd gnd cell_6t
Xbit_r134_c98 bl_98 br_98 wl_134 vdd gnd cell_6t
Xbit_r135_c98 bl_98 br_98 wl_135 vdd gnd cell_6t
Xbit_r136_c98 bl_98 br_98 wl_136 vdd gnd cell_6t
Xbit_r137_c98 bl_98 br_98 wl_137 vdd gnd cell_6t
Xbit_r138_c98 bl_98 br_98 wl_138 vdd gnd cell_6t
Xbit_r139_c98 bl_98 br_98 wl_139 vdd gnd cell_6t
Xbit_r140_c98 bl_98 br_98 wl_140 vdd gnd cell_6t
Xbit_r141_c98 bl_98 br_98 wl_141 vdd gnd cell_6t
Xbit_r142_c98 bl_98 br_98 wl_142 vdd gnd cell_6t
Xbit_r143_c98 bl_98 br_98 wl_143 vdd gnd cell_6t
Xbit_r144_c98 bl_98 br_98 wl_144 vdd gnd cell_6t
Xbit_r145_c98 bl_98 br_98 wl_145 vdd gnd cell_6t
Xbit_r146_c98 bl_98 br_98 wl_146 vdd gnd cell_6t
Xbit_r147_c98 bl_98 br_98 wl_147 vdd gnd cell_6t
Xbit_r148_c98 bl_98 br_98 wl_148 vdd gnd cell_6t
Xbit_r149_c98 bl_98 br_98 wl_149 vdd gnd cell_6t
Xbit_r150_c98 bl_98 br_98 wl_150 vdd gnd cell_6t
Xbit_r151_c98 bl_98 br_98 wl_151 vdd gnd cell_6t
Xbit_r152_c98 bl_98 br_98 wl_152 vdd gnd cell_6t
Xbit_r153_c98 bl_98 br_98 wl_153 vdd gnd cell_6t
Xbit_r154_c98 bl_98 br_98 wl_154 vdd gnd cell_6t
Xbit_r155_c98 bl_98 br_98 wl_155 vdd gnd cell_6t
Xbit_r156_c98 bl_98 br_98 wl_156 vdd gnd cell_6t
Xbit_r157_c98 bl_98 br_98 wl_157 vdd gnd cell_6t
Xbit_r158_c98 bl_98 br_98 wl_158 vdd gnd cell_6t
Xbit_r159_c98 bl_98 br_98 wl_159 vdd gnd cell_6t
Xbit_r160_c98 bl_98 br_98 wl_160 vdd gnd cell_6t
Xbit_r161_c98 bl_98 br_98 wl_161 vdd gnd cell_6t
Xbit_r162_c98 bl_98 br_98 wl_162 vdd gnd cell_6t
Xbit_r163_c98 bl_98 br_98 wl_163 vdd gnd cell_6t
Xbit_r164_c98 bl_98 br_98 wl_164 vdd gnd cell_6t
Xbit_r165_c98 bl_98 br_98 wl_165 vdd gnd cell_6t
Xbit_r166_c98 bl_98 br_98 wl_166 vdd gnd cell_6t
Xbit_r167_c98 bl_98 br_98 wl_167 vdd gnd cell_6t
Xbit_r168_c98 bl_98 br_98 wl_168 vdd gnd cell_6t
Xbit_r169_c98 bl_98 br_98 wl_169 vdd gnd cell_6t
Xbit_r170_c98 bl_98 br_98 wl_170 vdd gnd cell_6t
Xbit_r171_c98 bl_98 br_98 wl_171 vdd gnd cell_6t
Xbit_r172_c98 bl_98 br_98 wl_172 vdd gnd cell_6t
Xbit_r173_c98 bl_98 br_98 wl_173 vdd gnd cell_6t
Xbit_r174_c98 bl_98 br_98 wl_174 vdd gnd cell_6t
Xbit_r175_c98 bl_98 br_98 wl_175 vdd gnd cell_6t
Xbit_r176_c98 bl_98 br_98 wl_176 vdd gnd cell_6t
Xbit_r177_c98 bl_98 br_98 wl_177 vdd gnd cell_6t
Xbit_r178_c98 bl_98 br_98 wl_178 vdd gnd cell_6t
Xbit_r179_c98 bl_98 br_98 wl_179 vdd gnd cell_6t
Xbit_r180_c98 bl_98 br_98 wl_180 vdd gnd cell_6t
Xbit_r181_c98 bl_98 br_98 wl_181 vdd gnd cell_6t
Xbit_r182_c98 bl_98 br_98 wl_182 vdd gnd cell_6t
Xbit_r183_c98 bl_98 br_98 wl_183 vdd gnd cell_6t
Xbit_r184_c98 bl_98 br_98 wl_184 vdd gnd cell_6t
Xbit_r185_c98 bl_98 br_98 wl_185 vdd gnd cell_6t
Xbit_r186_c98 bl_98 br_98 wl_186 vdd gnd cell_6t
Xbit_r187_c98 bl_98 br_98 wl_187 vdd gnd cell_6t
Xbit_r188_c98 bl_98 br_98 wl_188 vdd gnd cell_6t
Xbit_r189_c98 bl_98 br_98 wl_189 vdd gnd cell_6t
Xbit_r190_c98 bl_98 br_98 wl_190 vdd gnd cell_6t
Xbit_r191_c98 bl_98 br_98 wl_191 vdd gnd cell_6t
Xbit_r192_c98 bl_98 br_98 wl_192 vdd gnd cell_6t
Xbit_r193_c98 bl_98 br_98 wl_193 vdd gnd cell_6t
Xbit_r194_c98 bl_98 br_98 wl_194 vdd gnd cell_6t
Xbit_r195_c98 bl_98 br_98 wl_195 vdd gnd cell_6t
Xbit_r196_c98 bl_98 br_98 wl_196 vdd gnd cell_6t
Xbit_r197_c98 bl_98 br_98 wl_197 vdd gnd cell_6t
Xbit_r198_c98 bl_98 br_98 wl_198 vdd gnd cell_6t
Xbit_r199_c98 bl_98 br_98 wl_199 vdd gnd cell_6t
Xbit_r200_c98 bl_98 br_98 wl_200 vdd gnd cell_6t
Xbit_r201_c98 bl_98 br_98 wl_201 vdd gnd cell_6t
Xbit_r202_c98 bl_98 br_98 wl_202 vdd gnd cell_6t
Xbit_r203_c98 bl_98 br_98 wl_203 vdd gnd cell_6t
Xbit_r204_c98 bl_98 br_98 wl_204 vdd gnd cell_6t
Xbit_r205_c98 bl_98 br_98 wl_205 vdd gnd cell_6t
Xbit_r206_c98 bl_98 br_98 wl_206 vdd gnd cell_6t
Xbit_r207_c98 bl_98 br_98 wl_207 vdd gnd cell_6t
Xbit_r208_c98 bl_98 br_98 wl_208 vdd gnd cell_6t
Xbit_r209_c98 bl_98 br_98 wl_209 vdd gnd cell_6t
Xbit_r210_c98 bl_98 br_98 wl_210 vdd gnd cell_6t
Xbit_r211_c98 bl_98 br_98 wl_211 vdd gnd cell_6t
Xbit_r212_c98 bl_98 br_98 wl_212 vdd gnd cell_6t
Xbit_r213_c98 bl_98 br_98 wl_213 vdd gnd cell_6t
Xbit_r214_c98 bl_98 br_98 wl_214 vdd gnd cell_6t
Xbit_r215_c98 bl_98 br_98 wl_215 vdd gnd cell_6t
Xbit_r216_c98 bl_98 br_98 wl_216 vdd gnd cell_6t
Xbit_r217_c98 bl_98 br_98 wl_217 vdd gnd cell_6t
Xbit_r218_c98 bl_98 br_98 wl_218 vdd gnd cell_6t
Xbit_r219_c98 bl_98 br_98 wl_219 vdd gnd cell_6t
Xbit_r220_c98 bl_98 br_98 wl_220 vdd gnd cell_6t
Xbit_r221_c98 bl_98 br_98 wl_221 vdd gnd cell_6t
Xbit_r222_c98 bl_98 br_98 wl_222 vdd gnd cell_6t
Xbit_r223_c98 bl_98 br_98 wl_223 vdd gnd cell_6t
Xbit_r224_c98 bl_98 br_98 wl_224 vdd gnd cell_6t
Xbit_r225_c98 bl_98 br_98 wl_225 vdd gnd cell_6t
Xbit_r226_c98 bl_98 br_98 wl_226 vdd gnd cell_6t
Xbit_r227_c98 bl_98 br_98 wl_227 vdd gnd cell_6t
Xbit_r228_c98 bl_98 br_98 wl_228 vdd gnd cell_6t
Xbit_r229_c98 bl_98 br_98 wl_229 vdd gnd cell_6t
Xbit_r230_c98 bl_98 br_98 wl_230 vdd gnd cell_6t
Xbit_r231_c98 bl_98 br_98 wl_231 vdd gnd cell_6t
Xbit_r232_c98 bl_98 br_98 wl_232 vdd gnd cell_6t
Xbit_r233_c98 bl_98 br_98 wl_233 vdd gnd cell_6t
Xbit_r234_c98 bl_98 br_98 wl_234 vdd gnd cell_6t
Xbit_r235_c98 bl_98 br_98 wl_235 vdd gnd cell_6t
Xbit_r236_c98 bl_98 br_98 wl_236 vdd gnd cell_6t
Xbit_r237_c98 bl_98 br_98 wl_237 vdd gnd cell_6t
Xbit_r238_c98 bl_98 br_98 wl_238 vdd gnd cell_6t
Xbit_r239_c98 bl_98 br_98 wl_239 vdd gnd cell_6t
Xbit_r240_c98 bl_98 br_98 wl_240 vdd gnd cell_6t
Xbit_r241_c98 bl_98 br_98 wl_241 vdd gnd cell_6t
Xbit_r242_c98 bl_98 br_98 wl_242 vdd gnd cell_6t
Xbit_r243_c98 bl_98 br_98 wl_243 vdd gnd cell_6t
Xbit_r244_c98 bl_98 br_98 wl_244 vdd gnd cell_6t
Xbit_r245_c98 bl_98 br_98 wl_245 vdd gnd cell_6t
Xbit_r246_c98 bl_98 br_98 wl_246 vdd gnd cell_6t
Xbit_r247_c98 bl_98 br_98 wl_247 vdd gnd cell_6t
Xbit_r248_c98 bl_98 br_98 wl_248 vdd gnd cell_6t
Xbit_r249_c98 bl_98 br_98 wl_249 vdd gnd cell_6t
Xbit_r250_c98 bl_98 br_98 wl_250 vdd gnd cell_6t
Xbit_r251_c98 bl_98 br_98 wl_251 vdd gnd cell_6t
Xbit_r252_c98 bl_98 br_98 wl_252 vdd gnd cell_6t
Xbit_r253_c98 bl_98 br_98 wl_253 vdd gnd cell_6t
Xbit_r254_c98 bl_98 br_98 wl_254 vdd gnd cell_6t
Xbit_r255_c98 bl_98 br_98 wl_255 vdd gnd cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd cell_6t
Xbit_r1_c99 bl_99 br_99 wl_1 vdd gnd cell_6t
Xbit_r2_c99 bl_99 br_99 wl_2 vdd gnd cell_6t
Xbit_r3_c99 bl_99 br_99 wl_3 vdd gnd cell_6t
Xbit_r4_c99 bl_99 br_99 wl_4 vdd gnd cell_6t
Xbit_r5_c99 bl_99 br_99 wl_5 vdd gnd cell_6t
Xbit_r6_c99 bl_99 br_99 wl_6 vdd gnd cell_6t
Xbit_r7_c99 bl_99 br_99 wl_7 vdd gnd cell_6t
Xbit_r8_c99 bl_99 br_99 wl_8 vdd gnd cell_6t
Xbit_r9_c99 bl_99 br_99 wl_9 vdd gnd cell_6t
Xbit_r10_c99 bl_99 br_99 wl_10 vdd gnd cell_6t
Xbit_r11_c99 bl_99 br_99 wl_11 vdd gnd cell_6t
Xbit_r12_c99 bl_99 br_99 wl_12 vdd gnd cell_6t
Xbit_r13_c99 bl_99 br_99 wl_13 vdd gnd cell_6t
Xbit_r14_c99 bl_99 br_99 wl_14 vdd gnd cell_6t
Xbit_r15_c99 bl_99 br_99 wl_15 vdd gnd cell_6t
Xbit_r16_c99 bl_99 br_99 wl_16 vdd gnd cell_6t
Xbit_r17_c99 bl_99 br_99 wl_17 vdd gnd cell_6t
Xbit_r18_c99 bl_99 br_99 wl_18 vdd gnd cell_6t
Xbit_r19_c99 bl_99 br_99 wl_19 vdd gnd cell_6t
Xbit_r20_c99 bl_99 br_99 wl_20 vdd gnd cell_6t
Xbit_r21_c99 bl_99 br_99 wl_21 vdd gnd cell_6t
Xbit_r22_c99 bl_99 br_99 wl_22 vdd gnd cell_6t
Xbit_r23_c99 bl_99 br_99 wl_23 vdd gnd cell_6t
Xbit_r24_c99 bl_99 br_99 wl_24 vdd gnd cell_6t
Xbit_r25_c99 bl_99 br_99 wl_25 vdd gnd cell_6t
Xbit_r26_c99 bl_99 br_99 wl_26 vdd gnd cell_6t
Xbit_r27_c99 bl_99 br_99 wl_27 vdd gnd cell_6t
Xbit_r28_c99 bl_99 br_99 wl_28 vdd gnd cell_6t
Xbit_r29_c99 bl_99 br_99 wl_29 vdd gnd cell_6t
Xbit_r30_c99 bl_99 br_99 wl_30 vdd gnd cell_6t
Xbit_r31_c99 bl_99 br_99 wl_31 vdd gnd cell_6t
Xbit_r32_c99 bl_99 br_99 wl_32 vdd gnd cell_6t
Xbit_r33_c99 bl_99 br_99 wl_33 vdd gnd cell_6t
Xbit_r34_c99 bl_99 br_99 wl_34 vdd gnd cell_6t
Xbit_r35_c99 bl_99 br_99 wl_35 vdd gnd cell_6t
Xbit_r36_c99 bl_99 br_99 wl_36 vdd gnd cell_6t
Xbit_r37_c99 bl_99 br_99 wl_37 vdd gnd cell_6t
Xbit_r38_c99 bl_99 br_99 wl_38 vdd gnd cell_6t
Xbit_r39_c99 bl_99 br_99 wl_39 vdd gnd cell_6t
Xbit_r40_c99 bl_99 br_99 wl_40 vdd gnd cell_6t
Xbit_r41_c99 bl_99 br_99 wl_41 vdd gnd cell_6t
Xbit_r42_c99 bl_99 br_99 wl_42 vdd gnd cell_6t
Xbit_r43_c99 bl_99 br_99 wl_43 vdd gnd cell_6t
Xbit_r44_c99 bl_99 br_99 wl_44 vdd gnd cell_6t
Xbit_r45_c99 bl_99 br_99 wl_45 vdd gnd cell_6t
Xbit_r46_c99 bl_99 br_99 wl_46 vdd gnd cell_6t
Xbit_r47_c99 bl_99 br_99 wl_47 vdd gnd cell_6t
Xbit_r48_c99 bl_99 br_99 wl_48 vdd gnd cell_6t
Xbit_r49_c99 bl_99 br_99 wl_49 vdd gnd cell_6t
Xbit_r50_c99 bl_99 br_99 wl_50 vdd gnd cell_6t
Xbit_r51_c99 bl_99 br_99 wl_51 vdd gnd cell_6t
Xbit_r52_c99 bl_99 br_99 wl_52 vdd gnd cell_6t
Xbit_r53_c99 bl_99 br_99 wl_53 vdd gnd cell_6t
Xbit_r54_c99 bl_99 br_99 wl_54 vdd gnd cell_6t
Xbit_r55_c99 bl_99 br_99 wl_55 vdd gnd cell_6t
Xbit_r56_c99 bl_99 br_99 wl_56 vdd gnd cell_6t
Xbit_r57_c99 bl_99 br_99 wl_57 vdd gnd cell_6t
Xbit_r58_c99 bl_99 br_99 wl_58 vdd gnd cell_6t
Xbit_r59_c99 bl_99 br_99 wl_59 vdd gnd cell_6t
Xbit_r60_c99 bl_99 br_99 wl_60 vdd gnd cell_6t
Xbit_r61_c99 bl_99 br_99 wl_61 vdd gnd cell_6t
Xbit_r62_c99 bl_99 br_99 wl_62 vdd gnd cell_6t
Xbit_r63_c99 bl_99 br_99 wl_63 vdd gnd cell_6t
Xbit_r64_c99 bl_99 br_99 wl_64 vdd gnd cell_6t
Xbit_r65_c99 bl_99 br_99 wl_65 vdd gnd cell_6t
Xbit_r66_c99 bl_99 br_99 wl_66 vdd gnd cell_6t
Xbit_r67_c99 bl_99 br_99 wl_67 vdd gnd cell_6t
Xbit_r68_c99 bl_99 br_99 wl_68 vdd gnd cell_6t
Xbit_r69_c99 bl_99 br_99 wl_69 vdd gnd cell_6t
Xbit_r70_c99 bl_99 br_99 wl_70 vdd gnd cell_6t
Xbit_r71_c99 bl_99 br_99 wl_71 vdd gnd cell_6t
Xbit_r72_c99 bl_99 br_99 wl_72 vdd gnd cell_6t
Xbit_r73_c99 bl_99 br_99 wl_73 vdd gnd cell_6t
Xbit_r74_c99 bl_99 br_99 wl_74 vdd gnd cell_6t
Xbit_r75_c99 bl_99 br_99 wl_75 vdd gnd cell_6t
Xbit_r76_c99 bl_99 br_99 wl_76 vdd gnd cell_6t
Xbit_r77_c99 bl_99 br_99 wl_77 vdd gnd cell_6t
Xbit_r78_c99 bl_99 br_99 wl_78 vdd gnd cell_6t
Xbit_r79_c99 bl_99 br_99 wl_79 vdd gnd cell_6t
Xbit_r80_c99 bl_99 br_99 wl_80 vdd gnd cell_6t
Xbit_r81_c99 bl_99 br_99 wl_81 vdd gnd cell_6t
Xbit_r82_c99 bl_99 br_99 wl_82 vdd gnd cell_6t
Xbit_r83_c99 bl_99 br_99 wl_83 vdd gnd cell_6t
Xbit_r84_c99 bl_99 br_99 wl_84 vdd gnd cell_6t
Xbit_r85_c99 bl_99 br_99 wl_85 vdd gnd cell_6t
Xbit_r86_c99 bl_99 br_99 wl_86 vdd gnd cell_6t
Xbit_r87_c99 bl_99 br_99 wl_87 vdd gnd cell_6t
Xbit_r88_c99 bl_99 br_99 wl_88 vdd gnd cell_6t
Xbit_r89_c99 bl_99 br_99 wl_89 vdd gnd cell_6t
Xbit_r90_c99 bl_99 br_99 wl_90 vdd gnd cell_6t
Xbit_r91_c99 bl_99 br_99 wl_91 vdd gnd cell_6t
Xbit_r92_c99 bl_99 br_99 wl_92 vdd gnd cell_6t
Xbit_r93_c99 bl_99 br_99 wl_93 vdd gnd cell_6t
Xbit_r94_c99 bl_99 br_99 wl_94 vdd gnd cell_6t
Xbit_r95_c99 bl_99 br_99 wl_95 vdd gnd cell_6t
Xbit_r96_c99 bl_99 br_99 wl_96 vdd gnd cell_6t
Xbit_r97_c99 bl_99 br_99 wl_97 vdd gnd cell_6t
Xbit_r98_c99 bl_99 br_99 wl_98 vdd gnd cell_6t
Xbit_r99_c99 bl_99 br_99 wl_99 vdd gnd cell_6t
Xbit_r100_c99 bl_99 br_99 wl_100 vdd gnd cell_6t
Xbit_r101_c99 bl_99 br_99 wl_101 vdd gnd cell_6t
Xbit_r102_c99 bl_99 br_99 wl_102 vdd gnd cell_6t
Xbit_r103_c99 bl_99 br_99 wl_103 vdd gnd cell_6t
Xbit_r104_c99 bl_99 br_99 wl_104 vdd gnd cell_6t
Xbit_r105_c99 bl_99 br_99 wl_105 vdd gnd cell_6t
Xbit_r106_c99 bl_99 br_99 wl_106 vdd gnd cell_6t
Xbit_r107_c99 bl_99 br_99 wl_107 vdd gnd cell_6t
Xbit_r108_c99 bl_99 br_99 wl_108 vdd gnd cell_6t
Xbit_r109_c99 bl_99 br_99 wl_109 vdd gnd cell_6t
Xbit_r110_c99 bl_99 br_99 wl_110 vdd gnd cell_6t
Xbit_r111_c99 bl_99 br_99 wl_111 vdd gnd cell_6t
Xbit_r112_c99 bl_99 br_99 wl_112 vdd gnd cell_6t
Xbit_r113_c99 bl_99 br_99 wl_113 vdd gnd cell_6t
Xbit_r114_c99 bl_99 br_99 wl_114 vdd gnd cell_6t
Xbit_r115_c99 bl_99 br_99 wl_115 vdd gnd cell_6t
Xbit_r116_c99 bl_99 br_99 wl_116 vdd gnd cell_6t
Xbit_r117_c99 bl_99 br_99 wl_117 vdd gnd cell_6t
Xbit_r118_c99 bl_99 br_99 wl_118 vdd gnd cell_6t
Xbit_r119_c99 bl_99 br_99 wl_119 vdd gnd cell_6t
Xbit_r120_c99 bl_99 br_99 wl_120 vdd gnd cell_6t
Xbit_r121_c99 bl_99 br_99 wl_121 vdd gnd cell_6t
Xbit_r122_c99 bl_99 br_99 wl_122 vdd gnd cell_6t
Xbit_r123_c99 bl_99 br_99 wl_123 vdd gnd cell_6t
Xbit_r124_c99 bl_99 br_99 wl_124 vdd gnd cell_6t
Xbit_r125_c99 bl_99 br_99 wl_125 vdd gnd cell_6t
Xbit_r126_c99 bl_99 br_99 wl_126 vdd gnd cell_6t
Xbit_r127_c99 bl_99 br_99 wl_127 vdd gnd cell_6t
Xbit_r128_c99 bl_99 br_99 wl_128 vdd gnd cell_6t
Xbit_r129_c99 bl_99 br_99 wl_129 vdd gnd cell_6t
Xbit_r130_c99 bl_99 br_99 wl_130 vdd gnd cell_6t
Xbit_r131_c99 bl_99 br_99 wl_131 vdd gnd cell_6t
Xbit_r132_c99 bl_99 br_99 wl_132 vdd gnd cell_6t
Xbit_r133_c99 bl_99 br_99 wl_133 vdd gnd cell_6t
Xbit_r134_c99 bl_99 br_99 wl_134 vdd gnd cell_6t
Xbit_r135_c99 bl_99 br_99 wl_135 vdd gnd cell_6t
Xbit_r136_c99 bl_99 br_99 wl_136 vdd gnd cell_6t
Xbit_r137_c99 bl_99 br_99 wl_137 vdd gnd cell_6t
Xbit_r138_c99 bl_99 br_99 wl_138 vdd gnd cell_6t
Xbit_r139_c99 bl_99 br_99 wl_139 vdd gnd cell_6t
Xbit_r140_c99 bl_99 br_99 wl_140 vdd gnd cell_6t
Xbit_r141_c99 bl_99 br_99 wl_141 vdd gnd cell_6t
Xbit_r142_c99 bl_99 br_99 wl_142 vdd gnd cell_6t
Xbit_r143_c99 bl_99 br_99 wl_143 vdd gnd cell_6t
Xbit_r144_c99 bl_99 br_99 wl_144 vdd gnd cell_6t
Xbit_r145_c99 bl_99 br_99 wl_145 vdd gnd cell_6t
Xbit_r146_c99 bl_99 br_99 wl_146 vdd gnd cell_6t
Xbit_r147_c99 bl_99 br_99 wl_147 vdd gnd cell_6t
Xbit_r148_c99 bl_99 br_99 wl_148 vdd gnd cell_6t
Xbit_r149_c99 bl_99 br_99 wl_149 vdd gnd cell_6t
Xbit_r150_c99 bl_99 br_99 wl_150 vdd gnd cell_6t
Xbit_r151_c99 bl_99 br_99 wl_151 vdd gnd cell_6t
Xbit_r152_c99 bl_99 br_99 wl_152 vdd gnd cell_6t
Xbit_r153_c99 bl_99 br_99 wl_153 vdd gnd cell_6t
Xbit_r154_c99 bl_99 br_99 wl_154 vdd gnd cell_6t
Xbit_r155_c99 bl_99 br_99 wl_155 vdd gnd cell_6t
Xbit_r156_c99 bl_99 br_99 wl_156 vdd gnd cell_6t
Xbit_r157_c99 bl_99 br_99 wl_157 vdd gnd cell_6t
Xbit_r158_c99 bl_99 br_99 wl_158 vdd gnd cell_6t
Xbit_r159_c99 bl_99 br_99 wl_159 vdd gnd cell_6t
Xbit_r160_c99 bl_99 br_99 wl_160 vdd gnd cell_6t
Xbit_r161_c99 bl_99 br_99 wl_161 vdd gnd cell_6t
Xbit_r162_c99 bl_99 br_99 wl_162 vdd gnd cell_6t
Xbit_r163_c99 bl_99 br_99 wl_163 vdd gnd cell_6t
Xbit_r164_c99 bl_99 br_99 wl_164 vdd gnd cell_6t
Xbit_r165_c99 bl_99 br_99 wl_165 vdd gnd cell_6t
Xbit_r166_c99 bl_99 br_99 wl_166 vdd gnd cell_6t
Xbit_r167_c99 bl_99 br_99 wl_167 vdd gnd cell_6t
Xbit_r168_c99 bl_99 br_99 wl_168 vdd gnd cell_6t
Xbit_r169_c99 bl_99 br_99 wl_169 vdd gnd cell_6t
Xbit_r170_c99 bl_99 br_99 wl_170 vdd gnd cell_6t
Xbit_r171_c99 bl_99 br_99 wl_171 vdd gnd cell_6t
Xbit_r172_c99 bl_99 br_99 wl_172 vdd gnd cell_6t
Xbit_r173_c99 bl_99 br_99 wl_173 vdd gnd cell_6t
Xbit_r174_c99 bl_99 br_99 wl_174 vdd gnd cell_6t
Xbit_r175_c99 bl_99 br_99 wl_175 vdd gnd cell_6t
Xbit_r176_c99 bl_99 br_99 wl_176 vdd gnd cell_6t
Xbit_r177_c99 bl_99 br_99 wl_177 vdd gnd cell_6t
Xbit_r178_c99 bl_99 br_99 wl_178 vdd gnd cell_6t
Xbit_r179_c99 bl_99 br_99 wl_179 vdd gnd cell_6t
Xbit_r180_c99 bl_99 br_99 wl_180 vdd gnd cell_6t
Xbit_r181_c99 bl_99 br_99 wl_181 vdd gnd cell_6t
Xbit_r182_c99 bl_99 br_99 wl_182 vdd gnd cell_6t
Xbit_r183_c99 bl_99 br_99 wl_183 vdd gnd cell_6t
Xbit_r184_c99 bl_99 br_99 wl_184 vdd gnd cell_6t
Xbit_r185_c99 bl_99 br_99 wl_185 vdd gnd cell_6t
Xbit_r186_c99 bl_99 br_99 wl_186 vdd gnd cell_6t
Xbit_r187_c99 bl_99 br_99 wl_187 vdd gnd cell_6t
Xbit_r188_c99 bl_99 br_99 wl_188 vdd gnd cell_6t
Xbit_r189_c99 bl_99 br_99 wl_189 vdd gnd cell_6t
Xbit_r190_c99 bl_99 br_99 wl_190 vdd gnd cell_6t
Xbit_r191_c99 bl_99 br_99 wl_191 vdd gnd cell_6t
Xbit_r192_c99 bl_99 br_99 wl_192 vdd gnd cell_6t
Xbit_r193_c99 bl_99 br_99 wl_193 vdd gnd cell_6t
Xbit_r194_c99 bl_99 br_99 wl_194 vdd gnd cell_6t
Xbit_r195_c99 bl_99 br_99 wl_195 vdd gnd cell_6t
Xbit_r196_c99 bl_99 br_99 wl_196 vdd gnd cell_6t
Xbit_r197_c99 bl_99 br_99 wl_197 vdd gnd cell_6t
Xbit_r198_c99 bl_99 br_99 wl_198 vdd gnd cell_6t
Xbit_r199_c99 bl_99 br_99 wl_199 vdd gnd cell_6t
Xbit_r200_c99 bl_99 br_99 wl_200 vdd gnd cell_6t
Xbit_r201_c99 bl_99 br_99 wl_201 vdd gnd cell_6t
Xbit_r202_c99 bl_99 br_99 wl_202 vdd gnd cell_6t
Xbit_r203_c99 bl_99 br_99 wl_203 vdd gnd cell_6t
Xbit_r204_c99 bl_99 br_99 wl_204 vdd gnd cell_6t
Xbit_r205_c99 bl_99 br_99 wl_205 vdd gnd cell_6t
Xbit_r206_c99 bl_99 br_99 wl_206 vdd gnd cell_6t
Xbit_r207_c99 bl_99 br_99 wl_207 vdd gnd cell_6t
Xbit_r208_c99 bl_99 br_99 wl_208 vdd gnd cell_6t
Xbit_r209_c99 bl_99 br_99 wl_209 vdd gnd cell_6t
Xbit_r210_c99 bl_99 br_99 wl_210 vdd gnd cell_6t
Xbit_r211_c99 bl_99 br_99 wl_211 vdd gnd cell_6t
Xbit_r212_c99 bl_99 br_99 wl_212 vdd gnd cell_6t
Xbit_r213_c99 bl_99 br_99 wl_213 vdd gnd cell_6t
Xbit_r214_c99 bl_99 br_99 wl_214 vdd gnd cell_6t
Xbit_r215_c99 bl_99 br_99 wl_215 vdd gnd cell_6t
Xbit_r216_c99 bl_99 br_99 wl_216 vdd gnd cell_6t
Xbit_r217_c99 bl_99 br_99 wl_217 vdd gnd cell_6t
Xbit_r218_c99 bl_99 br_99 wl_218 vdd gnd cell_6t
Xbit_r219_c99 bl_99 br_99 wl_219 vdd gnd cell_6t
Xbit_r220_c99 bl_99 br_99 wl_220 vdd gnd cell_6t
Xbit_r221_c99 bl_99 br_99 wl_221 vdd gnd cell_6t
Xbit_r222_c99 bl_99 br_99 wl_222 vdd gnd cell_6t
Xbit_r223_c99 bl_99 br_99 wl_223 vdd gnd cell_6t
Xbit_r224_c99 bl_99 br_99 wl_224 vdd gnd cell_6t
Xbit_r225_c99 bl_99 br_99 wl_225 vdd gnd cell_6t
Xbit_r226_c99 bl_99 br_99 wl_226 vdd gnd cell_6t
Xbit_r227_c99 bl_99 br_99 wl_227 vdd gnd cell_6t
Xbit_r228_c99 bl_99 br_99 wl_228 vdd gnd cell_6t
Xbit_r229_c99 bl_99 br_99 wl_229 vdd gnd cell_6t
Xbit_r230_c99 bl_99 br_99 wl_230 vdd gnd cell_6t
Xbit_r231_c99 bl_99 br_99 wl_231 vdd gnd cell_6t
Xbit_r232_c99 bl_99 br_99 wl_232 vdd gnd cell_6t
Xbit_r233_c99 bl_99 br_99 wl_233 vdd gnd cell_6t
Xbit_r234_c99 bl_99 br_99 wl_234 vdd gnd cell_6t
Xbit_r235_c99 bl_99 br_99 wl_235 vdd gnd cell_6t
Xbit_r236_c99 bl_99 br_99 wl_236 vdd gnd cell_6t
Xbit_r237_c99 bl_99 br_99 wl_237 vdd gnd cell_6t
Xbit_r238_c99 bl_99 br_99 wl_238 vdd gnd cell_6t
Xbit_r239_c99 bl_99 br_99 wl_239 vdd gnd cell_6t
Xbit_r240_c99 bl_99 br_99 wl_240 vdd gnd cell_6t
Xbit_r241_c99 bl_99 br_99 wl_241 vdd gnd cell_6t
Xbit_r242_c99 bl_99 br_99 wl_242 vdd gnd cell_6t
Xbit_r243_c99 bl_99 br_99 wl_243 vdd gnd cell_6t
Xbit_r244_c99 bl_99 br_99 wl_244 vdd gnd cell_6t
Xbit_r245_c99 bl_99 br_99 wl_245 vdd gnd cell_6t
Xbit_r246_c99 bl_99 br_99 wl_246 vdd gnd cell_6t
Xbit_r247_c99 bl_99 br_99 wl_247 vdd gnd cell_6t
Xbit_r248_c99 bl_99 br_99 wl_248 vdd gnd cell_6t
Xbit_r249_c99 bl_99 br_99 wl_249 vdd gnd cell_6t
Xbit_r250_c99 bl_99 br_99 wl_250 vdd gnd cell_6t
Xbit_r251_c99 bl_99 br_99 wl_251 vdd gnd cell_6t
Xbit_r252_c99 bl_99 br_99 wl_252 vdd gnd cell_6t
Xbit_r253_c99 bl_99 br_99 wl_253 vdd gnd cell_6t
Xbit_r254_c99 bl_99 br_99 wl_254 vdd gnd cell_6t
Xbit_r255_c99 bl_99 br_99 wl_255 vdd gnd cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd cell_6t
Xbit_r1_c100 bl_100 br_100 wl_1 vdd gnd cell_6t
Xbit_r2_c100 bl_100 br_100 wl_2 vdd gnd cell_6t
Xbit_r3_c100 bl_100 br_100 wl_3 vdd gnd cell_6t
Xbit_r4_c100 bl_100 br_100 wl_4 vdd gnd cell_6t
Xbit_r5_c100 bl_100 br_100 wl_5 vdd gnd cell_6t
Xbit_r6_c100 bl_100 br_100 wl_6 vdd gnd cell_6t
Xbit_r7_c100 bl_100 br_100 wl_7 vdd gnd cell_6t
Xbit_r8_c100 bl_100 br_100 wl_8 vdd gnd cell_6t
Xbit_r9_c100 bl_100 br_100 wl_9 vdd gnd cell_6t
Xbit_r10_c100 bl_100 br_100 wl_10 vdd gnd cell_6t
Xbit_r11_c100 bl_100 br_100 wl_11 vdd gnd cell_6t
Xbit_r12_c100 bl_100 br_100 wl_12 vdd gnd cell_6t
Xbit_r13_c100 bl_100 br_100 wl_13 vdd gnd cell_6t
Xbit_r14_c100 bl_100 br_100 wl_14 vdd gnd cell_6t
Xbit_r15_c100 bl_100 br_100 wl_15 vdd gnd cell_6t
Xbit_r16_c100 bl_100 br_100 wl_16 vdd gnd cell_6t
Xbit_r17_c100 bl_100 br_100 wl_17 vdd gnd cell_6t
Xbit_r18_c100 bl_100 br_100 wl_18 vdd gnd cell_6t
Xbit_r19_c100 bl_100 br_100 wl_19 vdd gnd cell_6t
Xbit_r20_c100 bl_100 br_100 wl_20 vdd gnd cell_6t
Xbit_r21_c100 bl_100 br_100 wl_21 vdd gnd cell_6t
Xbit_r22_c100 bl_100 br_100 wl_22 vdd gnd cell_6t
Xbit_r23_c100 bl_100 br_100 wl_23 vdd gnd cell_6t
Xbit_r24_c100 bl_100 br_100 wl_24 vdd gnd cell_6t
Xbit_r25_c100 bl_100 br_100 wl_25 vdd gnd cell_6t
Xbit_r26_c100 bl_100 br_100 wl_26 vdd gnd cell_6t
Xbit_r27_c100 bl_100 br_100 wl_27 vdd gnd cell_6t
Xbit_r28_c100 bl_100 br_100 wl_28 vdd gnd cell_6t
Xbit_r29_c100 bl_100 br_100 wl_29 vdd gnd cell_6t
Xbit_r30_c100 bl_100 br_100 wl_30 vdd gnd cell_6t
Xbit_r31_c100 bl_100 br_100 wl_31 vdd gnd cell_6t
Xbit_r32_c100 bl_100 br_100 wl_32 vdd gnd cell_6t
Xbit_r33_c100 bl_100 br_100 wl_33 vdd gnd cell_6t
Xbit_r34_c100 bl_100 br_100 wl_34 vdd gnd cell_6t
Xbit_r35_c100 bl_100 br_100 wl_35 vdd gnd cell_6t
Xbit_r36_c100 bl_100 br_100 wl_36 vdd gnd cell_6t
Xbit_r37_c100 bl_100 br_100 wl_37 vdd gnd cell_6t
Xbit_r38_c100 bl_100 br_100 wl_38 vdd gnd cell_6t
Xbit_r39_c100 bl_100 br_100 wl_39 vdd gnd cell_6t
Xbit_r40_c100 bl_100 br_100 wl_40 vdd gnd cell_6t
Xbit_r41_c100 bl_100 br_100 wl_41 vdd gnd cell_6t
Xbit_r42_c100 bl_100 br_100 wl_42 vdd gnd cell_6t
Xbit_r43_c100 bl_100 br_100 wl_43 vdd gnd cell_6t
Xbit_r44_c100 bl_100 br_100 wl_44 vdd gnd cell_6t
Xbit_r45_c100 bl_100 br_100 wl_45 vdd gnd cell_6t
Xbit_r46_c100 bl_100 br_100 wl_46 vdd gnd cell_6t
Xbit_r47_c100 bl_100 br_100 wl_47 vdd gnd cell_6t
Xbit_r48_c100 bl_100 br_100 wl_48 vdd gnd cell_6t
Xbit_r49_c100 bl_100 br_100 wl_49 vdd gnd cell_6t
Xbit_r50_c100 bl_100 br_100 wl_50 vdd gnd cell_6t
Xbit_r51_c100 bl_100 br_100 wl_51 vdd gnd cell_6t
Xbit_r52_c100 bl_100 br_100 wl_52 vdd gnd cell_6t
Xbit_r53_c100 bl_100 br_100 wl_53 vdd gnd cell_6t
Xbit_r54_c100 bl_100 br_100 wl_54 vdd gnd cell_6t
Xbit_r55_c100 bl_100 br_100 wl_55 vdd gnd cell_6t
Xbit_r56_c100 bl_100 br_100 wl_56 vdd gnd cell_6t
Xbit_r57_c100 bl_100 br_100 wl_57 vdd gnd cell_6t
Xbit_r58_c100 bl_100 br_100 wl_58 vdd gnd cell_6t
Xbit_r59_c100 bl_100 br_100 wl_59 vdd gnd cell_6t
Xbit_r60_c100 bl_100 br_100 wl_60 vdd gnd cell_6t
Xbit_r61_c100 bl_100 br_100 wl_61 vdd gnd cell_6t
Xbit_r62_c100 bl_100 br_100 wl_62 vdd gnd cell_6t
Xbit_r63_c100 bl_100 br_100 wl_63 vdd gnd cell_6t
Xbit_r64_c100 bl_100 br_100 wl_64 vdd gnd cell_6t
Xbit_r65_c100 bl_100 br_100 wl_65 vdd gnd cell_6t
Xbit_r66_c100 bl_100 br_100 wl_66 vdd gnd cell_6t
Xbit_r67_c100 bl_100 br_100 wl_67 vdd gnd cell_6t
Xbit_r68_c100 bl_100 br_100 wl_68 vdd gnd cell_6t
Xbit_r69_c100 bl_100 br_100 wl_69 vdd gnd cell_6t
Xbit_r70_c100 bl_100 br_100 wl_70 vdd gnd cell_6t
Xbit_r71_c100 bl_100 br_100 wl_71 vdd gnd cell_6t
Xbit_r72_c100 bl_100 br_100 wl_72 vdd gnd cell_6t
Xbit_r73_c100 bl_100 br_100 wl_73 vdd gnd cell_6t
Xbit_r74_c100 bl_100 br_100 wl_74 vdd gnd cell_6t
Xbit_r75_c100 bl_100 br_100 wl_75 vdd gnd cell_6t
Xbit_r76_c100 bl_100 br_100 wl_76 vdd gnd cell_6t
Xbit_r77_c100 bl_100 br_100 wl_77 vdd gnd cell_6t
Xbit_r78_c100 bl_100 br_100 wl_78 vdd gnd cell_6t
Xbit_r79_c100 bl_100 br_100 wl_79 vdd gnd cell_6t
Xbit_r80_c100 bl_100 br_100 wl_80 vdd gnd cell_6t
Xbit_r81_c100 bl_100 br_100 wl_81 vdd gnd cell_6t
Xbit_r82_c100 bl_100 br_100 wl_82 vdd gnd cell_6t
Xbit_r83_c100 bl_100 br_100 wl_83 vdd gnd cell_6t
Xbit_r84_c100 bl_100 br_100 wl_84 vdd gnd cell_6t
Xbit_r85_c100 bl_100 br_100 wl_85 vdd gnd cell_6t
Xbit_r86_c100 bl_100 br_100 wl_86 vdd gnd cell_6t
Xbit_r87_c100 bl_100 br_100 wl_87 vdd gnd cell_6t
Xbit_r88_c100 bl_100 br_100 wl_88 vdd gnd cell_6t
Xbit_r89_c100 bl_100 br_100 wl_89 vdd gnd cell_6t
Xbit_r90_c100 bl_100 br_100 wl_90 vdd gnd cell_6t
Xbit_r91_c100 bl_100 br_100 wl_91 vdd gnd cell_6t
Xbit_r92_c100 bl_100 br_100 wl_92 vdd gnd cell_6t
Xbit_r93_c100 bl_100 br_100 wl_93 vdd gnd cell_6t
Xbit_r94_c100 bl_100 br_100 wl_94 vdd gnd cell_6t
Xbit_r95_c100 bl_100 br_100 wl_95 vdd gnd cell_6t
Xbit_r96_c100 bl_100 br_100 wl_96 vdd gnd cell_6t
Xbit_r97_c100 bl_100 br_100 wl_97 vdd gnd cell_6t
Xbit_r98_c100 bl_100 br_100 wl_98 vdd gnd cell_6t
Xbit_r99_c100 bl_100 br_100 wl_99 vdd gnd cell_6t
Xbit_r100_c100 bl_100 br_100 wl_100 vdd gnd cell_6t
Xbit_r101_c100 bl_100 br_100 wl_101 vdd gnd cell_6t
Xbit_r102_c100 bl_100 br_100 wl_102 vdd gnd cell_6t
Xbit_r103_c100 bl_100 br_100 wl_103 vdd gnd cell_6t
Xbit_r104_c100 bl_100 br_100 wl_104 vdd gnd cell_6t
Xbit_r105_c100 bl_100 br_100 wl_105 vdd gnd cell_6t
Xbit_r106_c100 bl_100 br_100 wl_106 vdd gnd cell_6t
Xbit_r107_c100 bl_100 br_100 wl_107 vdd gnd cell_6t
Xbit_r108_c100 bl_100 br_100 wl_108 vdd gnd cell_6t
Xbit_r109_c100 bl_100 br_100 wl_109 vdd gnd cell_6t
Xbit_r110_c100 bl_100 br_100 wl_110 vdd gnd cell_6t
Xbit_r111_c100 bl_100 br_100 wl_111 vdd gnd cell_6t
Xbit_r112_c100 bl_100 br_100 wl_112 vdd gnd cell_6t
Xbit_r113_c100 bl_100 br_100 wl_113 vdd gnd cell_6t
Xbit_r114_c100 bl_100 br_100 wl_114 vdd gnd cell_6t
Xbit_r115_c100 bl_100 br_100 wl_115 vdd gnd cell_6t
Xbit_r116_c100 bl_100 br_100 wl_116 vdd gnd cell_6t
Xbit_r117_c100 bl_100 br_100 wl_117 vdd gnd cell_6t
Xbit_r118_c100 bl_100 br_100 wl_118 vdd gnd cell_6t
Xbit_r119_c100 bl_100 br_100 wl_119 vdd gnd cell_6t
Xbit_r120_c100 bl_100 br_100 wl_120 vdd gnd cell_6t
Xbit_r121_c100 bl_100 br_100 wl_121 vdd gnd cell_6t
Xbit_r122_c100 bl_100 br_100 wl_122 vdd gnd cell_6t
Xbit_r123_c100 bl_100 br_100 wl_123 vdd gnd cell_6t
Xbit_r124_c100 bl_100 br_100 wl_124 vdd gnd cell_6t
Xbit_r125_c100 bl_100 br_100 wl_125 vdd gnd cell_6t
Xbit_r126_c100 bl_100 br_100 wl_126 vdd gnd cell_6t
Xbit_r127_c100 bl_100 br_100 wl_127 vdd gnd cell_6t
Xbit_r128_c100 bl_100 br_100 wl_128 vdd gnd cell_6t
Xbit_r129_c100 bl_100 br_100 wl_129 vdd gnd cell_6t
Xbit_r130_c100 bl_100 br_100 wl_130 vdd gnd cell_6t
Xbit_r131_c100 bl_100 br_100 wl_131 vdd gnd cell_6t
Xbit_r132_c100 bl_100 br_100 wl_132 vdd gnd cell_6t
Xbit_r133_c100 bl_100 br_100 wl_133 vdd gnd cell_6t
Xbit_r134_c100 bl_100 br_100 wl_134 vdd gnd cell_6t
Xbit_r135_c100 bl_100 br_100 wl_135 vdd gnd cell_6t
Xbit_r136_c100 bl_100 br_100 wl_136 vdd gnd cell_6t
Xbit_r137_c100 bl_100 br_100 wl_137 vdd gnd cell_6t
Xbit_r138_c100 bl_100 br_100 wl_138 vdd gnd cell_6t
Xbit_r139_c100 bl_100 br_100 wl_139 vdd gnd cell_6t
Xbit_r140_c100 bl_100 br_100 wl_140 vdd gnd cell_6t
Xbit_r141_c100 bl_100 br_100 wl_141 vdd gnd cell_6t
Xbit_r142_c100 bl_100 br_100 wl_142 vdd gnd cell_6t
Xbit_r143_c100 bl_100 br_100 wl_143 vdd gnd cell_6t
Xbit_r144_c100 bl_100 br_100 wl_144 vdd gnd cell_6t
Xbit_r145_c100 bl_100 br_100 wl_145 vdd gnd cell_6t
Xbit_r146_c100 bl_100 br_100 wl_146 vdd gnd cell_6t
Xbit_r147_c100 bl_100 br_100 wl_147 vdd gnd cell_6t
Xbit_r148_c100 bl_100 br_100 wl_148 vdd gnd cell_6t
Xbit_r149_c100 bl_100 br_100 wl_149 vdd gnd cell_6t
Xbit_r150_c100 bl_100 br_100 wl_150 vdd gnd cell_6t
Xbit_r151_c100 bl_100 br_100 wl_151 vdd gnd cell_6t
Xbit_r152_c100 bl_100 br_100 wl_152 vdd gnd cell_6t
Xbit_r153_c100 bl_100 br_100 wl_153 vdd gnd cell_6t
Xbit_r154_c100 bl_100 br_100 wl_154 vdd gnd cell_6t
Xbit_r155_c100 bl_100 br_100 wl_155 vdd gnd cell_6t
Xbit_r156_c100 bl_100 br_100 wl_156 vdd gnd cell_6t
Xbit_r157_c100 bl_100 br_100 wl_157 vdd gnd cell_6t
Xbit_r158_c100 bl_100 br_100 wl_158 vdd gnd cell_6t
Xbit_r159_c100 bl_100 br_100 wl_159 vdd gnd cell_6t
Xbit_r160_c100 bl_100 br_100 wl_160 vdd gnd cell_6t
Xbit_r161_c100 bl_100 br_100 wl_161 vdd gnd cell_6t
Xbit_r162_c100 bl_100 br_100 wl_162 vdd gnd cell_6t
Xbit_r163_c100 bl_100 br_100 wl_163 vdd gnd cell_6t
Xbit_r164_c100 bl_100 br_100 wl_164 vdd gnd cell_6t
Xbit_r165_c100 bl_100 br_100 wl_165 vdd gnd cell_6t
Xbit_r166_c100 bl_100 br_100 wl_166 vdd gnd cell_6t
Xbit_r167_c100 bl_100 br_100 wl_167 vdd gnd cell_6t
Xbit_r168_c100 bl_100 br_100 wl_168 vdd gnd cell_6t
Xbit_r169_c100 bl_100 br_100 wl_169 vdd gnd cell_6t
Xbit_r170_c100 bl_100 br_100 wl_170 vdd gnd cell_6t
Xbit_r171_c100 bl_100 br_100 wl_171 vdd gnd cell_6t
Xbit_r172_c100 bl_100 br_100 wl_172 vdd gnd cell_6t
Xbit_r173_c100 bl_100 br_100 wl_173 vdd gnd cell_6t
Xbit_r174_c100 bl_100 br_100 wl_174 vdd gnd cell_6t
Xbit_r175_c100 bl_100 br_100 wl_175 vdd gnd cell_6t
Xbit_r176_c100 bl_100 br_100 wl_176 vdd gnd cell_6t
Xbit_r177_c100 bl_100 br_100 wl_177 vdd gnd cell_6t
Xbit_r178_c100 bl_100 br_100 wl_178 vdd gnd cell_6t
Xbit_r179_c100 bl_100 br_100 wl_179 vdd gnd cell_6t
Xbit_r180_c100 bl_100 br_100 wl_180 vdd gnd cell_6t
Xbit_r181_c100 bl_100 br_100 wl_181 vdd gnd cell_6t
Xbit_r182_c100 bl_100 br_100 wl_182 vdd gnd cell_6t
Xbit_r183_c100 bl_100 br_100 wl_183 vdd gnd cell_6t
Xbit_r184_c100 bl_100 br_100 wl_184 vdd gnd cell_6t
Xbit_r185_c100 bl_100 br_100 wl_185 vdd gnd cell_6t
Xbit_r186_c100 bl_100 br_100 wl_186 vdd gnd cell_6t
Xbit_r187_c100 bl_100 br_100 wl_187 vdd gnd cell_6t
Xbit_r188_c100 bl_100 br_100 wl_188 vdd gnd cell_6t
Xbit_r189_c100 bl_100 br_100 wl_189 vdd gnd cell_6t
Xbit_r190_c100 bl_100 br_100 wl_190 vdd gnd cell_6t
Xbit_r191_c100 bl_100 br_100 wl_191 vdd gnd cell_6t
Xbit_r192_c100 bl_100 br_100 wl_192 vdd gnd cell_6t
Xbit_r193_c100 bl_100 br_100 wl_193 vdd gnd cell_6t
Xbit_r194_c100 bl_100 br_100 wl_194 vdd gnd cell_6t
Xbit_r195_c100 bl_100 br_100 wl_195 vdd gnd cell_6t
Xbit_r196_c100 bl_100 br_100 wl_196 vdd gnd cell_6t
Xbit_r197_c100 bl_100 br_100 wl_197 vdd gnd cell_6t
Xbit_r198_c100 bl_100 br_100 wl_198 vdd gnd cell_6t
Xbit_r199_c100 bl_100 br_100 wl_199 vdd gnd cell_6t
Xbit_r200_c100 bl_100 br_100 wl_200 vdd gnd cell_6t
Xbit_r201_c100 bl_100 br_100 wl_201 vdd gnd cell_6t
Xbit_r202_c100 bl_100 br_100 wl_202 vdd gnd cell_6t
Xbit_r203_c100 bl_100 br_100 wl_203 vdd gnd cell_6t
Xbit_r204_c100 bl_100 br_100 wl_204 vdd gnd cell_6t
Xbit_r205_c100 bl_100 br_100 wl_205 vdd gnd cell_6t
Xbit_r206_c100 bl_100 br_100 wl_206 vdd gnd cell_6t
Xbit_r207_c100 bl_100 br_100 wl_207 vdd gnd cell_6t
Xbit_r208_c100 bl_100 br_100 wl_208 vdd gnd cell_6t
Xbit_r209_c100 bl_100 br_100 wl_209 vdd gnd cell_6t
Xbit_r210_c100 bl_100 br_100 wl_210 vdd gnd cell_6t
Xbit_r211_c100 bl_100 br_100 wl_211 vdd gnd cell_6t
Xbit_r212_c100 bl_100 br_100 wl_212 vdd gnd cell_6t
Xbit_r213_c100 bl_100 br_100 wl_213 vdd gnd cell_6t
Xbit_r214_c100 bl_100 br_100 wl_214 vdd gnd cell_6t
Xbit_r215_c100 bl_100 br_100 wl_215 vdd gnd cell_6t
Xbit_r216_c100 bl_100 br_100 wl_216 vdd gnd cell_6t
Xbit_r217_c100 bl_100 br_100 wl_217 vdd gnd cell_6t
Xbit_r218_c100 bl_100 br_100 wl_218 vdd gnd cell_6t
Xbit_r219_c100 bl_100 br_100 wl_219 vdd gnd cell_6t
Xbit_r220_c100 bl_100 br_100 wl_220 vdd gnd cell_6t
Xbit_r221_c100 bl_100 br_100 wl_221 vdd gnd cell_6t
Xbit_r222_c100 bl_100 br_100 wl_222 vdd gnd cell_6t
Xbit_r223_c100 bl_100 br_100 wl_223 vdd gnd cell_6t
Xbit_r224_c100 bl_100 br_100 wl_224 vdd gnd cell_6t
Xbit_r225_c100 bl_100 br_100 wl_225 vdd gnd cell_6t
Xbit_r226_c100 bl_100 br_100 wl_226 vdd gnd cell_6t
Xbit_r227_c100 bl_100 br_100 wl_227 vdd gnd cell_6t
Xbit_r228_c100 bl_100 br_100 wl_228 vdd gnd cell_6t
Xbit_r229_c100 bl_100 br_100 wl_229 vdd gnd cell_6t
Xbit_r230_c100 bl_100 br_100 wl_230 vdd gnd cell_6t
Xbit_r231_c100 bl_100 br_100 wl_231 vdd gnd cell_6t
Xbit_r232_c100 bl_100 br_100 wl_232 vdd gnd cell_6t
Xbit_r233_c100 bl_100 br_100 wl_233 vdd gnd cell_6t
Xbit_r234_c100 bl_100 br_100 wl_234 vdd gnd cell_6t
Xbit_r235_c100 bl_100 br_100 wl_235 vdd gnd cell_6t
Xbit_r236_c100 bl_100 br_100 wl_236 vdd gnd cell_6t
Xbit_r237_c100 bl_100 br_100 wl_237 vdd gnd cell_6t
Xbit_r238_c100 bl_100 br_100 wl_238 vdd gnd cell_6t
Xbit_r239_c100 bl_100 br_100 wl_239 vdd gnd cell_6t
Xbit_r240_c100 bl_100 br_100 wl_240 vdd gnd cell_6t
Xbit_r241_c100 bl_100 br_100 wl_241 vdd gnd cell_6t
Xbit_r242_c100 bl_100 br_100 wl_242 vdd gnd cell_6t
Xbit_r243_c100 bl_100 br_100 wl_243 vdd gnd cell_6t
Xbit_r244_c100 bl_100 br_100 wl_244 vdd gnd cell_6t
Xbit_r245_c100 bl_100 br_100 wl_245 vdd gnd cell_6t
Xbit_r246_c100 bl_100 br_100 wl_246 vdd gnd cell_6t
Xbit_r247_c100 bl_100 br_100 wl_247 vdd gnd cell_6t
Xbit_r248_c100 bl_100 br_100 wl_248 vdd gnd cell_6t
Xbit_r249_c100 bl_100 br_100 wl_249 vdd gnd cell_6t
Xbit_r250_c100 bl_100 br_100 wl_250 vdd gnd cell_6t
Xbit_r251_c100 bl_100 br_100 wl_251 vdd gnd cell_6t
Xbit_r252_c100 bl_100 br_100 wl_252 vdd gnd cell_6t
Xbit_r253_c100 bl_100 br_100 wl_253 vdd gnd cell_6t
Xbit_r254_c100 bl_100 br_100 wl_254 vdd gnd cell_6t
Xbit_r255_c100 bl_100 br_100 wl_255 vdd gnd cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd cell_6t
Xbit_r1_c101 bl_101 br_101 wl_1 vdd gnd cell_6t
Xbit_r2_c101 bl_101 br_101 wl_2 vdd gnd cell_6t
Xbit_r3_c101 bl_101 br_101 wl_3 vdd gnd cell_6t
Xbit_r4_c101 bl_101 br_101 wl_4 vdd gnd cell_6t
Xbit_r5_c101 bl_101 br_101 wl_5 vdd gnd cell_6t
Xbit_r6_c101 bl_101 br_101 wl_6 vdd gnd cell_6t
Xbit_r7_c101 bl_101 br_101 wl_7 vdd gnd cell_6t
Xbit_r8_c101 bl_101 br_101 wl_8 vdd gnd cell_6t
Xbit_r9_c101 bl_101 br_101 wl_9 vdd gnd cell_6t
Xbit_r10_c101 bl_101 br_101 wl_10 vdd gnd cell_6t
Xbit_r11_c101 bl_101 br_101 wl_11 vdd gnd cell_6t
Xbit_r12_c101 bl_101 br_101 wl_12 vdd gnd cell_6t
Xbit_r13_c101 bl_101 br_101 wl_13 vdd gnd cell_6t
Xbit_r14_c101 bl_101 br_101 wl_14 vdd gnd cell_6t
Xbit_r15_c101 bl_101 br_101 wl_15 vdd gnd cell_6t
Xbit_r16_c101 bl_101 br_101 wl_16 vdd gnd cell_6t
Xbit_r17_c101 bl_101 br_101 wl_17 vdd gnd cell_6t
Xbit_r18_c101 bl_101 br_101 wl_18 vdd gnd cell_6t
Xbit_r19_c101 bl_101 br_101 wl_19 vdd gnd cell_6t
Xbit_r20_c101 bl_101 br_101 wl_20 vdd gnd cell_6t
Xbit_r21_c101 bl_101 br_101 wl_21 vdd gnd cell_6t
Xbit_r22_c101 bl_101 br_101 wl_22 vdd gnd cell_6t
Xbit_r23_c101 bl_101 br_101 wl_23 vdd gnd cell_6t
Xbit_r24_c101 bl_101 br_101 wl_24 vdd gnd cell_6t
Xbit_r25_c101 bl_101 br_101 wl_25 vdd gnd cell_6t
Xbit_r26_c101 bl_101 br_101 wl_26 vdd gnd cell_6t
Xbit_r27_c101 bl_101 br_101 wl_27 vdd gnd cell_6t
Xbit_r28_c101 bl_101 br_101 wl_28 vdd gnd cell_6t
Xbit_r29_c101 bl_101 br_101 wl_29 vdd gnd cell_6t
Xbit_r30_c101 bl_101 br_101 wl_30 vdd gnd cell_6t
Xbit_r31_c101 bl_101 br_101 wl_31 vdd gnd cell_6t
Xbit_r32_c101 bl_101 br_101 wl_32 vdd gnd cell_6t
Xbit_r33_c101 bl_101 br_101 wl_33 vdd gnd cell_6t
Xbit_r34_c101 bl_101 br_101 wl_34 vdd gnd cell_6t
Xbit_r35_c101 bl_101 br_101 wl_35 vdd gnd cell_6t
Xbit_r36_c101 bl_101 br_101 wl_36 vdd gnd cell_6t
Xbit_r37_c101 bl_101 br_101 wl_37 vdd gnd cell_6t
Xbit_r38_c101 bl_101 br_101 wl_38 vdd gnd cell_6t
Xbit_r39_c101 bl_101 br_101 wl_39 vdd gnd cell_6t
Xbit_r40_c101 bl_101 br_101 wl_40 vdd gnd cell_6t
Xbit_r41_c101 bl_101 br_101 wl_41 vdd gnd cell_6t
Xbit_r42_c101 bl_101 br_101 wl_42 vdd gnd cell_6t
Xbit_r43_c101 bl_101 br_101 wl_43 vdd gnd cell_6t
Xbit_r44_c101 bl_101 br_101 wl_44 vdd gnd cell_6t
Xbit_r45_c101 bl_101 br_101 wl_45 vdd gnd cell_6t
Xbit_r46_c101 bl_101 br_101 wl_46 vdd gnd cell_6t
Xbit_r47_c101 bl_101 br_101 wl_47 vdd gnd cell_6t
Xbit_r48_c101 bl_101 br_101 wl_48 vdd gnd cell_6t
Xbit_r49_c101 bl_101 br_101 wl_49 vdd gnd cell_6t
Xbit_r50_c101 bl_101 br_101 wl_50 vdd gnd cell_6t
Xbit_r51_c101 bl_101 br_101 wl_51 vdd gnd cell_6t
Xbit_r52_c101 bl_101 br_101 wl_52 vdd gnd cell_6t
Xbit_r53_c101 bl_101 br_101 wl_53 vdd gnd cell_6t
Xbit_r54_c101 bl_101 br_101 wl_54 vdd gnd cell_6t
Xbit_r55_c101 bl_101 br_101 wl_55 vdd gnd cell_6t
Xbit_r56_c101 bl_101 br_101 wl_56 vdd gnd cell_6t
Xbit_r57_c101 bl_101 br_101 wl_57 vdd gnd cell_6t
Xbit_r58_c101 bl_101 br_101 wl_58 vdd gnd cell_6t
Xbit_r59_c101 bl_101 br_101 wl_59 vdd gnd cell_6t
Xbit_r60_c101 bl_101 br_101 wl_60 vdd gnd cell_6t
Xbit_r61_c101 bl_101 br_101 wl_61 vdd gnd cell_6t
Xbit_r62_c101 bl_101 br_101 wl_62 vdd gnd cell_6t
Xbit_r63_c101 bl_101 br_101 wl_63 vdd gnd cell_6t
Xbit_r64_c101 bl_101 br_101 wl_64 vdd gnd cell_6t
Xbit_r65_c101 bl_101 br_101 wl_65 vdd gnd cell_6t
Xbit_r66_c101 bl_101 br_101 wl_66 vdd gnd cell_6t
Xbit_r67_c101 bl_101 br_101 wl_67 vdd gnd cell_6t
Xbit_r68_c101 bl_101 br_101 wl_68 vdd gnd cell_6t
Xbit_r69_c101 bl_101 br_101 wl_69 vdd gnd cell_6t
Xbit_r70_c101 bl_101 br_101 wl_70 vdd gnd cell_6t
Xbit_r71_c101 bl_101 br_101 wl_71 vdd gnd cell_6t
Xbit_r72_c101 bl_101 br_101 wl_72 vdd gnd cell_6t
Xbit_r73_c101 bl_101 br_101 wl_73 vdd gnd cell_6t
Xbit_r74_c101 bl_101 br_101 wl_74 vdd gnd cell_6t
Xbit_r75_c101 bl_101 br_101 wl_75 vdd gnd cell_6t
Xbit_r76_c101 bl_101 br_101 wl_76 vdd gnd cell_6t
Xbit_r77_c101 bl_101 br_101 wl_77 vdd gnd cell_6t
Xbit_r78_c101 bl_101 br_101 wl_78 vdd gnd cell_6t
Xbit_r79_c101 bl_101 br_101 wl_79 vdd gnd cell_6t
Xbit_r80_c101 bl_101 br_101 wl_80 vdd gnd cell_6t
Xbit_r81_c101 bl_101 br_101 wl_81 vdd gnd cell_6t
Xbit_r82_c101 bl_101 br_101 wl_82 vdd gnd cell_6t
Xbit_r83_c101 bl_101 br_101 wl_83 vdd gnd cell_6t
Xbit_r84_c101 bl_101 br_101 wl_84 vdd gnd cell_6t
Xbit_r85_c101 bl_101 br_101 wl_85 vdd gnd cell_6t
Xbit_r86_c101 bl_101 br_101 wl_86 vdd gnd cell_6t
Xbit_r87_c101 bl_101 br_101 wl_87 vdd gnd cell_6t
Xbit_r88_c101 bl_101 br_101 wl_88 vdd gnd cell_6t
Xbit_r89_c101 bl_101 br_101 wl_89 vdd gnd cell_6t
Xbit_r90_c101 bl_101 br_101 wl_90 vdd gnd cell_6t
Xbit_r91_c101 bl_101 br_101 wl_91 vdd gnd cell_6t
Xbit_r92_c101 bl_101 br_101 wl_92 vdd gnd cell_6t
Xbit_r93_c101 bl_101 br_101 wl_93 vdd gnd cell_6t
Xbit_r94_c101 bl_101 br_101 wl_94 vdd gnd cell_6t
Xbit_r95_c101 bl_101 br_101 wl_95 vdd gnd cell_6t
Xbit_r96_c101 bl_101 br_101 wl_96 vdd gnd cell_6t
Xbit_r97_c101 bl_101 br_101 wl_97 vdd gnd cell_6t
Xbit_r98_c101 bl_101 br_101 wl_98 vdd gnd cell_6t
Xbit_r99_c101 bl_101 br_101 wl_99 vdd gnd cell_6t
Xbit_r100_c101 bl_101 br_101 wl_100 vdd gnd cell_6t
Xbit_r101_c101 bl_101 br_101 wl_101 vdd gnd cell_6t
Xbit_r102_c101 bl_101 br_101 wl_102 vdd gnd cell_6t
Xbit_r103_c101 bl_101 br_101 wl_103 vdd gnd cell_6t
Xbit_r104_c101 bl_101 br_101 wl_104 vdd gnd cell_6t
Xbit_r105_c101 bl_101 br_101 wl_105 vdd gnd cell_6t
Xbit_r106_c101 bl_101 br_101 wl_106 vdd gnd cell_6t
Xbit_r107_c101 bl_101 br_101 wl_107 vdd gnd cell_6t
Xbit_r108_c101 bl_101 br_101 wl_108 vdd gnd cell_6t
Xbit_r109_c101 bl_101 br_101 wl_109 vdd gnd cell_6t
Xbit_r110_c101 bl_101 br_101 wl_110 vdd gnd cell_6t
Xbit_r111_c101 bl_101 br_101 wl_111 vdd gnd cell_6t
Xbit_r112_c101 bl_101 br_101 wl_112 vdd gnd cell_6t
Xbit_r113_c101 bl_101 br_101 wl_113 vdd gnd cell_6t
Xbit_r114_c101 bl_101 br_101 wl_114 vdd gnd cell_6t
Xbit_r115_c101 bl_101 br_101 wl_115 vdd gnd cell_6t
Xbit_r116_c101 bl_101 br_101 wl_116 vdd gnd cell_6t
Xbit_r117_c101 bl_101 br_101 wl_117 vdd gnd cell_6t
Xbit_r118_c101 bl_101 br_101 wl_118 vdd gnd cell_6t
Xbit_r119_c101 bl_101 br_101 wl_119 vdd gnd cell_6t
Xbit_r120_c101 bl_101 br_101 wl_120 vdd gnd cell_6t
Xbit_r121_c101 bl_101 br_101 wl_121 vdd gnd cell_6t
Xbit_r122_c101 bl_101 br_101 wl_122 vdd gnd cell_6t
Xbit_r123_c101 bl_101 br_101 wl_123 vdd gnd cell_6t
Xbit_r124_c101 bl_101 br_101 wl_124 vdd gnd cell_6t
Xbit_r125_c101 bl_101 br_101 wl_125 vdd gnd cell_6t
Xbit_r126_c101 bl_101 br_101 wl_126 vdd gnd cell_6t
Xbit_r127_c101 bl_101 br_101 wl_127 vdd gnd cell_6t
Xbit_r128_c101 bl_101 br_101 wl_128 vdd gnd cell_6t
Xbit_r129_c101 bl_101 br_101 wl_129 vdd gnd cell_6t
Xbit_r130_c101 bl_101 br_101 wl_130 vdd gnd cell_6t
Xbit_r131_c101 bl_101 br_101 wl_131 vdd gnd cell_6t
Xbit_r132_c101 bl_101 br_101 wl_132 vdd gnd cell_6t
Xbit_r133_c101 bl_101 br_101 wl_133 vdd gnd cell_6t
Xbit_r134_c101 bl_101 br_101 wl_134 vdd gnd cell_6t
Xbit_r135_c101 bl_101 br_101 wl_135 vdd gnd cell_6t
Xbit_r136_c101 bl_101 br_101 wl_136 vdd gnd cell_6t
Xbit_r137_c101 bl_101 br_101 wl_137 vdd gnd cell_6t
Xbit_r138_c101 bl_101 br_101 wl_138 vdd gnd cell_6t
Xbit_r139_c101 bl_101 br_101 wl_139 vdd gnd cell_6t
Xbit_r140_c101 bl_101 br_101 wl_140 vdd gnd cell_6t
Xbit_r141_c101 bl_101 br_101 wl_141 vdd gnd cell_6t
Xbit_r142_c101 bl_101 br_101 wl_142 vdd gnd cell_6t
Xbit_r143_c101 bl_101 br_101 wl_143 vdd gnd cell_6t
Xbit_r144_c101 bl_101 br_101 wl_144 vdd gnd cell_6t
Xbit_r145_c101 bl_101 br_101 wl_145 vdd gnd cell_6t
Xbit_r146_c101 bl_101 br_101 wl_146 vdd gnd cell_6t
Xbit_r147_c101 bl_101 br_101 wl_147 vdd gnd cell_6t
Xbit_r148_c101 bl_101 br_101 wl_148 vdd gnd cell_6t
Xbit_r149_c101 bl_101 br_101 wl_149 vdd gnd cell_6t
Xbit_r150_c101 bl_101 br_101 wl_150 vdd gnd cell_6t
Xbit_r151_c101 bl_101 br_101 wl_151 vdd gnd cell_6t
Xbit_r152_c101 bl_101 br_101 wl_152 vdd gnd cell_6t
Xbit_r153_c101 bl_101 br_101 wl_153 vdd gnd cell_6t
Xbit_r154_c101 bl_101 br_101 wl_154 vdd gnd cell_6t
Xbit_r155_c101 bl_101 br_101 wl_155 vdd gnd cell_6t
Xbit_r156_c101 bl_101 br_101 wl_156 vdd gnd cell_6t
Xbit_r157_c101 bl_101 br_101 wl_157 vdd gnd cell_6t
Xbit_r158_c101 bl_101 br_101 wl_158 vdd gnd cell_6t
Xbit_r159_c101 bl_101 br_101 wl_159 vdd gnd cell_6t
Xbit_r160_c101 bl_101 br_101 wl_160 vdd gnd cell_6t
Xbit_r161_c101 bl_101 br_101 wl_161 vdd gnd cell_6t
Xbit_r162_c101 bl_101 br_101 wl_162 vdd gnd cell_6t
Xbit_r163_c101 bl_101 br_101 wl_163 vdd gnd cell_6t
Xbit_r164_c101 bl_101 br_101 wl_164 vdd gnd cell_6t
Xbit_r165_c101 bl_101 br_101 wl_165 vdd gnd cell_6t
Xbit_r166_c101 bl_101 br_101 wl_166 vdd gnd cell_6t
Xbit_r167_c101 bl_101 br_101 wl_167 vdd gnd cell_6t
Xbit_r168_c101 bl_101 br_101 wl_168 vdd gnd cell_6t
Xbit_r169_c101 bl_101 br_101 wl_169 vdd gnd cell_6t
Xbit_r170_c101 bl_101 br_101 wl_170 vdd gnd cell_6t
Xbit_r171_c101 bl_101 br_101 wl_171 vdd gnd cell_6t
Xbit_r172_c101 bl_101 br_101 wl_172 vdd gnd cell_6t
Xbit_r173_c101 bl_101 br_101 wl_173 vdd gnd cell_6t
Xbit_r174_c101 bl_101 br_101 wl_174 vdd gnd cell_6t
Xbit_r175_c101 bl_101 br_101 wl_175 vdd gnd cell_6t
Xbit_r176_c101 bl_101 br_101 wl_176 vdd gnd cell_6t
Xbit_r177_c101 bl_101 br_101 wl_177 vdd gnd cell_6t
Xbit_r178_c101 bl_101 br_101 wl_178 vdd gnd cell_6t
Xbit_r179_c101 bl_101 br_101 wl_179 vdd gnd cell_6t
Xbit_r180_c101 bl_101 br_101 wl_180 vdd gnd cell_6t
Xbit_r181_c101 bl_101 br_101 wl_181 vdd gnd cell_6t
Xbit_r182_c101 bl_101 br_101 wl_182 vdd gnd cell_6t
Xbit_r183_c101 bl_101 br_101 wl_183 vdd gnd cell_6t
Xbit_r184_c101 bl_101 br_101 wl_184 vdd gnd cell_6t
Xbit_r185_c101 bl_101 br_101 wl_185 vdd gnd cell_6t
Xbit_r186_c101 bl_101 br_101 wl_186 vdd gnd cell_6t
Xbit_r187_c101 bl_101 br_101 wl_187 vdd gnd cell_6t
Xbit_r188_c101 bl_101 br_101 wl_188 vdd gnd cell_6t
Xbit_r189_c101 bl_101 br_101 wl_189 vdd gnd cell_6t
Xbit_r190_c101 bl_101 br_101 wl_190 vdd gnd cell_6t
Xbit_r191_c101 bl_101 br_101 wl_191 vdd gnd cell_6t
Xbit_r192_c101 bl_101 br_101 wl_192 vdd gnd cell_6t
Xbit_r193_c101 bl_101 br_101 wl_193 vdd gnd cell_6t
Xbit_r194_c101 bl_101 br_101 wl_194 vdd gnd cell_6t
Xbit_r195_c101 bl_101 br_101 wl_195 vdd gnd cell_6t
Xbit_r196_c101 bl_101 br_101 wl_196 vdd gnd cell_6t
Xbit_r197_c101 bl_101 br_101 wl_197 vdd gnd cell_6t
Xbit_r198_c101 bl_101 br_101 wl_198 vdd gnd cell_6t
Xbit_r199_c101 bl_101 br_101 wl_199 vdd gnd cell_6t
Xbit_r200_c101 bl_101 br_101 wl_200 vdd gnd cell_6t
Xbit_r201_c101 bl_101 br_101 wl_201 vdd gnd cell_6t
Xbit_r202_c101 bl_101 br_101 wl_202 vdd gnd cell_6t
Xbit_r203_c101 bl_101 br_101 wl_203 vdd gnd cell_6t
Xbit_r204_c101 bl_101 br_101 wl_204 vdd gnd cell_6t
Xbit_r205_c101 bl_101 br_101 wl_205 vdd gnd cell_6t
Xbit_r206_c101 bl_101 br_101 wl_206 vdd gnd cell_6t
Xbit_r207_c101 bl_101 br_101 wl_207 vdd gnd cell_6t
Xbit_r208_c101 bl_101 br_101 wl_208 vdd gnd cell_6t
Xbit_r209_c101 bl_101 br_101 wl_209 vdd gnd cell_6t
Xbit_r210_c101 bl_101 br_101 wl_210 vdd gnd cell_6t
Xbit_r211_c101 bl_101 br_101 wl_211 vdd gnd cell_6t
Xbit_r212_c101 bl_101 br_101 wl_212 vdd gnd cell_6t
Xbit_r213_c101 bl_101 br_101 wl_213 vdd gnd cell_6t
Xbit_r214_c101 bl_101 br_101 wl_214 vdd gnd cell_6t
Xbit_r215_c101 bl_101 br_101 wl_215 vdd gnd cell_6t
Xbit_r216_c101 bl_101 br_101 wl_216 vdd gnd cell_6t
Xbit_r217_c101 bl_101 br_101 wl_217 vdd gnd cell_6t
Xbit_r218_c101 bl_101 br_101 wl_218 vdd gnd cell_6t
Xbit_r219_c101 bl_101 br_101 wl_219 vdd gnd cell_6t
Xbit_r220_c101 bl_101 br_101 wl_220 vdd gnd cell_6t
Xbit_r221_c101 bl_101 br_101 wl_221 vdd gnd cell_6t
Xbit_r222_c101 bl_101 br_101 wl_222 vdd gnd cell_6t
Xbit_r223_c101 bl_101 br_101 wl_223 vdd gnd cell_6t
Xbit_r224_c101 bl_101 br_101 wl_224 vdd gnd cell_6t
Xbit_r225_c101 bl_101 br_101 wl_225 vdd gnd cell_6t
Xbit_r226_c101 bl_101 br_101 wl_226 vdd gnd cell_6t
Xbit_r227_c101 bl_101 br_101 wl_227 vdd gnd cell_6t
Xbit_r228_c101 bl_101 br_101 wl_228 vdd gnd cell_6t
Xbit_r229_c101 bl_101 br_101 wl_229 vdd gnd cell_6t
Xbit_r230_c101 bl_101 br_101 wl_230 vdd gnd cell_6t
Xbit_r231_c101 bl_101 br_101 wl_231 vdd gnd cell_6t
Xbit_r232_c101 bl_101 br_101 wl_232 vdd gnd cell_6t
Xbit_r233_c101 bl_101 br_101 wl_233 vdd gnd cell_6t
Xbit_r234_c101 bl_101 br_101 wl_234 vdd gnd cell_6t
Xbit_r235_c101 bl_101 br_101 wl_235 vdd gnd cell_6t
Xbit_r236_c101 bl_101 br_101 wl_236 vdd gnd cell_6t
Xbit_r237_c101 bl_101 br_101 wl_237 vdd gnd cell_6t
Xbit_r238_c101 bl_101 br_101 wl_238 vdd gnd cell_6t
Xbit_r239_c101 bl_101 br_101 wl_239 vdd gnd cell_6t
Xbit_r240_c101 bl_101 br_101 wl_240 vdd gnd cell_6t
Xbit_r241_c101 bl_101 br_101 wl_241 vdd gnd cell_6t
Xbit_r242_c101 bl_101 br_101 wl_242 vdd gnd cell_6t
Xbit_r243_c101 bl_101 br_101 wl_243 vdd gnd cell_6t
Xbit_r244_c101 bl_101 br_101 wl_244 vdd gnd cell_6t
Xbit_r245_c101 bl_101 br_101 wl_245 vdd gnd cell_6t
Xbit_r246_c101 bl_101 br_101 wl_246 vdd gnd cell_6t
Xbit_r247_c101 bl_101 br_101 wl_247 vdd gnd cell_6t
Xbit_r248_c101 bl_101 br_101 wl_248 vdd gnd cell_6t
Xbit_r249_c101 bl_101 br_101 wl_249 vdd gnd cell_6t
Xbit_r250_c101 bl_101 br_101 wl_250 vdd gnd cell_6t
Xbit_r251_c101 bl_101 br_101 wl_251 vdd gnd cell_6t
Xbit_r252_c101 bl_101 br_101 wl_252 vdd gnd cell_6t
Xbit_r253_c101 bl_101 br_101 wl_253 vdd gnd cell_6t
Xbit_r254_c101 bl_101 br_101 wl_254 vdd gnd cell_6t
Xbit_r255_c101 bl_101 br_101 wl_255 vdd gnd cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd cell_6t
Xbit_r1_c102 bl_102 br_102 wl_1 vdd gnd cell_6t
Xbit_r2_c102 bl_102 br_102 wl_2 vdd gnd cell_6t
Xbit_r3_c102 bl_102 br_102 wl_3 vdd gnd cell_6t
Xbit_r4_c102 bl_102 br_102 wl_4 vdd gnd cell_6t
Xbit_r5_c102 bl_102 br_102 wl_5 vdd gnd cell_6t
Xbit_r6_c102 bl_102 br_102 wl_6 vdd gnd cell_6t
Xbit_r7_c102 bl_102 br_102 wl_7 vdd gnd cell_6t
Xbit_r8_c102 bl_102 br_102 wl_8 vdd gnd cell_6t
Xbit_r9_c102 bl_102 br_102 wl_9 vdd gnd cell_6t
Xbit_r10_c102 bl_102 br_102 wl_10 vdd gnd cell_6t
Xbit_r11_c102 bl_102 br_102 wl_11 vdd gnd cell_6t
Xbit_r12_c102 bl_102 br_102 wl_12 vdd gnd cell_6t
Xbit_r13_c102 bl_102 br_102 wl_13 vdd gnd cell_6t
Xbit_r14_c102 bl_102 br_102 wl_14 vdd gnd cell_6t
Xbit_r15_c102 bl_102 br_102 wl_15 vdd gnd cell_6t
Xbit_r16_c102 bl_102 br_102 wl_16 vdd gnd cell_6t
Xbit_r17_c102 bl_102 br_102 wl_17 vdd gnd cell_6t
Xbit_r18_c102 bl_102 br_102 wl_18 vdd gnd cell_6t
Xbit_r19_c102 bl_102 br_102 wl_19 vdd gnd cell_6t
Xbit_r20_c102 bl_102 br_102 wl_20 vdd gnd cell_6t
Xbit_r21_c102 bl_102 br_102 wl_21 vdd gnd cell_6t
Xbit_r22_c102 bl_102 br_102 wl_22 vdd gnd cell_6t
Xbit_r23_c102 bl_102 br_102 wl_23 vdd gnd cell_6t
Xbit_r24_c102 bl_102 br_102 wl_24 vdd gnd cell_6t
Xbit_r25_c102 bl_102 br_102 wl_25 vdd gnd cell_6t
Xbit_r26_c102 bl_102 br_102 wl_26 vdd gnd cell_6t
Xbit_r27_c102 bl_102 br_102 wl_27 vdd gnd cell_6t
Xbit_r28_c102 bl_102 br_102 wl_28 vdd gnd cell_6t
Xbit_r29_c102 bl_102 br_102 wl_29 vdd gnd cell_6t
Xbit_r30_c102 bl_102 br_102 wl_30 vdd gnd cell_6t
Xbit_r31_c102 bl_102 br_102 wl_31 vdd gnd cell_6t
Xbit_r32_c102 bl_102 br_102 wl_32 vdd gnd cell_6t
Xbit_r33_c102 bl_102 br_102 wl_33 vdd gnd cell_6t
Xbit_r34_c102 bl_102 br_102 wl_34 vdd gnd cell_6t
Xbit_r35_c102 bl_102 br_102 wl_35 vdd gnd cell_6t
Xbit_r36_c102 bl_102 br_102 wl_36 vdd gnd cell_6t
Xbit_r37_c102 bl_102 br_102 wl_37 vdd gnd cell_6t
Xbit_r38_c102 bl_102 br_102 wl_38 vdd gnd cell_6t
Xbit_r39_c102 bl_102 br_102 wl_39 vdd gnd cell_6t
Xbit_r40_c102 bl_102 br_102 wl_40 vdd gnd cell_6t
Xbit_r41_c102 bl_102 br_102 wl_41 vdd gnd cell_6t
Xbit_r42_c102 bl_102 br_102 wl_42 vdd gnd cell_6t
Xbit_r43_c102 bl_102 br_102 wl_43 vdd gnd cell_6t
Xbit_r44_c102 bl_102 br_102 wl_44 vdd gnd cell_6t
Xbit_r45_c102 bl_102 br_102 wl_45 vdd gnd cell_6t
Xbit_r46_c102 bl_102 br_102 wl_46 vdd gnd cell_6t
Xbit_r47_c102 bl_102 br_102 wl_47 vdd gnd cell_6t
Xbit_r48_c102 bl_102 br_102 wl_48 vdd gnd cell_6t
Xbit_r49_c102 bl_102 br_102 wl_49 vdd gnd cell_6t
Xbit_r50_c102 bl_102 br_102 wl_50 vdd gnd cell_6t
Xbit_r51_c102 bl_102 br_102 wl_51 vdd gnd cell_6t
Xbit_r52_c102 bl_102 br_102 wl_52 vdd gnd cell_6t
Xbit_r53_c102 bl_102 br_102 wl_53 vdd gnd cell_6t
Xbit_r54_c102 bl_102 br_102 wl_54 vdd gnd cell_6t
Xbit_r55_c102 bl_102 br_102 wl_55 vdd gnd cell_6t
Xbit_r56_c102 bl_102 br_102 wl_56 vdd gnd cell_6t
Xbit_r57_c102 bl_102 br_102 wl_57 vdd gnd cell_6t
Xbit_r58_c102 bl_102 br_102 wl_58 vdd gnd cell_6t
Xbit_r59_c102 bl_102 br_102 wl_59 vdd gnd cell_6t
Xbit_r60_c102 bl_102 br_102 wl_60 vdd gnd cell_6t
Xbit_r61_c102 bl_102 br_102 wl_61 vdd gnd cell_6t
Xbit_r62_c102 bl_102 br_102 wl_62 vdd gnd cell_6t
Xbit_r63_c102 bl_102 br_102 wl_63 vdd gnd cell_6t
Xbit_r64_c102 bl_102 br_102 wl_64 vdd gnd cell_6t
Xbit_r65_c102 bl_102 br_102 wl_65 vdd gnd cell_6t
Xbit_r66_c102 bl_102 br_102 wl_66 vdd gnd cell_6t
Xbit_r67_c102 bl_102 br_102 wl_67 vdd gnd cell_6t
Xbit_r68_c102 bl_102 br_102 wl_68 vdd gnd cell_6t
Xbit_r69_c102 bl_102 br_102 wl_69 vdd gnd cell_6t
Xbit_r70_c102 bl_102 br_102 wl_70 vdd gnd cell_6t
Xbit_r71_c102 bl_102 br_102 wl_71 vdd gnd cell_6t
Xbit_r72_c102 bl_102 br_102 wl_72 vdd gnd cell_6t
Xbit_r73_c102 bl_102 br_102 wl_73 vdd gnd cell_6t
Xbit_r74_c102 bl_102 br_102 wl_74 vdd gnd cell_6t
Xbit_r75_c102 bl_102 br_102 wl_75 vdd gnd cell_6t
Xbit_r76_c102 bl_102 br_102 wl_76 vdd gnd cell_6t
Xbit_r77_c102 bl_102 br_102 wl_77 vdd gnd cell_6t
Xbit_r78_c102 bl_102 br_102 wl_78 vdd gnd cell_6t
Xbit_r79_c102 bl_102 br_102 wl_79 vdd gnd cell_6t
Xbit_r80_c102 bl_102 br_102 wl_80 vdd gnd cell_6t
Xbit_r81_c102 bl_102 br_102 wl_81 vdd gnd cell_6t
Xbit_r82_c102 bl_102 br_102 wl_82 vdd gnd cell_6t
Xbit_r83_c102 bl_102 br_102 wl_83 vdd gnd cell_6t
Xbit_r84_c102 bl_102 br_102 wl_84 vdd gnd cell_6t
Xbit_r85_c102 bl_102 br_102 wl_85 vdd gnd cell_6t
Xbit_r86_c102 bl_102 br_102 wl_86 vdd gnd cell_6t
Xbit_r87_c102 bl_102 br_102 wl_87 vdd gnd cell_6t
Xbit_r88_c102 bl_102 br_102 wl_88 vdd gnd cell_6t
Xbit_r89_c102 bl_102 br_102 wl_89 vdd gnd cell_6t
Xbit_r90_c102 bl_102 br_102 wl_90 vdd gnd cell_6t
Xbit_r91_c102 bl_102 br_102 wl_91 vdd gnd cell_6t
Xbit_r92_c102 bl_102 br_102 wl_92 vdd gnd cell_6t
Xbit_r93_c102 bl_102 br_102 wl_93 vdd gnd cell_6t
Xbit_r94_c102 bl_102 br_102 wl_94 vdd gnd cell_6t
Xbit_r95_c102 bl_102 br_102 wl_95 vdd gnd cell_6t
Xbit_r96_c102 bl_102 br_102 wl_96 vdd gnd cell_6t
Xbit_r97_c102 bl_102 br_102 wl_97 vdd gnd cell_6t
Xbit_r98_c102 bl_102 br_102 wl_98 vdd gnd cell_6t
Xbit_r99_c102 bl_102 br_102 wl_99 vdd gnd cell_6t
Xbit_r100_c102 bl_102 br_102 wl_100 vdd gnd cell_6t
Xbit_r101_c102 bl_102 br_102 wl_101 vdd gnd cell_6t
Xbit_r102_c102 bl_102 br_102 wl_102 vdd gnd cell_6t
Xbit_r103_c102 bl_102 br_102 wl_103 vdd gnd cell_6t
Xbit_r104_c102 bl_102 br_102 wl_104 vdd gnd cell_6t
Xbit_r105_c102 bl_102 br_102 wl_105 vdd gnd cell_6t
Xbit_r106_c102 bl_102 br_102 wl_106 vdd gnd cell_6t
Xbit_r107_c102 bl_102 br_102 wl_107 vdd gnd cell_6t
Xbit_r108_c102 bl_102 br_102 wl_108 vdd gnd cell_6t
Xbit_r109_c102 bl_102 br_102 wl_109 vdd gnd cell_6t
Xbit_r110_c102 bl_102 br_102 wl_110 vdd gnd cell_6t
Xbit_r111_c102 bl_102 br_102 wl_111 vdd gnd cell_6t
Xbit_r112_c102 bl_102 br_102 wl_112 vdd gnd cell_6t
Xbit_r113_c102 bl_102 br_102 wl_113 vdd gnd cell_6t
Xbit_r114_c102 bl_102 br_102 wl_114 vdd gnd cell_6t
Xbit_r115_c102 bl_102 br_102 wl_115 vdd gnd cell_6t
Xbit_r116_c102 bl_102 br_102 wl_116 vdd gnd cell_6t
Xbit_r117_c102 bl_102 br_102 wl_117 vdd gnd cell_6t
Xbit_r118_c102 bl_102 br_102 wl_118 vdd gnd cell_6t
Xbit_r119_c102 bl_102 br_102 wl_119 vdd gnd cell_6t
Xbit_r120_c102 bl_102 br_102 wl_120 vdd gnd cell_6t
Xbit_r121_c102 bl_102 br_102 wl_121 vdd gnd cell_6t
Xbit_r122_c102 bl_102 br_102 wl_122 vdd gnd cell_6t
Xbit_r123_c102 bl_102 br_102 wl_123 vdd gnd cell_6t
Xbit_r124_c102 bl_102 br_102 wl_124 vdd gnd cell_6t
Xbit_r125_c102 bl_102 br_102 wl_125 vdd gnd cell_6t
Xbit_r126_c102 bl_102 br_102 wl_126 vdd gnd cell_6t
Xbit_r127_c102 bl_102 br_102 wl_127 vdd gnd cell_6t
Xbit_r128_c102 bl_102 br_102 wl_128 vdd gnd cell_6t
Xbit_r129_c102 bl_102 br_102 wl_129 vdd gnd cell_6t
Xbit_r130_c102 bl_102 br_102 wl_130 vdd gnd cell_6t
Xbit_r131_c102 bl_102 br_102 wl_131 vdd gnd cell_6t
Xbit_r132_c102 bl_102 br_102 wl_132 vdd gnd cell_6t
Xbit_r133_c102 bl_102 br_102 wl_133 vdd gnd cell_6t
Xbit_r134_c102 bl_102 br_102 wl_134 vdd gnd cell_6t
Xbit_r135_c102 bl_102 br_102 wl_135 vdd gnd cell_6t
Xbit_r136_c102 bl_102 br_102 wl_136 vdd gnd cell_6t
Xbit_r137_c102 bl_102 br_102 wl_137 vdd gnd cell_6t
Xbit_r138_c102 bl_102 br_102 wl_138 vdd gnd cell_6t
Xbit_r139_c102 bl_102 br_102 wl_139 vdd gnd cell_6t
Xbit_r140_c102 bl_102 br_102 wl_140 vdd gnd cell_6t
Xbit_r141_c102 bl_102 br_102 wl_141 vdd gnd cell_6t
Xbit_r142_c102 bl_102 br_102 wl_142 vdd gnd cell_6t
Xbit_r143_c102 bl_102 br_102 wl_143 vdd gnd cell_6t
Xbit_r144_c102 bl_102 br_102 wl_144 vdd gnd cell_6t
Xbit_r145_c102 bl_102 br_102 wl_145 vdd gnd cell_6t
Xbit_r146_c102 bl_102 br_102 wl_146 vdd gnd cell_6t
Xbit_r147_c102 bl_102 br_102 wl_147 vdd gnd cell_6t
Xbit_r148_c102 bl_102 br_102 wl_148 vdd gnd cell_6t
Xbit_r149_c102 bl_102 br_102 wl_149 vdd gnd cell_6t
Xbit_r150_c102 bl_102 br_102 wl_150 vdd gnd cell_6t
Xbit_r151_c102 bl_102 br_102 wl_151 vdd gnd cell_6t
Xbit_r152_c102 bl_102 br_102 wl_152 vdd gnd cell_6t
Xbit_r153_c102 bl_102 br_102 wl_153 vdd gnd cell_6t
Xbit_r154_c102 bl_102 br_102 wl_154 vdd gnd cell_6t
Xbit_r155_c102 bl_102 br_102 wl_155 vdd gnd cell_6t
Xbit_r156_c102 bl_102 br_102 wl_156 vdd gnd cell_6t
Xbit_r157_c102 bl_102 br_102 wl_157 vdd gnd cell_6t
Xbit_r158_c102 bl_102 br_102 wl_158 vdd gnd cell_6t
Xbit_r159_c102 bl_102 br_102 wl_159 vdd gnd cell_6t
Xbit_r160_c102 bl_102 br_102 wl_160 vdd gnd cell_6t
Xbit_r161_c102 bl_102 br_102 wl_161 vdd gnd cell_6t
Xbit_r162_c102 bl_102 br_102 wl_162 vdd gnd cell_6t
Xbit_r163_c102 bl_102 br_102 wl_163 vdd gnd cell_6t
Xbit_r164_c102 bl_102 br_102 wl_164 vdd gnd cell_6t
Xbit_r165_c102 bl_102 br_102 wl_165 vdd gnd cell_6t
Xbit_r166_c102 bl_102 br_102 wl_166 vdd gnd cell_6t
Xbit_r167_c102 bl_102 br_102 wl_167 vdd gnd cell_6t
Xbit_r168_c102 bl_102 br_102 wl_168 vdd gnd cell_6t
Xbit_r169_c102 bl_102 br_102 wl_169 vdd gnd cell_6t
Xbit_r170_c102 bl_102 br_102 wl_170 vdd gnd cell_6t
Xbit_r171_c102 bl_102 br_102 wl_171 vdd gnd cell_6t
Xbit_r172_c102 bl_102 br_102 wl_172 vdd gnd cell_6t
Xbit_r173_c102 bl_102 br_102 wl_173 vdd gnd cell_6t
Xbit_r174_c102 bl_102 br_102 wl_174 vdd gnd cell_6t
Xbit_r175_c102 bl_102 br_102 wl_175 vdd gnd cell_6t
Xbit_r176_c102 bl_102 br_102 wl_176 vdd gnd cell_6t
Xbit_r177_c102 bl_102 br_102 wl_177 vdd gnd cell_6t
Xbit_r178_c102 bl_102 br_102 wl_178 vdd gnd cell_6t
Xbit_r179_c102 bl_102 br_102 wl_179 vdd gnd cell_6t
Xbit_r180_c102 bl_102 br_102 wl_180 vdd gnd cell_6t
Xbit_r181_c102 bl_102 br_102 wl_181 vdd gnd cell_6t
Xbit_r182_c102 bl_102 br_102 wl_182 vdd gnd cell_6t
Xbit_r183_c102 bl_102 br_102 wl_183 vdd gnd cell_6t
Xbit_r184_c102 bl_102 br_102 wl_184 vdd gnd cell_6t
Xbit_r185_c102 bl_102 br_102 wl_185 vdd gnd cell_6t
Xbit_r186_c102 bl_102 br_102 wl_186 vdd gnd cell_6t
Xbit_r187_c102 bl_102 br_102 wl_187 vdd gnd cell_6t
Xbit_r188_c102 bl_102 br_102 wl_188 vdd gnd cell_6t
Xbit_r189_c102 bl_102 br_102 wl_189 vdd gnd cell_6t
Xbit_r190_c102 bl_102 br_102 wl_190 vdd gnd cell_6t
Xbit_r191_c102 bl_102 br_102 wl_191 vdd gnd cell_6t
Xbit_r192_c102 bl_102 br_102 wl_192 vdd gnd cell_6t
Xbit_r193_c102 bl_102 br_102 wl_193 vdd gnd cell_6t
Xbit_r194_c102 bl_102 br_102 wl_194 vdd gnd cell_6t
Xbit_r195_c102 bl_102 br_102 wl_195 vdd gnd cell_6t
Xbit_r196_c102 bl_102 br_102 wl_196 vdd gnd cell_6t
Xbit_r197_c102 bl_102 br_102 wl_197 vdd gnd cell_6t
Xbit_r198_c102 bl_102 br_102 wl_198 vdd gnd cell_6t
Xbit_r199_c102 bl_102 br_102 wl_199 vdd gnd cell_6t
Xbit_r200_c102 bl_102 br_102 wl_200 vdd gnd cell_6t
Xbit_r201_c102 bl_102 br_102 wl_201 vdd gnd cell_6t
Xbit_r202_c102 bl_102 br_102 wl_202 vdd gnd cell_6t
Xbit_r203_c102 bl_102 br_102 wl_203 vdd gnd cell_6t
Xbit_r204_c102 bl_102 br_102 wl_204 vdd gnd cell_6t
Xbit_r205_c102 bl_102 br_102 wl_205 vdd gnd cell_6t
Xbit_r206_c102 bl_102 br_102 wl_206 vdd gnd cell_6t
Xbit_r207_c102 bl_102 br_102 wl_207 vdd gnd cell_6t
Xbit_r208_c102 bl_102 br_102 wl_208 vdd gnd cell_6t
Xbit_r209_c102 bl_102 br_102 wl_209 vdd gnd cell_6t
Xbit_r210_c102 bl_102 br_102 wl_210 vdd gnd cell_6t
Xbit_r211_c102 bl_102 br_102 wl_211 vdd gnd cell_6t
Xbit_r212_c102 bl_102 br_102 wl_212 vdd gnd cell_6t
Xbit_r213_c102 bl_102 br_102 wl_213 vdd gnd cell_6t
Xbit_r214_c102 bl_102 br_102 wl_214 vdd gnd cell_6t
Xbit_r215_c102 bl_102 br_102 wl_215 vdd gnd cell_6t
Xbit_r216_c102 bl_102 br_102 wl_216 vdd gnd cell_6t
Xbit_r217_c102 bl_102 br_102 wl_217 vdd gnd cell_6t
Xbit_r218_c102 bl_102 br_102 wl_218 vdd gnd cell_6t
Xbit_r219_c102 bl_102 br_102 wl_219 vdd gnd cell_6t
Xbit_r220_c102 bl_102 br_102 wl_220 vdd gnd cell_6t
Xbit_r221_c102 bl_102 br_102 wl_221 vdd gnd cell_6t
Xbit_r222_c102 bl_102 br_102 wl_222 vdd gnd cell_6t
Xbit_r223_c102 bl_102 br_102 wl_223 vdd gnd cell_6t
Xbit_r224_c102 bl_102 br_102 wl_224 vdd gnd cell_6t
Xbit_r225_c102 bl_102 br_102 wl_225 vdd gnd cell_6t
Xbit_r226_c102 bl_102 br_102 wl_226 vdd gnd cell_6t
Xbit_r227_c102 bl_102 br_102 wl_227 vdd gnd cell_6t
Xbit_r228_c102 bl_102 br_102 wl_228 vdd gnd cell_6t
Xbit_r229_c102 bl_102 br_102 wl_229 vdd gnd cell_6t
Xbit_r230_c102 bl_102 br_102 wl_230 vdd gnd cell_6t
Xbit_r231_c102 bl_102 br_102 wl_231 vdd gnd cell_6t
Xbit_r232_c102 bl_102 br_102 wl_232 vdd gnd cell_6t
Xbit_r233_c102 bl_102 br_102 wl_233 vdd gnd cell_6t
Xbit_r234_c102 bl_102 br_102 wl_234 vdd gnd cell_6t
Xbit_r235_c102 bl_102 br_102 wl_235 vdd gnd cell_6t
Xbit_r236_c102 bl_102 br_102 wl_236 vdd gnd cell_6t
Xbit_r237_c102 bl_102 br_102 wl_237 vdd gnd cell_6t
Xbit_r238_c102 bl_102 br_102 wl_238 vdd gnd cell_6t
Xbit_r239_c102 bl_102 br_102 wl_239 vdd gnd cell_6t
Xbit_r240_c102 bl_102 br_102 wl_240 vdd gnd cell_6t
Xbit_r241_c102 bl_102 br_102 wl_241 vdd gnd cell_6t
Xbit_r242_c102 bl_102 br_102 wl_242 vdd gnd cell_6t
Xbit_r243_c102 bl_102 br_102 wl_243 vdd gnd cell_6t
Xbit_r244_c102 bl_102 br_102 wl_244 vdd gnd cell_6t
Xbit_r245_c102 bl_102 br_102 wl_245 vdd gnd cell_6t
Xbit_r246_c102 bl_102 br_102 wl_246 vdd gnd cell_6t
Xbit_r247_c102 bl_102 br_102 wl_247 vdd gnd cell_6t
Xbit_r248_c102 bl_102 br_102 wl_248 vdd gnd cell_6t
Xbit_r249_c102 bl_102 br_102 wl_249 vdd gnd cell_6t
Xbit_r250_c102 bl_102 br_102 wl_250 vdd gnd cell_6t
Xbit_r251_c102 bl_102 br_102 wl_251 vdd gnd cell_6t
Xbit_r252_c102 bl_102 br_102 wl_252 vdd gnd cell_6t
Xbit_r253_c102 bl_102 br_102 wl_253 vdd gnd cell_6t
Xbit_r254_c102 bl_102 br_102 wl_254 vdd gnd cell_6t
Xbit_r255_c102 bl_102 br_102 wl_255 vdd gnd cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd cell_6t
Xbit_r1_c103 bl_103 br_103 wl_1 vdd gnd cell_6t
Xbit_r2_c103 bl_103 br_103 wl_2 vdd gnd cell_6t
Xbit_r3_c103 bl_103 br_103 wl_3 vdd gnd cell_6t
Xbit_r4_c103 bl_103 br_103 wl_4 vdd gnd cell_6t
Xbit_r5_c103 bl_103 br_103 wl_5 vdd gnd cell_6t
Xbit_r6_c103 bl_103 br_103 wl_6 vdd gnd cell_6t
Xbit_r7_c103 bl_103 br_103 wl_7 vdd gnd cell_6t
Xbit_r8_c103 bl_103 br_103 wl_8 vdd gnd cell_6t
Xbit_r9_c103 bl_103 br_103 wl_9 vdd gnd cell_6t
Xbit_r10_c103 bl_103 br_103 wl_10 vdd gnd cell_6t
Xbit_r11_c103 bl_103 br_103 wl_11 vdd gnd cell_6t
Xbit_r12_c103 bl_103 br_103 wl_12 vdd gnd cell_6t
Xbit_r13_c103 bl_103 br_103 wl_13 vdd gnd cell_6t
Xbit_r14_c103 bl_103 br_103 wl_14 vdd gnd cell_6t
Xbit_r15_c103 bl_103 br_103 wl_15 vdd gnd cell_6t
Xbit_r16_c103 bl_103 br_103 wl_16 vdd gnd cell_6t
Xbit_r17_c103 bl_103 br_103 wl_17 vdd gnd cell_6t
Xbit_r18_c103 bl_103 br_103 wl_18 vdd gnd cell_6t
Xbit_r19_c103 bl_103 br_103 wl_19 vdd gnd cell_6t
Xbit_r20_c103 bl_103 br_103 wl_20 vdd gnd cell_6t
Xbit_r21_c103 bl_103 br_103 wl_21 vdd gnd cell_6t
Xbit_r22_c103 bl_103 br_103 wl_22 vdd gnd cell_6t
Xbit_r23_c103 bl_103 br_103 wl_23 vdd gnd cell_6t
Xbit_r24_c103 bl_103 br_103 wl_24 vdd gnd cell_6t
Xbit_r25_c103 bl_103 br_103 wl_25 vdd gnd cell_6t
Xbit_r26_c103 bl_103 br_103 wl_26 vdd gnd cell_6t
Xbit_r27_c103 bl_103 br_103 wl_27 vdd gnd cell_6t
Xbit_r28_c103 bl_103 br_103 wl_28 vdd gnd cell_6t
Xbit_r29_c103 bl_103 br_103 wl_29 vdd gnd cell_6t
Xbit_r30_c103 bl_103 br_103 wl_30 vdd gnd cell_6t
Xbit_r31_c103 bl_103 br_103 wl_31 vdd gnd cell_6t
Xbit_r32_c103 bl_103 br_103 wl_32 vdd gnd cell_6t
Xbit_r33_c103 bl_103 br_103 wl_33 vdd gnd cell_6t
Xbit_r34_c103 bl_103 br_103 wl_34 vdd gnd cell_6t
Xbit_r35_c103 bl_103 br_103 wl_35 vdd gnd cell_6t
Xbit_r36_c103 bl_103 br_103 wl_36 vdd gnd cell_6t
Xbit_r37_c103 bl_103 br_103 wl_37 vdd gnd cell_6t
Xbit_r38_c103 bl_103 br_103 wl_38 vdd gnd cell_6t
Xbit_r39_c103 bl_103 br_103 wl_39 vdd gnd cell_6t
Xbit_r40_c103 bl_103 br_103 wl_40 vdd gnd cell_6t
Xbit_r41_c103 bl_103 br_103 wl_41 vdd gnd cell_6t
Xbit_r42_c103 bl_103 br_103 wl_42 vdd gnd cell_6t
Xbit_r43_c103 bl_103 br_103 wl_43 vdd gnd cell_6t
Xbit_r44_c103 bl_103 br_103 wl_44 vdd gnd cell_6t
Xbit_r45_c103 bl_103 br_103 wl_45 vdd gnd cell_6t
Xbit_r46_c103 bl_103 br_103 wl_46 vdd gnd cell_6t
Xbit_r47_c103 bl_103 br_103 wl_47 vdd gnd cell_6t
Xbit_r48_c103 bl_103 br_103 wl_48 vdd gnd cell_6t
Xbit_r49_c103 bl_103 br_103 wl_49 vdd gnd cell_6t
Xbit_r50_c103 bl_103 br_103 wl_50 vdd gnd cell_6t
Xbit_r51_c103 bl_103 br_103 wl_51 vdd gnd cell_6t
Xbit_r52_c103 bl_103 br_103 wl_52 vdd gnd cell_6t
Xbit_r53_c103 bl_103 br_103 wl_53 vdd gnd cell_6t
Xbit_r54_c103 bl_103 br_103 wl_54 vdd gnd cell_6t
Xbit_r55_c103 bl_103 br_103 wl_55 vdd gnd cell_6t
Xbit_r56_c103 bl_103 br_103 wl_56 vdd gnd cell_6t
Xbit_r57_c103 bl_103 br_103 wl_57 vdd gnd cell_6t
Xbit_r58_c103 bl_103 br_103 wl_58 vdd gnd cell_6t
Xbit_r59_c103 bl_103 br_103 wl_59 vdd gnd cell_6t
Xbit_r60_c103 bl_103 br_103 wl_60 vdd gnd cell_6t
Xbit_r61_c103 bl_103 br_103 wl_61 vdd gnd cell_6t
Xbit_r62_c103 bl_103 br_103 wl_62 vdd gnd cell_6t
Xbit_r63_c103 bl_103 br_103 wl_63 vdd gnd cell_6t
Xbit_r64_c103 bl_103 br_103 wl_64 vdd gnd cell_6t
Xbit_r65_c103 bl_103 br_103 wl_65 vdd gnd cell_6t
Xbit_r66_c103 bl_103 br_103 wl_66 vdd gnd cell_6t
Xbit_r67_c103 bl_103 br_103 wl_67 vdd gnd cell_6t
Xbit_r68_c103 bl_103 br_103 wl_68 vdd gnd cell_6t
Xbit_r69_c103 bl_103 br_103 wl_69 vdd gnd cell_6t
Xbit_r70_c103 bl_103 br_103 wl_70 vdd gnd cell_6t
Xbit_r71_c103 bl_103 br_103 wl_71 vdd gnd cell_6t
Xbit_r72_c103 bl_103 br_103 wl_72 vdd gnd cell_6t
Xbit_r73_c103 bl_103 br_103 wl_73 vdd gnd cell_6t
Xbit_r74_c103 bl_103 br_103 wl_74 vdd gnd cell_6t
Xbit_r75_c103 bl_103 br_103 wl_75 vdd gnd cell_6t
Xbit_r76_c103 bl_103 br_103 wl_76 vdd gnd cell_6t
Xbit_r77_c103 bl_103 br_103 wl_77 vdd gnd cell_6t
Xbit_r78_c103 bl_103 br_103 wl_78 vdd gnd cell_6t
Xbit_r79_c103 bl_103 br_103 wl_79 vdd gnd cell_6t
Xbit_r80_c103 bl_103 br_103 wl_80 vdd gnd cell_6t
Xbit_r81_c103 bl_103 br_103 wl_81 vdd gnd cell_6t
Xbit_r82_c103 bl_103 br_103 wl_82 vdd gnd cell_6t
Xbit_r83_c103 bl_103 br_103 wl_83 vdd gnd cell_6t
Xbit_r84_c103 bl_103 br_103 wl_84 vdd gnd cell_6t
Xbit_r85_c103 bl_103 br_103 wl_85 vdd gnd cell_6t
Xbit_r86_c103 bl_103 br_103 wl_86 vdd gnd cell_6t
Xbit_r87_c103 bl_103 br_103 wl_87 vdd gnd cell_6t
Xbit_r88_c103 bl_103 br_103 wl_88 vdd gnd cell_6t
Xbit_r89_c103 bl_103 br_103 wl_89 vdd gnd cell_6t
Xbit_r90_c103 bl_103 br_103 wl_90 vdd gnd cell_6t
Xbit_r91_c103 bl_103 br_103 wl_91 vdd gnd cell_6t
Xbit_r92_c103 bl_103 br_103 wl_92 vdd gnd cell_6t
Xbit_r93_c103 bl_103 br_103 wl_93 vdd gnd cell_6t
Xbit_r94_c103 bl_103 br_103 wl_94 vdd gnd cell_6t
Xbit_r95_c103 bl_103 br_103 wl_95 vdd gnd cell_6t
Xbit_r96_c103 bl_103 br_103 wl_96 vdd gnd cell_6t
Xbit_r97_c103 bl_103 br_103 wl_97 vdd gnd cell_6t
Xbit_r98_c103 bl_103 br_103 wl_98 vdd gnd cell_6t
Xbit_r99_c103 bl_103 br_103 wl_99 vdd gnd cell_6t
Xbit_r100_c103 bl_103 br_103 wl_100 vdd gnd cell_6t
Xbit_r101_c103 bl_103 br_103 wl_101 vdd gnd cell_6t
Xbit_r102_c103 bl_103 br_103 wl_102 vdd gnd cell_6t
Xbit_r103_c103 bl_103 br_103 wl_103 vdd gnd cell_6t
Xbit_r104_c103 bl_103 br_103 wl_104 vdd gnd cell_6t
Xbit_r105_c103 bl_103 br_103 wl_105 vdd gnd cell_6t
Xbit_r106_c103 bl_103 br_103 wl_106 vdd gnd cell_6t
Xbit_r107_c103 bl_103 br_103 wl_107 vdd gnd cell_6t
Xbit_r108_c103 bl_103 br_103 wl_108 vdd gnd cell_6t
Xbit_r109_c103 bl_103 br_103 wl_109 vdd gnd cell_6t
Xbit_r110_c103 bl_103 br_103 wl_110 vdd gnd cell_6t
Xbit_r111_c103 bl_103 br_103 wl_111 vdd gnd cell_6t
Xbit_r112_c103 bl_103 br_103 wl_112 vdd gnd cell_6t
Xbit_r113_c103 bl_103 br_103 wl_113 vdd gnd cell_6t
Xbit_r114_c103 bl_103 br_103 wl_114 vdd gnd cell_6t
Xbit_r115_c103 bl_103 br_103 wl_115 vdd gnd cell_6t
Xbit_r116_c103 bl_103 br_103 wl_116 vdd gnd cell_6t
Xbit_r117_c103 bl_103 br_103 wl_117 vdd gnd cell_6t
Xbit_r118_c103 bl_103 br_103 wl_118 vdd gnd cell_6t
Xbit_r119_c103 bl_103 br_103 wl_119 vdd gnd cell_6t
Xbit_r120_c103 bl_103 br_103 wl_120 vdd gnd cell_6t
Xbit_r121_c103 bl_103 br_103 wl_121 vdd gnd cell_6t
Xbit_r122_c103 bl_103 br_103 wl_122 vdd gnd cell_6t
Xbit_r123_c103 bl_103 br_103 wl_123 vdd gnd cell_6t
Xbit_r124_c103 bl_103 br_103 wl_124 vdd gnd cell_6t
Xbit_r125_c103 bl_103 br_103 wl_125 vdd gnd cell_6t
Xbit_r126_c103 bl_103 br_103 wl_126 vdd gnd cell_6t
Xbit_r127_c103 bl_103 br_103 wl_127 vdd gnd cell_6t
Xbit_r128_c103 bl_103 br_103 wl_128 vdd gnd cell_6t
Xbit_r129_c103 bl_103 br_103 wl_129 vdd gnd cell_6t
Xbit_r130_c103 bl_103 br_103 wl_130 vdd gnd cell_6t
Xbit_r131_c103 bl_103 br_103 wl_131 vdd gnd cell_6t
Xbit_r132_c103 bl_103 br_103 wl_132 vdd gnd cell_6t
Xbit_r133_c103 bl_103 br_103 wl_133 vdd gnd cell_6t
Xbit_r134_c103 bl_103 br_103 wl_134 vdd gnd cell_6t
Xbit_r135_c103 bl_103 br_103 wl_135 vdd gnd cell_6t
Xbit_r136_c103 bl_103 br_103 wl_136 vdd gnd cell_6t
Xbit_r137_c103 bl_103 br_103 wl_137 vdd gnd cell_6t
Xbit_r138_c103 bl_103 br_103 wl_138 vdd gnd cell_6t
Xbit_r139_c103 bl_103 br_103 wl_139 vdd gnd cell_6t
Xbit_r140_c103 bl_103 br_103 wl_140 vdd gnd cell_6t
Xbit_r141_c103 bl_103 br_103 wl_141 vdd gnd cell_6t
Xbit_r142_c103 bl_103 br_103 wl_142 vdd gnd cell_6t
Xbit_r143_c103 bl_103 br_103 wl_143 vdd gnd cell_6t
Xbit_r144_c103 bl_103 br_103 wl_144 vdd gnd cell_6t
Xbit_r145_c103 bl_103 br_103 wl_145 vdd gnd cell_6t
Xbit_r146_c103 bl_103 br_103 wl_146 vdd gnd cell_6t
Xbit_r147_c103 bl_103 br_103 wl_147 vdd gnd cell_6t
Xbit_r148_c103 bl_103 br_103 wl_148 vdd gnd cell_6t
Xbit_r149_c103 bl_103 br_103 wl_149 vdd gnd cell_6t
Xbit_r150_c103 bl_103 br_103 wl_150 vdd gnd cell_6t
Xbit_r151_c103 bl_103 br_103 wl_151 vdd gnd cell_6t
Xbit_r152_c103 bl_103 br_103 wl_152 vdd gnd cell_6t
Xbit_r153_c103 bl_103 br_103 wl_153 vdd gnd cell_6t
Xbit_r154_c103 bl_103 br_103 wl_154 vdd gnd cell_6t
Xbit_r155_c103 bl_103 br_103 wl_155 vdd gnd cell_6t
Xbit_r156_c103 bl_103 br_103 wl_156 vdd gnd cell_6t
Xbit_r157_c103 bl_103 br_103 wl_157 vdd gnd cell_6t
Xbit_r158_c103 bl_103 br_103 wl_158 vdd gnd cell_6t
Xbit_r159_c103 bl_103 br_103 wl_159 vdd gnd cell_6t
Xbit_r160_c103 bl_103 br_103 wl_160 vdd gnd cell_6t
Xbit_r161_c103 bl_103 br_103 wl_161 vdd gnd cell_6t
Xbit_r162_c103 bl_103 br_103 wl_162 vdd gnd cell_6t
Xbit_r163_c103 bl_103 br_103 wl_163 vdd gnd cell_6t
Xbit_r164_c103 bl_103 br_103 wl_164 vdd gnd cell_6t
Xbit_r165_c103 bl_103 br_103 wl_165 vdd gnd cell_6t
Xbit_r166_c103 bl_103 br_103 wl_166 vdd gnd cell_6t
Xbit_r167_c103 bl_103 br_103 wl_167 vdd gnd cell_6t
Xbit_r168_c103 bl_103 br_103 wl_168 vdd gnd cell_6t
Xbit_r169_c103 bl_103 br_103 wl_169 vdd gnd cell_6t
Xbit_r170_c103 bl_103 br_103 wl_170 vdd gnd cell_6t
Xbit_r171_c103 bl_103 br_103 wl_171 vdd gnd cell_6t
Xbit_r172_c103 bl_103 br_103 wl_172 vdd gnd cell_6t
Xbit_r173_c103 bl_103 br_103 wl_173 vdd gnd cell_6t
Xbit_r174_c103 bl_103 br_103 wl_174 vdd gnd cell_6t
Xbit_r175_c103 bl_103 br_103 wl_175 vdd gnd cell_6t
Xbit_r176_c103 bl_103 br_103 wl_176 vdd gnd cell_6t
Xbit_r177_c103 bl_103 br_103 wl_177 vdd gnd cell_6t
Xbit_r178_c103 bl_103 br_103 wl_178 vdd gnd cell_6t
Xbit_r179_c103 bl_103 br_103 wl_179 vdd gnd cell_6t
Xbit_r180_c103 bl_103 br_103 wl_180 vdd gnd cell_6t
Xbit_r181_c103 bl_103 br_103 wl_181 vdd gnd cell_6t
Xbit_r182_c103 bl_103 br_103 wl_182 vdd gnd cell_6t
Xbit_r183_c103 bl_103 br_103 wl_183 vdd gnd cell_6t
Xbit_r184_c103 bl_103 br_103 wl_184 vdd gnd cell_6t
Xbit_r185_c103 bl_103 br_103 wl_185 vdd gnd cell_6t
Xbit_r186_c103 bl_103 br_103 wl_186 vdd gnd cell_6t
Xbit_r187_c103 bl_103 br_103 wl_187 vdd gnd cell_6t
Xbit_r188_c103 bl_103 br_103 wl_188 vdd gnd cell_6t
Xbit_r189_c103 bl_103 br_103 wl_189 vdd gnd cell_6t
Xbit_r190_c103 bl_103 br_103 wl_190 vdd gnd cell_6t
Xbit_r191_c103 bl_103 br_103 wl_191 vdd gnd cell_6t
Xbit_r192_c103 bl_103 br_103 wl_192 vdd gnd cell_6t
Xbit_r193_c103 bl_103 br_103 wl_193 vdd gnd cell_6t
Xbit_r194_c103 bl_103 br_103 wl_194 vdd gnd cell_6t
Xbit_r195_c103 bl_103 br_103 wl_195 vdd gnd cell_6t
Xbit_r196_c103 bl_103 br_103 wl_196 vdd gnd cell_6t
Xbit_r197_c103 bl_103 br_103 wl_197 vdd gnd cell_6t
Xbit_r198_c103 bl_103 br_103 wl_198 vdd gnd cell_6t
Xbit_r199_c103 bl_103 br_103 wl_199 vdd gnd cell_6t
Xbit_r200_c103 bl_103 br_103 wl_200 vdd gnd cell_6t
Xbit_r201_c103 bl_103 br_103 wl_201 vdd gnd cell_6t
Xbit_r202_c103 bl_103 br_103 wl_202 vdd gnd cell_6t
Xbit_r203_c103 bl_103 br_103 wl_203 vdd gnd cell_6t
Xbit_r204_c103 bl_103 br_103 wl_204 vdd gnd cell_6t
Xbit_r205_c103 bl_103 br_103 wl_205 vdd gnd cell_6t
Xbit_r206_c103 bl_103 br_103 wl_206 vdd gnd cell_6t
Xbit_r207_c103 bl_103 br_103 wl_207 vdd gnd cell_6t
Xbit_r208_c103 bl_103 br_103 wl_208 vdd gnd cell_6t
Xbit_r209_c103 bl_103 br_103 wl_209 vdd gnd cell_6t
Xbit_r210_c103 bl_103 br_103 wl_210 vdd gnd cell_6t
Xbit_r211_c103 bl_103 br_103 wl_211 vdd gnd cell_6t
Xbit_r212_c103 bl_103 br_103 wl_212 vdd gnd cell_6t
Xbit_r213_c103 bl_103 br_103 wl_213 vdd gnd cell_6t
Xbit_r214_c103 bl_103 br_103 wl_214 vdd gnd cell_6t
Xbit_r215_c103 bl_103 br_103 wl_215 vdd gnd cell_6t
Xbit_r216_c103 bl_103 br_103 wl_216 vdd gnd cell_6t
Xbit_r217_c103 bl_103 br_103 wl_217 vdd gnd cell_6t
Xbit_r218_c103 bl_103 br_103 wl_218 vdd gnd cell_6t
Xbit_r219_c103 bl_103 br_103 wl_219 vdd gnd cell_6t
Xbit_r220_c103 bl_103 br_103 wl_220 vdd gnd cell_6t
Xbit_r221_c103 bl_103 br_103 wl_221 vdd gnd cell_6t
Xbit_r222_c103 bl_103 br_103 wl_222 vdd gnd cell_6t
Xbit_r223_c103 bl_103 br_103 wl_223 vdd gnd cell_6t
Xbit_r224_c103 bl_103 br_103 wl_224 vdd gnd cell_6t
Xbit_r225_c103 bl_103 br_103 wl_225 vdd gnd cell_6t
Xbit_r226_c103 bl_103 br_103 wl_226 vdd gnd cell_6t
Xbit_r227_c103 bl_103 br_103 wl_227 vdd gnd cell_6t
Xbit_r228_c103 bl_103 br_103 wl_228 vdd gnd cell_6t
Xbit_r229_c103 bl_103 br_103 wl_229 vdd gnd cell_6t
Xbit_r230_c103 bl_103 br_103 wl_230 vdd gnd cell_6t
Xbit_r231_c103 bl_103 br_103 wl_231 vdd gnd cell_6t
Xbit_r232_c103 bl_103 br_103 wl_232 vdd gnd cell_6t
Xbit_r233_c103 bl_103 br_103 wl_233 vdd gnd cell_6t
Xbit_r234_c103 bl_103 br_103 wl_234 vdd gnd cell_6t
Xbit_r235_c103 bl_103 br_103 wl_235 vdd gnd cell_6t
Xbit_r236_c103 bl_103 br_103 wl_236 vdd gnd cell_6t
Xbit_r237_c103 bl_103 br_103 wl_237 vdd gnd cell_6t
Xbit_r238_c103 bl_103 br_103 wl_238 vdd gnd cell_6t
Xbit_r239_c103 bl_103 br_103 wl_239 vdd gnd cell_6t
Xbit_r240_c103 bl_103 br_103 wl_240 vdd gnd cell_6t
Xbit_r241_c103 bl_103 br_103 wl_241 vdd gnd cell_6t
Xbit_r242_c103 bl_103 br_103 wl_242 vdd gnd cell_6t
Xbit_r243_c103 bl_103 br_103 wl_243 vdd gnd cell_6t
Xbit_r244_c103 bl_103 br_103 wl_244 vdd gnd cell_6t
Xbit_r245_c103 bl_103 br_103 wl_245 vdd gnd cell_6t
Xbit_r246_c103 bl_103 br_103 wl_246 vdd gnd cell_6t
Xbit_r247_c103 bl_103 br_103 wl_247 vdd gnd cell_6t
Xbit_r248_c103 bl_103 br_103 wl_248 vdd gnd cell_6t
Xbit_r249_c103 bl_103 br_103 wl_249 vdd gnd cell_6t
Xbit_r250_c103 bl_103 br_103 wl_250 vdd gnd cell_6t
Xbit_r251_c103 bl_103 br_103 wl_251 vdd gnd cell_6t
Xbit_r252_c103 bl_103 br_103 wl_252 vdd gnd cell_6t
Xbit_r253_c103 bl_103 br_103 wl_253 vdd gnd cell_6t
Xbit_r254_c103 bl_103 br_103 wl_254 vdd gnd cell_6t
Xbit_r255_c103 bl_103 br_103 wl_255 vdd gnd cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd cell_6t
Xbit_r1_c104 bl_104 br_104 wl_1 vdd gnd cell_6t
Xbit_r2_c104 bl_104 br_104 wl_2 vdd gnd cell_6t
Xbit_r3_c104 bl_104 br_104 wl_3 vdd gnd cell_6t
Xbit_r4_c104 bl_104 br_104 wl_4 vdd gnd cell_6t
Xbit_r5_c104 bl_104 br_104 wl_5 vdd gnd cell_6t
Xbit_r6_c104 bl_104 br_104 wl_6 vdd gnd cell_6t
Xbit_r7_c104 bl_104 br_104 wl_7 vdd gnd cell_6t
Xbit_r8_c104 bl_104 br_104 wl_8 vdd gnd cell_6t
Xbit_r9_c104 bl_104 br_104 wl_9 vdd gnd cell_6t
Xbit_r10_c104 bl_104 br_104 wl_10 vdd gnd cell_6t
Xbit_r11_c104 bl_104 br_104 wl_11 vdd gnd cell_6t
Xbit_r12_c104 bl_104 br_104 wl_12 vdd gnd cell_6t
Xbit_r13_c104 bl_104 br_104 wl_13 vdd gnd cell_6t
Xbit_r14_c104 bl_104 br_104 wl_14 vdd gnd cell_6t
Xbit_r15_c104 bl_104 br_104 wl_15 vdd gnd cell_6t
Xbit_r16_c104 bl_104 br_104 wl_16 vdd gnd cell_6t
Xbit_r17_c104 bl_104 br_104 wl_17 vdd gnd cell_6t
Xbit_r18_c104 bl_104 br_104 wl_18 vdd gnd cell_6t
Xbit_r19_c104 bl_104 br_104 wl_19 vdd gnd cell_6t
Xbit_r20_c104 bl_104 br_104 wl_20 vdd gnd cell_6t
Xbit_r21_c104 bl_104 br_104 wl_21 vdd gnd cell_6t
Xbit_r22_c104 bl_104 br_104 wl_22 vdd gnd cell_6t
Xbit_r23_c104 bl_104 br_104 wl_23 vdd gnd cell_6t
Xbit_r24_c104 bl_104 br_104 wl_24 vdd gnd cell_6t
Xbit_r25_c104 bl_104 br_104 wl_25 vdd gnd cell_6t
Xbit_r26_c104 bl_104 br_104 wl_26 vdd gnd cell_6t
Xbit_r27_c104 bl_104 br_104 wl_27 vdd gnd cell_6t
Xbit_r28_c104 bl_104 br_104 wl_28 vdd gnd cell_6t
Xbit_r29_c104 bl_104 br_104 wl_29 vdd gnd cell_6t
Xbit_r30_c104 bl_104 br_104 wl_30 vdd gnd cell_6t
Xbit_r31_c104 bl_104 br_104 wl_31 vdd gnd cell_6t
Xbit_r32_c104 bl_104 br_104 wl_32 vdd gnd cell_6t
Xbit_r33_c104 bl_104 br_104 wl_33 vdd gnd cell_6t
Xbit_r34_c104 bl_104 br_104 wl_34 vdd gnd cell_6t
Xbit_r35_c104 bl_104 br_104 wl_35 vdd gnd cell_6t
Xbit_r36_c104 bl_104 br_104 wl_36 vdd gnd cell_6t
Xbit_r37_c104 bl_104 br_104 wl_37 vdd gnd cell_6t
Xbit_r38_c104 bl_104 br_104 wl_38 vdd gnd cell_6t
Xbit_r39_c104 bl_104 br_104 wl_39 vdd gnd cell_6t
Xbit_r40_c104 bl_104 br_104 wl_40 vdd gnd cell_6t
Xbit_r41_c104 bl_104 br_104 wl_41 vdd gnd cell_6t
Xbit_r42_c104 bl_104 br_104 wl_42 vdd gnd cell_6t
Xbit_r43_c104 bl_104 br_104 wl_43 vdd gnd cell_6t
Xbit_r44_c104 bl_104 br_104 wl_44 vdd gnd cell_6t
Xbit_r45_c104 bl_104 br_104 wl_45 vdd gnd cell_6t
Xbit_r46_c104 bl_104 br_104 wl_46 vdd gnd cell_6t
Xbit_r47_c104 bl_104 br_104 wl_47 vdd gnd cell_6t
Xbit_r48_c104 bl_104 br_104 wl_48 vdd gnd cell_6t
Xbit_r49_c104 bl_104 br_104 wl_49 vdd gnd cell_6t
Xbit_r50_c104 bl_104 br_104 wl_50 vdd gnd cell_6t
Xbit_r51_c104 bl_104 br_104 wl_51 vdd gnd cell_6t
Xbit_r52_c104 bl_104 br_104 wl_52 vdd gnd cell_6t
Xbit_r53_c104 bl_104 br_104 wl_53 vdd gnd cell_6t
Xbit_r54_c104 bl_104 br_104 wl_54 vdd gnd cell_6t
Xbit_r55_c104 bl_104 br_104 wl_55 vdd gnd cell_6t
Xbit_r56_c104 bl_104 br_104 wl_56 vdd gnd cell_6t
Xbit_r57_c104 bl_104 br_104 wl_57 vdd gnd cell_6t
Xbit_r58_c104 bl_104 br_104 wl_58 vdd gnd cell_6t
Xbit_r59_c104 bl_104 br_104 wl_59 vdd gnd cell_6t
Xbit_r60_c104 bl_104 br_104 wl_60 vdd gnd cell_6t
Xbit_r61_c104 bl_104 br_104 wl_61 vdd gnd cell_6t
Xbit_r62_c104 bl_104 br_104 wl_62 vdd gnd cell_6t
Xbit_r63_c104 bl_104 br_104 wl_63 vdd gnd cell_6t
Xbit_r64_c104 bl_104 br_104 wl_64 vdd gnd cell_6t
Xbit_r65_c104 bl_104 br_104 wl_65 vdd gnd cell_6t
Xbit_r66_c104 bl_104 br_104 wl_66 vdd gnd cell_6t
Xbit_r67_c104 bl_104 br_104 wl_67 vdd gnd cell_6t
Xbit_r68_c104 bl_104 br_104 wl_68 vdd gnd cell_6t
Xbit_r69_c104 bl_104 br_104 wl_69 vdd gnd cell_6t
Xbit_r70_c104 bl_104 br_104 wl_70 vdd gnd cell_6t
Xbit_r71_c104 bl_104 br_104 wl_71 vdd gnd cell_6t
Xbit_r72_c104 bl_104 br_104 wl_72 vdd gnd cell_6t
Xbit_r73_c104 bl_104 br_104 wl_73 vdd gnd cell_6t
Xbit_r74_c104 bl_104 br_104 wl_74 vdd gnd cell_6t
Xbit_r75_c104 bl_104 br_104 wl_75 vdd gnd cell_6t
Xbit_r76_c104 bl_104 br_104 wl_76 vdd gnd cell_6t
Xbit_r77_c104 bl_104 br_104 wl_77 vdd gnd cell_6t
Xbit_r78_c104 bl_104 br_104 wl_78 vdd gnd cell_6t
Xbit_r79_c104 bl_104 br_104 wl_79 vdd gnd cell_6t
Xbit_r80_c104 bl_104 br_104 wl_80 vdd gnd cell_6t
Xbit_r81_c104 bl_104 br_104 wl_81 vdd gnd cell_6t
Xbit_r82_c104 bl_104 br_104 wl_82 vdd gnd cell_6t
Xbit_r83_c104 bl_104 br_104 wl_83 vdd gnd cell_6t
Xbit_r84_c104 bl_104 br_104 wl_84 vdd gnd cell_6t
Xbit_r85_c104 bl_104 br_104 wl_85 vdd gnd cell_6t
Xbit_r86_c104 bl_104 br_104 wl_86 vdd gnd cell_6t
Xbit_r87_c104 bl_104 br_104 wl_87 vdd gnd cell_6t
Xbit_r88_c104 bl_104 br_104 wl_88 vdd gnd cell_6t
Xbit_r89_c104 bl_104 br_104 wl_89 vdd gnd cell_6t
Xbit_r90_c104 bl_104 br_104 wl_90 vdd gnd cell_6t
Xbit_r91_c104 bl_104 br_104 wl_91 vdd gnd cell_6t
Xbit_r92_c104 bl_104 br_104 wl_92 vdd gnd cell_6t
Xbit_r93_c104 bl_104 br_104 wl_93 vdd gnd cell_6t
Xbit_r94_c104 bl_104 br_104 wl_94 vdd gnd cell_6t
Xbit_r95_c104 bl_104 br_104 wl_95 vdd gnd cell_6t
Xbit_r96_c104 bl_104 br_104 wl_96 vdd gnd cell_6t
Xbit_r97_c104 bl_104 br_104 wl_97 vdd gnd cell_6t
Xbit_r98_c104 bl_104 br_104 wl_98 vdd gnd cell_6t
Xbit_r99_c104 bl_104 br_104 wl_99 vdd gnd cell_6t
Xbit_r100_c104 bl_104 br_104 wl_100 vdd gnd cell_6t
Xbit_r101_c104 bl_104 br_104 wl_101 vdd gnd cell_6t
Xbit_r102_c104 bl_104 br_104 wl_102 vdd gnd cell_6t
Xbit_r103_c104 bl_104 br_104 wl_103 vdd gnd cell_6t
Xbit_r104_c104 bl_104 br_104 wl_104 vdd gnd cell_6t
Xbit_r105_c104 bl_104 br_104 wl_105 vdd gnd cell_6t
Xbit_r106_c104 bl_104 br_104 wl_106 vdd gnd cell_6t
Xbit_r107_c104 bl_104 br_104 wl_107 vdd gnd cell_6t
Xbit_r108_c104 bl_104 br_104 wl_108 vdd gnd cell_6t
Xbit_r109_c104 bl_104 br_104 wl_109 vdd gnd cell_6t
Xbit_r110_c104 bl_104 br_104 wl_110 vdd gnd cell_6t
Xbit_r111_c104 bl_104 br_104 wl_111 vdd gnd cell_6t
Xbit_r112_c104 bl_104 br_104 wl_112 vdd gnd cell_6t
Xbit_r113_c104 bl_104 br_104 wl_113 vdd gnd cell_6t
Xbit_r114_c104 bl_104 br_104 wl_114 vdd gnd cell_6t
Xbit_r115_c104 bl_104 br_104 wl_115 vdd gnd cell_6t
Xbit_r116_c104 bl_104 br_104 wl_116 vdd gnd cell_6t
Xbit_r117_c104 bl_104 br_104 wl_117 vdd gnd cell_6t
Xbit_r118_c104 bl_104 br_104 wl_118 vdd gnd cell_6t
Xbit_r119_c104 bl_104 br_104 wl_119 vdd gnd cell_6t
Xbit_r120_c104 bl_104 br_104 wl_120 vdd gnd cell_6t
Xbit_r121_c104 bl_104 br_104 wl_121 vdd gnd cell_6t
Xbit_r122_c104 bl_104 br_104 wl_122 vdd gnd cell_6t
Xbit_r123_c104 bl_104 br_104 wl_123 vdd gnd cell_6t
Xbit_r124_c104 bl_104 br_104 wl_124 vdd gnd cell_6t
Xbit_r125_c104 bl_104 br_104 wl_125 vdd gnd cell_6t
Xbit_r126_c104 bl_104 br_104 wl_126 vdd gnd cell_6t
Xbit_r127_c104 bl_104 br_104 wl_127 vdd gnd cell_6t
Xbit_r128_c104 bl_104 br_104 wl_128 vdd gnd cell_6t
Xbit_r129_c104 bl_104 br_104 wl_129 vdd gnd cell_6t
Xbit_r130_c104 bl_104 br_104 wl_130 vdd gnd cell_6t
Xbit_r131_c104 bl_104 br_104 wl_131 vdd gnd cell_6t
Xbit_r132_c104 bl_104 br_104 wl_132 vdd gnd cell_6t
Xbit_r133_c104 bl_104 br_104 wl_133 vdd gnd cell_6t
Xbit_r134_c104 bl_104 br_104 wl_134 vdd gnd cell_6t
Xbit_r135_c104 bl_104 br_104 wl_135 vdd gnd cell_6t
Xbit_r136_c104 bl_104 br_104 wl_136 vdd gnd cell_6t
Xbit_r137_c104 bl_104 br_104 wl_137 vdd gnd cell_6t
Xbit_r138_c104 bl_104 br_104 wl_138 vdd gnd cell_6t
Xbit_r139_c104 bl_104 br_104 wl_139 vdd gnd cell_6t
Xbit_r140_c104 bl_104 br_104 wl_140 vdd gnd cell_6t
Xbit_r141_c104 bl_104 br_104 wl_141 vdd gnd cell_6t
Xbit_r142_c104 bl_104 br_104 wl_142 vdd gnd cell_6t
Xbit_r143_c104 bl_104 br_104 wl_143 vdd gnd cell_6t
Xbit_r144_c104 bl_104 br_104 wl_144 vdd gnd cell_6t
Xbit_r145_c104 bl_104 br_104 wl_145 vdd gnd cell_6t
Xbit_r146_c104 bl_104 br_104 wl_146 vdd gnd cell_6t
Xbit_r147_c104 bl_104 br_104 wl_147 vdd gnd cell_6t
Xbit_r148_c104 bl_104 br_104 wl_148 vdd gnd cell_6t
Xbit_r149_c104 bl_104 br_104 wl_149 vdd gnd cell_6t
Xbit_r150_c104 bl_104 br_104 wl_150 vdd gnd cell_6t
Xbit_r151_c104 bl_104 br_104 wl_151 vdd gnd cell_6t
Xbit_r152_c104 bl_104 br_104 wl_152 vdd gnd cell_6t
Xbit_r153_c104 bl_104 br_104 wl_153 vdd gnd cell_6t
Xbit_r154_c104 bl_104 br_104 wl_154 vdd gnd cell_6t
Xbit_r155_c104 bl_104 br_104 wl_155 vdd gnd cell_6t
Xbit_r156_c104 bl_104 br_104 wl_156 vdd gnd cell_6t
Xbit_r157_c104 bl_104 br_104 wl_157 vdd gnd cell_6t
Xbit_r158_c104 bl_104 br_104 wl_158 vdd gnd cell_6t
Xbit_r159_c104 bl_104 br_104 wl_159 vdd gnd cell_6t
Xbit_r160_c104 bl_104 br_104 wl_160 vdd gnd cell_6t
Xbit_r161_c104 bl_104 br_104 wl_161 vdd gnd cell_6t
Xbit_r162_c104 bl_104 br_104 wl_162 vdd gnd cell_6t
Xbit_r163_c104 bl_104 br_104 wl_163 vdd gnd cell_6t
Xbit_r164_c104 bl_104 br_104 wl_164 vdd gnd cell_6t
Xbit_r165_c104 bl_104 br_104 wl_165 vdd gnd cell_6t
Xbit_r166_c104 bl_104 br_104 wl_166 vdd gnd cell_6t
Xbit_r167_c104 bl_104 br_104 wl_167 vdd gnd cell_6t
Xbit_r168_c104 bl_104 br_104 wl_168 vdd gnd cell_6t
Xbit_r169_c104 bl_104 br_104 wl_169 vdd gnd cell_6t
Xbit_r170_c104 bl_104 br_104 wl_170 vdd gnd cell_6t
Xbit_r171_c104 bl_104 br_104 wl_171 vdd gnd cell_6t
Xbit_r172_c104 bl_104 br_104 wl_172 vdd gnd cell_6t
Xbit_r173_c104 bl_104 br_104 wl_173 vdd gnd cell_6t
Xbit_r174_c104 bl_104 br_104 wl_174 vdd gnd cell_6t
Xbit_r175_c104 bl_104 br_104 wl_175 vdd gnd cell_6t
Xbit_r176_c104 bl_104 br_104 wl_176 vdd gnd cell_6t
Xbit_r177_c104 bl_104 br_104 wl_177 vdd gnd cell_6t
Xbit_r178_c104 bl_104 br_104 wl_178 vdd gnd cell_6t
Xbit_r179_c104 bl_104 br_104 wl_179 vdd gnd cell_6t
Xbit_r180_c104 bl_104 br_104 wl_180 vdd gnd cell_6t
Xbit_r181_c104 bl_104 br_104 wl_181 vdd gnd cell_6t
Xbit_r182_c104 bl_104 br_104 wl_182 vdd gnd cell_6t
Xbit_r183_c104 bl_104 br_104 wl_183 vdd gnd cell_6t
Xbit_r184_c104 bl_104 br_104 wl_184 vdd gnd cell_6t
Xbit_r185_c104 bl_104 br_104 wl_185 vdd gnd cell_6t
Xbit_r186_c104 bl_104 br_104 wl_186 vdd gnd cell_6t
Xbit_r187_c104 bl_104 br_104 wl_187 vdd gnd cell_6t
Xbit_r188_c104 bl_104 br_104 wl_188 vdd gnd cell_6t
Xbit_r189_c104 bl_104 br_104 wl_189 vdd gnd cell_6t
Xbit_r190_c104 bl_104 br_104 wl_190 vdd gnd cell_6t
Xbit_r191_c104 bl_104 br_104 wl_191 vdd gnd cell_6t
Xbit_r192_c104 bl_104 br_104 wl_192 vdd gnd cell_6t
Xbit_r193_c104 bl_104 br_104 wl_193 vdd gnd cell_6t
Xbit_r194_c104 bl_104 br_104 wl_194 vdd gnd cell_6t
Xbit_r195_c104 bl_104 br_104 wl_195 vdd gnd cell_6t
Xbit_r196_c104 bl_104 br_104 wl_196 vdd gnd cell_6t
Xbit_r197_c104 bl_104 br_104 wl_197 vdd gnd cell_6t
Xbit_r198_c104 bl_104 br_104 wl_198 vdd gnd cell_6t
Xbit_r199_c104 bl_104 br_104 wl_199 vdd gnd cell_6t
Xbit_r200_c104 bl_104 br_104 wl_200 vdd gnd cell_6t
Xbit_r201_c104 bl_104 br_104 wl_201 vdd gnd cell_6t
Xbit_r202_c104 bl_104 br_104 wl_202 vdd gnd cell_6t
Xbit_r203_c104 bl_104 br_104 wl_203 vdd gnd cell_6t
Xbit_r204_c104 bl_104 br_104 wl_204 vdd gnd cell_6t
Xbit_r205_c104 bl_104 br_104 wl_205 vdd gnd cell_6t
Xbit_r206_c104 bl_104 br_104 wl_206 vdd gnd cell_6t
Xbit_r207_c104 bl_104 br_104 wl_207 vdd gnd cell_6t
Xbit_r208_c104 bl_104 br_104 wl_208 vdd gnd cell_6t
Xbit_r209_c104 bl_104 br_104 wl_209 vdd gnd cell_6t
Xbit_r210_c104 bl_104 br_104 wl_210 vdd gnd cell_6t
Xbit_r211_c104 bl_104 br_104 wl_211 vdd gnd cell_6t
Xbit_r212_c104 bl_104 br_104 wl_212 vdd gnd cell_6t
Xbit_r213_c104 bl_104 br_104 wl_213 vdd gnd cell_6t
Xbit_r214_c104 bl_104 br_104 wl_214 vdd gnd cell_6t
Xbit_r215_c104 bl_104 br_104 wl_215 vdd gnd cell_6t
Xbit_r216_c104 bl_104 br_104 wl_216 vdd gnd cell_6t
Xbit_r217_c104 bl_104 br_104 wl_217 vdd gnd cell_6t
Xbit_r218_c104 bl_104 br_104 wl_218 vdd gnd cell_6t
Xbit_r219_c104 bl_104 br_104 wl_219 vdd gnd cell_6t
Xbit_r220_c104 bl_104 br_104 wl_220 vdd gnd cell_6t
Xbit_r221_c104 bl_104 br_104 wl_221 vdd gnd cell_6t
Xbit_r222_c104 bl_104 br_104 wl_222 vdd gnd cell_6t
Xbit_r223_c104 bl_104 br_104 wl_223 vdd gnd cell_6t
Xbit_r224_c104 bl_104 br_104 wl_224 vdd gnd cell_6t
Xbit_r225_c104 bl_104 br_104 wl_225 vdd gnd cell_6t
Xbit_r226_c104 bl_104 br_104 wl_226 vdd gnd cell_6t
Xbit_r227_c104 bl_104 br_104 wl_227 vdd gnd cell_6t
Xbit_r228_c104 bl_104 br_104 wl_228 vdd gnd cell_6t
Xbit_r229_c104 bl_104 br_104 wl_229 vdd gnd cell_6t
Xbit_r230_c104 bl_104 br_104 wl_230 vdd gnd cell_6t
Xbit_r231_c104 bl_104 br_104 wl_231 vdd gnd cell_6t
Xbit_r232_c104 bl_104 br_104 wl_232 vdd gnd cell_6t
Xbit_r233_c104 bl_104 br_104 wl_233 vdd gnd cell_6t
Xbit_r234_c104 bl_104 br_104 wl_234 vdd gnd cell_6t
Xbit_r235_c104 bl_104 br_104 wl_235 vdd gnd cell_6t
Xbit_r236_c104 bl_104 br_104 wl_236 vdd gnd cell_6t
Xbit_r237_c104 bl_104 br_104 wl_237 vdd gnd cell_6t
Xbit_r238_c104 bl_104 br_104 wl_238 vdd gnd cell_6t
Xbit_r239_c104 bl_104 br_104 wl_239 vdd gnd cell_6t
Xbit_r240_c104 bl_104 br_104 wl_240 vdd gnd cell_6t
Xbit_r241_c104 bl_104 br_104 wl_241 vdd gnd cell_6t
Xbit_r242_c104 bl_104 br_104 wl_242 vdd gnd cell_6t
Xbit_r243_c104 bl_104 br_104 wl_243 vdd gnd cell_6t
Xbit_r244_c104 bl_104 br_104 wl_244 vdd gnd cell_6t
Xbit_r245_c104 bl_104 br_104 wl_245 vdd gnd cell_6t
Xbit_r246_c104 bl_104 br_104 wl_246 vdd gnd cell_6t
Xbit_r247_c104 bl_104 br_104 wl_247 vdd gnd cell_6t
Xbit_r248_c104 bl_104 br_104 wl_248 vdd gnd cell_6t
Xbit_r249_c104 bl_104 br_104 wl_249 vdd gnd cell_6t
Xbit_r250_c104 bl_104 br_104 wl_250 vdd gnd cell_6t
Xbit_r251_c104 bl_104 br_104 wl_251 vdd gnd cell_6t
Xbit_r252_c104 bl_104 br_104 wl_252 vdd gnd cell_6t
Xbit_r253_c104 bl_104 br_104 wl_253 vdd gnd cell_6t
Xbit_r254_c104 bl_104 br_104 wl_254 vdd gnd cell_6t
Xbit_r255_c104 bl_104 br_104 wl_255 vdd gnd cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd cell_6t
Xbit_r1_c105 bl_105 br_105 wl_1 vdd gnd cell_6t
Xbit_r2_c105 bl_105 br_105 wl_2 vdd gnd cell_6t
Xbit_r3_c105 bl_105 br_105 wl_3 vdd gnd cell_6t
Xbit_r4_c105 bl_105 br_105 wl_4 vdd gnd cell_6t
Xbit_r5_c105 bl_105 br_105 wl_5 vdd gnd cell_6t
Xbit_r6_c105 bl_105 br_105 wl_6 vdd gnd cell_6t
Xbit_r7_c105 bl_105 br_105 wl_7 vdd gnd cell_6t
Xbit_r8_c105 bl_105 br_105 wl_8 vdd gnd cell_6t
Xbit_r9_c105 bl_105 br_105 wl_9 vdd gnd cell_6t
Xbit_r10_c105 bl_105 br_105 wl_10 vdd gnd cell_6t
Xbit_r11_c105 bl_105 br_105 wl_11 vdd gnd cell_6t
Xbit_r12_c105 bl_105 br_105 wl_12 vdd gnd cell_6t
Xbit_r13_c105 bl_105 br_105 wl_13 vdd gnd cell_6t
Xbit_r14_c105 bl_105 br_105 wl_14 vdd gnd cell_6t
Xbit_r15_c105 bl_105 br_105 wl_15 vdd gnd cell_6t
Xbit_r16_c105 bl_105 br_105 wl_16 vdd gnd cell_6t
Xbit_r17_c105 bl_105 br_105 wl_17 vdd gnd cell_6t
Xbit_r18_c105 bl_105 br_105 wl_18 vdd gnd cell_6t
Xbit_r19_c105 bl_105 br_105 wl_19 vdd gnd cell_6t
Xbit_r20_c105 bl_105 br_105 wl_20 vdd gnd cell_6t
Xbit_r21_c105 bl_105 br_105 wl_21 vdd gnd cell_6t
Xbit_r22_c105 bl_105 br_105 wl_22 vdd gnd cell_6t
Xbit_r23_c105 bl_105 br_105 wl_23 vdd gnd cell_6t
Xbit_r24_c105 bl_105 br_105 wl_24 vdd gnd cell_6t
Xbit_r25_c105 bl_105 br_105 wl_25 vdd gnd cell_6t
Xbit_r26_c105 bl_105 br_105 wl_26 vdd gnd cell_6t
Xbit_r27_c105 bl_105 br_105 wl_27 vdd gnd cell_6t
Xbit_r28_c105 bl_105 br_105 wl_28 vdd gnd cell_6t
Xbit_r29_c105 bl_105 br_105 wl_29 vdd gnd cell_6t
Xbit_r30_c105 bl_105 br_105 wl_30 vdd gnd cell_6t
Xbit_r31_c105 bl_105 br_105 wl_31 vdd gnd cell_6t
Xbit_r32_c105 bl_105 br_105 wl_32 vdd gnd cell_6t
Xbit_r33_c105 bl_105 br_105 wl_33 vdd gnd cell_6t
Xbit_r34_c105 bl_105 br_105 wl_34 vdd gnd cell_6t
Xbit_r35_c105 bl_105 br_105 wl_35 vdd gnd cell_6t
Xbit_r36_c105 bl_105 br_105 wl_36 vdd gnd cell_6t
Xbit_r37_c105 bl_105 br_105 wl_37 vdd gnd cell_6t
Xbit_r38_c105 bl_105 br_105 wl_38 vdd gnd cell_6t
Xbit_r39_c105 bl_105 br_105 wl_39 vdd gnd cell_6t
Xbit_r40_c105 bl_105 br_105 wl_40 vdd gnd cell_6t
Xbit_r41_c105 bl_105 br_105 wl_41 vdd gnd cell_6t
Xbit_r42_c105 bl_105 br_105 wl_42 vdd gnd cell_6t
Xbit_r43_c105 bl_105 br_105 wl_43 vdd gnd cell_6t
Xbit_r44_c105 bl_105 br_105 wl_44 vdd gnd cell_6t
Xbit_r45_c105 bl_105 br_105 wl_45 vdd gnd cell_6t
Xbit_r46_c105 bl_105 br_105 wl_46 vdd gnd cell_6t
Xbit_r47_c105 bl_105 br_105 wl_47 vdd gnd cell_6t
Xbit_r48_c105 bl_105 br_105 wl_48 vdd gnd cell_6t
Xbit_r49_c105 bl_105 br_105 wl_49 vdd gnd cell_6t
Xbit_r50_c105 bl_105 br_105 wl_50 vdd gnd cell_6t
Xbit_r51_c105 bl_105 br_105 wl_51 vdd gnd cell_6t
Xbit_r52_c105 bl_105 br_105 wl_52 vdd gnd cell_6t
Xbit_r53_c105 bl_105 br_105 wl_53 vdd gnd cell_6t
Xbit_r54_c105 bl_105 br_105 wl_54 vdd gnd cell_6t
Xbit_r55_c105 bl_105 br_105 wl_55 vdd gnd cell_6t
Xbit_r56_c105 bl_105 br_105 wl_56 vdd gnd cell_6t
Xbit_r57_c105 bl_105 br_105 wl_57 vdd gnd cell_6t
Xbit_r58_c105 bl_105 br_105 wl_58 vdd gnd cell_6t
Xbit_r59_c105 bl_105 br_105 wl_59 vdd gnd cell_6t
Xbit_r60_c105 bl_105 br_105 wl_60 vdd gnd cell_6t
Xbit_r61_c105 bl_105 br_105 wl_61 vdd gnd cell_6t
Xbit_r62_c105 bl_105 br_105 wl_62 vdd gnd cell_6t
Xbit_r63_c105 bl_105 br_105 wl_63 vdd gnd cell_6t
Xbit_r64_c105 bl_105 br_105 wl_64 vdd gnd cell_6t
Xbit_r65_c105 bl_105 br_105 wl_65 vdd gnd cell_6t
Xbit_r66_c105 bl_105 br_105 wl_66 vdd gnd cell_6t
Xbit_r67_c105 bl_105 br_105 wl_67 vdd gnd cell_6t
Xbit_r68_c105 bl_105 br_105 wl_68 vdd gnd cell_6t
Xbit_r69_c105 bl_105 br_105 wl_69 vdd gnd cell_6t
Xbit_r70_c105 bl_105 br_105 wl_70 vdd gnd cell_6t
Xbit_r71_c105 bl_105 br_105 wl_71 vdd gnd cell_6t
Xbit_r72_c105 bl_105 br_105 wl_72 vdd gnd cell_6t
Xbit_r73_c105 bl_105 br_105 wl_73 vdd gnd cell_6t
Xbit_r74_c105 bl_105 br_105 wl_74 vdd gnd cell_6t
Xbit_r75_c105 bl_105 br_105 wl_75 vdd gnd cell_6t
Xbit_r76_c105 bl_105 br_105 wl_76 vdd gnd cell_6t
Xbit_r77_c105 bl_105 br_105 wl_77 vdd gnd cell_6t
Xbit_r78_c105 bl_105 br_105 wl_78 vdd gnd cell_6t
Xbit_r79_c105 bl_105 br_105 wl_79 vdd gnd cell_6t
Xbit_r80_c105 bl_105 br_105 wl_80 vdd gnd cell_6t
Xbit_r81_c105 bl_105 br_105 wl_81 vdd gnd cell_6t
Xbit_r82_c105 bl_105 br_105 wl_82 vdd gnd cell_6t
Xbit_r83_c105 bl_105 br_105 wl_83 vdd gnd cell_6t
Xbit_r84_c105 bl_105 br_105 wl_84 vdd gnd cell_6t
Xbit_r85_c105 bl_105 br_105 wl_85 vdd gnd cell_6t
Xbit_r86_c105 bl_105 br_105 wl_86 vdd gnd cell_6t
Xbit_r87_c105 bl_105 br_105 wl_87 vdd gnd cell_6t
Xbit_r88_c105 bl_105 br_105 wl_88 vdd gnd cell_6t
Xbit_r89_c105 bl_105 br_105 wl_89 vdd gnd cell_6t
Xbit_r90_c105 bl_105 br_105 wl_90 vdd gnd cell_6t
Xbit_r91_c105 bl_105 br_105 wl_91 vdd gnd cell_6t
Xbit_r92_c105 bl_105 br_105 wl_92 vdd gnd cell_6t
Xbit_r93_c105 bl_105 br_105 wl_93 vdd gnd cell_6t
Xbit_r94_c105 bl_105 br_105 wl_94 vdd gnd cell_6t
Xbit_r95_c105 bl_105 br_105 wl_95 vdd gnd cell_6t
Xbit_r96_c105 bl_105 br_105 wl_96 vdd gnd cell_6t
Xbit_r97_c105 bl_105 br_105 wl_97 vdd gnd cell_6t
Xbit_r98_c105 bl_105 br_105 wl_98 vdd gnd cell_6t
Xbit_r99_c105 bl_105 br_105 wl_99 vdd gnd cell_6t
Xbit_r100_c105 bl_105 br_105 wl_100 vdd gnd cell_6t
Xbit_r101_c105 bl_105 br_105 wl_101 vdd gnd cell_6t
Xbit_r102_c105 bl_105 br_105 wl_102 vdd gnd cell_6t
Xbit_r103_c105 bl_105 br_105 wl_103 vdd gnd cell_6t
Xbit_r104_c105 bl_105 br_105 wl_104 vdd gnd cell_6t
Xbit_r105_c105 bl_105 br_105 wl_105 vdd gnd cell_6t
Xbit_r106_c105 bl_105 br_105 wl_106 vdd gnd cell_6t
Xbit_r107_c105 bl_105 br_105 wl_107 vdd gnd cell_6t
Xbit_r108_c105 bl_105 br_105 wl_108 vdd gnd cell_6t
Xbit_r109_c105 bl_105 br_105 wl_109 vdd gnd cell_6t
Xbit_r110_c105 bl_105 br_105 wl_110 vdd gnd cell_6t
Xbit_r111_c105 bl_105 br_105 wl_111 vdd gnd cell_6t
Xbit_r112_c105 bl_105 br_105 wl_112 vdd gnd cell_6t
Xbit_r113_c105 bl_105 br_105 wl_113 vdd gnd cell_6t
Xbit_r114_c105 bl_105 br_105 wl_114 vdd gnd cell_6t
Xbit_r115_c105 bl_105 br_105 wl_115 vdd gnd cell_6t
Xbit_r116_c105 bl_105 br_105 wl_116 vdd gnd cell_6t
Xbit_r117_c105 bl_105 br_105 wl_117 vdd gnd cell_6t
Xbit_r118_c105 bl_105 br_105 wl_118 vdd gnd cell_6t
Xbit_r119_c105 bl_105 br_105 wl_119 vdd gnd cell_6t
Xbit_r120_c105 bl_105 br_105 wl_120 vdd gnd cell_6t
Xbit_r121_c105 bl_105 br_105 wl_121 vdd gnd cell_6t
Xbit_r122_c105 bl_105 br_105 wl_122 vdd gnd cell_6t
Xbit_r123_c105 bl_105 br_105 wl_123 vdd gnd cell_6t
Xbit_r124_c105 bl_105 br_105 wl_124 vdd gnd cell_6t
Xbit_r125_c105 bl_105 br_105 wl_125 vdd gnd cell_6t
Xbit_r126_c105 bl_105 br_105 wl_126 vdd gnd cell_6t
Xbit_r127_c105 bl_105 br_105 wl_127 vdd gnd cell_6t
Xbit_r128_c105 bl_105 br_105 wl_128 vdd gnd cell_6t
Xbit_r129_c105 bl_105 br_105 wl_129 vdd gnd cell_6t
Xbit_r130_c105 bl_105 br_105 wl_130 vdd gnd cell_6t
Xbit_r131_c105 bl_105 br_105 wl_131 vdd gnd cell_6t
Xbit_r132_c105 bl_105 br_105 wl_132 vdd gnd cell_6t
Xbit_r133_c105 bl_105 br_105 wl_133 vdd gnd cell_6t
Xbit_r134_c105 bl_105 br_105 wl_134 vdd gnd cell_6t
Xbit_r135_c105 bl_105 br_105 wl_135 vdd gnd cell_6t
Xbit_r136_c105 bl_105 br_105 wl_136 vdd gnd cell_6t
Xbit_r137_c105 bl_105 br_105 wl_137 vdd gnd cell_6t
Xbit_r138_c105 bl_105 br_105 wl_138 vdd gnd cell_6t
Xbit_r139_c105 bl_105 br_105 wl_139 vdd gnd cell_6t
Xbit_r140_c105 bl_105 br_105 wl_140 vdd gnd cell_6t
Xbit_r141_c105 bl_105 br_105 wl_141 vdd gnd cell_6t
Xbit_r142_c105 bl_105 br_105 wl_142 vdd gnd cell_6t
Xbit_r143_c105 bl_105 br_105 wl_143 vdd gnd cell_6t
Xbit_r144_c105 bl_105 br_105 wl_144 vdd gnd cell_6t
Xbit_r145_c105 bl_105 br_105 wl_145 vdd gnd cell_6t
Xbit_r146_c105 bl_105 br_105 wl_146 vdd gnd cell_6t
Xbit_r147_c105 bl_105 br_105 wl_147 vdd gnd cell_6t
Xbit_r148_c105 bl_105 br_105 wl_148 vdd gnd cell_6t
Xbit_r149_c105 bl_105 br_105 wl_149 vdd gnd cell_6t
Xbit_r150_c105 bl_105 br_105 wl_150 vdd gnd cell_6t
Xbit_r151_c105 bl_105 br_105 wl_151 vdd gnd cell_6t
Xbit_r152_c105 bl_105 br_105 wl_152 vdd gnd cell_6t
Xbit_r153_c105 bl_105 br_105 wl_153 vdd gnd cell_6t
Xbit_r154_c105 bl_105 br_105 wl_154 vdd gnd cell_6t
Xbit_r155_c105 bl_105 br_105 wl_155 vdd gnd cell_6t
Xbit_r156_c105 bl_105 br_105 wl_156 vdd gnd cell_6t
Xbit_r157_c105 bl_105 br_105 wl_157 vdd gnd cell_6t
Xbit_r158_c105 bl_105 br_105 wl_158 vdd gnd cell_6t
Xbit_r159_c105 bl_105 br_105 wl_159 vdd gnd cell_6t
Xbit_r160_c105 bl_105 br_105 wl_160 vdd gnd cell_6t
Xbit_r161_c105 bl_105 br_105 wl_161 vdd gnd cell_6t
Xbit_r162_c105 bl_105 br_105 wl_162 vdd gnd cell_6t
Xbit_r163_c105 bl_105 br_105 wl_163 vdd gnd cell_6t
Xbit_r164_c105 bl_105 br_105 wl_164 vdd gnd cell_6t
Xbit_r165_c105 bl_105 br_105 wl_165 vdd gnd cell_6t
Xbit_r166_c105 bl_105 br_105 wl_166 vdd gnd cell_6t
Xbit_r167_c105 bl_105 br_105 wl_167 vdd gnd cell_6t
Xbit_r168_c105 bl_105 br_105 wl_168 vdd gnd cell_6t
Xbit_r169_c105 bl_105 br_105 wl_169 vdd gnd cell_6t
Xbit_r170_c105 bl_105 br_105 wl_170 vdd gnd cell_6t
Xbit_r171_c105 bl_105 br_105 wl_171 vdd gnd cell_6t
Xbit_r172_c105 bl_105 br_105 wl_172 vdd gnd cell_6t
Xbit_r173_c105 bl_105 br_105 wl_173 vdd gnd cell_6t
Xbit_r174_c105 bl_105 br_105 wl_174 vdd gnd cell_6t
Xbit_r175_c105 bl_105 br_105 wl_175 vdd gnd cell_6t
Xbit_r176_c105 bl_105 br_105 wl_176 vdd gnd cell_6t
Xbit_r177_c105 bl_105 br_105 wl_177 vdd gnd cell_6t
Xbit_r178_c105 bl_105 br_105 wl_178 vdd gnd cell_6t
Xbit_r179_c105 bl_105 br_105 wl_179 vdd gnd cell_6t
Xbit_r180_c105 bl_105 br_105 wl_180 vdd gnd cell_6t
Xbit_r181_c105 bl_105 br_105 wl_181 vdd gnd cell_6t
Xbit_r182_c105 bl_105 br_105 wl_182 vdd gnd cell_6t
Xbit_r183_c105 bl_105 br_105 wl_183 vdd gnd cell_6t
Xbit_r184_c105 bl_105 br_105 wl_184 vdd gnd cell_6t
Xbit_r185_c105 bl_105 br_105 wl_185 vdd gnd cell_6t
Xbit_r186_c105 bl_105 br_105 wl_186 vdd gnd cell_6t
Xbit_r187_c105 bl_105 br_105 wl_187 vdd gnd cell_6t
Xbit_r188_c105 bl_105 br_105 wl_188 vdd gnd cell_6t
Xbit_r189_c105 bl_105 br_105 wl_189 vdd gnd cell_6t
Xbit_r190_c105 bl_105 br_105 wl_190 vdd gnd cell_6t
Xbit_r191_c105 bl_105 br_105 wl_191 vdd gnd cell_6t
Xbit_r192_c105 bl_105 br_105 wl_192 vdd gnd cell_6t
Xbit_r193_c105 bl_105 br_105 wl_193 vdd gnd cell_6t
Xbit_r194_c105 bl_105 br_105 wl_194 vdd gnd cell_6t
Xbit_r195_c105 bl_105 br_105 wl_195 vdd gnd cell_6t
Xbit_r196_c105 bl_105 br_105 wl_196 vdd gnd cell_6t
Xbit_r197_c105 bl_105 br_105 wl_197 vdd gnd cell_6t
Xbit_r198_c105 bl_105 br_105 wl_198 vdd gnd cell_6t
Xbit_r199_c105 bl_105 br_105 wl_199 vdd gnd cell_6t
Xbit_r200_c105 bl_105 br_105 wl_200 vdd gnd cell_6t
Xbit_r201_c105 bl_105 br_105 wl_201 vdd gnd cell_6t
Xbit_r202_c105 bl_105 br_105 wl_202 vdd gnd cell_6t
Xbit_r203_c105 bl_105 br_105 wl_203 vdd gnd cell_6t
Xbit_r204_c105 bl_105 br_105 wl_204 vdd gnd cell_6t
Xbit_r205_c105 bl_105 br_105 wl_205 vdd gnd cell_6t
Xbit_r206_c105 bl_105 br_105 wl_206 vdd gnd cell_6t
Xbit_r207_c105 bl_105 br_105 wl_207 vdd gnd cell_6t
Xbit_r208_c105 bl_105 br_105 wl_208 vdd gnd cell_6t
Xbit_r209_c105 bl_105 br_105 wl_209 vdd gnd cell_6t
Xbit_r210_c105 bl_105 br_105 wl_210 vdd gnd cell_6t
Xbit_r211_c105 bl_105 br_105 wl_211 vdd gnd cell_6t
Xbit_r212_c105 bl_105 br_105 wl_212 vdd gnd cell_6t
Xbit_r213_c105 bl_105 br_105 wl_213 vdd gnd cell_6t
Xbit_r214_c105 bl_105 br_105 wl_214 vdd gnd cell_6t
Xbit_r215_c105 bl_105 br_105 wl_215 vdd gnd cell_6t
Xbit_r216_c105 bl_105 br_105 wl_216 vdd gnd cell_6t
Xbit_r217_c105 bl_105 br_105 wl_217 vdd gnd cell_6t
Xbit_r218_c105 bl_105 br_105 wl_218 vdd gnd cell_6t
Xbit_r219_c105 bl_105 br_105 wl_219 vdd gnd cell_6t
Xbit_r220_c105 bl_105 br_105 wl_220 vdd gnd cell_6t
Xbit_r221_c105 bl_105 br_105 wl_221 vdd gnd cell_6t
Xbit_r222_c105 bl_105 br_105 wl_222 vdd gnd cell_6t
Xbit_r223_c105 bl_105 br_105 wl_223 vdd gnd cell_6t
Xbit_r224_c105 bl_105 br_105 wl_224 vdd gnd cell_6t
Xbit_r225_c105 bl_105 br_105 wl_225 vdd gnd cell_6t
Xbit_r226_c105 bl_105 br_105 wl_226 vdd gnd cell_6t
Xbit_r227_c105 bl_105 br_105 wl_227 vdd gnd cell_6t
Xbit_r228_c105 bl_105 br_105 wl_228 vdd gnd cell_6t
Xbit_r229_c105 bl_105 br_105 wl_229 vdd gnd cell_6t
Xbit_r230_c105 bl_105 br_105 wl_230 vdd gnd cell_6t
Xbit_r231_c105 bl_105 br_105 wl_231 vdd gnd cell_6t
Xbit_r232_c105 bl_105 br_105 wl_232 vdd gnd cell_6t
Xbit_r233_c105 bl_105 br_105 wl_233 vdd gnd cell_6t
Xbit_r234_c105 bl_105 br_105 wl_234 vdd gnd cell_6t
Xbit_r235_c105 bl_105 br_105 wl_235 vdd gnd cell_6t
Xbit_r236_c105 bl_105 br_105 wl_236 vdd gnd cell_6t
Xbit_r237_c105 bl_105 br_105 wl_237 vdd gnd cell_6t
Xbit_r238_c105 bl_105 br_105 wl_238 vdd gnd cell_6t
Xbit_r239_c105 bl_105 br_105 wl_239 vdd gnd cell_6t
Xbit_r240_c105 bl_105 br_105 wl_240 vdd gnd cell_6t
Xbit_r241_c105 bl_105 br_105 wl_241 vdd gnd cell_6t
Xbit_r242_c105 bl_105 br_105 wl_242 vdd gnd cell_6t
Xbit_r243_c105 bl_105 br_105 wl_243 vdd gnd cell_6t
Xbit_r244_c105 bl_105 br_105 wl_244 vdd gnd cell_6t
Xbit_r245_c105 bl_105 br_105 wl_245 vdd gnd cell_6t
Xbit_r246_c105 bl_105 br_105 wl_246 vdd gnd cell_6t
Xbit_r247_c105 bl_105 br_105 wl_247 vdd gnd cell_6t
Xbit_r248_c105 bl_105 br_105 wl_248 vdd gnd cell_6t
Xbit_r249_c105 bl_105 br_105 wl_249 vdd gnd cell_6t
Xbit_r250_c105 bl_105 br_105 wl_250 vdd gnd cell_6t
Xbit_r251_c105 bl_105 br_105 wl_251 vdd gnd cell_6t
Xbit_r252_c105 bl_105 br_105 wl_252 vdd gnd cell_6t
Xbit_r253_c105 bl_105 br_105 wl_253 vdd gnd cell_6t
Xbit_r254_c105 bl_105 br_105 wl_254 vdd gnd cell_6t
Xbit_r255_c105 bl_105 br_105 wl_255 vdd gnd cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd cell_6t
Xbit_r1_c106 bl_106 br_106 wl_1 vdd gnd cell_6t
Xbit_r2_c106 bl_106 br_106 wl_2 vdd gnd cell_6t
Xbit_r3_c106 bl_106 br_106 wl_3 vdd gnd cell_6t
Xbit_r4_c106 bl_106 br_106 wl_4 vdd gnd cell_6t
Xbit_r5_c106 bl_106 br_106 wl_5 vdd gnd cell_6t
Xbit_r6_c106 bl_106 br_106 wl_6 vdd gnd cell_6t
Xbit_r7_c106 bl_106 br_106 wl_7 vdd gnd cell_6t
Xbit_r8_c106 bl_106 br_106 wl_8 vdd gnd cell_6t
Xbit_r9_c106 bl_106 br_106 wl_9 vdd gnd cell_6t
Xbit_r10_c106 bl_106 br_106 wl_10 vdd gnd cell_6t
Xbit_r11_c106 bl_106 br_106 wl_11 vdd gnd cell_6t
Xbit_r12_c106 bl_106 br_106 wl_12 vdd gnd cell_6t
Xbit_r13_c106 bl_106 br_106 wl_13 vdd gnd cell_6t
Xbit_r14_c106 bl_106 br_106 wl_14 vdd gnd cell_6t
Xbit_r15_c106 bl_106 br_106 wl_15 vdd gnd cell_6t
Xbit_r16_c106 bl_106 br_106 wl_16 vdd gnd cell_6t
Xbit_r17_c106 bl_106 br_106 wl_17 vdd gnd cell_6t
Xbit_r18_c106 bl_106 br_106 wl_18 vdd gnd cell_6t
Xbit_r19_c106 bl_106 br_106 wl_19 vdd gnd cell_6t
Xbit_r20_c106 bl_106 br_106 wl_20 vdd gnd cell_6t
Xbit_r21_c106 bl_106 br_106 wl_21 vdd gnd cell_6t
Xbit_r22_c106 bl_106 br_106 wl_22 vdd gnd cell_6t
Xbit_r23_c106 bl_106 br_106 wl_23 vdd gnd cell_6t
Xbit_r24_c106 bl_106 br_106 wl_24 vdd gnd cell_6t
Xbit_r25_c106 bl_106 br_106 wl_25 vdd gnd cell_6t
Xbit_r26_c106 bl_106 br_106 wl_26 vdd gnd cell_6t
Xbit_r27_c106 bl_106 br_106 wl_27 vdd gnd cell_6t
Xbit_r28_c106 bl_106 br_106 wl_28 vdd gnd cell_6t
Xbit_r29_c106 bl_106 br_106 wl_29 vdd gnd cell_6t
Xbit_r30_c106 bl_106 br_106 wl_30 vdd gnd cell_6t
Xbit_r31_c106 bl_106 br_106 wl_31 vdd gnd cell_6t
Xbit_r32_c106 bl_106 br_106 wl_32 vdd gnd cell_6t
Xbit_r33_c106 bl_106 br_106 wl_33 vdd gnd cell_6t
Xbit_r34_c106 bl_106 br_106 wl_34 vdd gnd cell_6t
Xbit_r35_c106 bl_106 br_106 wl_35 vdd gnd cell_6t
Xbit_r36_c106 bl_106 br_106 wl_36 vdd gnd cell_6t
Xbit_r37_c106 bl_106 br_106 wl_37 vdd gnd cell_6t
Xbit_r38_c106 bl_106 br_106 wl_38 vdd gnd cell_6t
Xbit_r39_c106 bl_106 br_106 wl_39 vdd gnd cell_6t
Xbit_r40_c106 bl_106 br_106 wl_40 vdd gnd cell_6t
Xbit_r41_c106 bl_106 br_106 wl_41 vdd gnd cell_6t
Xbit_r42_c106 bl_106 br_106 wl_42 vdd gnd cell_6t
Xbit_r43_c106 bl_106 br_106 wl_43 vdd gnd cell_6t
Xbit_r44_c106 bl_106 br_106 wl_44 vdd gnd cell_6t
Xbit_r45_c106 bl_106 br_106 wl_45 vdd gnd cell_6t
Xbit_r46_c106 bl_106 br_106 wl_46 vdd gnd cell_6t
Xbit_r47_c106 bl_106 br_106 wl_47 vdd gnd cell_6t
Xbit_r48_c106 bl_106 br_106 wl_48 vdd gnd cell_6t
Xbit_r49_c106 bl_106 br_106 wl_49 vdd gnd cell_6t
Xbit_r50_c106 bl_106 br_106 wl_50 vdd gnd cell_6t
Xbit_r51_c106 bl_106 br_106 wl_51 vdd gnd cell_6t
Xbit_r52_c106 bl_106 br_106 wl_52 vdd gnd cell_6t
Xbit_r53_c106 bl_106 br_106 wl_53 vdd gnd cell_6t
Xbit_r54_c106 bl_106 br_106 wl_54 vdd gnd cell_6t
Xbit_r55_c106 bl_106 br_106 wl_55 vdd gnd cell_6t
Xbit_r56_c106 bl_106 br_106 wl_56 vdd gnd cell_6t
Xbit_r57_c106 bl_106 br_106 wl_57 vdd gnd cell_6t
Xbit_r58_c106 bl_106 br_106 wl_58 vdd gnd cell_6t
Xbit_r59_c106 bl_106 br_106 wl_59 vdd gnd cell_6t
Xbit_r60_c106 bl_106 br_106 wl_60 vdd gnd cell_6t
Xbit_r61_c106 bl_106 br_106 wl_61 vdd gnd cell_6t
Xbit_r62_c106 bl_106 br_106 wl_62 vdd gnd cell_6t
Xbit_r63_c106 bl_106 br_106 wl_63 vdd gnd cell_6t
Xbit_r64_c106 bl_106 br_106 wl_64 vdd gnd cell_6t
Xbit_r65_c106 bl_106 br_106 wl_65 vdd gnd cell_6t
Xbit_r66_c106 bl_106 br_106 wl_66 vdd gnd cell_6t
Xbit_r67_c106 bl_106 br_106 wl_67 vdd gnd cell_6t
Xbit_r68_c106 bl_106 br_106 wl_68 vdd gnd cell_6t
Xbit_r69_c106 bl_106 br_106 wl_69 vdd gnd cell_6t
Xbit_r70_c106 bl_106 br_106 wl_70 vdd gnd cell_6t
Xbit_r71_c106 bl_106 br_106 wl_71 vdd gnd cell_6t
Xbit_r72_c106 bl_106 br_106 wl_72 vdd gnd cell_6t
Xbit_r73_c106 bl_106 br_106 wl_73 vdd gnd cell_6t
Xbit_r74_c106 bl_106 br_106 wl_74 vdd gnd cell_6t
Xbit_r75_c106 bl_106 br_106 wl_75 vdd gnd cell_6t
Xbit_r76_c106 bl_106 br_106 wl_76 vdd gnd cell_6t
Xbit_r77_c106 bl_106 br_106 wl_77 vdd gnd cell_6t
Xbit_r78_c106 bl_106 br_106 wl_78 vdd gnd cell_6t
Xbit_r79_c106 bl_106 br_106 wl_79 vdd gnd cell_6t
Xbit_r80_c106 bl_106 br_106 wl_80 vdd gnd cell_6t
Xbit_r81_c106 bl_106 br_106 wl_81 vdd gnd cell_6t
Xbit_r82_c106 bl_106 br_106 wl_82 vdd gnd cell_6t
Xbit_r83_c106 bl_106 br_106 wl_83 vdd gnd cell_6t
Xbit_r84_c106 bl_106 br_106 wl_84 vdd gnd cell_6t
Xbit_r85_c106 bl_106 br_106 wl_85 vdd gnd cell_6t
Xbit_r86_c106 bl_106 br_106 wl_86 vdd gnd cell_6t
Xbit_r87_c106 bl_106 br_106 wl_87 vdd gnd cell_6t
Xbit_r88_c106 bl_106 br_106 wl_88 vdd gnd cell_6t
Xbit_r89_c106 bl_106 br_106 wl_89 vdd gnd cell_6t
Xbit_r90_c106 bl_106 br_106 wl_90 vdd gnd cell_6t
Xbit_r91_c106 bl_106 br_106 wl_91 vdd gnd cell_6t
Xbit_r92_c106 bl_106 br_106 wl_92 vdd gnd cell_6t
Xbit_r93_c106 bl_106 br_106 wl_93 vdd gnd cell_6t
Xbit_r94_c106 bl_106 br_106 wl_94 vdd gnd cell_6t
Xbit_r95_c106 bl_106 br_106 wl_95 vdd gnd cell_6t
Xbit_r96_c106 bl_106 br_106 wl_96 vdd gnd cell_6t
Xbit_r97_c106 bl_106 br_106 wl_97 vdd gnd cell_6t
Xbit_r98_c106 bl_106 br_106 wl_98 vdd gnd cell_6t
Xbit_r99_c106 bl_106 br_106 wl_99 vdd gnd cell_6t
Xbit_r100_c106 bl_106 br_106 wl_100 vdd gnd cell_6t
Xbit_r101_c106 bl_106 br_106 wl_101 vdd gnd cell_6t
Xbit_r102_c106 bl_106 br_106 wl_102 vdd gnd cell_6t
Xbit_r103_c106 bl_106 br_106 wl_103 vdd gnd cell_6t
Xbit_r104_c106 bl_106 br_106 wl_104 vdd gnd cell_6t
Xbit_r105_c106 bl_106 br_106 wl_105 vdd gnd cell_6t
Xbit_r106_c106 bl_106 br_106 wl_106 vdd gnd cell_6t
Xbit_r107_c106 bl_106 br_106 wl_107 vdd gnd cell_6t
Xbit_r108_c106 bl_106 br_106 wl_108 vdd gnd cell_6t
Xbit_r109_c106 bl_106 br_106 wl_109 vdd gnd cell_6t
Xbit_r110_c106 bl_106 br_106 wl_110 vdd gnd cell_6t
Xbit_r111_c106 bl_106 br_106 wl_111 vdd gnd cell_6t
Xbit_r112_c106 bl_106 br_106 wl_112 vdd gnd cell_6t
Xbit_r113_c106 bl_106 br_106 wl_113 vdd gnd cell_6t
Xbit_r114_c106 bl_106 br_106 wl_114 vdd gnd cell_6t
Xbit_r115_c106 bl_106 br_106 wl_115 vdd gnd cell_6t
Xbit_r116_c106 bl_106 br_106 wl_116 vdd gnd cell_6t
Xbit_r117_c106 bl_106 br_106 wl_117 vdd gnd cell_6t
Xbit_r118_c106 bl_106 br_106 wl_118 vdd gnd cell_6t
Xbit_r119_c106 bl_106 br_106 wl_119 vdd gnd cell_6t
Xbit_r120_c106 bl_106 br_106 wl_120 vdd gnd cell_6t
Xbit_r121_c106 bl_106 br_106 wl_121 vdd gnd cell_6t
Xbit_r122_c106 bl_106 br_106 wl_122 vdd gnd cell_6t
Xbit_r123_c106 bl_106 br_106 wl_123 vdd gnd cell_6t
Xbit_r124_c106 bl_106 br_106 wl_124 vdd gnd cell_6t
Xbit_r125_c106 bl_106 br_106 wl_125 vdd gnd cell_6t
Xbit_r126_c106 bl_106 br_106 wl_126 vdd gnd cell_6t
Xbit_r127_c106 bl_106 br_106 wl_127 vdd gnd cell_6t
Xbit_r128_c106 bl_106 br_106 wl_128 vdd gnd cell_6t
Xbit_r129_c106 bl_106 br_106 wl_129 vdd gnd cell_6t
Xbit_r130_c106 bl_106 br_106 wl_130 vdd gnd cell_6t
Xbit_r131_c106 bl_106 br_106 wl_131 vdd gnd cell_6t
Xbit_r132_c106 bl_106 br_106 wl_132 vdd gnd cell_6t
Xbit_r133_c106 bl_106 br_106 wl_133 vdd gnd cell_6t
Xbit_r134_c106 bl_106 br_106 wl_134 vdd gnd cell_6t
Xbit_r135_c106 bl_106 br_106 wl_135 vdd gnd cell_6t
Xbit_r136_c106 bl_106 br_106 wl_136 vdd gnd cell_6t
Xbit_r137_c106 bl_106 br_106 wl_137 vdd gnd cell_6t
Xbit_r138_c106 bl_106 br_106 wl_138 vdd gnd cell_6t
Xbit_r139_c106 bl_106 br_106 wl_139 vdd gnd cell_6t
Xbit_r140_c106 bl_106 br_106 wl_140 vdd gnd cell_6t
Xbit_r141_c106 bl_106 br_106 wl_141 vdd gnd cell_6t
Xbit_r142_c106 bl_106 br_106 wl_142 vdd gnd cell_6t
Xbit_r143_c106 bl_106 br_106 wl_143 vdd gnd cell_6t
Xbit_r144_c106 bl_106 br_106 wl_144 vdd gnd cell_6t
Xbit_r145_c106 bl_106 br_106 wl_145 vdd gnd cell_6t
Xbit_r146_c106 bl_106 br_106 wl_146 vdd gnd cell_6t
Xbit_r147_c106 bl_106 br_106 wl_147 vdd gnd cell_6t
Xbit_r148_c106 bl_106 br_106 wl_148 vdd gnd cell_6t
Xbit_r149_c106 bl_106 br_106 wl_149 vdd gnd cell_6t
Xbit_r150_c106 bl_106 br_106 wl_150 vdd gnd cell_6t
Xbit_r151_c106 bl_106 br_106 wl_151 vdd gnd cell_6t
Xbit_r152_c106 bl_106 br_106 wl_152 vdd gnd cell_6t
Xbit_r153_c106 bl_106 br_106 wl_153 vdd gnd cell_6t
Xbit_r154_c106 bl_106 br_106 wl_154 vdd gnd cell_6t
Xbit_r155_c106 bl_106 br_106 wl_155 vdd gnd cell_6t
Xbit_r156_c106 bl_106 br_106 wl_156 vdd gnd cell_6t
Xbit_r157_c106 bl_106 br_106 wl_157 vdd gnd cell_6t
Xbit_r158_c106 bl_106 br_106 wl_158 vdd gnd cell_6t
Xbit_r159_c106 bl_106 br_106 wl_159 vdd gnd cell_6t
Xbit_r160_c106 bl_106 br_106 wl_160 vdd gnd cell_6t
Xbit_r161_c106 bl_106 br_106 wl_161 vdd gnd cell_6t
Xbit_r162_c106 bl_106 br_106 wl_162 vdd gnd cell_6t
Xbit_r163_c106 bl_106 br_106 wl_163 vdd gnd cell_6t
Xbit_r164_c106 bl_106 br_106 wl_164 vdd gnd cell_6t
Xbit_r165_c106 bl_106 br_106 wl_165 vdd gnd cell_6t
Xbit_r166_c106 bl_106 br_106 wl_166 vdd gnd cell_6t
Xbit_r167_c106 bl_106 br_106 wl_167 vdd gnd cell_6t
Xbit_r168_c106 bl_106 br_106 wl_168 vdd gnd cell_6t
Xbit_r169_c106 bl_106 br_106 wl_169 vdd gnd cell_6t
Xbit_r170_c106 bl_106 br_106 wl_170 vdd gnd cell_6t
Xbit_r171_c106 bl_106 br_106 wl_171 vdd gnd cell_6t
Xbit_r172_c106 bl_106 br_106 wl_172 vdd gnd cell_6t
Xbit_r173_c106 bl_106 br_106 wl_173 vdd gnd cell_6t
Xbit_r174_c106 bl_106 br_106 wl_174 vdd gnd cell_6t
Xbit_r175_c106 bl_106 br_106 wl_175 vdd gnd cell_6t
Xbit_r176_c106 bl_106 br_106 wl_176 vdd gnd cell_6t
Xbit_r177_c106 bl_106 br_106 wl_177 vdd gnd cell_6t
Xbit_r178_c106 bl_106 br_106 wl_178 vdd gnd cell_6t
Xbit_r179_c106 bl_106 br_106 wl_179 vdd gnd cell_6t
Xbit_r180_c106 bl_106 br_106 wl_180 vdd gnd cell_6t
Xbit_r181_c106 bl_106 br_106 wl_181 vdd gnd cell_6t
Xbit_r182_c106 bl_106 br_106 wl_182 vdd gnd cell_6t
Xbit_r183_c106 bl_106 br_106 wl_183 vdd gnd cell_6t
Xbit_r184_c106 bl_106 br_106 wl_184 vdd gnd cell_6t
Xbit_r185_c106 bl_106 br_106 wl_185 vdd gnd cell_6t
Xbit_r186_c106 bl_106 br_106 wl_186 vdd gnd cell_6t
Xbit_r187_c106 bl_106 br_106 wl_187 vdd gnd cell_6t
Xbit_r188_c106 bl_106 br_106 wl_188 vdd gnd cell_6t
Xbit_r189_c106 bl_106 br_106 wl_189 vdd gnd cell_6t
Xbit_r190_c106 bl_106 br_106 wl_190 vdd gnd cell_6t
Xbit_r191_c106 bl_106 br_106 wl_191 vdd gnd cell_6t
Xbit_r192_c106 bl_106 br_106 wl_192 vdd gnd cell_6t
Xbit_r193_c106 bl_106 br_106 wl_193 vdd gnd cell_6t
Xbit_r194_c106 bl_106 br_106 wl_194 vdd gnd cell_6t
Xbit_r195_c106 bl_106 br_106 wl_195 vdd gnd cell_6t
Xbit_r196_c106 bl_106 br_106 wl_196 vdd gnd cell_6t
Xbit_r197_c106 bl_106 br_106 wl_197 vdd gnd cell_6t
Xbit_r198_c106 bl_106 br_106 wl_198 vdd gnd cell_6t
Xbit_r199_c106 bl_106 br_106 wl_199 vdd gnd cell_6t
Xbit_r200_c106 bl_106 br_106 wl_200 vdd gnd cell_6t
Xbit_r201_c106 bl_106 br_106 wl_201 vdd gnd cell_6t
Xbit_r202_c106 bl_106 br_106 wl_202 vdd gnd cell_6t
Xbit_r203_c106 bl_106 br_106 wl_203 vdd gnd cell_6t
Xbit_r204_c106 bl_106 br_106 wl_204 vdd gnd cell_6t
Xbit_r205_c106 bl_106 br_106 wl_205 vdd gnd cell_6t
Xbit_r206_c106 bl_106 br_106 wl_206 vdd gnd cell_6t
Xbit_r207_c106 bl_106 br_106 wl_207 vdd gnd cell_6t
Xbit_r208_c106 bl_106 br_106 wl_208 vdd gnd cell_6t
Xbit_r209_c106 bl_106 br_106 wl_209 vdd gnd cell_6t
Xbit_r210_c106 bl_106 br_106 wl_210 vdd gnd cell_6t
Xbit_r211_c106 bl_106 br_106 wl_211 vdd gnd cell_6t
Xbit_r212_c106 bl_106 br_106 wl_212 vdd gnd cell_6t
Xbit_r213_c106 bl_106 br_106 wl_213 vdd gnd cell_6t
Xbit_r214_c106 bl_106 br_106 wl_214 vdd gnd cell_6t
Xbit_r215_c106 bl_106 br_106 wl_215 vdd gnd cell_6t
Xbit_r216_c106 bl_106 br_106 wl_216 vdd gnd cell_6t
Xbit_r217_c106 bl_106 br_106 wl_217 vdd gnd cell_6t
Xbit_r218_c106 bl_106 br_106 wl_218 vdd gnd cell_6t
Xbit_r219_c106 bl_106 br_106 wl_219 vdd gnd cell_6t
Xbit_r220_c106 bl_106 br_106 wl_220 vdd gnd cell_6t
Xbit_r221_c106 bl_106 br_106 wl_221 vdd gnd cell_6t
Xbit_r222_c106 bl_106 br_106 wl_222 vdd gnd cell_6t
Xbit_r223_c106 bl_106 br_106 wl_223 vdd gnd cell_6t
Xbit_r224_c106 bl_106 br_106 wl_224 vdd gnd cell_6t
Xbit_r225_c106 bl_106 br_106 wl_225 vdd gnd cell_6t
Xbit_r226_c106 bl_106 br_106 wl_226 vdd gnd cell_6t
Xbit_r227_c106 bl_106 br_106 wl_227 vdd gnd cell_6t
Xbit_r228_c106 bl_106 br_106 wl_228 vdd gnd cell_6t
Xbit_r229_c106 bl_106 br_106 wl_229 vdd gnd cell_6t
Xbit_r230_c106 bl_106 br_106 wl_230 vdd gnd cell_6t
Xbit_r231_c106 bl_106 br_106 wl_231 vdd gnd cell_6t
Xbit_r232_c106 bl_106 br_106 wl_232 vdd gnd cell_6t
Xbit_r233_c106 bl_106 br_106 wl_233 vdd gnd cell_6t
Xbit_r234_c106 bl_106 br_106 wl_234 vdd gnd cell_6t
Xbit_r235_c106 bl_106 br_106 wl_235 vdd gnd cell_6t
Xbit_r236_c106 bl_106 br_106 wl_236 vdd gnd cell_6t
Xbit_r237_c106 bl_106 br_106 wl_237 vdd gnd cell_6t
Xbit_r238_c106 bl_106 br_106 wl_238 vdd gnd cell_6t
Xbit_r239_c106 bl_106 br_106 wl_239 vdd gnd cell_6t
Xbit_r240_c106 bl_106 br_106 wl_240 vdd gnd cell_6t
Xbit_r241_c106 bl_106 br_106 wl_241 vdd gnd cell_6t
Xbit_r242_c106 bl_106 br_106 wl_242 vdd gnd cell_6t
Xbit_r243_c106 bl_106 br_106 wl_243 vdd gnd cell_6t
Xbit_r244_c106 bl_106 br_106 wl_244 vdd gnd cell_6t
Xbit_r245_c106 bl_106 br_106 wl_245 vdd gnd cell_6t
Xbit_r246_c106 bl_106 br_106 wl_246 vdd gnd cell_6t
Xbit_r247_c106 bl_106 br_106 wl_247 vdd gnd cell_6t
Xbit_r248_c106 bl_106 br_106 wl_248 vdd gnd cell_6t
Xbit_r249_c106 bl_106 br_106 wl_249 vdd gnd cell_6t
Xbit_r250_c106 bl_106 br_106 wl_250 vdd gnd cell_6t
Xbit_r251_c106 bl_106 br_106 wl_251 vdd gnd cell_6t
Xbit_r252_c106 bl_106 br_106 wl_252 vdd gnd cell_6t
Xbit_r253_c106 bl_106 br_106 wl_253 vdd gnd cell_6t
Xbit_r254_c106 bl_106 br_106 wl_254 vdd gnd cell_6t
Xbit_r255_c106 bl_106 br_106 wl_255 vdd gnd cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd cell_6t
Xbit_r1_c107 bl_107 br_107 wl_1 vdd gnd cell_6t
Xbit_r2_c107 bl_107 br_107 wl_2 vdd gnd cell_6t
Xbit_r3_c107 bl_107 br_107 wl_3 vdd gnd cell_6t
Xbit_r4_c107 bl_107 br_107 wl_4 vdd gnd cell_6t
Xbit_r5_c107 bl_107 br_107 wl_5 vdd gnd cell_6t
Xbit_r6_c107 bl_107 br_107 wl_6 vdd gnd cell_6t
Xbit_r7_c107 bl_107 br_107 wl_7 vdd gnd cell_6t
Xbit_r8_c107 bl_107 br_107 wl_8 vdd gnd cell_6t
Xbit_r9_c107 bl_107 br_107 wl_9 vdd gnd cell_6t
Xbit_r10_c107 bl_107 br_107 wl_10 vdd gnd cell_6t
Xbit_r11_c107 bl_107 br_107 wl_11 vdd gnd cell_6t
Xbit_r12_c107 bl_107 br_107 wl_12 vdd gnd cell_6t
Xbit_r13_c107 bl_107 br_107 wl_13 vdd gnd cell_6t
Xbit_r14_c107 bl_107 br_107 wl_14 vdd gnd cell_6t
Xbit_r15_c107 bl_107 br_107 wl_15 vdd gnd cell_6t
Xbit_r16_c107 bl_107 br_107 wl_16 vdd gnd cell_6t
Xbit_r17_c107 bl_107 br_107 wl_17 vdd gnd cell_6t
Xbit_r18_c107 bl_107 br_107 wl_18 vdd gnd cell_6t
Xbit_r19_c107 bl_107 br_107 wl_19 vdd gnd cell_6t
Xbit_r20_c107 bl_107 br_107 wl_20 vdd gnd cell_6t
Xbit_r21_c107 bl_107 br_107 wl_21 vdd gnd cell_6t
Xbit_r22_c107 bl_107 br_107 wl_22 vdd gnd cell_6t
Xbit_r23_c107 bl_107 br_107 wl_23 vdd gnd cell_6t
Xbit_r24_c107 bl_107 br_107 wl_24 vdd gnd cell_6t
Xbit_r25_c107 bl_107 br_107 wl_25 vdd gnd cell_6t
Xbit_r26_c107 bl_107 br_107 wl_26 vdd gnd cell_6t
Xbit_r27_c107 bl_107 br_107 wl_27 vdd gnd cell_6t
Xbit_r28_c107 bl_107 br_107 wl_28 vdd gnd cell_6t
Xbit_r29_c107 bl_107 br_107 wl_29 vdd gnd cell_6t
Xbit_r30_c107 bl_107 br_107 wl_30 vdd gnd cell_6t
Xbit_r31_c107 bl_107 br_107 wl_31 vdd gnd cell_6t
Xbit_r32_c107 bl_107 br_107 wl_32 vdd gnd cell_6t
Xbit_r33_c107 bl_107 br_107 wl_33 vdd gnd cell_6t
Xbit_r34_c107 bl_107 br_107 wl_34 vdd gnd cell_6t
Xbit_r35_c107 bl_107 br_107 wl_35 vdd gnd cell_6t
Xbit_r36_c107 bl_107 br_107 wl_36 vdd gnd cell_6t
Xbit_r37_c107 bl_107 br_107 wl_37 vdd gnd cell_6t
Xbit_r38_c107 bl_107 br_107 wl_38 vdd gnd cell_6t
Xbit_r39_c107 bl_107 br_107 wl_39 vdd gnd cell_6t
Xbit_r40_c107 bl_107 br_107 wl_40 vdd gnd cell_6t
Xbit_r41_c107 bl_107 br_107 wl_41 vdd gnd cell_6t
Xbit_r42_c107 bl_107 br_107 wl_42 vdd gnd cell_6t
Xbit_r43_c107 bl_107 br_107 wl_43 vdd gnd cell_6t
Xbit_r44_c107 bl_107 br_107 wl_44 vdd gnd cell_6t
Xbit_r45_c107 bl_107 br_107 wl_45 vdd gnd cell_6t
Xbit_r46_c107 bl_107 br_107 wl_46 vdd gnd cell_6t
Xbit_r47_c107 bl_107 br_107 wl_47 vdd gnd cell_6t
Xbit_r48_c107 bl_107 br_107 wl_48 vdd gnd cell_6t
Xbit_r49_c107 bl_107 br_107 wl_49 vdd gnd cell_6t
Xbit_r50_c107 bl_107 br_107 wl_50 vdd gnd cell_6t
Xbit_r51_c107 bl_107 br_107 wl_51 vdd gnd cell_6t
Xbit_r52_c107 bl_107 br_107 wl_52 vdd gnd cell_6t
Xbit_r53_c107 bl_107 br_107 wl_53 vdd gnd cell_6t
Xbit_r54_c107 bl_107 br_107 wl_54 vdd gnd cell_6t
Xbit_r55_c107 bl_107 br_107 wl_55 vdd gnd cell_6t
Xbit_r56_c107 bl_107 br_107 wl_56 vdd gnd cell_6t
Xbit_r57_c107 bl_107 br_107 wl_57 vdd gnd cell_6t
Xbit_r58_c107 bl_107 br_107 wl_58 vdd gnd cell_6t
Xbit_r59_c107 bl_107 br_107 wl_59 vdd gnd cell_6t
Xbit_r60_c107 bl_107 br_107 wl_60 vdd gnd cell_6t
Xbit_r61_c107 bl_107 br_107 wl_61 vdd gnd cell_6t
Xbit_r62_c107 bl_107 br_107 wl_62 vdd gnd cell_6t
Xbit_r63_c107 bl_107 br_107 wl_63 vdd gnd cell_6t
Xbit_r64_c107 bl_107 br_107 wl_64 vdd gnd cell_6t
Xbit_r65_c107 bl_107 br_107 wl_65 vdd gnd cell_6t
Xbit_r66_c107 bl_107 br_107 wl_66 vdd gnd cell_6t
Xbit_r67_c107 bl_107 br_107 wl_67 vdd gnd cell_6t
Xbit_r68_c107 bl_107 br_107 wl_68 vdd gnd cell_6t
Xbit_r69_c107 bl_107 br_107 wl_69 vdd gnd cell_6t
Xbit_r70_c107 bl_107 br_107 wl_70 vdd gnd cell_6t
Xbit_r71_c107 bl_107 br_107 wl_71 vdd gnd cell_6t
Xbit_r72_c107 bl_107 br_107 wl_72 vdd gnd cell_6t
Xbit_r73_c107 bl_107 br_107 wl_73 vdd gnd cell_6t
Xbit_r74_c107 bl_107 br_107 wl_74 vdd gnd cell_6t
Xbit_r75_c107 bl_107 br_107 wl_75 vdd gnd cell_6t
Xbit_r76_c107 bl_107 br_107 wl_76 vdd gnd cell_6t
Xbit_r77_c107 bl_107 br_107 wl_77 vdd gnd cell_6t
Xbit_r78_c107 bl_107 br_107 wl_78 vdd gnd cell_6t
Xbit_r79_c107 bl_107 br_107 wl_79 vdd gnd cell_6t
Xbit_r80_c107 bl_107 br_107 wl_80 vdd gnd cell_6t
Xbit_r81_c107 bl_107 br_107 wl_81 vdd gnd cell_6t
Xbit_r82_c107 bl_107 br_107 wl_82 vdd gnd cell_6t
Xbit_r83_c107 bl_107 br_107 wl_83 vdd gnd cell_6t
Xbit_r84_c107 bl_107 br_107 wl_84 vdd gnd cell_6t
Xbit_r85_c107 bl_107 br_107 wl_85 vdd gnd cell_6t
Xbit_r86_c107 bl_107 br_107 wl_86 vdd gnd cell_6t
Xbit_r87_c107 bl_107 br_107 wl_87 vdd gnd cell_6t
Xbit_r88_c107 bl_107 br_107 wl_88 vdd gnd cell_6t
Xbit_r89_c107 bl_107 br_107 wl_89 vdd gnd cell_6t
Xbit_r90_c107 bl_107 br_107 wl_90 vdd gnd cell_6t
Xbit_r91_c107 bl_107 br_107 wl_91 vdd gnd cell_6t
Xbit_r92_c107 bl_107 br_107 wl_92 vdd gnd cell_6t
Xbit_r93_c107 bl_107 br_107 wl_93 vdd gnd cell_6t
Xbit_r94_c107 bl_107 br_107 wl_94 vdd gnd cell_6t
Xbit_r95_c107 bl_107 br_107 wl_95 vdd gnd cell_6t
Xbit_r96_c107 bl_107 br_107 wl_96 vdd gnd cell_6t
Xbit_r97_c107 bl_107 br_107 wl_97 vdd gnd cell_6t
Xbit_r98_c107 bl_107 br_107 wl_98 vdd gnd cell_6t
Xbit_r99_c107 bl_107 br_107 wl_99 vdd gnd cell_6t
Xbit_r100_c107 bl_107 br_107 wl_100 vdd gnd cell_6t
Xbit_r101_c107 bl_107 br_107 wl_101 vdd gnd cell_6t
Xbit_r102_c107 bl_107 br_107 wl_102 vdd gnd cell_6t
Xbit_r103_c107 bl_107 br_107 wl_103 vdd gnd cell_6t
Xbit_r104_c107 bl_107 br_107 wl_104 vdd gnd cell_6t
Xbit_r105_c107 bl_107 br_107 wl_105 vdd gnd cell_6t
Xbit_r106_c107 bl_107 br_107 wl_106 vdd gnd cell_6t
Xbit_r107_c107 bl_107 br_107 wl_107 vdd gnd cell_6t
Xbit_r108_c107 bl_107 br_107 wl_108 vdd gnd cell_6t
Xbit_r109_c107 bl_107 br_107 wl_109 vdd gnd cell_6t
Xbit_r110_c107 bl_107 br_107 wl_110 vdd gnd cell_6t
Xbit_r111_c107 bl_107 br_107 wl_111 vdd gnd cell_6t
Xbit_r112_c107 bl_107 br_107 wl_112 vdd gnd cell_6t
Xbit_r113_c107 bl_107 br_107 wl_113 vdd gnd cell_6t
Xbit_r114_c107 bl_107 br_107 wl_114 vdd gnd cell_6t
Xbit_r115_c107 bl_107 br_107 wl_115 vdd gnd cell_6t
Xbit_r116_c107 bl_107 br_107 wl_116 vdd gnd cell_6t
Xbit_r117_c107 bl_107 br_107 wl_117 vdd gnd cell_6t
Xbit_r118_c107 bl_107 br_107 wl_118 vdd gnd cell_6t
Xbit_r119_c107 bl_107 br_107 wl_119 vdd gnd cell_6t
Xbit_r120_c107 bl_107 br_107 wl_120 vdd gnd cell_6t
Xbit_r121_c107 bl_107 br_107 wl_121 vdd gnd cell_6t
Xbit_r122_c107 bl_107 br_107 wl_122 vdd gnd cell_6t
Xbit_r123_c107 bl_107 br_107 wl_123 vdd gnd cell_6t
Xbit_r124_c107 bl_107 br_107 wl_124 vdd gnd cell_6t
Xbit_r125_c107 bl_107 br_107 wl_125 vdd gnd cell_6t
Xbit_r126_c107 bl_107 br_107 wl_126 vdd gnd cell_6t
Xbit_r127_c107 bl_107 br_107 wl_127 vdd gnd cell_6t
Xbit_r128_c107 bl_107 br_107 wl_128 vdd gnd cell_6t
Xbit_r129_c107 bl_107 br_107 wl_129 vdd gnd cell_6t
Xbit_r130_c107 bl_107 br_107 wl_130 vdd gnd cell_6t
Xbit_r131_c107 bl_107 br_107 wl_131 vdd gnd cell_6t
Xbit_r132_c107 bl_107 br_107 wl_132 vdd gnd cell_6t
Xbit_r133_c107 bl_107 br_107 wl_133 vdd gnd cell_6t
Xbit_r134_c107 bl_107 br_107 wl_134 vdd gnd cell_6t
Xbit_r135_c107 bl_107 br_107 wl_135 vdd gnd cell_6t
Xbit_r136_c107 bl_107 br_107 wl_136 vdd gnd cell_6t
Xbit_r137_c107 bl_107 br_107 wl_137 vdd gnd cell_6t
Xbit_r138_c107 bl_107 br_107 wl_138 vdd gnd cell_6t
Xbit_r139_c107 bl_107 br_107 wl_139 vdd gnd cell_6t
Xbit_r140_c107 bl_107 br_107 wl_140 vdd gnd cell_6t
Xbit_r141_c107 bl_107 br_107 wl_141 vdd gnd cell_6t
Xbit_r142_c107 bl_107 br_107 wl_142 vdd gnd cell_6t
Xbit_r143_c107 bl_107 br_107 wl_143 vdd gnd cell_6t
Xbit_r144_c107 bl_107 br_107 wl_144 vdd gnd cell_6t
Xbit_r145_c107 bl_107 br_107 wl_145 vdd gnd cell_6t
Xbit_r146_c107 bl_107 br_107 wl_146 vdd gnd cell_6t
Xbit_r147_c107 bl_107 br_107 wl_147 vdd gnd cell_6t
Xbit_r148_c107 bl_107 br_107 wl_148 vdd gnd cell_6t
Xbit_r149_c107 bl_107 br_107 wl_149 vdd gnd cell_6t
Xbit_r150_c107 bl_107 br_107 wl_150 vdd gnd cell_6t
Xbit_r151_c107 bl_107 br_107 wl_151 vdd gnd cell_6t
Xbit_r152_c107 bl_107 br_107 wl_152 vdd gnd cell_6t
Xbit_r153_c107 bl_107 br_107 wl_153 vdd gnd cell_6t
Xbit_r154_c107 bl_107 br_107 wl_154 vdd gnd cell_6t
Xbit_r155_c107 bl_107 br_107 wl_155 vdd gnd cell_6t
Xbit_r156_c107 bl_107 br_107 wl_156 vdd gnd cell_6t
Xbit_r157_c107 bl_107 br_107 wl_157 vdd gnd cell_6t
Xbit_r158_c107 bl_107 br_107 wl_158 vdd gnd cell_6t
Xbit_r159_c107 bl_107 br_107 wl_159 vdd gnd cell_6t
Xbit_r160_c107 bl_107 br_107 wl_160 vdd gnd cell_6t
Xbit_r161_c107 bl_107 br_107 wl_161 vdd gnd cell_6t
Xbit_r162_c107 bl_107 br_107 wl_162 vdd gnd cell_6t
Xbit_r163_c107 bl_107 br_107 wl_163 vdd gnd cell_6t
Xbit_r164_c107 bl_107 br_107 wl_164 vdd gnd cell_6t
Xbit_r165_c107 bl_107 br_107 wl_165 vdd gnd cell_6t
Xbit_r166_c107 bl_107 br_107 wl_166 vdd gnd cell_6t
Xbit_r167_c107 bl_107 br_107 wl_167 vdd gnd cell_6t
Xbit_r168_c107 bl_107 br_107 wl_168 vdd gnd cell_6t
Xbit_r169_c107 bl_107 br_107 wl_169 vdd gnd cell_6t
Xbit_r170_c107 bl_107 br_107 wl_170 vdd gnd cell_6t
Xbit_r171_c107 bl_107 br_107 wl_171 vdd gnd cell_6t
Xbit_r172_c107 bl_107 br_107 wl_172 vdd gnd cell_6t
Xbit_r173_c107 bl_107 br_107 wl_173 vdd gnd cell_6t
Xbit_r174_c107 bl_107 br_107 wl_174 vdd gnd cell_6t
Xbit_r175_c107 bl_107 br_107 wl_175 vdd gnd cell_6t
Xbit_r176_c107 bl_107 br_107 wl_176 vdd gnd cell_6t
Xbit_r177_c107 bl_107 br_107 wl_177 vdd gnd cell_6t
Xbit_r178_c107 bl_107 br_107 wl_178 vdd gnd cell_6t
Xbit_r179_c107 bl_107 br_107 wl_179 vdd gnd cell_6t
Xbit_r180_c107 bl_107 br_107 wl_180 vdd gnd cell_6t
Xbit_r181_c107 bl_107 br_107 wl_181 vdd gnd cell_6t
Xbit_r182_c107 bl_107 br_107 wl_182 vdd gnd cell_6t
Xbit_r183_c107 bl_107 br_107 wl_183 vdd gnd cell_6t
Xbit_r184_c107 bl_107 br_107 wl_184 vdd gnd cell_6t
Xbit_r185_c107 bl_107 br_107 wl_185 vdd gnd cell_6t
Xbit_r186_c107 bl_107 br_107 wl_186 vdd gnd cell_6t
Xbit_r187_c107 bl_107 br_107 wl_187 vdd gnd cell_6t
Xbit_r188_c107 bl_107 br_107 wl_188 vdd gnd cell_6t
Xbit_r189_c107 bl_107 br_107 wl_189 vdd gnd cell_6t
Xbit_r190_c107 bl_107 br_107 wl_190 vdd gnd cell_6t
Xbit_r191_c107 bl_107 br_107 wl_191 vdd gnd cell_6t
Xbit_r192_c107 bl_107 br_107 wl_192 vdd gnd cell_6t
Xbit_r193_c107 bl_107 br_107 wl_193 vdd gnd cell_6t
Xbit_r194_c107 bl_107 br_107 wl_194 vdd gnd cell_6t
Xbit_r195_c107 bl_107 br_107 wl_195 vdd gnd cell_6t
Xbit_r196_c107 bl_107 br_107 wl_196 vdd gnd cell_6t
Xbit_r197_c107 bl_107 br_107 wl_197 vdd gnd cell_6t
Xbit_r198_c107 bl_107 br_107 wl_198 vdd gnd cell_6t
Xbit_r199_c107 bl_107 br_107 wl_199 vdd gnd cell_6t
Xbit_r200_c107 bl_107 br_107 wl_200 vdd gnd cell_6t
Xbit_r201_c107 bl_107 br_107 wl_201 vdd gnd cell_6t
Xbit_r202_c107 bl_107 br_107 wl_202 vdd gnd cell_6t
Xbit_r203_c107 bl_107 br_107 wl_203 vdd gnd cell_6t
Xbit_r204_c107 bl_107 br_107 wl_204 vdd gnd cell_6t
Xbit_r205_c107 bl_107 br_107 wl_205 vdd gnd cell_6t
Xbit_r206_c107 bl_107 br_107 wl_206 vdd gnd cell_6t
Xbit_r207_c107 bl_107 br_107 wl_207 vdd gnd cell_6t
Xbit_r208_c107 bl_107 br_107 wl_208 vdd gnd cell_6t
Xbit_r209_c107 bl_107 br_107 wl_209 vdd gnd cell_6t
Xbit_r210_c107 bl_107 br_107 wl_210 vdd gnd cell_6t
Xbit_r211_c107 bl_107 br_107 wl_211 vdd gnd cell_6t
Xbit_r212_c107 bl_107 br_107 wl_212 vdd gnd cell_6t
Xbit_r213_c107 bl_107 br_107 wl_213 vdd gnd cell_6t
Xbit_r214_c107 bl_107 br_107 wl_214 vdd gnd cell_6t
Xbit_r215_c107 bl_107 br_107 wl_215 vdd gnd cell_6t
Xbit_r216_c107 bl_107 br_107 wl_216 vdd gnd cell_6t
Xbit_r217_c107 bl_107 br_107 wl_217 vdd gnd cell_6t
Xbit_r218_c107 bl_107 br_107 wl_218 vdd gnd cell_6t
Xbit_r219_c107 bl_107 br_107 wl_219 vdd gnd cell_6t
Xbit_r220_c107 bl_107 br_107 wl_220 vdd gnd cell_6t
Xbit_r221_c107 bl_107 br_107 wl_221 vdd gnd cell_6t
Xbit_r222_c107 bl_107 br_107 wl_222 vdd gnd cell_6t
Xbit_r223_c107 bl_107 br_107 wl_223 vdd gnd cell_6t
Xbit_r224_c107 bl_107 br_107 wl_224 vdd gnd cell_6t
Xbit_r225_c107 bl_107 br_107 wl_225 vdd gnd cell_6t
Xbit_r226_c107 bl_107 br_107 wl_226 vdd gnd cell_6t
Xbit_r227_c107 bl_107 br_107 wl_227 vdd gnd cell_6t
Xbit_r228_c107 bl_107 br_107 wl_228 vdd gnd cell_6t
Xbit_r229_c107 bl_107 br_107 wl_229 vdd gnd cell_6t
Xbit_r230_c107 bl_107 br_107 wl_230 vdd gnd cell_6t
Xbit_r231_c107 bl_107 br_107 wl_231 vdd gnd cell_6t
Xbit_r232_c107 bl_107 br_107 wl_232 vdd gnd cell_6t
Xbit_r233_c107 bl_107 br_107 wl_233 vdd gnd cell_6t
Xbit_r234_c107 bl_107 br_107 wl_234 vdd gnd cell_6t
Xbit_r235_c107 bl_107 br_107 wl_235 vdd gnd cell_6t
Xbit_r236_c107 bl_107 br_107 wl_236 vdd gnd cell_6t
Xbit_r237_c107 bl_107 br_107 wl_237 vdd gnd cell_6t
Xbit_r238_c107 bl_107 br_107 wl_238 vdd gnd cell_6t
Xbit_r239_c107 bl_107 br_107 wl_239 vdd gnd cell_6t
Xbit_r240_c107 bl_107 br_107 wl_240 vdd gnd cell_6t
Xbit_r241_c107 bl_107 br_107 wl_241 vdd gnd cell_6t
Xbit_r242_c107 bl_107 br_107 wl_242 vdd gnd cell_6t
Xbit_r243_c107 bl_107 br_107 wl_243 vdd gnd cell_6t
Xbit_r244_c107 bl_107 br_107 wl_244 vdd gnd cell_6t
Xbit_r245_c107 bl_107 br_107 wl_245 vdd gnd cell_6t
Xbit_r246_c107 bl_107 br_107 wl_246 vdd gnd cell_6t
Xbit_r247_c107 bl_107 br_107 wl_247 vdd gnd cell_6t
Xbit_r248_c107 bl_107 br_107 wl_248 vdd gnd cell_6t
Xbit_r249_c107 bl_107 br_107 wl_249 vdd gnd cell_6t
Xbit_r250_c107 bl_107 br_107 wl_250 vdd gnd cell_6t
Xbit_r251_c107 bl_107 br_107 wl_251 vdd gnd cell_6t
Xbit_r252_c107 bl_107 br_107 wl_252 vdd gnd cell_6t
Xbit_r253_c107 bl_107 br_107 wl_253 vdd gnd cell_6t
Xbit_r254_c107 bl_107 br_107 wl_254 vdd gnd cell_6t
Xbit_r255_c107 bl_107 br_107 wl_255 vdd gnd cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd cell_6t
Xbit_r1_c108 bl_108 br_108 wl_1 vdd gnd cell_6t
Xbit_r2_c108 bl_108 br_108 wl_2 vdd gnd cell_6t
Xbit_r3_c108 bl_108 br_108 wl_3 vdd gnd cell_6t
Xbit_r4_c108 bl_108 br_108 wl_4 vdd gnd cell_6t
Xbit_r5_c108 bl_108 br_108 wl_5 vdd gnd cell_6t
Xbit_r6_c108 bl_108 br_108 wl_6 vdd gnd cell_6t
Xbit_r7_c108 bl_108 br_108 wl_7 vdd gnd cell_6t
Xbit_r8_c108 bl_108 br_108 wl_8 vdd gnd cell_6t
Xbit_r9_c108 bl_108 br_108 wl_9 vdd gnd cell_6t
Xbit_r10_c108 bl_108 br_108 wl_10 vdd gnd cell_6t
Xbit_r11_c108 bl_108 br_108 wl_11 vdd gnd cell_6t
Xbit_r12_c108 bl_108 br_108 wl_12 vdd gnd cell_6t
Xbit_r13_c108 bl_108 br_108 wl_13 vdd gnd cell_6t
Xbit_r14_c108 bl_108 br_108 wl_14 vdd gnd cell_6t
Xbit_r15_c108 bl_108 br_108 wl_15 vdd gnd cell_6t
Xbit_r16_c108 bl_108 br_108 wl_16 vdd gnd cell_6t
Xbit_r17_c108 bl_108 br_108 wl_17 vdd gnd cell_6t
Xbit_r18_c108 bl_108 br_108 wl_18 vdd gnd cell_6t
Xbit_r19_c108 bl_108 br_108 wl_19 vdd gnd cell_6t
Xbit_r20_c108 bl_108 br_108 wl_20 vdd gnd cell_6t
Xbit_r21_c108 bl_108 br_108 wl_21 vdd gnd cell_6t
Xbit_r22_c108 bl_108 br_108 wl_22 vdd gnd cell_6t
Xbit_r23_c108 bl_108 br_108 wl_23 vdd gnd cell_6t
Xbit_r24_c108 bl_108 br_108 wl_24 vdd gnd cell_6t
Xbit_r25_c108 bl_108 br_108 wl_25 vdd gnd cell_6t
Xbit_r26_c108 bl_108 br_108 wl_26 vdd gnd cell_6t
Xbit_r27_c108 bl_108 br_108 wl_27 vdd gnd cell_6t
Xbit_r28_c108 bl_108 br_108 wl_28 vdd gnd cell_6t
Xbit_r29_c108 bl_108 br_108 wl_29 vdd gnd cell_6t
Xbit_r30_c108 bl_108 br_108 wl_30 vdd gnd cell_6t
Xbit_r31_c108 bl_108 br_108 wl_31 vdd gnd cell_6t
Xbit_r32_c108 bl_108 br_108 wl_32 vdd gnd cell_6t
Xbit_r33_c108 bl_108 br_108 wl_33 vdd gnd cell_6t
Xbit_r34_c108 bl_108 br_108 wl_34 vdd gnd cell_6t
Xbit_r35_c108 bl_108 br_108 wl_35 vdd gnd cell_6t
Xbit_r36_c108 bl_108 br_108 wl_36 vdd gnd cell_6t
Xbit_r37_c108 bl_108 br_108 wl_37 vdd gnd cell_6t
Xbit_r38_c108 bl_108 br_108 wl_38 vdd gnd cell_6t
Xbit_r39_c108 bl_108 br_108 wl_39 vdd gnd cell_6t
Xbit_r40_c108 bl_108 br_108 wl_40 vdd gnd cell_6t
Xbit_r41_c108 bl_108 br_108 wl_41 vdd gnd cell_6t
Xbit_r42_c108 bl_108 br_108 wl_42 vdd gnd cell_6t
Xbit_r43_c108 bl_108 br_108 wl_43 vdd gnd cell_6t
Xbit_r44_c108 bl_108 br_108 wl_44 vdd gnd cell_6t
Xbit_r45_c108 bl_108 br_108 wl_45 vdd gnd cell_6t
Xbit_r46_c108 bl_108 br_108 wl_46 vdd gnd cell_6t
Xbit_r47_c108 bl_108 br_108 wl_47 vdd gnd cell_6t
Xbit_r48_c108 bl_108 br_108 wl_48 vdd gnd cell_6t
Xbit_r49_c108 bl_108 br_108 wl_49 vdd gnd cell_6t
Xbit_r50_c108 bl_108 br_108 wl_50 vdd gnd cell_6t
Xbit_r51_c108 bl_108 br_108 wl_51 vdd gnd cell_6t
Xbit_r52_c108 bl_108 br_108 wl_52 vdd gnd cell_6t
Xbit_r53_c108 bl_108 br_108 wl_53 vdd gnd cell_6t
Xbit_r54_c108 bl_108 br_108 wl_54 vdd gnd cell_6t
Xbit_r55_c108 bl_108 br_108 wl_55 vdd gnd cell_6t
Xbit_r56_c108 bl_108 br_108 wl_56 vdd gnd cell_6t
Xbit_r57_c108 bl_108 br_108 wl_57 vdd gnd cell_6t
Xbit_r58_c108 bl_108 br_108 wl_58 vdd gnd cell_6t
Xbit_r59_c108 bl_108 br_108 wl_59 vdd gnd cell_6t
Xbit_r60_c108 bl_108 br_108 wl_60 vdd gnd cell_6t
Xbit_r61_c108 bl_108 br_108 wl_61 vdd gnd cell_6t
Xbit_r62_c108 bl_108 br_108 wl_62 vdd gnd cell_6t
Xbit_r63_c108 bl_108 br_108 wl_63 vdd gnd cell_6t
Xbit_r64_c108 bl_108 br_108 wl_64 vdd gnd cell_6t
Xbit_r65_c108 bl_108 br_108 wl_65 vdd gnd cell_6t
Xbit_r66_c108 bl_108 br_108 wl_66 vdd gnd cell_6t
Xbit_r67_c108 bl_108 br_108 wl_67 vdd gnd cell_6t
Xbit_r68_c108 bl_108 br_108 wl_68 vdd gnd cell_6t
Xbit_r69_c108 bl_108 br_108 wl_69 vdd gnd cell_6t
Xbit_r70_c108 bl_108 br_108 wl_70 vdd gnd cell_6t
Xbit_r71_c108 bl_108 br_108 wl_71 vdd gnd cell_6t
Xbit_r72_c108 bl_108 br_108 wl_72 vdd gnd cell_6t
Xbit_r73_c108 bl_108 br_108 wl_73 vdd gnd cell_6t
Xbit_r74_c108 bl_108 br_108 wl_74 vdd gnd cell_6t
Xbit_r75_c108 bl_108 br_108 wl_75 vdd gnd cell_6t
Xbit_r76_c108 bl_108 br_108 wl_76 vdd gnd cell_6t
Xbit_r77_c108 bl_108 br_108 wl_77 vdd gnd cell_6t
Xbit_r78_c108 bl_108 br_108 wl_78 vdd gnd cell_6t
Xbit_r79_c108 bl_108 br_108 wl_79 vdd gnd cell_6t
Xbit_r80_c108 bl_108 br_108 wl_80 vdd gnd cell_6t
Xbit_r81_c108 bl_108 br_108 wl_81 vdd gnd cell_6t
Xbit_r82_c108 bl_108 br_108 wl_82 vdd gnd cell_6t
Xbit_r83_c108 bl_108 br_108 wl_83 vdd gnd cell_6t
Xbit_r84_c108 bl_108 br_108 wl_84 vdd gnd cell_6t
Xbit_r85_c108 bl_108 br_108 wl_85 vdd gnd cell_6t
Xbit_r86_c108 bl_108 br_108 wl_86 vdd gnd cell_6t
Xbit_r87_c108 bl_108 br_108 wl_87 vdd gnd cell_6t
Xbit_r88_c108 bl_108 br_108 wl_88 vdd gnd cell_6t
Xbit_r89_c108 bl_108 br_108 wl_89 vdd gnd cell_6t
Xbit_r90_c108 bl_108 br_108 wl_90 vdd gnd cell_6t
Xbit_r91_c108 bl_108 br_108 wl_91 vdd gnd cell_6t
Xbit_r92_c108 bl_108 br_108 wl_92 vdd gnd cell_6t
Xbit_r93_c108 bl_108 br_108 wl_93 vdd gnd cell_6t
Xbit_r94_c108 bl_108 br_108 wl_94 vdd gnd cell_6t
Xbit_r95_c108 bl_108 br_108 wl_95 vdd gnd cell_6t
Xbit_r96_c108 bl_108 br_108 wl_96 vdd gnd cell_6t
Xbit_r97_c108 bl_108 br_108 wl_97 vdd gnd cell_6t
Xbit_r98_c108 bl_108 br_108 wl_98 vdd gnd cell_6t
Xbit_r99_c108 bl_108 br_108 wl_99 vdd gnd cell_6t
Xbit_r100_c108 bl_108 br_108 wl_100 vdd gnd cell_6t
Xbit_r101_c108 bl_108 br_108 wl_101 vdd gnd cell_6t
Xbit_r102_c108 bl_108 br_108 wl_102 vdd gnd cell_6t
Xbit_r103_c108 bl_108 br_108 wl_103 vdd gnd cell_6t
Xbit_r104_c108 bl_108 br_108 wl_104 vdd gnd cell_6t
Xbit_r105_c108 bl_108 br_108 wl_105 vdd gnd cell_6t
Xbit_r106_c108 bl_108 br_108 wl_106 vdd gnd cell_6t
Xbit_r107_c108 bl_108 br_108 wl_107 vdd gnd cell_6t
Xbit_r108_c108 bl_108 br_108 wl_108 vdd gnd cell_6t
Xbit_r109_c108 bl_108 br_108 wl_109 vdd gnd cell_6t
Xbit_r110_c108 bl_108 br_108 wl_110 vdd gnd cell_6t
Xbit_r111_c108 bl_108 br_108 wl_111 vdd gnd cell_6t
Xbit_r112_c108 bl_108 br_108 wl_112 vdd gnd cell_6t
Xbit_r113_c108 bl_108 br_108 wl_113 vdd gnd cell_6t
Xbit_r114_c108 bl_108 br_108 wl_114 vdd gnd cell_6t
Xbit_r115_c108 bl_108 br_108 wl_115 vdd gnd cell_6t
Xbit_r116_c108 bl_108 br_108 wl_116 vdd gnd cell_6t
Xbit_r117_c108 bl_108 br_108 wl_117 vdd gnd cell_6t
Xbit_r118_c108 bl_108 br_108 wl_118 vdd gnd cell_6t
Xbit_r119_c108 bl_108 br_108 wl_119 vdd gnd cell_6t
Xbit_r120_c108 bl_108 br_108 wl_120 vdd gnd cell_6t
Xbit_r121_c108 bl_108 br_108 wl_121 vdd gnd cell_6t
Xbit_r122_c108 bl_108 br_108 wl_122 vdd gnd cell_6t
Xbit_r123_c108 bl_108 br_108 wl_123 vdd gnd cell_6t
Xbit_r124_c108 bl_108 br_108 wl_124 vdd gnd cell_6t
Xbit_r125_c108 bl_108 br_108 wl_125 vdd gnd cell_6t
Xbit_r126_c108 bl_108 br_108 wl_126 vdd gnd cell_6t
Xbit_r127_c108 bl_108 br_108 wl_127 vdd gnd cell_6t
Xbit_r128_c108 bl_108 br_108 wl_128 vdd gnd cell_6t
Xbit_r129_c108 bl_108 br_108 wl_129 vdd gnd cell_6t
Xbit_r130_c108 bl_108 br_108 wl_130 vdd gnd cell_6t
Xbit_r131_c108 bl_108 br_108 wl_131 vdd gnd cell_6t
Xbit_r132_c108 bl_108 br_108 wl_132 vdd gnd cell_6t
Xbit_r133_c108 bl_108 br_108 wl_133 vdd gnd cell_6t
Xbit_r134_c108 bl_108 br_108 wl_134 vdd gnd cell_6t
Xbit_r135_c108 bl_108 br_108 wl_135 vdd gnd cell_6t
Xbit_r136_c108 bl_108 br_108 wl_136 vdd gnd cell_6t
Xbit_r137_c108 bl_108 br_108 wl_137 vdd gnd cell_6t
Xbit_r138_c108 bl_108 br_108 wl_138 vdd gnd cell_6t
Xbit_r139_c108 bl_108 br_108 wl_139 vdd gnd cell_6t
Xbit_r140_c108 bl_108 br_108 wl_140 vdd gnd cell_6t
Xbit_r141_c108 bl_108 br_108 wl_141 vdd gnd cell_6t
Xbit_r142_c108 bl_108 br_108 wl_142 vdd gnd cell_6t
Xbit_r143_c108 bl_108 br_108 wl_143 vdd gnd cell_6t
Xbit_r144_c108 bl_108 br_108 wl_144 vdd gnd cell_6t
Xbit_r145_c108 bl_108 br_108 wl_145 vdd gnd cell_6t
Xbit_r146_c108 bl_108 br_108 wl_146 vdd gnd cell_6t
Xbit_r147_c108 bl_108 br_108 wl_147 vdd gnd cell_6t
Xbit_r148_c108 bl_108 br_108 wl_148 vdd gnd cell_6t
Xbit_r149_c108 bl_108 br_108 wl_149 vdd gnd cell_6t
Xbit_r150_c108 bl_108 br_108 wl_150 vdd gnd cell_6t
Xbit_r151_c108 bl_108 br_108 wl_151 vdd gnd cell_6t
Xbit_r152_c108 bl_108 br_108 wl_152 vdd gnd cell_6t
Xbit_r153_c108 bl_108 br_108 wl_153 vdd gnd cell_6t
Xbit_r154_c108 bl_108 br_108 wl_154 vdd gnd cell_6t
Xbit_r155_c108 bl_108 br_108 wl_155 vdd gnd cell_6t
Xbit_r156_c108 bl_108 br_108 wl_156 vdd gnd cell_6t
Xbit_r157_c108 bl_108 br_108 wl_157 vdd gnd cell_6t
Xbit_r158_c108 bl_108 br_108 wl_158 vdd gnd cell_6t
Xbit_r159_c108 bl_108 br_108 wl_159 vdd gnd cell_6t
Xbit_r160_c108 bl_108 br_108 wl_160 vdd gnd cell_6t
Xbit_r161_c108 bl_108 br_108 wl_161 vdd gnd cell_6t
Xbit_r162_c108 bl_108 br_108 wl_162 vdd gnd cell_6t
Xbit_r163_c108 bl_108 br_108 wl_163 vdd gnd cell_6t
Xbit_r164_c108 bl_108 br_108 wl_164 vdd gnd cell_6t
Xbit_r165_c108 bl_108 br_108 wl_165 vdd gnd cell_6t
Xbit_r166_c108 bl_108 br_108 wl_166 vdd gnd cell_6t
Xbit_r167_c108 bl_108 br_108 wl_167 vdd gnd cell_6t
Xbit_r168_c108 bl_108 br_108 wl_168 vdd gnd cell_6t
Xbit_r169_c108 bl_108 br_108 wl_169 vdd gnd cell_6t
Xbit_r170_c108 bl_108 br_108 wl_170 vdd gnd cell_6t
Xbit_r171_c108 bl_108 br_108 wl_171 vdd gnd cell_6t
Xbit_r172_c108 bl_108 br_108 wl_172 vdd gnd cell_6t
Xbit_r173_c108 bl_108 br_108 wl_173 vdd gnd cell_6t
Xbit_r174_c108 bl_108 br_108 wl_174 vdd gnd cell_6t
Xbit_r175_c108 bl_108 br_108 wl_175 vdd gnd cell_6t
Xbit_r176_c108 bl_108 br_108 wl_176 vdd gnd cell_6t
Xbit_r177_c108 bl_108 br_108 wl_177 vdd gnd cell_6t
Xbit_r178_c108 bl_108 br_108 wl_178 vdd gnd cell_6t
Xbit_r179_c108 bl_108 br_108 wl_179 vdd gnd cell_6t
Xbit_r180_c108 bl_108 br_108 wl_180 vdd gnd cell_6t
Xbit_r181_c108 bl_108 br_108 wl_181 vdd gnd cell_6t
Xbit_r182_c108 bl_108 br_108 wl_182 vdd gnd cell_6t
Xbit_r183_c108 bl_108 br_108 wl_183 vdd gnd cell_6t
Xbit_r184_c108 bl_108 br_108 wl_184 vdd gnd cell_6t
Xbit_r185_c108 bl_108 br_108 wl_185 vdd gnd cell_6t
Xbit_r186_c108 bl_108 br_108 wl_186 vdd gnd cell_6t
Xbit_r187_c108 bl_108 br_108 wl_187 vdd gnd cell_6t
Xbit_r188_c108 bl_108 br_108 wl_188 vdd gnd cell_6t
Xbit_r189_c108 bl_108 br_108 wl_189 vdd gnd cell_6t
Xbit_r190_c108 bl_108 br_108 wl_190 vdd gnd cell_6t
Xbit_r191_c108 bl_108 br_108 wl_191 vdd gnd cell_6t
Xbit_r192_c108 bl_108 br_108 wl_192 vdd gnd cell_6t
Xbit_r193_c108 bl_108 br_108 wl_193 vdd gnd cell_6t
Xbit_r194_c108 bl_108 br_108 wl_194 vdd gnd cell_6t
Xbit_r195_c108 bl_108 br_108 wl_195 vdd gnd cell_6t
Xbit_r196_c108 bl_108 br_108 wl_196 vdd gnd cell_6t
Xbit_r197_c108 bl_108 br_108 wl_197 vdd gnd cell_6t
Xbit_r198_c108 bl_108 br_108 wl_198 vdd gnd cell_6t
Xbit_r199_c108 bl_108 br_108 wl_199 vdd gnd cell_6t
Xbit_r200_c108 bl_108 br_108 wl_200 vdd gnd cell_6t
Xbit_r201_c108 bl_108 br_108 wl_201 vdd gnd cell_6t
Xbit_r202_c108 bl_108 br_108 wl_202 vdd gnd cell_6t
Xbit_r203_c108 bl_108 br_108 wl_203 vdd gnd cell_6t
Xbit_r204_c108 bl_108 br_108 wl_204 vdd gnd cell_6t
Xbit_r205_c108 bl_108 br_108 wl_205 vdd gnd cell_6t
Xbit_r206_c108 bl_108 br_108 wl_206 vdd gnd cell_6t
Xbit_r207_c108 bl_108 br_108 wl_207 vdd gnd cell_6t
Xbit_r208_c108 bl_108 br_108 wl_208 vdd gnd cell_6t
Xbit_r209_c108 bl_108 br_108 wl_209 vdd gnd cell_6t
Xbit_r210_c108 bl_108 br_108 wl_210 vdd gnd cell_6t
Xbit_r211_c108 bl_108 br_108 wl_211 vdd gnd cell_6t
Xbit_r212_c108 bl_108 br_108 wl_212 vdd gnd cell_6t
Xbit_r213_c108 bl_108 br_108 wl_213 vdd gnd cell_6t
Xbit_r214_c108 bl_108 br_108 wl_214 vdd gnd cell_6t
Xbit_r215_c108 bl_108 br_108 wl_215 vdd gnd cell_6t
Xbit_r216_c108 bl_108 br_108 wl_216 vdd gnd cell_6t
Xbit_r217_c108 bl_108 br_108 wl_217 vdd gnd cell_6t
Xbit_r218_c108 bl_108 br_108 wl_218 vdd gnd cell_6t
Xbit_r219_c108 bl_108 br_108 wl_219 vdd gnd cell_6t
Xbit_r220_c108 bl_108 br_108 wl_220 vdd gnd cell_6t
Xbit_r221_c108 bl_108 br_108 wl_221 vdd gnd cell_6t
Xbit_r222_c108 bl_108 br_108 wl_222 vdd gnd cell_6t
Xbit_r223_c108 bl_108 br_108 wl_223 vdd gnd cell_6t
Xbit_r224_c108 bl_108 br_108 wl_224 vdd gnd cell_6t
Xbit_r225_c108 bl_108 br_108 wl_225 vdd gnd cell_6t
Xbit_r226_c108 bl_108 br_108 wl_226 vdd gnd cell_6t
Xbit_r227_c108 bl_108 br_108 wl_227 vdd gnd cell_6t
Xbit_r228_c108 bl_108 br_108 wl_228 vdd gnd cell_6t
Xbit_r229_c108 bl_108 br_108 wl_229 vdd gnd cell_6t
Xbit_r230_c108 bl_108 br_108 wl_230 vdd gnd cell_6t
Xbit_r231_c108 bl_108 br_108 wl_231 vdd gnd cell_6t
Xbit_r232_c108 bl_108 br_108 wl_232 vdd gnd cell_6t
Xbit_r233_c108 bl_108 br_108 wl_233 vdd gnd cell_6t
Xbit_r234_c108 bl_108 br_108 wl_234 vdd gnd cell_6t
Xbit_r235_c108 bl_108 br_108 wl_235 vdd gnd cell_6t
Xbit_r236_c108 bl_108 br_108 wl_236 vdd gnd cell_6t
Xbit_r237_c108 bl_108 br_108 wl_237 vdd gnd cell_6t
Xbit_r238_c108 bl_108 br_108 wl_238 vdd gnd cell_6t
Xbit_r239_c108 bl_108 br_108 wl_239 vdd gnd cell_6t
Xbit_r240_c108 bl_108 br_108 wl_240 vdd gnd cell_6t
Xbit_r241_c108 bl_108 br_108 wl_241 vdd gnd cell_6t
Xbit_r242_c108 bl_108 br_108 wl_242 vdd gnd cell_6t
Xbit_r243_c108 bl_108 br_108 wl_243 vdd gnd cell_6t
Xbit_r244_c108 bl_108 br_108 wl_244 vdd gnd cell_6t
Xbit_r245_c108 bl_108 br_108 wl_245 vdd gnd cell_6t
Xbit_r246_c108 bl_108 br_108 wl_246 vdd gnd cell_6t
Xbit_r247_c108 bl_108 br_108 wl_247 vdd gnd cell_6t
Xbit_r248_c108 bl_108 br_108 wl_248 vdd gnd cell_6t
Xbit_r249_c108 bl_108 br_108 wl_249 vdd gnd cell_6t
Xbit_r250_c108 bl_108 br_108 wl_250 vdd gnd cell_6t
Xbit_r251_c108 bl_108 br_108 wl_251 vdd gnd cell_6t
Xbit_r252_c108 bl_108 br_108 wl_252 vdd gnd cell_6t
Xbit_r253_c108 bl_108 br_108 wl_253 vdd gnd cell_6t
Xbit_r254_c108 bl_108 br_108 wl_254 vdd gnd cell_6t
Xbit_r255_c108 bl_108 br_108 wl_255 vdd gnd cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd cell_6t
Xbit_r1_c109 bl_109 br_109 wl_1 vdd gnd cell_6t
Xbit_r2_c109 bl_109 br_109 wl_2 vdd gnd cell_6t
Xbit_r3_c109 bl_109 br_109 wl_3 vdd gnd cell_6t
Xbit_r4_c109 bl_109 br_109 wl_4 vdd gnd cell_6t
Xbit_r5_c109 bl_109 br_109 wl_5 vdd gnd cell_6t
Xbit_r6_c109 bl_109 br_109 wl_6 vdd gnd cell_6t
Xbit_r7_c109 bl_109 br_109 wl_7 vdd gnd cell_6t
Xbit_r8_c109 bl_109 br_109 wl_8 vdd gnd cell_6t
Xbit_r9_c109 bl_109 br_109 wl_9 vdd gnd cell_6t
Xbit_r10_c109 bl_109 br_109 wl_10 vdd gnd cell_6t
Xbit_r11_c109 bl_109 br_109 wl_11 vdd gnd cell_6t
Xbit_r12_c109 bl_109 br_109 wl_12 vdd gnd cell_6t
Xbit_r13_c109 bl_109 br_109 wl_13 vdd gnd cell_6t
Xbit_r14_c109 bl_109 br_109 wl_14 vdd gnd cell_6t
Xbit_r15_c109 bl_109 br_109 wl_15 vdd gnd cell_6t
Xbit_r16_c109 bl_109 br_109 wl_16 vdd gnd cell_6t
Xbit_r17_c109 bl_109 br_109 wl_17 vdd gnd cell_6t
Xbit_r18_c109 bl_109 br_109 wl_18 vdd gnd cell_6t
Xbit_r19_c109 bl_109 br_109 wl_19 vdd gnd cell_6t
Xbit_r20_c109 bl_109 br_109 wl_20 vdd gnd cell_6t
Xbit_r21_c109 bl_109 br_109 wl_21 vdd gnd cell_6t
Xbit_r22_c109 bl_109 br_109 wl_22 vdd gnd cell_6t
Xbit_r23_c109 bl_109 br_109 wl_23 vdd gnd cell_6t
Xbit_r24_c109 bl_109 br_109 wl_24 vdd gnd cell_6t
Xbit_r25_c109 bl_109 br_109 wl_25 vdd gnd cell_6t
Xbit_r26_c109 bl_109 br_109 wl_26 vdd gnd cell_6t
Xbit_r27_c109 bl_109 br_109 wl_27 vdd gnd cell_6t
Xbit_r28_c109 bl_109 br_109 wl_28 vdd gnd cell_6t
Xbit_r29_c109 bl_109 br_109 wl_29 vdd gnd cell_6t
Xbit_r30_c109 bl_109 br_109 wl_30 vdd gnd cell_6t
Xbit_r31_c109 bl_109 br_109 wl_31 vdd gnd cell_6t
Xbit_r32_c109 bl_109 br_109 wl_32 vdd gnd cell_6t
Xbit_r33_c109 bl_109 br_109 wl_33 vdd gnd cell_6t
Xbit_r34_c109 bl_109 br_109 wl_34 vdd gnd cell_6t
Xbit_r35_c109 bl_109 br_109 wl_35 vdd gnd cell_6t
Xbit_r36_c109 bl_109 br_109 wl_36 vdd gnd cell_6t
Xbit_r37_c109 bl_109 br_109 wl_37 vdd gnd cell_6t
Xbit_r38_c109 bl_109 br_109 wl_38 vdd gnd cell_6t
Xbit_r39_c109 bl_109 br_109 wl_39 vdd gnd cell_6t
Xbit_r40_c109 bl_109 br_109 wl_40 vdd gnd cell_6t
Xbit_r41_c109 bl_109 br_109 wl_41 vdd gnd cell_6t
Xbit_r42_c109 bl_109 br_109 wl_42 vdd gnd cell_6t
Xbit_r43_c109 bl_109 br_109 wl_43 vdd gnd cell_6t
Xbit_r44_c109 bl_109 br_109 wl_44 vdd gnd cell_6t
Xbit_r45_c109 bl_109 br_109 wl_45 vdd gnd cell_6t
Xbit_r46_c109 bl_109 br_109 wl_46 vdd gnd cell_6t
Xbit_r47_c109 bl_109 br_109 wl_47 vdd gnd cell_6t
Xbit_r48_c109 bl_109 br_109 wl_48 vdd gnd cell_6t
Xbit_r49_c109 bl_109 br_109 wl_49 vdd gnd cell_6t
Xbit_r50_c109 bl_109 br_109 wl_50 vdd gnd cell_6t
Xbit_r51_c109 bl_109 br_109 wl_51 vdd gnd cell_6t
Xbit_r52_c109 bl_109 br_109 wl_52 vdd gnd cell_6t
Xbit_r53_c109 bl_109 br_109 wl_53 vdd gnd cell_6t
Xbit_r54_c109 bl_109 br_109 wl_54 vdd gnd cell_6t
Xbit_r55_c109 bl_109 br_109 wl_55 vdd gnd cell_6t
Xbit_r56_c109 bl_109 br_109 wl_56 vdd gnd cell_6t
Xbit_r57_c109 bl_109 br_109 wl_57 vdd gnd cell_6t
Xbit_r58_c109 bl_109 br_109 wl_58 vdd gnd cell_6t
Xbit_r59_c109 bl_109 br_109 wl_59 vdd gnd cell_6t
Xbit_r60_c109 bl_109 br_109 wl_60 vdd gnd cell_6t
Xbit_r61_c109 bl_109 br_109 wl_61 vdd gnd cell_6t
Xbit_r62_c109 bl_109 br_109 wl_62 vdd gnd cell_6t
Xbit_r63_c109 bl_109 br_109 wl_63 vdd gnd cell_6t
Xbit_r64_c109 bl_109 br_109 wl_64 vdd gnd cell_6t
Xbit_r65_c109 bl_109 br_109 wl_65 vdd gnd cell_6t
Xbit_r66_c109 bl_109 br_109 wl_66 vdd gnd cell_6t
Xbit_r67_c109 bl_109 br_109 wl_67 vdd gnd cell_6t
Xbit_r68_c109 bl_109 br_109 wl_68 vdd gnd cell_6t
Xbit_r69_c109 bl_109 br_109 wl_69 vdd gnd cell_6t
Xbit_r70_c109 bl_109 br_109 wl_70 vdd gnd cell_6t
Xbit_r71_c109 bl_109 br_109 wl_71 vdd gnd cell_6t
Xbit_r72_c109 bl_109 br_109 wl_72 vdd gnd cell_6t
Xbit_r73_c109 bl_109 br_109 wl_73 vdd gnd cell_6t
Xbit_r74_c109 bl_109 br_109 wl_74 vdd gnd cell_6t
Xbit_r75_c109 bl_109 br_109 wl_75 vdd gnd cell_6t
Xbit_r76_c109 bl_109 br_109 wl_76 vdd gnd cell_6t
Xbit_r77_c109 bl_109 br_109 wl_77 vdd gnd cell_6t
Xbit_r78_c109 bl_109 br_109 wl_78 vdd gnd cell_6t
Xbit_r79_c109 bl_109 br_109 wl_79 vdd gnd cell_6t
Xbit_r80_c109 bl_109 br_109 wl_80 vdd gnd cell_6t
Xbit_r81_c109 bl_109 br_109 wl_81 vdd gnd cell_6t
Xbit_r82_c109 bl_109 br_109 wl_82 vdd gnd cell_6t
Xbit_r83_c109 bl_109 br_109 wl_83 vdd gnd cell_6t
Xbit_r84_c109 bl_109 br_109 wl_84 vdd gnd cell_6t
Xbit_r85_c109 bl_109 br_109 wl_85 vdd gnd cell_6t
Xbit_r86_c109 bl_109 br_109 wl_86 vdd gnd cell_6t
Xbit_r87_c109 bl_109 br_109 wl_87 vdd gnd cell_6t
Xbit_r88_c109 bl_109 br_109 wl_88 vdd gnd cell_6t
Xbit_r89_c109 bl_109 br_109 wl_89 vdd gnd cell_6t
Xbit_r90_c109 bl_109 br_109 wl_90 vdd gnd cell_6t
Xbit_r91_c109 bl_109 br_109 wl_91 vdd gnd cell_6t
Xbit_r92_c109 bl_109 br_109 wl_92 vdd gnd cell_6t
Xbit_r93_c109 bl_109 br_109 wl_93 vdd gnd cell_6t
Xbit_r94_c109 bl_109 br_109 wl_94 vdd gnd cell_6t
Xbit_r95_c109 bl_109 br_109 wl_95 vdd gnd cell_6t
Xbit_r96_c109 bl_109 br_109 wl_96 vdd gnd cell_6t
Xbit_r97_c109 bl_109 br_109 wl_97 vdd gnd cell_6t
Xbit_r98_c109 bl_109 br_109 wl_98 vdd gnd cell_6t
Xbit_r99_c109 bl_109 br_109 wl_99 vdd gnd cell_6t
Xbit_r100_c109 bl_109 br_109 wl_100 vdd gnd cell_6t
Xbit_r101_c109 bl_109 br_109 wl_101 vdd gnd cell_6t
Xbit_r102_c109 bl_109 br_109 wl_102 vdd gnd cell_6t
Xbit_r103_c109 bl_109 br_109 wl_103 vdd gnd cell_6t
Xbit_r104_c109 bl_109 br_109 wl_104 vdd gnd cell_6t
Xbit_r105_c109 bl_109 br_109 wl_105 vdd gnd cell_6t
Xbit_r106_c109 bl_109 br_109 wl_106 vdd gnd cell_6t
Xbit_r107_c109 bl_109 br_109 wl_107 vdd gnd cell_6t
Xbit_r108_c109 bl_109 br_109 wl_108 vdd gnd cell_6t
Xbit_r109_c109 bl_109 br_109 wl_109 vdd gnd cell_6t
Xbit_r110_c109 bl_109 br_109 wl_110 vdd gnd cell_6t
Xbit_r111_c109 bl_109 br_109 wl_111 vdd gnd cell_6t
Xbit_r112_c109 bl_109 br_109 wl_112 vdd gnd cell_6t
Xbit_r113_c109 bl_109 br_109 wl_113 vdd gnd cell_6t
Xbit_r114_c109 bl_109 br_109 wl_114 vdd gnd cell_6t
Xbit_r115_c109 bl_109 br_109 wl_115 vdd gnd cell_6t
Xbit_r116_c109 bl_109 br_109 wl_116 vdd gnd cell_6t
Xbit_r117_c109 bl_109 br_109 wl_117 vdd gnd cell_6t
Xbit_r118_c109 bl_109 br_109 wl_118 vdd gnd cell_6t
Xbit_r119_c109 bl_109 br_109 wl_119 vdd gnd cell_6t
Xbit_r120_c109 bl_109 br_109 wl_120 vdd gnd cell_6t
Xbit_r121_c109 bl_109 br_109 wl_121 vdd gnd cell_6t
Xbit_r122_c109 bl_109 br_109 wl_122 vdd gnd cell_6t
Xbit_r123_c109 bl_109 br_109 wl_123 vdd gnd cell_6t
Xbit_r124_c109 bl_109 br_109 wl_124 vdd gnd cell_6t
Xbit_r125_c109 bl_109 br_109 wl_125 vdd gnd cell_6t
Xbit_r126_c109 bl_109 br_109 wl_126 vdd gnd cell_6t
Xbit_r127_c109 bl_109 br_109 wl_127 vdd gnd cell_6t
Xbit_r128_c109 bl_109 br_109 wl_128 vdd gnd cell_6t
Xbit_r129_c109 bl_109 br_109 wl_129 vdd gnd cell_6t
Xbit_r130_c109 bl_109 br_109 wl_130 vdd gnd cell_6t
Xbit_r131_c109 bl_109 br_109 wl_131 vdd gnd cell_6t
Xbit_r132_c109 bl_109 br_109 wl_132 vdd gnd cell_6t
Xbit_r133_c109 bl_109 br_109 wl_133 vdd gnd cell_6t
Xbit_r134_c109 bl_109 br_109 wl_134 vdd gnd cell_6t
Xbit_r135_c109 bl_109 br_109 wl_135 vdd gnd cell_6t
Xbit_r136_c109 bl_109 br_109 wl_136 vdd gnd cell_6t
Xbit_r137_c109 bl_109 br_109 wl_137 vdd gnd cell_6t
Xbit_r138_c109 bl_109 br_109 wl_138 vdd gnd cell_6t
Xbit_r139_c109 bl_109 br_109 wl_139 vdd gnd cell_6t
Xbit_r140_c109 bl_109 br_109 wl_140 vdd gnd cell_6t
Xbit_r141_c109 bl_109 br_109 wl_141 vdd gnd cell_6t
Xbit_r142_c109 bl_109 br_109 wl_142 vdd gnd cell_6t
Xbit_r143_c109 bl_109 br_109 wl_143 vdd gnd cell_6t
Xbit_r144_c109 bl_109 br_109 wl_144 vdd gnd cell_6t
Xbit_r145_c109 bl_109 br_109 wl_145 vdd gnd cell_6t
Xbit_r146_c109 bl_109 br_109 wl_146 vdd gnd cell_6t
Xbit_r147_c109 bl_109 br_109 wl_147 vdd gnd cell_6t
Xbit_r148_c109 bl_109 br_109 wl_148 vdd gnd cell_6t
Xbit_r149_c109 bl_109 br_109 wl_149 vdd gnd cell_6t
Xbit_r150_c109 bl_109 br_109 wl_150 vdd gnd cell_6t
Xbit_r151_c109 bl_109 br_109 wl_151 vdd gnd cell_6t
Xbit_r152_c109 bl_109 br_109 wl_152 vdd gnd cell_6t
Xbit_r153_c109 bl_109 br_109 wl_153 vdd gnd cell_6t
Xbit_r154_c109 bl_109 br_109 wl_154 vdd gnd cell_6t
Xbit_r155_c109 bl_109 br_109 wl_155 vdd gnd cell_6t
Xbit_r156_c109 bl_109 br_109 wl_156 vdd gnd cell_6t
Xbit_r157_c109 bl_109 br_109 wl_157 vdd gnd cell_6t
Xbit_r158_c109 bl_109 br_109 wl_158 vdd gnd cell_6t
Xbit_r159_c109 bl_109 br_109 wl_159 vdd gnd cell_6t
Xbit_r160_c109 bl_109 br_109 wl_160 vdd gnd cell_6t
Xbit_r161_c109 bl_109 br_109 wl_161 vdd gnd cell_6t
Xbit_r162_c109 bl_109 br_109 wl_162 vdd gnd cell_6t
Xbit_r163_c109 bl_109 br_109 wl_163 vdd gnd cell_6t
Xbit_r164_c109 bl_109 br_109 wl_164 vdd gnd cell_6t
Xbit_r165_c109 bl_109 br_109 wl_165 vdd gnd cell_6t
Xbit_r166_c109 bl_109 br_109 wl_166 vdd gnd cell_6t
Xbit_r167_c109 bl_109 br_109 wl_167 vdd gnd cell_6t
Xbit_r168_c109 bl_109 br_109 wl_168 vdd gnd cell_6t
Xbit_r169_c109 bl_109 br_109 wl_169 vdd gnd cell_6t
Xbit_r170_c109 bl_109 br_109 wl_170 vdd gnd cell_6t
Xbit_r171_c109 bl_109 br_109 wl_171 vdd gnd cell_6t
Xbit_r172_c109 bl_109 br_109 wl_172 vdd gnd cell_6t
Xbit_r173_c109 bl_109 br_109 wl_173 vdd gnd cell_6t
Xbit_r174_c109 bl_109 br_109 wl_174 vdd gnd cell_6t
Xbit_r175_c109 bl_109 br_109 wl_175 vdd gnd cell_6t
Xbit_r176_c109 bl_109 br_109 wl_176 vdd gnd cell_6t
Xbit_r177_c109 bl_109 br_109 wl_177 vdd gnd cell_6t
Xbit_r178_c109 bl_109 br_109 wl_178 vdd gnd cell_6t
Xbit_r179_c109 bl_109 br_109 wl_179 vdd gnd cell_6t
Xbit_r180_c109 bl_109 br_109 wl_180 vdd gnd cell_6t
Xbit_r181_c109 bl_109 br_109 wl_181 vdd gnd cell_6t
Xbit_r182_c109 bl_109 br_109 wl_182 vdd gnd cell_6t
Xbit_r183_c109 bl_109 br_109 wl_183 vdd gnd cell_6t
Xbit_r184_c109 bl_109 br_109 wl_184 vdd gnd cell_6t
Xbit_r185_c109 bl_109 br_109 wl_185 vdd gnd cell_6t
Xbit_r186_c109 bl_109 br_109 wl_186 vdd gnd cell_6t
Xbit_r187_c109 bl_109 br_109 wl_187 vdd gnd cell_6t
Xbit_r188_c109 bl_109 br_109 wl_188 vdd gnd cell_6t
Xbit_r189_c109 bl_109 br_109 wl_189 vdd gnd cell_6t
Xbit_r190_c109 bl_109 br_109 wl_190 vdd gnd cell_6t
Xbit_r191_c109 bl_109 br_109 wl_191 vdd gnd cell_6t
Xbit_r192_c109 bl_109 br_109 wl_192 vdd gnd cell_6t
Xbit_r193_c109 bl_109 br_109 wl_193 vdd gnd cell_6t
Xbit_r194_c109 bl_109 br_109 wl_194 vdd gnd cell_6t
Xbit_r195_c109 bl_109 br_109 wl_195 vdd gnd cell_6t
Xbit_r196_c109 bl_109 br_109 wl_196 vdd gnd cell_6t
Xbit_r197_c109 bl_109 br_109 wl_197 vdd gnd cell_6t
Xbit_r198_c109 bl_109 br_109 wl_198 vdd gnd cell_6t
Xbit_r199_c109 bl_109 br_109 wl_199 vdd gnd cell_6t
Xbit_r200_c109 bl_109 br_109 wl_200 vdd gnd cell_6t
Xbit_r201_c109 bl_109 br_109 wl_201 vdd gnd cell_6t
Xbit_r202_c109 bl_109 br_109 wl_202 vdd gnd cell_6t
Xbit_r203_c109 bl_109 br_109 wl_203 vdd gnd cell_6t
Xbit_r204_c109 bl_109 br_109 wl_204 vdd gnd cell_6t
Xbit_r205_c109 bl_109 br_109 wl_205 vdd gnd cell_6t
Xbit_r206_c109 bl_109 br_109 wl_206 vdd gnd cell_6t
Xbit_r207_c109 bl_109 br_109 wl_207 vdd gnd cell_6t
Xbit_r208_c109 bl_109 br_109 wl_208 vdd gnd cell_6t
Xbit_r209_c109 bl_109 br_109 wl_209 vdd gnd cell_6t
Xbit_r210_c109 bl_109 br_109 wl_210 vdd gnd cell_6t
Xbit_r211_c109 bl_109 br_109 wl_211 vdd gnd cell_6t
Xbit_r212_c109 bl_109 br_109 wl_212 vdd gnd cell_6t
Xbit_r213_c109 bl_109 br_109 wl_213 vdd gnd cell_6t
Xbit_r214_c109 bl_109 br_109 wl_214 vdd gnd cell_6t
Xbit_r215_c109 bl_109 br_109 wl_215 vdd gnd cell_6t
Xbit_r216_c109 bl_109 br_109 wl_216 vdd gnd cell_6t
Xbit_r217_c109 bl_109 br_109 wl_217 vdd gnd cell_6t
Xbit_r218_c109 bl_109 br_109 wl_218 vdd gnd cell_6t
Xbit_r219_c109 bl_109 br_109 wl_219 vdd gnd cell_6t
Xbit_r220_c109 bl_109 br_109 wl_220 vdd gnd cell_6t
Xbit_r221_c109 bl_109 br_109 wl_221 vdd gnd cell_6t
Xbit_r222_c109 bl_109 br_109 wl_222 vdd gnd cell_6t
Xbit_r223_c109 bl_109 br_109 wl_223 vdd gnd cell_6t
Xbit_r224_c109 bl_109 br_109 wl_224 vdd gnd cell_6t
Xbit_r225_c109 bl_109 br_109 wl_225 vdd gnd cell_6t
Xbit_r226_c109 bl_109 br_109 wl_226 vdd gnd cell_6t
Xbit_r227_c109 bl_109 br_109 wl_227 vdd gnd cell_6t
Xbit_r228_c109 bl_109 br_109 wl_228 vdd gnd cell_6t
Xbit_r229_c109 bl_109 br_109 wl_229 vdd gnd cell_6t
Xbit_r230_c109 bl_109 br_109 wl_230 vdd gnd cell_6t
Xbit_r231_c109 bl_109 br_109 wl_231 vdd gnd cell_6t
Xbit_r232_c109 bl_109 br_109 wl_232 vdd gnd cell_6t
Xbit_r233_c109 bl_109 br_109 wl_233 vdd gnd cell_6t
Xbit_r234_c109 bl_109 br_109 wl_234 vdd gnd cell_6t
Xbit_r235_c109 bl_109 br_109 wl_235 vdd gnd cell_6t
Xbit_r236_c109 bl_109 br_109 wl_236 vdd gnd cell_6t
Xbit_r237_c109 bl_109 br_109 wl_237 vdd gnd cell_6t
Xbit_r238_c109 bl_109 br_109 wl_238 vdd gnd cell_6t
Xbit_r239_c109 bl_109 br_109 wl_239 vdd gnd cell_6t
Xbit_r240_c109 bl_109 br_109 wl_240 vdd gnd cell_6t
Xbit_r241_c109 bl_109 br_109 wl_241 vdd gnd cell_6t
Xbit_r242_c109 bl_109 br_109 wl_242 vdd gnd cell_6t
Xbit_r243_c109 bl_109 br_109 wl_243 vdd gnd cell_6t
Xbit_r244_c109 bl_109 br_109 wl_244 vdd gnd cell_6t
Xbit_r245_c109 bl_109 br_109 wl_245 vdd gnd cell_6t
Xbit_r246_c109 bl_109 br_109 wl_246 vdd gnd cell_6t
Xbit_r247_c109 bl_109 br_109 wl_247 vdd gnd cell_6t
Xbit_r248_c109 bl_109 br_109 wl_248 vdd gnd cell_6t
Xbit_r249_c109 bl_109 br_109 wl_249 vdd gnd cell_6t
Xbit_r250_c109 bl_109 br_109 wl_250 vdd gnd cell_6t
Xbit_r251_c109 bl_109 br_109 wl_251 vdd gnd cell_6t
Xbit_r252_c109 bl_109 br_109 wl_252 vdd gnd cell_6t
Xbit_r253_c109 bl_109 br_109 wl_253 vdd gnd cell_6t
Xbit_r254_c109 bl_109 br_109 wl_254 vdd gnd cell_6t
Xbit_r255_c109 bl_109 br_109 wl_255 vdd gnd cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd cell_6t
Xbit_r1_c110 bl_110 br_110 wl_1 vdd gnd cell_6t
Xbit_r2_c110 bl_110 br_110 wl_2 vdd gnd cell_6t
Xbit_r3_c110 bl_110 br_110 wl_3 vdd gnd cell_6t
Xbit_r4_c110 bl_110 br_110 wl_4 vdd gnd cell_6t
Xbit_r5_c110 bl_110 br_110 wl_5 vdd gnd cell_6t
Xbit_r6_c110 bl_110 br_110 wl_6 vdd gnd cell_6t
Xbit_r7_c110 bl_110 br_110 wl_7 vdd gnd cell_6t
Xbit_r8_c110 bl_110 br_110 wl_8 vdd gnd cell_6t
Xbit_r9_c110 bl_110 br_110 wl_9 vdd gnd cell_6t
Xbit_r10_c110 bl_110 br_110 wl_10 vdd gnd cell_6t
Xbit_r11_c110 bl_110 br_110 wl_11 vdd gnd cell_6t
Xbit_r12_c110 bl_110 br_110 wl_12 vdd gnd cell_6t
Xbit_r13_c110 bl_110 br_110 wl_13 vdd gnd cell_6t
Xbit_r14_c110 bl_110 br_110 wl_14 vdd gnd cell_6t
Xbit_r15_c110 bl_110 br_110 wl_15 vdd gnd cell_6t
Xbit_r16_c110 bl_110 br_110 wl_16 vdd gnd cell_6t
Xbit_r17_c110 bl_110 br_110 wl_17 vdd gnd cell_6t
Xbit_r18_c110 bl_110 br_110 wl_18 vdd gnd cell_6t
Xbit_r19_c110 bl_110 br_110 wl_19 vdd gnd cell_6t
Xbit_r20_c110 bl_110 br_110 wl_20 vdd gnd cell_6t
Xbit_r21_c110 bl_110 br_110 wl_21 vdd gnd cell_6t
Xbit_r22_c110 bl_110 br_110 wl_22 vdd gnd cell_6t
Xbit_r23_c110 bl_110 br_110 wl_23 vdd gnd cell_6t
Xbit_r24_c110 bl_110 br_110 wl_24 vdd gnd cell_6t
Xbit_r25_c110 bl_110 br_110 wl_25 vdd gnd cell_6t
Xbit_r26_c110 bl_110 br_110 wl_26 vdd gnd cell_6t
Xbit_r27_c110 bl_110 br_110 wl_27 vdd gnd cell_6t
Xbit_r28_c110 bl_110 br_110 wl_28 vdd gnd cell_6t
Xbit_r29_c110 bl_110 br_110 wl_29 vdd gnd cell_6t
Xbit_r30_c110 bl_110 br_110 wl_30 vdd gnd cell_6t
Xbit_r31_c110 bl_110 br_110 wl_31 vdd gnd cell_6t
Xbit_r32_c110 bl_110 br_110 wl_32 vdd gnd cell_6t
Xbit_r33_c110 bl_110 br_110 wl_33 vdd gnd cell_6t
Xbit_r34_c110 bl_110 br_110 wl_34 vdd gnd cell_6t
Xbit_r35_c110 bl_110 br_110 wl_35 vdd gnd cell_6t
Xbit_r36_c110 bl_110 br_110 wl_36 vdd gnd cell_6t
Xbit_r37_c110 bl_110 br_110 wl_37 vdd gnd cell_6t
Xbit_r38_c110 bl_110 br_110 wl_38 vdd gnd cell_6t
Xbit_r39_c110 bl_110 br_110 wl_39 vdd gnd cell_6t
Xbit_r40_c110 bl_110 br_110 wl_40 vdd gnd cell_6t
Xbit_r41_c110 bl_110 br_110 wl_41 vdd gnd cell_6t
Xbit_r42_c110 bl_110 br_110 wl_42 vdd gnd cell_6t
Xbit_r43_c110 bl_110 br_110 wl_43 vdd gnd cell_6t
Xbit_r44_c110 bl_110 br_110 wl_44 vdd gnd cell_6t
Xbit_r45_c110 bl_110 br_110 wl_45 vdd gnd cell_6t
Xbit_r46_c110 bl_110 br_110 wl_46 vdd gnd cell_6t
Xbit_r47_c110 bl_110 br_110 wl_47 vdd gnd cell_6t
Xbit_r48_c110 bl_110 br_110 wl_48 vdd gnd cell_6t
Xbit_r49_c110 bl_110 br_110 wl_49 vdd gnd cell_6t
Xbit_r50_c110 bl_110 br_110 wl_50 vdd gnd cell_6t
Xbit_r51_c110 bl_110 br_110 wl_51 vdd gnd cell_6t
Xbit_r52_c110 bl_110 br_110 wl_52 vdd gnd cell_6t
Xbit_r53_c110 bl_110 br_110 wl_53 vdd gnd cell_6t
Xbit_r54_c110 bl_110 br_110 wl_54 vdd gnd cell_6t
Xbit_r55_c110 bl_110 br_110 wl_55 vdd gnd cell_6t
Xbit_r56_c110 bl_110 br_110 wl_56 vdd gnd cell_6t
Xbit_r57_c110 bl_110 br_110 wl_57 vdd gnd cell_6t
Xbit_r58_c110 bl_110 br_110 wl_58 vdd gnd cell_6t
Xbit_r59_c110 bl_110 br_110 wl_59 vdd gnd cell_6t
Xbit_r60_c110 bl_110 br_110 wl_60 vdd gnd cell_6t
Xbit_r61_c110 bl_110 br_110 wl_61 vdd gnd cell_6t
Xbit_r62_c110 bl_110 br_110 wl_62 vdd gnd cell_6t
Xbit_r63_c110 bl_110 br_110 wl_63 vdd gnd cell_6t
Xbit_r64_c110 bl_110 br_110 wl_64 vdd gnd cell_6t
Xbit_r65_c110 bl_110 br_110 wl_65 vdd gnd cell_6t
Xbit_r66_c110 bl_110 br_110 wl_66 vdd gnd cell_6t
Xbit_r67_c110 bl_110 br_110 wl_67 vdd gnd cell_6t
Xbit_r68_c110 bl_110 br_110 wl_68 vdd gnd cell_6t
Xbit_r69_c110 bl_110 br_110 wl_69 vdd gnd cell_6t
Xbit_r70_c110 bl_110 br_110 wl_70 vdd gnd cell_6t
Xbit_r71_c110 bl_110 br_110 wl_71 vdd gnd cell_6t
Xbit_r72_c110 bl_110 br_110 wl_72 vdd gnd cell_6t
Xbit_r73_c110 bl_110 br_110 wl_73 vdd gnd cell_6t
Xbit_r74_c110 bl_110 br_110 wl_74 vdd gnd cell_6t
Xbit_r75_c110 bl_110 br_110 wl_75 vdd gnd cell_6t
Xbit_r76_c110 bl_110 br_110 wl_76 vdd gnd cell_6t
Xbit_r77_c110 bl_110 br_110 wl_77 vdd gnd cell_6t
Xbit_r78_c110 bl_110 br_110 wl_78 vdd gnd cell_6t
Xbit_r79_c110 bl_110 br_110 wl_79 vdd gnd cell_6t
Xbit_r80_c110 bl_110 br_110 wl_80 vdd gnd cell_6t
Xbit_r81_c110 bl_110 br_110 wl_81 vdd gnd cell_6t
Xbit_r82_c110 bl_110 br_110 wl_82 vdd gnd cell_6t
Xbit_r83_c110 bl_110 br_110 wl_83 vdd gnd cell_6t
Xbit_r84_c110 bl_110 br_110 wl_84 vdd gnd cell_6t
Xbit_r85_c110 bl_110 br_110 wl_85 vdd gnd cell_6t
Xbit_r86_c110 bl_110 br_110 wl_86 vdd gnd cell_6t
Xbit_r87_c110 bl_110 br_110 wl_87 vdd gnd cell_6t
Xbit_r88_c110 bl_110 br_110 wl_88 vdd gnd cell_6t
Xbit_r89_c110 bl_110 br_110 wl_89 vdd gnd cell_6t
Xbit_r90_c110 bl_110 br_110 wl_90 vdd gnd cell_6t
Xbit_r91_c110 bl_110 br_110 wl_91 vdd gnd cell_6t
Xbit_r92_c110 bl_110 br_110 wl_92 vdd gnd cell_6t
Xbit_r93_c110 bl_110 br_110 wl_93 vdd gnd cell_6t
Xbit_r94_c110 bl_110 br_110 wl_94 vdd gnd cell_6t
Xbit_r95_c110 bl_110 br_110 wl_95 vdd gnd cell_6t
Xbit_r96_c110 bl_110 br_110 wl_96 vdd gnd cell_6t
Xbit_r97_c110 bl_110 br_110 wl_97 vdd gnd cell_6t
Xbit_r98_c110 bl_110 br_110 wl_98 vdd gnd cell_6t
Xbit_r99_c110 bl_110 br_110 wl_99 vdd gnd cell_6t
Xbit_r100_c110 bl_110 br_110 wl_100 vdd gnd cell_6t
Xbit_r101_c110 bl_110 br_110 wl_101 vdd gnd cell_6t
Xbit_r102_c110 bl_110 br_110 wl_102 vdd gnd cell_6t
Xbit_r103_c110 bl_110 br_110 wl_103 vdd gnd cell_6t
Xbit_r104_c110 bl_110 br_110 wl_104 vdd gnd cell_6t
Xbit_r105_c110 bl_110 br_110 wl_105 vdd gnd cell_6t
Xbit_r106_c110 bl_110 br_110 wl_106 vdd gnd cell_6t
Xbit_r107_c110 bl_110 br_110 wl_107 vdd gnd cell_6t
Xbit_r108_c110 bl_110 br_110 wl_108 vdd gnd cell_6t
Xbit_r109_c110 bl_110 br_110 wl_109 vdd gnd cell_6t
Xbit_r110_c110 bl_110 br_110 wl_110 vdd gnd cell_6t
Xbit_r111_c110 bl_110 br_110 wl_111 vdd gnd cell_6t
Xbit_r112_c110 bl_110 br_110 wl_112 vdd gnd cell_6t
Xbit_r113_c110 bl_110 br_110 wl_113 vdd gnd cell_6t
Xbit_r114_c110 bl_110 br_110 wl_114 vdd gnd cell_6t
Xbit_r115_c110 bl_110 br_110 wl_115 vdd gnd cell_6t
Xbit_r116_c110 bl_110 br_110 wl_116 vdd gnd cell_6t
Xbit_r117_c110 bl_110 br_110 wl_117 vdd gnd cell_6t
Xbit_r118_c110 bl_110 br_110 wl_118 vdd gnd cell_6t
Xbit_r119_c110 bl_110 br_110 wl_119 vdd gnd cell_6t
Xbit_r120_c110 bl_110 br_110 wl_120 vdd gnd cell_6t
Xbit_r121_c110 bl_110 br_110 wl_121 vdd gnd cell_6t
Xbit_r122_c110 bl_110 br_110 wl_122 vdd gnd cell_6t
Xbit_r123_c110 bl_110 br_110 wl_123 vdd gnd cell_6t
Xbit_r124_c110 bl_110 br_110 wl_124 vdd gnd cell_6t
Xbit_r125_c110 bl_110 br_110 wl_125 vdd gnd cell_6t
Xbit_r126_c110 bl_110 br_110 wl_126 vdd gnd cell_6t
Xbit_r127_c110 bl_110 br_110 wl_127 vdd gnd cell_6t
Xbit_r128_c110 bl_110 br_110 wl_128 vdd gnd cell_6t
Xbit_r129_c110 bl_110 br_110 wl_129 vdd gnd cell_6t
Xbit_r130_c110 bl_110 br_110 wl_130 vdd gnd cell_6t
Xbit_r131_c110 bl_110 br_110 wl_131 vdd gnd cell_6t
Xbit_r132_c110 bl_110 br_110 wl_132 vdd gnd cell_6t
Xbit_r133_c110 bl_110 br_110 wl_133 vdd gnd cell_6t
Xbit_r134_c110 bl_110 br_110 wl_134 vdd gnd cell_6t
Xbit_r135_c110 bl_110 br_110 wl_135 vdd gnd cell_6t
Xbit_r136_c110 bl_110 br_110 wl_136 vdd gnd cell_6t
Xbit_r137_c110 bl_110 br_110 wl_137 vdd gnd cell_6t
Xbit_r138_c110 bl_110 br_110 wl_138 vdd gnd cell_6t
Xbit_r139_c110 bl_110 br_110 wl_139 vdd gnd cell_6t
Xbit_r140_c110 bl_110 br_110 wl_140 vdd gnd cell_6t
Xbit_r141_c110 bl_110 br_110 wl_141 vdd gnd cell_6t
Xbit_r142_c110 bl_110 br_110 wl_142 vdd gnd cell_6t
Xbit_r143_c110 bl_110 br_110 wl_143 vdd gnd cell_6t
Xbit_r144_c110 bl_110 br_110 wl_144 vdd gnd cell_6t
Xbit_r145_c110 bl_110 br_110 wl_145 vdd gnd cell_6t
Xbit_r146_c110 bl_110 br_110 wl_146 vdd gnd cell_6t
Xbit_r147_c110 bl_110 br_110 wl_147 vdd gnd cell_6t
Xbit_r148_c110 bl_110 br_110 wl_148 vdd gnd cell_6t
Xbit_r149_c110 bl_110 br_110 wl_149 vdd gnd cell_6t
Xbit_r150_c110 bl_110 br_110 wl_150 vdd gnd cell_6t
Xbit_r151_c110 bl_110 br_110 wl_151 vdd gnd cell_6t
Xbit_r152_c110 bl_110 br_110 wl_152 vdd gnd cell_6t
Xbit_r153_c110 bl_110 br_110 wl_153 vdd gnd cell_6t
Xbit_r154_c110 bl_110 br_110 wl_154 vdd gnd cell_6t
Xbit_r155_c110 bl_110 br_110 wl_155 vdd gnd cell_6t
Xbit_r156_c110 bl_110 br_110 wl_156 vdd gnd cell_6t
Xbit_r157_c110 bl_110 br_110 wl_157 vdd gnd cell_6t
Xbit_r158_c110 bl_110 br_110 wl_158 vdd gnd cell_6t
Xbit_r159_c110 bl_110 br_110 wl_159 vdd gnd cell_6t
Xbit_r160_c110 bl_110 br_110 wl_160 vdd gnd cell_6t
Xbit_r161_c110 bl_110 br_110 wl_161 vdd gnd cell_6t
Xbit_r162_c110 bl_110 br_110 wl_162 vdd gnd cell_6t
Xbit_r163_c110 bl_110 br_110 wl_163 vdd gnd cell_6t
Xbit_r164_c110 bl_110 br_110 wl_164 vdd gnd cell_6t
Xbit_r165_c110 bl_110 br_110 wl_165 vdd gnd cell_6t
Xbit_r166_c110 bl_110 br_110 wl_166 vdd gnd cell_6t
Xbit_r167_c110 bl_110 br_110 wl_167 vdd gnd cell_6t
Xbit_r168_c110 bl_110 br_110 wl_168 vdd gnd cell_6t
Xbit_r169_c110 bl_110 br_110 wl_169 vdd gnd cell_6t
Xbit_r170_c110 bl_110 br_110 wl_170 vdd gnd cell_6t
Xbit_r171_c110 bl_110 br_110 wl_171 vdd gnd cell_6t
Xbit_r172_c110 bl_110 br_110 wl_172 vdd gnd cell_6t
Xbit_r173_c110 bl_110 br_110 wl_173 vdd gnd cell_6t
Xbit_r174_c110 bl_110 br_110 wl_174 vdd gnd cell_6t
Xbit_r175_c110 bl_110 br_110 wl_175 vdd gnd cell_6t
Xbit_r176_c110 bl_110 br_110 wl_176 vdd gnd cell_6t
Xbit_r177_c110 bl_110 br_110 wl_177 vdd gnd cell_6t
Xbit_r178_c110 bl_110 br_110 wl_178 vdd gnd cell_6t
Xbit_r179_c110 bl_110 br_110 wl_179 vdd gnd cell_6t
Xbit_r180_c110 bl_110 br_110 wl_180 vdd gnd cell_6t
Xbit_r181_c110 bl_110 br_110 wl_181 vdd gnd cell_6t
Xbit_r182_c110 bl_110 br_110 wl_182 vdd gnd cell_6t
Xbit_r183_c110 bl_110 br_110 wl_183 vdd gnd cell_6t
Xbit_r184_c110 bl_110 br_110 wl_184 vdd gnd cell_6t
Xbit_r185_c110 bl_110 br_110 wl_185 vdd gnd cell_6t
Xbit_r186_c110 bl_110 br_110 wl_186 vdd gnd cell_6t
Xbit_r187_c110 bl_110 br_110 wl_187 vdd gnd cell_6t
Xbit_r188_c110 bl_110 br_110 wl_188 vdd gnd cell_6t
Xbit_r189_c110 bl_110 br_110 wl_189 vdd gnd cell_6t
Xbit_r190_c110 bl_110 br_110 wl_190 vdd gnd cell_6t
Xbit_r191_c110 bl_110 br_110 wl_191 vdd gnd cell_6t
Xbit_r192_c110 bl_110 br_110 wl_192 vdd gnd cell_6t
Xbit_r193_c110 bl_110 br_110 wl_193 vdd gnd cell_6t
Xbit_r194_c110 bl_110 br_110 wl_194 vdd gnd cell_6t
Xbit_r195_c110 bl_110 br_110 wl_195 vdd gnd cell_6t
Xbit_r196_c110 bl_110 br_110 wl_196 vdd gnd cell_6t
Xbit_r197_c110 bl_110 br_110 wl_197 vdd gnd cell_6t
Xbit_r198_c110 bl_110 br_110 wl_198 vdd gnd cell_6t
Xbit_r199_c110 bl_110 br_110 wl_199 vdd gnd cell_6t
Xbit_r200_c110 bl_110 br_110 wl_200 vdd gnd cell_6t
Xbit_r201_c110 bl_110 br_110 wl_201 vdd gnd cell_6t
Xbit_r202_c110 bl_110 br_110 wl_202 vdd gnd cell_6t
Xbit_r203_c110 bl_110 br_110 wl_203 vdd gnd cell_6t
Xbit_r204_c110 bl_110 br_110 wl_204 vdd gnd cell_6t
Xbit_r205_c110 bl_110 br_110 wl_205 vdd gnd cell_6t
Xbit_r206_c110 bl_110 br_110 wl_206 vdd gnd cell_6t
Xbit_r207_c110 bl_110 br_110 wl_207 vdd gnd cell_6t
Xbit_r208_c110 bl_110 br_110 wl_208 vdd gnd cell_6t
Xbit_r209_c110 bl_110 br_110 wl_209 vdd gnd cell_6t
Xbit_r210_c110 bl_110 br_110 wl_210 vdd gnd cell_6t
Xbit_r211_c110 bl_110 br_110 wl_211 vdd gnd cell_6t
Xbit_r212_c110 bl_110 br_110 wl_212 vdd gnd cell_6t
Xbit_r213_c110 bl_110 br_110 wl_213 vdd gnd cell_6t
Xbit_r214_c110 bl_110 br_110 wl_214 vdd gnd cell_6t
Xbit_r215_c110 bl_110 br_110 wl_215 vdd gnd cell_6t
Xbit_r216_c110 bl_110 br_110 wl_216 vdd gnd cell_6t
Xbit_r217_c110 bl_110 br_110 wl_217 vdd gnd cell_6t
Xbit_r218_c110 bl_110 br_110 wl_218 vdd gnd cell_6t
Xbit_r219_c110 bl_110 br_110 wl_219 vdd gnd cell_6t
Xbit_r220_c110 bl_110 br_110 wl_220 vdd gnd cell_6t
Xbit_r221_c110 bl_110 br_110 wl_221 vdd gnd cell_6t
Xbit_r222_c110 bl_110 br_110 wl_222 vdd gnd cell_6t
Xbit_r223_c110 bl_110 br_110 wl_223 vdd gnd cell_6t
Xbit_r224_c110 bl_110 br_110 wl_224 vdd gnd cell_6t
Xbit_r225_c110 bl_110 br_110 wl_225 vdd gnd cell_6t
Xbit_r226_c110 bl_110 br_110 wl_226 vdd gnd cell_6t
Xbit_r227_c110 bl_110 br_110 wl_227 vdd gnd cell_6t
Xbit_r228_c110 bl_110 br_110 wl_228 vdd gnd cell_6t
Xbit_r229_c110 bl_110 br_110 wl_229 vdd gnd cell_6t
Xbit_r230_c110 bl_110 br_110 wl_230 vdd gnd cell_6t
Xbit_r231_c110 bl_110 br_110 wl_231 vdd gnd cell_6t
Xbit_r232_c110 bl_110 br_110 wl_232 vdd gnd cell_6t
Xbit_r233_c110 bl_110 br_110 wl_233 vdd gnd cell_6t
Xbit_r234_c110 bl_110 br_110 wl_234 vdd gnd cell_6t
Xbit_r235_c110 bl_110 br_110 wl_235 vdd gnd cell_6t
Xbit_r236_c110 bl_110 br_110 wl_236 vdd gnd cell_6t
Xbit_r237_c110 bl_110 br_110 wl_237 vdd gnd cell_6t
Xbit_r238_c110 bl_110 br_110 wl_238 vdd gnd cell_6t
Xbit_r239_c110 bl_110 br_110 wl_239 vdd gnd cell_6t
Xbit_r240_c110 bl_110 br_110 wl_240 vdd gnd cell_6t
Xbit_r241_c110 bl_110 br_110 wl_241 vdd gnd cell_6t
Xbit_r242_c110 bl_110 br_110 wl_242 vdd gnd cell_6t
Xbit_r243_c110 bl_110 br_110 wl_243 vdd gnd cell_6t
Xbit_r244_c110 bl_110 br_110 wl_244 vdd gnd cell_6t
Xbit_r245_c110 bl_110 br_110 wl_245 vdd gnd cell_6t
Xbit_r246_c110 bl_110 br_110 wl_246 vdd gnd cell_6t
Xbit_r247_c110 bl_110 br_110 wl_247 vdd gnd cell_6t
Xbit_r248_c110 bl_110 br_110 wl_248 vdd gnd cell_6t
Xbit_r249_c110 bl_110 br_110 wl_249 vdd gnd cell_6t
Xbit_r250_c110 bl_110 br_110 wl_250 vdd gnd cell_6t
Xbit_r251_c110 bl_110 br_110 wl_251 vdd gnd cell_6t
Xbit_r252_c110 bl_110 br_110 wl_252 vdd gnd cell_6t
Xbit_r253_c110 bl_110 br_110 wl_253 vdd gnd cell_6t
Xbit_r254_c110 bl_110 br_110 wl_254 vdd gnd cell_6t
Xbit_r255_c110 bl_110 br_110 wl_255 vdd gnd cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd cell_6t
Xbit_r1_c111 bl_111 br_111 wl_1 vdd gnd cell_6t
Xbit_r2_c111 bl_111 br_111 wl_2 vdd gnd cell_6t
Xbit_r3_c111 bl_111 br_111 wl_3 vdd gnd cell_6t
Xbit_r4_c111 bl_111 br_111 wl_4 vdd gnd cell_6t
Xbit_r5_c111 bl_111 br_111 wl_5 vdd gnd cell_6t
Xbit_r6_c111 bl_111 br_111 wl_6 vdd gnd cell_6t
Xbit_r7_c111 bl_111 br_111 wl_7 vdd gnd cell_6t
Xbit_r8_c111 bl_111 br_111 wl_8 vdd gnd cell_6t
Xbit_r9_c111 bl_111 br_111 wl_9 vdd gnd cell_6t
Xbit_r10_c111 bl_111 br_111 wl_10 vdd gnd cell_6t
Xbit_r11_c111 bl_111 br_111 wl_11 vdd gnd cell_6t
Xbit_r12_c111 bl_111 br_111 wl_12 vdd gnd cell_6t
Xbit_r13_c111 bl_111 br_111 wl_13 vdd gnd cell_6t
Xbit_r14_c111 bl_111 br_111 wl_14 vdd gnd cell_6t
Xbit_r15_c111 bl_111 br_111 wl_15 vdd gnd cell_6t
Xbit_r16_c111 bl_111 br_111 wl_16 vdd gnd cell_6t
Xbit_r17_c111 bl_111 br_111 wl_17 vdd gnd cell_6t
Xbit_r18_c111 bl_111 br_111 wl_18 vdd gnd cell_6t
Xbit_r19_c111 bl_111 br_111 wl_19 vdd gnd cell_6t
Xbit_r20_c111 bl_111 br_111 wl_20 vdd gnd cell_6t
Xbit_r21_c111 bl_111 br_111 wl_21 vdd gnd cell_6t
Xbit_r22_c111 bl_111 br_111 wl_22 vdd gnd cell_6t
Xbit_r23_c111 bl_111 br_111 wl_23 vdd gnd cell_6t
Xbit_r24_c111 bl_111 br_111 wl_24 vdd gnd cell_6t
Xbit_r25_c111 bl_111 br_111 wl_25 vdd gnd cell_6t
Xbit_r26_c111 bl_111 br_111 wl_26 vdd gnd cell_6t
Xbit_r27_c111 bl_111 br_111 wl_27 vdd gnd cell_6t
Xbit_r28_c111 bl_111 br_111 wl_28 vdd gnd cell_6t
Xbit_r29_c111 bl_111 br_111 wl_29 vdd gnd cell_6t
Xbit_r30_c111 bl_111 br_111 wl_30 vdd gnd cell_6t
Xbit_r31_c111 bl_111 br_111 wl_31 vdd gnd cell_6t
Xbit_r32_c111 bl_111 br_111 wl_32 vdd gnd cell_6t
Xbit_r33_c111 bl_111 br_111 wl_33 vdd gnd cell_6t
Xbit_r34_c111 bl_111 br_111 wl_34 vdd gnd cell_6t
Xbit_r35_c111 bl_111 br_111 wl_35 vdd gnd cell_6t
Xbit_r36_c111 bl_111 br_111 wl_36 vdd gnd cell_6t
Xbit_r37_c111 bl_111 br_111 wl_37 vdd gnd cell_6t
Xbit_r38_c111 bl_111 br_111 wl_38 vdd gnd cell_6t
Xbit_r39_c111 bl_111 br_111 wl_39 vdd gnd cell_6t
Xbit_r40_c111 bl_111 br_111 wl_40 vdd gnd cell_6t
Xbit_r41_c111 bl_111 br_111 wl_41 vdd gnd cell_6t
Xbit_r42_c111 bl_111 br_111 wl_42 vdd gnd cell_6t
Xbit_r43_c111 bl_111 br_111 wl_43 vdd gnd cell_6t
Xbit_r44_c111 bl_111 br_111 wl_44 vdd gnd cell_6t
Xbit_r45_c111 bl_111 br_111 wl_45 vdd gnd cell_6t
Xbit_r46_c111 bl_111 br_111 wl_46 vdd gnd cell_6t
Xbit_r47_c111 bl_111 br_111 wl_47 vdd gnd cell_6t
Xbit_r48_c111 bl_111 br_111 wl_48 vdd gnd cell_6t
Xbit_r49_c111 bl_111 br_111 wl_49 vdd gnd cell_6t
Xbit_r50_c111 bl_111 br_111 wl_50 vdd gnd cell_6t
Xbit_r51_c111 bl_111 br_111 wl_51 vdd gnd cell_6t
Xbit_r52_c111 bl_111 br_111 wl_52 vdd gnd cell_6t
Xbit_r53_c111 bl_111 br_111 wl_53 vdd gnd cell_6t
Xbit_r54_c111 bl_111 br_111 wl_54 vdd gnd cell_6t
Xbit_r55_c111 bl_111 br_111 wl_55 vdd gnd cell_6t
Xbit_r56_c111 bl_111 br_111 wl_56 vdd gnd cell_6t
Xbit_r57_c111 bl_111 br_111 wl_57 vdd gnd cell_6t
Xbit_r58_c111 bl_111 br_111 wl_58 vdd gnd cell_6t
Xbit_r59_c111 bl_111 br_111 wl_59 vdd gnd cell_6t
Xbit_r60_c111 bl_111 br_111 wl_60 vdd gnd cell_6t
Xbit_r61_c111 bl_111 br_111 wl_61 vdd gnd cell_6t
Xbit_r62_c111 bl_111 br_111 wl_62 vdd gnd cell_6t
Xbit_r63_c111 bl_111 br_111 wl_63 vdd gnd cell_6t
Xbit_r64_c111 bl_111 br_111 wl_64 vdd gnd cell_6t
Xbit_r65_c111 bl_111 br_111 wl_65 vdd gnd cell_6t
Xbit_r66_c111 bl_111 br_111 wl_66 vdd gnd cell_6t
Xbit_r67_c111 bl_111 br_111 wl_67 vdd gnd cell_6t
Xbit_r68_c111 bl_111 br_111 wl_68 vdd gnd cell_6t
Xbit_r69_c111 bl_111 br_111 wl_69 vdd gnd cell_6t
Xbit_r70_c111 bl_111 br_111 wl_70 vdd gnd cell_6t
Xbit_r71_c111 bl_111 br_111 wl_71 vdd gnd cell_6t
Xbit_r72_c111 bl_111 br_111 wl_72 vdd gnd cell_6t
Xbit_r73_c111 bl_111 br_111 wl_73 vdd gnd cell_6t
Xbit_r74_c111 bl_111 br_111 wl_74 vdd gnd cell_6t
Xbit_r75_c111 bl_111 br_111 wl_75 vdd gnd cell_6t
Xbit_r76_c111 bl_111 br_111 wl_76 vdd gnd cell_6t
Xbit_r77_c111 bl_111 br_111 wl_77 vdd gnd cell_6t
Xbit_r78_c111 bl_111 br_111 wl_78 vdd gnd cell_6t
Xbit_r79_c111 bl_111 br_111 wl_79 vdd gnd cell_6t
Xbit_r80_c111 bl_111 br_111 wl_80 vdd gnd cell_6t
Xbit_r81_c111 bl_111 br_111 wl_81 vdd gnd cell_6t
Xbit_r82_c111 bl_111 br_111 wl_82 vdd gnd cell_6t
Xbit_r83_c111 bl_111 br_111 wl_83 vdd gnd cell_6t
Xbit_r84_c111 bl_111 br_111 wl_84 vdd gnd cell_6t
Xbit_r85_c111 bl_111 br_111 wl_85 vdd gnd cell_6t
Xbit_r86_c111 bl_111 br_111 wl_86 vdd gnd cell_6t
Xbit_r87_c111 bl_111 br_111 wl_87 vdd gnd cell_6t
Xbit_r88_c111 bl_111 br_111 wl_88 vdd gnd cell_6t
Xbit_r89_c111 bl_111 br_111 wl_89 vdd gnd cell_6t
Xbit_r90_c111 bl_111 br_111 wl_90 vdd gnd cell_6t
Xbit_r91_c111 bl_111 br_111 wl_91 vdd gnd cell_6t
Xbit_r92_c111 bl_111 br_111 wl_92 vdd gnd cell_6t
Xbit_r93_c111 bl_111 br_111 wl_93 vdd gnd cell_6t
Xbit_r94_c111 bl_111 br_111 wl_94 vdd gnd cell_6t
Xbit_r95_c111 bl_111 br_111 wl_95 vdd gnd cell_6t
Xbit_r96_c111 bl_111 br_111 wl_96 vdd gnd cell_6t
Xbit_r97_c111 bl_111 br_111 wl_97 vdd gnd cell_6t
Xbit_r98_c111 bl_111 br_111 wl_98 vdd gnd cell_6t
Xbit_r99_c111 bl_111 br_111 wl_99 vdd gnd cell_6t
Xbit_r100_c111 bl_111 br_111 wl_100 vdd gnd cell_6t
Xbit_r101_c111 bl_111 br_111 wl_101 vdd gnd cell_6t
Xbit_r102_c111 bl_111 br_111 wl_102 vdd gnd cell_6t
Xbit_r103_c111 bl_111 br_111 wl_103 vdd gnd cell_6t
Xbit_r104_c111 bl_111 br_111 wl_104 vdd gnd cell_6t
Xbit_r105_c111 bl_111 br_111 wl_105 vdd gnd cell_6t
Xbit_r106_c111 bl_111 br_111 wl_106 vdd gnd cell_6t
Xbit_r107_c111 bl_111 br_111 wl_107 vdd gnd cell_6t
Xbit_r108_c111 bl_111 br_111 wl_108 vdd gnd cell_6t
Xbit_r109_c111 bl_111 br_111 wl_109 vdd gnd cell_6t
Xbit_r110_c111 bl_111 br_111 wl_110 vdd gnd cell_6t
Xbit_r111_c111 bl_111 br_111 wl_111 vdd gnd cell_6t
Xbit_r112_c111 bl_111 br_111 wl_112 vdd gnd cell_6t
Xbit_r113_c111 bl_111 br_111 wl_113 vdd gnd cell_6t
Xbit_r114_c111 bl_111 br_111 wl_114 vdd gnd cell_6t
Xbit_r115_c111 bl_111 br_111 wl_115 vdd gnd cell_6t
Xbit_r116_c111 bl_111 br_111 wl_116 vdd gnd cell_6t
Xbit_r117_c111 bl_111 br_111 wl_117 vdd gnd cell_6t
Xbit_r118_c111 bl_111 br_111 wl_118 vdd gnd cell_6t
Xbit_r119_c111 bl_111 br_111 wl_119 vdd gnd cell_6t
Xbit_r120_c111 bl_111 br_111 wl_120 vdd gnd cell_6t
Xbit_r121_c111 bl_111 br_111 wl_121 vdd gnd cell_6t
Xbit_r122_c111 bl_111 br_111 wl_122 vdd gnd cell_6t
Xbit_r123_c111 bl_111 br_111 wl_123 vdd gnd cell_6t
Xbit_r124_c111 bl_111 br_111 wl_124 vdd gnd cell_6t
Xbit_r125_c111 bl_111 br_111 wl_125 vdd gnd cell_6t
Xbit_r126_c111 bl_111 br_111 wl_126 vdd gnd cell_6t
Xbit_r127_c111 bl_111 br_111 wl_127 vdd gnd cell_6t
Xbit_r128_c111 bl_111 br_111 wl_128 vdd gnd cell_6t
Xbit_r129_c111 bl_111 br_111 wl_129 vdd gnd cell_6t
Xbit_r130_c111 bl_111 br_111 wl_130 vdd gnd cell_6t
Xbit_r131_c111 bl_111 br_111 wl_131 vdd gnd cell_6t
Xbit_r132_c111 bl_111 br_111 wl_132 vdd gnd cell_6t
Xbit_r133_c111 bl_111 br_111 wl_133 vdd gnd cell_6t
Xbit_r134_c111 bl_111 br_111 wl_134 vdd gnd cell_6t
Xbit_r135_c111 bl_111 br_111 wl_135 vdd gnd cell_6t
Xbit_r136_c111 bl_111 br_111 wl_136 vdd gnd cell_6t
Xbit_r137_c111 bl_111 br_111 wl_137 vdd gnd cell_6t
Xbit_r138_c111 bl_111 br_111 wl_138 vdd gnd cell_6t
Xbit_r139_c111 bl_111 br_111 wl_139 vdd gnd cell_6t
Xbit_r140_c111 bl_111 br_111 wl_140 vdd gnd cell_6t
Xbit_r141_c111 bl_111 br_111 wl_141 vdd gnd cell_6t
Xbit_r142_c111 bl_111 br_111 wl_142 vdd gnd cell_6t
Xbit_r143_c111 bl_111 br_111 wl_143 vdd gnd cell_6t
Xbit_r144_c111 bl_111 br_111 wl_144 vdd gnd cell_6t
Xbit_r145_c111 bl_111 br_111 wl_145 vdd gnd cell_6t
Xbit_r146_c111 bl_111 br_111 wl_146 vdd gnd cell_6t
Xbit_r147_c111 bl_111 br_111 wl_147 vdd gnd cell_6t
Xbit_r148_c111 bl_111 br_111 wl_148 vdd gnd cell_6t
Xbit_r149_c111 bl_111 br_111 wl_149 vdd gnd cell_6t
Xbit_r150_c111 bl_111 br_111 wl_150 vdd gnd cell_6t
Xbit_r151_c111 bl_111 br_111 wl_151 vdd gnd cell_6t
Xbit_r152_c111 bl_111 br_111 wl_152 vdd gnd cell_6t
Xbit_r153_c111 bl_111 br_111 wl_153 vdd gnd cell_6t
Xbit_r154_c111 bl_111 br_111 wl_154 vdd gnd cell_6t
Xbit_r155_c111 bl_111 br_111 wl_155 vdd gnd cell_6t
Xbit_r156_c111 bl_111 br_111 wl_156 vdd gnd cell_6t
Xbit_r157_c111 bl_111 br_111 wl_157 vdd gnd cell_6t
Xbit_r158_c111 bl_111 br_111 wl_158 vdd gnd cell_6t
Xbit_r159_c111 bl_111 br_111 wl_159 vdd gnd cell_6t
Xbit_r160_c111 bl_111 br_111 wl_160 vdd gnd cell_6t
Xbit_r161_c111 bl_111 br_111 wl_161 vdd gnd cell_6t
Xbit_r162_c111 bl_111 br_111 wl_162 vdd gnd cell_6t
Xbit_r163_c111 bl_111 br_111 wl_163 vdd gnd cell_6t
Xbit_r164_c111 bl_111 br_111 wl_164 vdd gnd cell_6t
Xbit_r165_c111 bl_111 br_111 wl_165 vdd gnd cell_6t
Xbit_r166_c111 bl_111 br_111 wl_166 vdd gnd cell_6t
Xbit_r167_c111 bl_111 br_111 wl_167 vdd gnd cell_6t
Xbit_r168_c111 bl_111 br_111 wl_168 vdd gnd cell_6t
Xbit_r169_c111 bl_111 br_111 wl_169 vdd gnd cell_6t
Xbit_r170_c111 bl_111 br_111 wl_170 vdd gnd cell_6t
Xbit_r171_c111 bl_111 br_111 wl_171 vdd gnd cell_6t
Xbit_r172_c111 bl_111 br_111 wl_172 vdd gnd cell_6t
Xbit_r173_c111 bl_111 br_111 wl_173 vdd gnd cell_6t
Xbit_r174_c111 bl_111 br_111 wl_174 vdd gnd cell_6t
Xbit_r175_c111 bl_111 br_111 wl_175 vdd gnd cell_6t
Xbit_r176_c111 bl_111 br_111 wl_176 vdd gnd cell_6t
Xbit_r177_c111 bl_111 br_111 wl_177 vdd gnd cell_6t
Xbit_r178_c111 bl_111 br_111 wl_178 vdd gnd cell_6t
Xbit_r179_c111 bl_111 br_111 wl_179 vdd gnd cell_6t
Xbit_r180_c111 bl_111 br_111 wl_180 vdd gnd cell_6t
Xbit_r181_c111 bl_111 br_111 wl_181 vdd gnd cell_6t
Xbit_r182_c111 bl_111 br_111 wl_182 vdd gnd cell_6t
Xbit_r183_c111 bl_111 br_111 wl_183 vdd gnd cell_6t
Xbit_r184_c111 bl_111 br_111 wl_184 vdd gnd cell_6t
Xbit_r185_c111 bl_111 br_111 wl_185 vdd gnd cell_6t
Xbit_r186_c111 bl_111 br_111 wl_186 vdd gnd cell_6t
Xbit_r187_c111 bl_111 br_111 wl_187 vdd gnd cell_6t
Xbit_r188_c111 bl_111 br_111 wl_188 vdd gnd cell_6t
Xbit_r189_c111 bl_111 br_111 wl_189 vdd gnd cell_6t
Xbit_r190_c111 bl_111 br_111 wl_190 vdd gnd cell_6t
Xbit_r191_c111 bl_111 br_111 wl_191 vdd gnd cell_6t
Xbit_r192_c111 bl_111 br_111 wl_192 vdd gnd cell_6t
Xbit_r193_c111 bl_111 br_111 wl_193 vdd gnd cell_6t
Xbit_r194_c111 bl_111 br_111 wl_194 vdd gnd cell_6t
Xbit_r195_c111 bl_111 br_111 wl_195 vdd gnd cell_6t
Xbit_r196_c111 bl_111 br_111 wl_196 vdd gnd cell_6t
Xbit_r197_c111 bl_111 br_111 wl_197 vdd gnd cell_6t
Xbit_r198_c111 bl_111 br_111 wl_198 vdd gnd cell_6t
Xbit_r199_c111 bl_111 br_111 wl_199 vdd gnd cell_6t
Xbit_r200_c111 bl_111 br_111 wl_200 vdd gnd cell_6t
Xbit_r201_c111 bl_111 br_111 wl_201 vdd gnd cell_6t
Xbit_r202_c111 bl_111 br_111 wl_202 vdd gnd cell_6t
Xbit_r203_c111 bl_111 br_111 wl_203 vdd gnd cell_6t
Xbit_r204_c111 bl_111 br_111 wl_204 vdd gnd cell_6t
Xbit_r205_c111 bl_111 br_111 wl_205 vdd gnd cell_6t
Xbit_r206_c111 bl_111 br_111 wl_206 vdd gnd cell_6t
Xbit_r207_c111 bl_111 br_111 wl_207 vdd gnd cell_6t
Xbit_r208_c111 bl_111 br_111 wl_208 vdd gnd cell_6t
Xbit_r209_c111 bl_111 br_111 wl_209 vdd gnd cell_6t
Xbit_r210_c111 bl_111 br_111 wl_210 vdd gnd cell_6t
Xbit_r211_c111 bl_111 br_111 wl_211 vdd gnd cell_6t
Xbit_r212_c111 bl_111 br_111 wl_212 vdd gnd cell_6t
Xbit_r213_c111 bl_111 br_111 wl_213 vdd gnd cell_6t
Xbit_r214_c111 bl_111 br_111 wl_214 vdd gnd cell_6t
Xbit_r215_c111 bl_111 br_111 wl_215 vdd gnd cell_6t
Xbit_r216_c111 bl_111 br_111 wl_216 vdd gnd cell_6t
Xbit_r217_c111 bl_111 br_111 wl_217 vdd gnd cell_6t
Xbit_r218_c111 bl_111 br_111 wl_218 vdd gnd cell_6t
Xbit_r219_c111 bl_111 br_111 wl_219 vdd gnd cell_6t
Xbit_r220_c111 bl_111 br_111 wl_220 vdd gnd cell_6t
Xbit_r221_c111 bl_111 br_111 wl_221 vdd gnd cell_6t
Xbit_r222_c111 bl_111 br_111 wl_222 vdd gnd cell_6t
Xbit_r223_c111 bl_111 br_111 wl_223 vdd gnd cell_6t
Xbit_r224_c111 bl_111 br_111 wl_224 vdd gnd cell_6t
Xbit_r225_c111 bl_111 br_111 wl_225 vdd gnd cell_6t
Xbit_r226_c111 bl_111 br_111 wl_226 vdd gnd cell_6t
Xbit_r227_c111 bl_111 br_111 wl_227 vdd gnd cell_6t
Xbit_r228_c111 bl_111 br_111 wl_228 vdd gnd cell_6t
Xbit_r229_c111 bl_111 br_111 wl_229 vdd gnd cell_6t
Xbit_r230_c111 bl_111 br_111 wl_230 vdd gnd cell_6t
Xbit_r231_c111 bl_111 br_111 wl_231 vdd gnd cell_6t
Xbit_r232_c111 bl_111 br_111 wl_232 vdd gnd cell_6t
Xbit_r233_c111 bl_111 br_111 wl_233 vdd gnd cell_6t
Xbit_r234_c111 bl_111 br_111 wl_234 vdd gnd cell_6t
Xbit_r235_c111 bl_111 br_111 wl_235 vdd gnd cell_6t
Xbit_r236_c111 bl_111 br_111 wl_236 vdd gnd cell_6t
Xbit_r237_c111 bl_111 br_111 wl_237 vdd gnd cell_6t
Xbit_r238_c111 bl_111 br_111 wl_238 vdd gnd cell_6t
Xbit_r239_c111 bl_111 br_111 wl_239 vdd gnd cell_6t
Xbit_r240_c111 bl_111 br_111 wl_240 vdd gnd cell_6t
Xbit_r241_c111 bl_111 br_111 wl_241 vdd gnd cell_6t
Xbit_r242_c111 bl_111 br_111 wl_242 vdd gnd cell_6t
Xbit_r243_c111 bl_111 br_111 wl_243 vdd gnd cell_6t
Xbit_r244_c111 bl_111 br_111 wl_244 vdd gnd cell_6t
Xbit_r245_c111 bl_111 br_111 wl_245 vdd gnd cell_6t
Xbit_r246_c111 bl_111 br_111 wl_246 vdd gnd cell_6t
Xbit_r247_c111 bl_111 br_111 wl_247 vdd gnd cell_6t
Xbit_r248_c111 bl_111 br_111 wl_248 vdd gnd cell_6t
Xbit_r249_c111 bl_111 br_111 wl_249 vdd gnd cell_6t
Xbit_r250_c111 bl_111 br_111 wl_250 vdd gnd cell_6t
Xbit_r251_c111 bl_111 br_111 wl_251 vdd gnd cell_6t
Xbit_r252_c111 bl_111 br_111 wl_252 vdd gnd cell_6t
Xbit_r253_c111 bl_111 br_111 wl_253 vdd gnd cell_6t
Xbit_r254_c111 bl_111 br_111 wl_254 vdd gnd cell_6t
Xbit_r255_c111 bl_111 br_111 wl_255 vdd gnd cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd cell_6t
Xbit_r1_c112 bl_112 br_112 wl_1 vdd gnd cell_6t
Xbit_r2_c112 bl_112 br_112 wl_2 vdd gnd cell_6t
Xbit_r3_c112 bl_112 br_112 wl_3 vdd gnd cell_6t
Xbit_r4_c112 bl_112 br_112 wl_4 vdd gnd cell_6t
Xbit_r5_c112 bl_112 br_112 wl_5 vdd gnd cell_6t
Xbit_r6_c112 bl_112 br_112 wl_6 vdd gnd cell_6t
Xbit_r7_c112 bl_112 br_112 wl_7 vdd gnd cell_6t
Xbit_r8_c112 bl_112 br_112 wl_8 vdd gnd cell_6t
Xbit_r9_c112 bl_112 br_112 wl_9 vdd gnd cell_6t
Xbit_r10_c112 bl_112 br_112 wl_10 vdd gnd cell_6t
Xbit_r11_c112 bl_112 br_112 wl_11 vdd gnd cell_6t
Xbit_r12_c112 bl_112 br_112 wl_12 vdd gnd cell_6t
Xbit_r13_c112 bl_112 br_112 wl_13 vdd gnd cell_6t
Xbit_r14_c112 bl_112 br_112 wl_14 vdd gnd cell_6t
Xbit_r15_c112 bl_112 br_112 wl_15 vdd gnd cell_6t
Xbit_r16_c112 bl_112 br_112 wl_16 vdd gnd cell_6t
Xbit_r17_c112 bl_112 br_112 wl_17 vdd gnd cell_6t
Xbit_r18_c112 bl_112 br_112 wl_18 vdd gnd cell_6t
Xbit_r19_c112 bl_112 br_112 wl_19 vdd gnd cell_6t
Xbit_r20_c112 bl_112 br_112 wl_20 vdd gnd cell_6t
Xbit_r21_c112 bl_112 br_112 wl_21 vdd gnd cell_6t
Xbit_r22_c112 bl_112 br_112 wl_22 vdd gnd cell_6t
Xbit_r23_c112 bl_112 br_112 wl_23 vdd gnd cell_6t
Xbit_r24_c112 bl_112 br_112 wl_24 vdd gnd cell_6t
Xbit_r25_c112 bl_112 br_112 wl_25 vdd gnd cell_6t
Xbit_r26_c112 bl_112 br_112 wl_26 vdd gnd cell_6t
Xbit_r27_c112 bl_112 br_112 wl_27 vdd gnd cell_6t
Xbit_r28_c112 bl_112 br_112 wl_28 vdd gnd cell_6t
Xbit_r29_c112 bl_112 br_112 wl_29 vdd gnd cell_6t
Xbit_r30_c112 bl_112 br_112 wl_30 vdd gnd cell_6t
Xbit_r31_c112 bl_112 br_112 wl_31 vdd gnd cell_6t
Xbit_r32_c112 bl_112 br_112 wl_32 vdd gnd cell_6t
Xbit_r33_c112 bl_112 br_112 wl_33 vdd gnd cell_6t
Xbit_r34_c112 bl_112 br_112 wl_34 vdd gnd cell_6t
Xbit_r35_c112 bl_112 br_112 wl_35 vdd gnd cell_6t
Xbit_r36_c112 bl_112 br_112 wl_36 vdd gnd cell_6t
Xbit_r37_c112 bl_112 br_112 wl_37 vdd gnd cell_6t
Xbit_r38_c112 bl_112 br_112 wl_38 vdd gnd cell_6t
Xbit_r39_c112 bl_112 br_112 wl_39 vdd gnd cell_6t
Xbit_r40_c112 bl_112 br_112 wl_40 vdd gnd cell_6t
Xbit_r41_c112 bl_112 br_112 wl_41 vdd gnd cell_6t
Xbit_r42_c112 bl_112 br_112 wl_42 vdd gnd cell_6t
Xbit_r43_c112 bl_112 br_112 wl_43 vdd gnd cell_6t
Xbit_r44_c112 bl_112 br_112 wl_44 vdd gnd cell_6t
Xbit_r45_c112 bl_112 br_112 wl_45 vdd gnd cell_6t
Xbit_r46_c112 bl_112 br_112 wl_46 vdd gnd cell_6t
Xbit_r47_c112 bl_112 br_112 wl_47 vdd gnd cell_6t
Xbit_r48_c112 bl_112 br_112 wl_48 vdd gnd cell_6t
Xbit_r49_c112 bl_112 br_112 wl_49 vdd gnd cell_6t
Xbit_r50_c112 bl_112 br_112 wl_50 vdd gnd cell_6t
Xbit_r51_c112 bl_112 br_112 wl_51 vdd gnd cell_6t
Xbit_r52_c112 bl_112 br_112 wl_52 vdd gnd cell_6t
Xbit_r53_c112 bl_112 br_112 wl_53 vdd gnd cell_6t
Xbit_r54_c112 bl_112 br_112 wl_54 vdd gnd cell_6t
Xbit_r55_c112 bl_112 br_112 wl_55 vdd gnd cell_6t
Xbit_r56_c112 bl_112 br_112 wl_56 vdd gnd cell_6t
Xbit_r57_c112 bl_112 br_112 wl_57 vdd gnd cell_6t
Xbit_r58_c112 bl_112 br_112 wl_58 vdd gnd cell_6t
Xbit_r59_c112 bl_112 br_112 wl_59 vdd gnd cell_6t
Xbit_r60_c112 bl_112 br_112 wl_60 vdd gnd cell_6t
Xbit_r61_c112 bl_112 br_112 wl_61 vdd gnd cell_6t
Xbit_r62_c112 bl_112 br_112 wl_62 vdd gnd cell_6t
Xbit_r63_c112 bl_112 br_112 wl_63 vdd gnd cell_6t
Xbit_r64_c112 bl_112 br_112 wl_64 vdd gnd cell_6t
Xbit_r65_c112 bl_112 br_112 wl_65 vdd gnd cell_6t
Xbit_r66_c112 bl_112 br_112 wl_66 vdd gnd cell_6t
Xbit_r67_c112 bl_112 br_112 wl_67 vdd gnd cell_6t
Xbit_r68_c112 bl_112 br_112 wl_68 vdd gnd cell_6t
Xbit_r69_c112 bl_112 br_112 wl_69 vdd gnd cell_6t
Xbit_r70_c112 bl_112 br_112 wl_70 vdd gnd cell_6t
Xbit_r71_c112 bl_112 br_112 wl_71 vdd gnd cell_6t
Xbit_r72_c112 bl_112 br_112 wl_72 vdd gnd cell_6t
Xbit_r73_c112 bl_112 br_112 wl_73 vdd gnd cell_6t
Xbit_r74_c112 bl_112 br_112 wl_74 vdd gnd cell_6t
Xbit_r75_c112 bl_112 br_112 wl_75 vdd gnd cell_6t
Xbit_r76_c112 bl_112 br_112 wl_76 vdd gnd cell_6t
Xbit_r77_c112 bl_112 br_112 wl_77 vdd gnd cell_6t
Xbit_r78_c112 bl_112 br_112 wl_78 vdd gnd cell_6t
Xbit_r79_c112 bl_112 br_112 wl_79 vdd gnd cell_6t
Xbit_r80_c112 bl_112 br_112 wl_80 vdd gnd cell_6t
Xbit_r81_c112 bl_112 br_112 wl_81 vdd gnd cell_6t
Xbit_r82_c112 bl_112 br_112 wl_82 vdd gnd cell_6t
Xbit_r83_c112 bl_112 br_112 wl_83 vdd gnd cell_6t
Xbit_r84_c112 bl_112 br_112 wl_84 vdd gnd cell_6t
Xbit_r85_c112 bl_112 br_112 wl_85 vdd gnd cell_6t
Xbit_r86_c112 bl_112 br_112 wl_86 vdd gnd cell_6t
Xbit_r87_c112 bl_112 br_112 wl_87 vdd gnd cell_6t
Xbit_r88_c112 bl_112 br_112 wl_88 vdd gnd cell_6t
Xbit_r89_c112 bl_112 br_112 wl_89 vdd gnd cell_6t
Xbit_r90_c112 bl_112 br_112 wl_90 vdd gnd cell_6t
Xbit_r91_c112 bl_112 br_112 wl_91 vdd gnd cell_6t
Xbit_r92_c112 bl_112 br_112 wl_92 vdd gnd cell_6t
Xbit_r93_c112 bl_112 br_112 wl_93 vdd gnd cell_6t
Xbit_r94_c112 bl_112 br_112 wl_94 vdd gnd cell_6t
Xbit_r95_c112 bl_112 br_112 wl_95 vdd gnd cell_6t
Xbit_r96_c112 bl_112 br_112 wl_96 vdd gnd cell_6t
Xbit_r97_c112 bl_112 br_112 wl_97 vdd gnd cell_6t
Xbit_r98_c112 bl_112 br_112 wl_98 vdd gnd cell_6t
Xbit_r99_c112 bl_112 br_112 wl_99 vdd gnd cell_6t
Xbit_r100_c112 bl_112 br_112 wl_100 vdd gnd cell_6t
Xbit_r101_c112 bl_112 br_112 wl_101 vdd gnd cell_6t
Xbit_r102_c112 bl_112 br_112 wl_102 vdd gnd cell_6t
Xbit_r103_c112 bl_112 br_112 wl_103 vdd gnd cell_6t
Xbit_r104_c112 bl_112 br_112 wl_104 vdd gnd cell_6t
Xbit_r105_c112 bl_112 br_112 wl_105 vdd gnd cell_6t
Xbit_r106_c112 bl_112 br_112 wl_106 vdd gnd cell_6t
Xbit_r107_c112 bl_112 br_112 wl_107 vdd gnd cell_6t
Xbit_r108_c112 bl_112 br_112 wl_108 vdd gnd cell_6t
Xbit_r109_c112 bl_112 br_112 wl_109 vdd gnd cell_6t
Xbit_r110_c112 bl_112 br_112 wl_110 vdd gnd cell_6t
Xbit_r111_c112 bl_112 br_112 wl_111 vdd gnd cell_6t
Xbit_r112_c112 bl_112 br_112 wl_112 vdd gnd cell_6t
Xbit_r113_c112 bl_112 br_112 wl_113 vdd gnd cell_6t
Xbit_r114_c112 bl_112 br_112 wl_114 vdd gnd cell_6t
Xbit_r115_c112 bl_112 br_112 wl_115 vdd gnd cell_6t
Xbit_r116_c112 bl_112 br_112 wl_116 vdd gnd cell_6t
Xbit_r117_c112 bl_112 br_112 wl_117 vdd gnd cell_6t
Xbit_r118_c112 bl_112 br_112 wl_118 vdd gnd cell_6t
Xbit_r119_c112 bl_112 br_112 wl_119 vdd gnd cell_6t
Xbit_r120_c112 bl_112 br_112 wl_120 vdd gnd cell_6t
Xbit_r121_c112 bl_112 br_112 wl_121 vdd gnd cell_6t
Xbit_r122_c112 bl_112 br_112 wl_122 vdd gnd cell_6t
Xbit_r123_c112 bl_112 br_112 wl_123 vdd gnd cell_6t
Xbit_r124_c112 bl_112 br_112 wl_124 vdd gnd cell_6t
Xbit_r125_c112 bl_112 br_112 wl_125 vdd gnd cell_6t
Xbit_r126_c112 bl_112 br_112 wl_126 vdd gnd cell_6t
Xbit_r127_c112 bl_112 br_112 wl_127 vdd gnd cell_6t
Xbit_r128_c112 bl_112 br_112 wl_128 vdd gnd cell_6t
Xbit_r129_c112 bl_112 br_112 wl_129 vdd gnd cell_6t
Xbit_r130_c112 bl_112 br_112 wl_130 vdd gnd cell_6t
Xbit_r131_c112 bl_112 br_112 wl_131 vdd gnd cell_6t
Xbit_r132_c112 bl_112 br_112 wl_132 vdd gnd cell_6t
Xbit_r133_c112 bl_112 br_112 wl_133 vdd gnd cell_6t
Xbit_r134_c112 bl_112 br_112 wl_134 vdd gnd cell_6t
Xbit_r135_c112 bl_112 br_112 wl_135 vdd gnd cell_6t
Xbit_r136_c112 bl_112 br_112 wl_136 vdd gnd cell_6t
Xbit_r137_c112 bl_112 br_112 wl_137 vdd gnd cell_6t
Xbit_r138_c112 bl_112 br_112 wl_138 vdd gnd cell_6t
Xbit_r139_c112 bl_112 br_112 wl_139 vdd gnd cell_6t
Xbit_r140_c112 bl_112 br_112 wl_140 vdd gnd cell_6t
Xbit_r141_c112 bl_112 br_112 wl_141 vdd gnd cell_6t
Xbit_r142_c112 bl_112 br_112 wl_142 vdd gnd cell_6t
Xbit_r143_c112 bl_112 br_112 wl_143 vdd gnd cell_6t
Xbit_r144_c112 bl_112 br_112 wl_144 vdd gnd cell_6t
Xbit_r145_c112 bl_112 br_112 wl_145 vdd gnd cell_6t
Xbit_r146_c112 bl_112 br_112 wl_146 vdd gnd cell_6t
Xbit_r147_c112 bl_112 br_112 wl_147 vdd gnd cell_6t
Xbit_r148_c112 bl_112 br_112 wl_148 vdd gnd cell_6t
Xbit_r149_c112 bl_112 br_112 wl_149 vdd gnd cell_6t
Xbit_r150_c112 bl_112 br_112 wl_150 vdd gnd cell_6t
Xbit_r151_c112 bl_112 br_112 wl_151 vdd gnd cell_6t
Xbit_r152_c112 bl_112 br_112 wl_152 vdd gnd cell_6t
Xbit_r153_c112 bl_112 br_112 wl_153 vdd gnd cell_6t
Xbit_r154_c112 bl_112 br_112 wl_154 vdd gnd cell_6t
Xbit_r155_c112 bl_112 br_112 wl_155 vdd gnd cell_6t
Xbit_r156_c112 bl_112 br_112 wl_156 vdd gnd cell_6t
Xbit_r157_c112 bl_112 br_112 wl_157 vdd gnd cell_6t
Xbit_r158_c112 bl_112 br_112 wl_158 vdd gnd cell_6t
Xbit_r159_c112 bl_112 br_112 wl_159 vdd gnd cell_6t
Xbit_r160_c112 bl_112 br_112 wl_160 vdd gnd cell_6t
Xbit_r161_c112 bl_112 br_112 wl_161 vdd gnd cell_6t
Xbit_r162_c112 bl_112 br_112 wl_162 vdd gnd cell_6t
Xbit_r163_c112 bl_112 br_112 wl_163 vdd gnd cell_6t
Xbit_r164_c112 bl_112 br_112 wl_164 vdd gnd cell_6t
Xbit_r165_c112 bl_112 br_112 wl_165 vdd gnd cell_6t
Xbit_r166_c112 bl_112 br_112 wl_166 vdd gnd cell_6t
Xbit_r167_c112 bl_112 br_112 wl_167 vdd gnd cell_6t
Xbit_r168_c112 bl_112 br_112 wl_168 vdd gnd cell_6t
Xbit_r169_c112 bl_112 br_112 wl_169 vdd gnd cell_6t
Xbit_r170_c112 bl_112 br_112 wl_170 vdd gnd cell_6t
Xbit_r171_c112 bl_112 br_112 wl_171 vdd gnd cell_6t
Xbit_r172_c112 bl_112 br_112 wl_172 vdd gnd cell_6t
Xbit_r173_c112 bl_112 br_112 wl_173 vdd gnd cell_6t
Xbit_r174_c112 bl_112 br_112 wl_174 vdd gnd cell_6t
Xbit_r175_c112 bl_112 br_112 wl_175 vdd gnd cell_6t
Xbit_r176_c112 bl_112 br_112 wl_176 vdd gnd cell_6t
Xbit_r177_c112 bl_112 br_112 wl_177 vdd gnd cell_6t
Xbit_r178_c112 bl_112 br_112 wl_178 vdd gnd cell_6t
Xbit_r179_c112 bl_112 br_112 wl_179 vdd gnd cell_6t
Xbit_r180_c112 bl_112 br_112 wl_180 vdd gnd cell_6t
Xbit_r181_c112 bl_112 br_112 wl_181 vdd gnd cell_6t
Xbit_r182_c112 bl_112 br_112 wl_182 vdd gnd cell_6t
Xbit_r183_c112 bl_112 br_112 wl_183 vdd gnd cell_6t
Xbit_r184_c112 bl_112 br_112 wl_184 vdd gnd cell_6t
Xbit_r185_c112 bl_112 br_112 wl_185 vdd gnd cell_6t
Xbit_r186_c112 bl_112 br_112 wl_186 vdd gnd cell_6t
Xbit_r187_c112 bl_112 br_112 wl_187 vdd gnd cell_6t
Xbit_r188_c112 bl_112 br_112 wl_188 vdd gnd cell_6t
Xbit_r189_c112 bl_112 br_112 wl_189 vdd gnd cell_6t
Xbit_r190_c112 bl_112 br_112 wl_190 vdd gnd cell_6t
Xbit_r191_c112 bl_112 br_112 wl_191 vdd gnd cell_6t
Xbit_r192_c112 bl_112 br_112 wl_192 vdd gnd cell_6t
Xbit_r193_c112 bl_112 br_112 wl_193 vdd gnd cell_6t
Xbit_r194_c112 bl_112 br_112 wl_194 vdd gnd cell_6t
Xbit_r195_c112 bl_112 br_112 wl_195 vdd gnd cell_6t
Xbit_r196_c112 bl_112 br_112 wl_196 vdd gnd cell_6t
Xbit_r197_c112 bl_112 br_112 wl_197 vdd gnd cell_6t
Xbit_r198_c112 bl_112 br_112 wl_198 vdd gnd cell_6t
Xbit_r199_c112 bl_112 br_112 wl_199 vdd gnd cell_6t
Xbit_r200_c112 bl_112 br_112 wl_200 vdd gnd cell_6t
Xbit_r201_c112 bl_112 br_112 wl_201 vdd gnd cell_6t
Xbit_r202_c112 bl_112 br_112 wl_202 vdd gnd cell_6t
Xbit_r203_c112 bl_112 br_112 wl_203 vdd gnd cell_6t
Xbit_r204_c112 bl_112 br_112 wl_204 vdd gnd cell_6t
Xbit_r205_c112 bl_112 br_112 wl_205 vdd gnd cell_6t
Xbit_r206_c112 bl_112 br_112 wl_206 vdd gnd cell_6t
Xbit_r207_c112 bl_112 br_112 wl_207 vdd gnd cell_6t
Xbit_r208_c112 bl_112 br_112 wl_208 vdd gnd cell_6t
Xbit_r209_c112 bl_112 br_112 wl_209 vdd gnd cell_6t
Xbit_r210_c112 bl_112 br_112 wl_210 vdd gnd cell_6t
Xbit_r211_c112 bl_112 br_112 wl_211 vdd gnd cell_6t
Xbit_r212_c112 bl_112 br_112 wl_212 vdd gnd cell_6t
Xbit_r213_c112 bl_112 br_112 wl_213 vdd gnd cell_6t
Xbit_r214_c112 bl_112 br_112 wl_214 vdd gnd cell_6t
Xbit_r215_c112 bl_112 br_112 wl_215 vdd gnd cell_6t
Xbit_r216_c112 bl_112 br_112 wl_216 vdd gnd cell_6t
Xbit_r217_c112 bl_112 br_112 wl_217 vdd gnd cell_6t
Xbit_r218_c112 bl_112 br_112 wl_218 vdd gnd cell_6t
Xbit_r219_c112 bl_112 br_112 wl_219 vdd gnd cell_6t
Xbit_r220_c112 bl_112 br_112 wl_220 vdd gnd cell_6t
Xbit_r221_c112 bl_112 br_112 wl_221 vdd gnd cell_6t
Xbit_r222_c112 bl_112 br_112 wl_222 vdd gnd cell_6t
Xbit_r223_c112 bl_112 br_112 wl_223 vdd gnd cell_6t
Xbit_r224_c112 bl_112 br_112 wl_224 vdd gnd cell_6t
Xbit_r225_c112 bl_112 br_112 wl_225 vdd gnd cell_6t
Xbit_r226_c112 bl_112 br_112 wl_226 vdd gnd cell_6t
Xbit_r227_c112 bl_112 br_112 wl_227 vdd gnd cell_6t
Xbit_r228_c112 bl_112 br_112 wl_228 vdd gnd cell_6t
Xbit_r229_c112 bl_112 br_112 wl_229 vdd gnd cell_6t
Xbit_r230_c112 bl_112 br_112 wl_230 vdd gnd cell_6t
Xbit_r231_c112 bl_112 br_112 wl_231 vdd gnd cell_6t
Xbit_r232_c112 bl_112 br_112 wl_232 vdd gnd cell_6t
Xbit_r233_c112 bl_112 br_112 wl_233 vdd gnd cell_6t
Xbit_r234_c112 bl_112 br_112 wl_234 vdd gnd cell_6t
Xbit_r235_c112 bl_112 br_112 wl_235 vdd gnd cell_6t
Xbit_r236_c112 bl_112 br_112 wl_236 vdd gnd cell_6t
Xbit_r237_c112 bl_112 br_112 wl_237 vdd gnd cell_6t
Xbit_r238_c112 bl_112 br_112 wl_238 vdd gnd cell_6t
Xbit_r239_c112 bl_112 br_112 wl_239 vdd gnd cell_6t
Xbit_r240_c112 bl_112 br_112 wl_240 vdd gnd cell_6t
Xbit_r241_c112 bl_112 br_112 wl_241 vdd gnd cell_6t
Xbit_r242_c112 bl_112 br_112 wl_242 vdd gnd cell_6t
Xbit_r243_c112 bl_112 br_112 wl_243 vdd gnd cell_6t
Xbit_r244_c112 bl_112 br_112 wl_244 vdd gnd cell_6t
Xbit_r245_c112 bl_112 br_112 wl_245 vdd gnd cell_6t
Xbit_r246_c112 bl_112 br_112 wl_246 vdd gnd cell_6t
Xbit_r247_c112 bl_112 br_112 wl_247 vdd gnd cell_6t
Xbit_r248_c112 bl_112 br_112 wl_248 vdd gnd cell_6t
Xbit_r249_c112 bl_112 br_112 wl_249 vdd gnd cell_6t
Xbit_r250_c112 bl_112 br_112 wl_250 vdd gnd cell_6t
Xbit_r251_c112 bl_112 br_112 wl_251 vdd gnd cell_6t
Xbit_r252_c112 bl_112 br_112 wl_252 vdd gnd cell_6t
Xbit_r253_c112 bl_112 br_112 wl_253 vdd gnd cell_6t
Xbit_r254_c112 bl_112 br_112 wl_254 vdd gnd cell_6t
Xbit_r255_c112 bl_112 br_112 wl_255 vdd gnd cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd cell_6t
Xbit_r1_c113 bl_113 br_113 wl_1 vdd gnd cell_6t
Xbit_r2_c113 bl_113 br_113 wl_2 vdd gnd cell_6t
Xbit_r3_c113 bl_113 br_113 wl_3 vdd gnd cell_6t
Xbit_r4_c113 bl_113 br_113 wl_4 vdd gnd cell_6t
Xbit_r5_c113 bl_113 br_113 wl_5 vdd gnd cell_6t
Xbit_r6_c113 bl_113 br_113 wl_6 vdd gnd cell_6t
Xbit_r7_c113 bl_113 br_113 wl_7 vdd gnd cell_6t
Xbit_r8_c113 bl_113 br_113 wl_8 vdd gnd cell_6t
Xbit_r9_c113 bl_113 br_113 wl_9 vdd gnd cell_6t
Xbit_r10_c113 bl_113 br_113 wl_10 vdd gnd cell_6t
Xbit_r11_c113 bl_113 br_113 wl_11 vdd gnd cell_6t
Xbit_r12_c113 bl_113 br_113 wl_12 vdd gnd cell_6t
Xbit_r13_c113 bl_113 br_113 wl_13 vdd gnd cell_6t
Xbit_r14_c113 bl_113 br_113 wl_14 vdd gnd cell_6t
Xbit_r15_c113 bl_113 br_113 wl_15 vdd gnd cell_6t
Xbit_r16_c113 bl_113 br_113 wl_16 vdd gnd cell_6t
Xbit_r17_c113 bl_113 br_113 wl_17 vdd gnd cell_6t
Xbit_r18_c113 bl_113 br_113 wl_18 vdd gnd cell_6t
Xbit_r19_c113 bl_113 br_113 wl_19 vdd gnd cell_6t
Xbit_r20_c113 bl_113 br_113 wl_20 vdd gnd cell_6t
Xbit_r21_c113 bl_113 br_113 wl_21 vdd gnd cell_6t
Xbit_r22_c113 bl_113 br_113 wl_22 vdd gnd cell_6t
Xbit_r23_c113 bl_113 br_113 wl_23 vdd gnd cell_6t
Xbit_r24_c113 bl_113 br_113 wl_24 vdd gnd cell_6t
Xbit_r25_c113 bl_113 br_113 wl_25 vdd gnd cell_6t
Xbit_r26_c113 bl_113 br_113 wl_26 vdd gnd cell_6t
Xbit_r27_c113 bl_113 br_113 wl_27 vdd gnd cell_6t
Xbit_r28_c113 bl_113 br_113 wl_28 vdd gnd cell_6t
Xbit_r29_c113 bl_113 br_113 wl_29 vdd gnd cell_6t
Xbit_r30_c113 bl_113 br_113 wl_30 vdd gnd cell_6t
Xbit_r31_c113 bl_113 br_113 wl_31 vdd gnd cell_6t
Xbit_r32_c113 bl_113 br_113 wl_32 vdd gnd cell_6t
Xbit_r33_c113 bl_113 br_113 wl_33 vdd gnd cell_6t
Xbit_r34_c113 bl_113 br_113 wl_34 vdd gnd cell_6t
Xbit_r35_c113 bl_113 br_113 wl_35 vdd gnd cell_6t
Xbit_r36_c113 bl_113 br_113 wl_36 vdd gnd cell_6t
Xbit_r37_c113 bl_113 br_113 wl_37 vdd gnd cell_6t
Xbit_r38_c113 bl_113 br_113 wl_38 vdd gnd cell_6t
Xbit_r39_c113 bl_113 br_113 wl_39 vdd gnd cell_6t
Xbit_r40_c113 bl_113 br_113 wl_40 vdd gnd cell_6t
Xbit_r41_c113 bl_113 br_113 wl_41 vdd gnd cell_6t
Xbit_r42_c113 bl_113 br_113 wl_42 vdd gnd cell_6t
Xbit_r43_c113 bl_113 br_113 wl_43 vdd gnd cell_6t
Xbit_r44_c113 bl_113 br_113 wl_44 vdd gnd cell_6t
Xbit_r45_c113 bl_113 br_113 wl_45 vdd gnd cell_6t
Xbit_r46_c113 bl_113 br_113 wl_46 vdd gnd cell_6t
Xbit_r47_c113 bl_113 br_113 wl_47 vdd gnd cell_6t
Xbit_r48_c113 bl_113 br_113 wl_48 vdd gnd cell_6t
Xbit_r49_c113 bl_113 br_113 wl_49 vdd gnd cell_6t
Xbit_r50_c113 bl_113 br_113 wl_50 vdd gnd cell_6t
Xbit_r51_c113 bl_113 br_113 wl_51 vdd gnd cell_6t
Xbit_r52_c113 bl_113 br_113 wl_52 vdd gnd cell_6t
Xbit_r53_c113 bl_113 br_113 wl_53 vdd gnd cell_6t
Xbit_r54_c113 bl_113 br_113 wl_54 vdd gnd cell_6t
Xbit_r55_c113 bl_113 br_113 wl_55 vdd gnd cell_6t
Xbit_r56_c113 bl_113 br_113 wl_56 vdd gnd cell_6t
Xbit_r57_c113 bl_113 br_113 wl_57 vdd gnd cell_6t
Xbit_r58_c113 bl_113 br_113 wl_58 vdd gnd cell_6t
Xbit_r59_c113 bl_113 br_113 wl_59 vdd gnd cell_6t
Xbit_r60_c113 bl_113 br_113 wl_60 vdd gnd cell_6t
Xbit_r61_c113 bl_113 br_113 wl_61 vdd gnd cell_6t
Xbit_r62_c113 bl_113 br_113 wl_62 vdd gnd cell_6t
Xbit_r63_c113 bl_113 br_113 wl_63 vdd gnd cell_6t
Xbit_r64_c113 bl_113 br_113 wl_64 vdd gnd cell_6t
Xbit_r65_c113 bl_113 br_113 wl_65 vdd gnd cell_6t
Xbit_r66_c113 bl_113 br_113 wl_66 vdd gnd cell_6t
Xbit_r67_c113 bl_113 br_113 wl_67 vdd gnd cell_6t
Xbit_r68_c113 bl_113 br_113 wl_68 vdd gnd cell_6t
Xbit_r69_c113 bl_113 br_113 wl_69 vdd gnd cell_6t
Xbit_r70_c113 bl_113 br_113 wl_70 vdd gnd cell_6t
Xbit_r71_c113 bl_113 br_113 wl_71 vdd gnd cell_6t
Xbit_r72_c113 bl_113 br_113 wl_72 vdd gnd cell_6t
Xbit_r73_c113 bl_113 br_113 wl_73 vdd gnd cell_6t
Xbit_r74_c113 bl_113 br_113 wl_74 vdd gnd cell_6t
Xbit_r75_c113 bl_113 br_113 wl_75 vdd gnd cell_6t
Xbit_r76_c113 bl_113 br_113 wl_76 vdd gnd cell_6t
Xbit_r77_c113 bl_113 br_113 wl_77 vdd gnd cell_6t
Xbit_r78_c113 bl_113 br_113 wl_78 vdd gnd cell_6t
Xbit_r79_c113 bl_113 br_113 wl_79 vdd gnd cell_6t
Xbit_r80_c113 bl_113 br_113 wl_80 vdd gnd cell_6t
Xbit_r81_c113 bl_113 br_113 wl_81 vdd gnd cell_6t
Xbit_r82_c113 bl_113 br_113 wl_82 vdd gnd cell_6t
Xbit_r83_c113 bl_113 br_113 wl_83 vdd gnd cell_6t
Xbit_r84_c113 bl_113 br_113 wl_84 vdd gnd cell_6t
Xbit_r85_c113 bl_113 br_113 wl_85 vdd gnd cell_6t
Xbit_r86_c113 bl_113 br_113 wl_86 vdd gnd cell_6t
Xbit_r87_c113 bl_113 br_113 wl_87 vdd gnd cell_6t
Xbit_r88_c113 bl_113 br_113 wl_88 vdd gnd cell_6t
Xbit_r89_c113 bl_113 br_113 wl_89 vdd gnd cell_6t
Xbit_r90_c113 bl_113 br_113 wl_90 vdd gnd cell_6t
Xbit_r91_c113 bl_113 br_113 wl_91 vdd gnd cell_6t
Xbit_r92_c113 bl_113 br_113 wl_92 vdd gnd cell_6t
Xbit_r93_c113 bl_113 br_113 wl_93 vdd gnd cell_6t
Xbit_r94_c113 bl_113 br_113 wl_94 vdd gnd cell_6t
Xbit_r95_c113 bl_113 br_113 wl_95 vdd gnd cell_6t
Xbit_r96_c113 bl_113 br_113 wl_96 vdd gnd cell_6t
Xbit_r97_c113 bl_113 br_113 wl_97 vdd gnd cell_6t
Xbit_r98_c113 bl_113 br_113 wl_98 vdd gnd cell_6t
Xbit_r99_c113 bl_113 br_113 wl_99 vdd gnd cell_6t
Xbit_r100_c113 bl_113 br_113 wl_100 vdd gnd cell_6t
Xbit_r101_c113 bl_113 br_113 wl_101 vdd gnd cell_6t
Xbit_r102_c113 bl_113 br_113 wl_102 vdd gnd cell_6t
Xbit_r103_c113 bl_113 br_113 wl_103 vdd gnd cell_6t
Xbit_r104_c113 bl_113 br_113 wl_104 vdd gnd cell_6t
Xbit_r105_c113 bl_113 br_113 wl_105 vdd gnd cell_6t
Xbit_r106_c113 bl_113 br_113 wl_106 vdd gnd cell_6t
Xbit_r107_c113 bl_113 br_113 wl_107 vdd gnd cell_6t
Xbit_r108_c113 bl_113 br_113 wl_108 vdd gnd cell_6t
Xbit_r109_c113 bl_113 br_113 wl_109 vdd gnd cell_6t
Xbit_r110_c113 bl_113 br_113 wl_110 vdd gnd cell_6t
Xbit_r111_c113 bl_113 br_113 wl_111 vdd gnd cell_6t
Xbit_r112_c113 bl_113 br_113 wl_112 vdd gnd cell_6t
Xbit_r113_c113 bl_113 br_113 wl_113 vdd gnd cell_6t
Xbit_r114_c113 bl_113 br_113 wl_114 vdd gnd cell_6t
Xbit_r115_c113 bl_113 br_113 wl_115 vdd gnd cell_6t
Xbit_r116_c113 bl_113 br_113 wl_116 vdd gnd cell_6t
Xbit_r117_c113 bl_113 br_113 wl_117 vdd gnd cell_6t
Xbit_r118_c113 bl_113 br_113 wl_118 vdd gnd cell_6t
Xbit_r119_c113 bl_113 br_113 wl_119 vdd gnd cell_6t
Xbit_r120_c113 bl_113 br_113 wl_120 vdd gnd cell_6t
Xbit_r121_c113 bl_113 br_113 wl_121 vdd gnd cell_6t
Xbit_r122_c113 bl_113 br_113 wl_122 vdd gnd cell_6t
Xbit_r123_c113 bl_113 br_113 wl_123 vdd gnd cell_6t
Xbit_r124_c113 bl_113 br_113 wl_124 vdd gnd cell_6t
Xbit_r125_c113 bl_113 br_113 wl_125 vdd gnd cell_6t
Xbit_r126_c113 bl_113 br_113 wl_126 vdd gnd cell_6t
Xbit_r127_c113 bl_113 br_113 wl_127 vdd gnd cell_6t
Xbit_r128_c113 bl_113 br_113 wl_128 vdd gnd cell_6t
Xbit_r129_c113 bl_113 br_113 wl_129 vdd gnd cell_6t
Xbit_r130_c113 bl_113 br_113 wl_130 vdd gnd cell_6t
Xbit_r131_c113 bl_113 br_113 wl_131 vdd gnd cell_6t
Xbit_r132_c113 bl_113 br_113 wl_132 vdd gnd cell_6t
Xbit_r133_c113 bl_113 br_113 wl_133 vdd gnd cell_6t
Xbit_r134_c113 bl_113 br_113 wl_134 vdd gnd cell_6t
Xbit_r135_c113 bl_113 br_113 wl_135 vdd gnd cell_6t
Xbit_r136_c113 bl_113 br_113 wl_136 vdd gnd cell_6t
Xbit_r137_c113 bl_113 br_113 wl_137 vdd gnd cell_6t
Xbit_r138_c113 bl_113 br_113 wl_138 vdd gnd cell_6t
Xbit_r139_c113 bl_113 br_113 wl_139 vdd gnd cell_6t
Xbit_r140_c113 bl_113 br_113 wl_140 vdd gnd cell_6t
Xbit_r141_c113 bl_113 br_113 wl_141 vdd gnd cell_6t
Xbit_r142_c113 bl_113 br_113 wl_142 vdd gnd cell_6t
Xbit_r143_c113 bl_113 br_113 wl_143 vdd gnd cell_6t
Xbit_r144_c113 bl_113 br_113 wl_144 vdd gnd cell_6t
Xbit_r145_c113 bl_113 br_113 wl_145 vdd gnd cell_6t
Xbit_r146_c113 bl_113 br_113 wl_146 vdd gnd cell_6t
Xbit_r147_c113 bl_113 br_113 wl_147 vdd gnd cell_6t
Xbit_r148_c113 bl_113 br_113 wl_148 vdd gnd cell_6t
Xbit_r149_c113 bl_113 br_113 wl_149 vdd gnd cell_6t
Xbit_r150_c113 bl_113 br_113 wl_150 vdd gnd cell_6t
Xbit_r151_c113 bl_113 br_113 wl_151 vdd gnd cell_6t
Xbit_r152_c113 bl_113 br_113 wl_152 vdd gnd cell_6t
Xbit_r153_c113 bl_113 br_113 wl_153 vdd gnd cell_6t
Xbit_r154_c113 bl_113 br_113 wl_154 vdd gnd cell_6t
Xbit_r155_c113 bl_113 br_113 wl_155 vdd gnd cell_6t
Xbit_r156_c113 bl_113 br_113 wl_156 vdd gnd cell_6t
Xbit_r157_c113 bl_113 br_113 wl_157 vdd gnd cell_6t
Xbit_r158_c113 bl_113 br_113 wl_158 vdd gnd cell_6t
Xbit_r159_c113 bl_113 br_113 wl_159 vdd gnd cell_6t
Xbit_r160_c113 bl_113 br_113 wl_160 vdd gnd cell_6t
Xbit_r161_c113 bl_113 br_113 wl_161 vdd gnd cell_6t
Xbit_r162_c113 bl_113 br_113 wl_162 vdd gnd cell_6t
Xbit_r163_c113 bl_113 br_113 wl_163 vdd gnd cell_6t
Xbit_r164_c113 bl_113 br_113 wl_164 vdd gnd cell_6t
Xbit_r165_c113 bl_113 br_113 wl_165 vdd gnd cell_6t
Xbit_r166_c113 bl_113 br_113 wl_166 vdd gnd cell_6t
Xbit_r167_c113 bl_113 br_113 wl_167 vdd gnd cell_6t
Xbit_r168_c113 bl_113 br_113 wl_168 vdd gnd cell_6t
Xbit_r169_c113 bl_113 br_113 wl_169 vdd gnd cell_6t
Xbit_r170_c113 bl_113 br_113 wl_170 vdd gnd cell_6t
Xbit_r171_c113 bl_113 br_113 wl_171 vdd gnd cell_6t
Xbit_r172_c113 bl_113 br_113 wl_172 vdd gnd cell_6t
Xbit_r173_c113 bl_113 br_113 wl_173 vdd gnd cell_6t
Xbit_r174_c113 bl_113 br_113 wl_174 vdd gnd cell_6t
Xbit_r175_c113 bl_113 br_113 wl_175 vdd gnd cell_6t
Xbit_r176_c113 bl_113 br_113 wl_176 vdd gnd cell_6t
Xbit_r177_c113 bl_113 br_113 wl_177 vdd gnd cell_6t
Xbit_r178_c113 bl_113 br_113 wl_178 vdd gnd cell_6t
Xbit_r179_c113 bl_113 br_113 wl_179 vdd gnd cell_6t
Xbit_r180_c113 bl_113 br_113 wl_180 vdd gnd cell_6t
Xbit_r181_c113 bl_113 br_113 wl_181 vdd gnd cell_6t
Xbit_r182_c113 bl_113 br_113 wl_182 vdd gnd cell_6t
Xbit_r183_c113 bl_113 br_113 wl_183 vdd gnd cell_6t
Xbit_r184_c113 bl_113 br_113 wl_184 vdd gnd cell_6t
Xbit_r185_c113 bl_113 br_113 wl_185 vdd gnd cell_6t
Xbit_r186_c113 bl_113 br_113 wl_186 vdd gnd cell_6t
Xbit_r187_c113 bl_113 br_113 wl_187 vdd gnd cell_6t
Xbit_r188_c113 bl_113 br_113 wl_188 vdd gnd cell_6t
Xbit_r189_c113 bl_113 br_113 wl_189 vdd gnd cell_6t
Xbit_r190_c113 bl_113 br_113 wl_190 vdd gnd cell_6t
Xbit_r191_c113 bl_113 br_113 wl_191 vdd gnd cell_6t
Xbit_r192_c113 bl_113 br_113 wl_192 vdd gnd cell_6t
Xbit_r193_c113 bl_113 br_113 wl_193 vdd gnd cell_6t
Xbit_r194_c113 bl_113 br_113 wl_194 vdd gnd cell_6t
Xbit_r195_c113 bl_113 br_113 wl_195 vdd gnd cell_6t
Xbit_r196_c113 bl_113 br_113 wl_196 vdd gnd cell_6t
Xbit_r197_c113 bl_113 br_113 wl_197 vdd gnd cell_6t
Xbit_r198_c113 bl_113 br_113 wl_198 vdd gnd cell_6t
Xbit_r199_c113 bl_113 br_113 wl_199 vdd gnd cell_6t
Xbit_r200_c113 bl_113 br_113 wl_200 vdd gnd cell_6t
Xbit_r201_c113 bl_113 br_113 wl_201 vdd gnd cell_6t
Xbit_r202_c113 bl_113 br_113 wl_202 vdd gnd cell_6t
Xbit_r203_c113 bl_113 br_113 wl_203 vdd gnd cell_6t
Xbit_r204_c113 bl_113 br_113 wl_204 vdd gnd cell_6t
Xbit_r205_c113 bl_113 br_113 wl_205 vdd gnd cell_6t
Xbit_r206_c113 bl_113 br_113 wl_206 vdd gnd cell_6t
Xbit_r207_c113 bl_113 br_113 wl_207 vdd gnd cell_6t
Xbit_r208_c113 bl_113 br_113 wl_208 vdd gnd cell_6t
Xbit_r209_c113 bl_113 br_113 wl_209 vdd gnd cell_6t
Xbit_r210_c113 bl_113 br_113 wl_210 vdd gnd cell_6t
Xbit_r211_c113 bl_113 br_113 wl_211 vdd gnd cell_6t
Xbit_r212_c113 bl_113 br_113 wl_212 vdd gnd cell_6t
Xbit_r213_c113 bl_113 br_113 wl_213 vdd gnd cell_6t
Xbit_r214_c113 bl_113 br_113 wl_214 vdd gnd cell_6t
Xbit_r215_c113 bl_113 br_113 wl_215 vdd gnd cell_6t
Xbit_r216_c113 bl_113 br_113 wl_216 vdd gnd cell_6t
Xbit_r217_c113 bl_113 br_113 wl_217 vdd gnd cell_6t
Xbit_r218_c113 bl_113 br_113 wl_218 vdd gnd cell_6t
Xbit_r219_c113 bl_113 br_113 wl_219 vdd gnd cell_6t
Xbit_r220_c113 bl_113 br_113 wl_220 vdd gnd cell_6t
Xbit_r221_c113 bl_113 br_113 wl_221 vdd gnd cell_6t
Xbit_r222_c113 bl_113 br_113 wl_222 vdd gnd cell_6t
Xbit_r223_c113 bl_113 br_113 wl_223 vdd gnd cell_6t
Xbit_r224_c113 bl_113 br_113 wl_224 vdd gnd cell_6t
Xbit_r225_c113 bl_113 br_113 wl_225 vdd gnd cell_6t
Xbit_r226_c113 bl_113 br_113 wl_226 vdd gnd cell_6t
Xbit_r227_c113 bl_113 br_113 wl_227 vdd gnd cell_6t
Xbit_r228_c113 bl_113 br_113 wl_228 vdd gnd cell_6t
Xbit_r229_c113 bl_113 br_113 wl_229 vdd gnd cell_6t
Xbit_r230_c113 bl_113 br_113 wl_230 vdd gnd cell_6t
Xbit_r231_c113 bl_113 br_113 wl_231 vdd gnd cell_6t
Xbit_r232_c113 bl_113 br_113 wl_232 vdd gnd cell_6t
Xbit_r233_c113 bl_113 br_113 wl_233 vdd gnd cell_6t
Xbit_r234_c113 bl_113 br_113 wl_234 vdd gnd cell_6t
Xbit_r235_c113 bl_113 br_113 wl_235 vdd gnd cell_6t
Xbit_r236_c113 bl_113 br_113 wl_236 vdd gnd cell_6t
Xbit_r237_c113 bl_113 br_113 wl_237 vdd gnd cell_6t
Xbit_r238_c113 bl_113 br_113 wl_238 vdd gnd cell_6t
Xbit_r239_c113 bl_113 br_113 wl_239 vdd gnd cell_6t
Xbit_r240_c113 bl_113 br_113 wl_240 vdd gnd cell_6t
Xbit_r241_c113 bl_113 br_113 wl_241 vdd gnd cell_6t
Xbit_r242_c113 bl_113 br_113 wl_242 vdd gnd cell_6t
Xbit_r243_c113 bl_113 br_113 wl_243 vdd gnd cell_6t
Xbit_r244_c113 bl_113 br_113 wl_244 vdd gnd cell_6t
Xbit_r245_c113 bl_113 br_113 wl_245 vdd gnd cell_6t
Xbit_r246_c113 bl_113 br_113 wl_246 vdd gnd cell_6t
Xbit_r247_c113 bl_113 br_113 wl_247 vdd gnd cell_6t
Xbit_r248_c113 bl_113 br_113 wl_248 vdd gnd cell_6t
Xbit_r249_c113 bl_113 br_113 wl_249 vdd gnd cell_6t
Xbit_r250_c113 bl_113 br_113 wl_250 vdd gnd cell_6t
Xbit_r251_c113 bl_113 br_113 wl_251 vdd gnd cell_6t
Xbit_r252_c113 bl_113 br_113 wl_252 vdd gnd cell_6t
Xbit_r253_c113 bl_113 br_113 wl_253 vdd gnd cell_6t
Xbit_r254_c113 bl_113 br_113 wl_254 vdd gnd cell_6t
Xbit_r255_c113 bl_113 br_113 wl_255 vdd gnd cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd cell_6t
Xbit_r1_c114 bl_114 br_114 wl_1 vdd gnd cell_6t
Xbit_r2_c114 bl_114 br_114 wl_2 vdd gnd cell_6t
Xbit_r3_c114 bl_114 br_114 wl_3 vdd gnd cell_6t
Xbit_r4_c114 bl_114 br_114 wl_4 vdd gnd cell_6t
Xbit_r5_c114 bl_114 br_114 wl_5 vdd gnd cell_6t
Xbit_r6_c114 bl_114 br_114 wl_6 vdd gnd cell_6t
Xbit_r7_c114 bl_114 br_114 wl_7 vdd gnd cell_6t
Xbit_r8_c114 bl_114 br_114 wl_8 vdd gnd cell_6t
Xbit_r9_c114 bl_114 br_114 wl_9 vdd gnd cell_6t
Xbit_r10_c114 bl_114 br_114 wl_10 vdd gnd cell_6t
Xbit_r11_c114 bl_114 br_114 wl_11 vdd gnd cell_6t
Xbit_r12_c114 bl_114 br_114 wl_12 vdd gnd cell_6t
Xbit_r13_c114 bl_114 br_114 wl_13 vdd gnd cell_6t
Xbit_r14_c114 bl_114 br_114 wl_14 vdd gnd cell_6t
Xbit_r15_c114 bl_114 br_114 wl_15 vdd gnd cell_6t
Xbit_r16_c114 bl_114 br_114 wl_16 vdd gnd cell_6t
Xbit_r17_c114 bl_114 br_114 wl_17 vdd gnd cell_6t
Xbit_r18_c114 bl_114 br_114 wl_18 vdd gnd cell_6t
Xbit_r19_c114 bl_114 br_114 wl_19 vdd gnd cell_6t
Xbit_r20_c114 bl_114 br_114 wl_20 vdd gnd cell_6t
Xbit_r21_c114 bl_114 br_114 wl_21 vdd gnd cell_6t
Xbit_r22_c114 bl_114 br_114 wl_22 vdd gnd cell_6t
Xbit_r23_c114 bl_114 br_114 wl_23 vdd gnd cell_6t
Xbit_r24_c114 bl_114 br_114 wl_24 vdd gnd cell_6t
Xbit_r25_c114 bl_114 br_114 wl_25 vdd gnd cell_6t
Xbit_r26_c114 bl_114 br_114 wl_26 vdd gnd cell_6t
Xbit_r27_c114 bl_114 br_114 wl_27 vdd gnd cell_6t
Xbit_r28_c114 bl_114 br_114 wl_28 vdd gnd cell_6t
Xbit_r29_c114 bl_114 br_114 wl_29 vdd gnd cell_6t
Xbit_r30_c114 bl_114 br_114 wl_30 vdd gnd cell_6t
Xbit_r31_c114 bl_114 br_114 wl_31 vdd gnd cell_6t
Xbit_r32_c114 bl_114 br_114 wl_32 vdd gnd cell_6t
Xbit_r33_c114 bl_114 br_114 wl_33 vdd gnd cell_6t
Xbit_r34_c114 bl_114 br_114 wl_34 vdd gnd cell_6t
Xbit_r35_c114 bl_114 br_114 wl_35 vdd gnd cell_6t
Xbit_r36_c114 bl_114 br_114 wl_36 vdd gnd cell_6t
Xbit_r37_c114 bl_114 br_114 wl_37 vdd gnd cell_6t
Xbit_r38_c114 bl_114 br_114 wl_38 vdd gnd cell_6t
Xbit_r39_c114 bl_114 br_114 wl_39 vdd gnd cell_6t
Xbit_r40_c114 bl_114 br_114 wl_40 vdd gnd cell_6t
Xbit_r41_c114 bl_114 br_114 wl_41 vdd gnd cell_6t
Xbit_r42_c114 bl_114 br_114 wl_42 vdd gnd cell_6t
Xbit_r43_c114 bl_114 br_114 wl_43 vdd gnd cell_6t
Xbit_r44_c114 bl_114 br_114 wl_44 vdd gnd cell_6t
Xbit_r45_c114 bl_114 br_114 wl_45 vdd gnd cell_6t
Xbit_r46_c114 bl_114 br_114 wl_46 vdd gnd cell_6t
Xbit_r47_c114 bl_114 br_114 wl_47 vdd gnd cell_6t
Xbit_r48_c114 bl_114 br_114 wl_48 vdd gnd cell_6t
Xbit_r49_c114 bl_114 br_114 wl_49 vdd gnd cell_6t
Xbit_r50_c114 bl_114 br_114 wl_50 vdd gnd cell_6t
Xbit_r51_c114 bl_114 br_114 wl_51 vdd gnd cell_6t
Xbit_r52_c114 bl_114 br_114 wl_52 vdd gnd cell_6t
Xbit_r53_c114 bl_114 br_114 wl_53 vdd gnd cell_6t
Xbit_r54_c114 bl_114 br_114 wl_54 vdd gnd cell_6t
Xbit_r55_c114 bl_114 br_114 wl_55 vdd gnd cell_6t
Xbit_r56_c114 bl_114 br_114 wl_56 vdd gnd cell_6t
Xbit_r57_c114 bl_114 br_114 wl_57 vdd gnd cell_6t
Xbit_r58_c114 bl_114 br_114 wl_58 vdd gnd cell_6t
Xbit_r59_c114 bl_114 br_114 wl_59 vdd gnd cell_6t
Xbit_r60_c114 bl_114 br_114 wl_60 vdd gnd cell_6t
Xbit_r61_c114 bl_114 br_114 wl_61 vdd gnd cell_6t
Xbit_r62_c114 bl_114 br_114 wl_62 vdd gnd cell_6t
Xbit_r63_c114 bl_114 br_114 wl_63 vdd gnd cell_6t
Xbit_r64_c114 bl_114 br_114 wl_64 vdd gnd cell_6t
Xbit_r65_c114 bl_114 br_114 wl_65 vdd gnd cell_6t
Xbit_r66_c114 bl_114 br_114 wl_66 vdd gnd cell_6t
Xbit_r67_c114 bl_114 br_114 wl_67 vdd gnd cell_6t
Xbit_r68_c114 bl_114 br_114 wl_68 vdd gnd cell_6t
Xbit_r69_c114 bl_114 br_114 wl_69 vdd gnd cell_6t
Xbit_r70_c114 bl_114 br_114 wl_70 vdd gnd cell_6t
Xbit_r71_c114 bl_114 br_114 wl_71 vdd gnd cell_6t
Xbit_r72_c114 bl_114 br_114 wl_72 vdd gnd cell_6t
Xbit_r73_c114 bl_114 br_114 wl_73 vdd gnd cell_6t
Xbit_r74_c114 bl_114 br_114 wl_74 vdd gnd cell_6t
Xbit_r75_c114 bl_114 br_114 wl_75 vdd gnd cell_6t
Xbit_r76_c114 bl_114 br_114 wl_76 vdd gnd cell_6t
Xbit_r77_c114 bl_114 br_114 wl_77 vdd gnd cell_6t
Xbit_r78_c114 bl_114 br_114 wl_78 vdd gnd cell_6t
Xbit_r79_c114 bl_114 br_114 wl_79 vdd gnd cell_6t
Xbit_r80_c114 bl_114 br_114 wl_80 vdd gnd cell_6t
Xbit_r81_c114 bl_114 br_114 wl_81 vdd gnd cell_6t
Xbit_r82_c114 bl_114 br_114 wl_82 vdd gnd cell_6t
Xbit_r83_c114 bl_114 br_114 wl_83 vdd gnd cell_6t
Xbit_r84_c114 bl_114 br_114 wl_84 vdd gnd cell_6t
Xbit_r85_c114 bl_114 br_114 wl_85 vdd gnd cell_6t
Xbit_r86_c114 bl_114 br_114 wl_86 vdd gnd cell_6t
Xbit_r87_c114 bl_114 br_114 wl_87 vdd gnd cell_6t
Xbit_r88_c114 bl_114 br_114 wl_88 vdd gnd cell_6t
Xbit_r89_c114 bl_114 br_114 wl_89 vdd gnd cell_6t
Xbit_r90_c114 bl_114 br_114 wl_90 vdd gnd cell_6t
Xbit_r91_c114 bl_114 br_114 wl_91 vdd gnd cell_6t
Xbit_r92_c114 bl_114 br_114 wl_92 vdd gnd cell_6t
Xbit_r93_c114 bl_114 br_114 wl_93 vdd gnd cell_6t
Xbit_r94_c114 bl_114 br_114 wl_94 vdd gnd cell_6t
Xbit_r95_c114 bl_114 br_114 wl_95 vdd gnd cell_6t
Xbit_r96_c114 bl_114 br_114 wl_96 vdd gnd cell_6t
Xbit_r97_c114 bl_114 br_114 wl_97 vdd gnd cell_6t
Xbit_r98_c114 bl_114 br_114 wl_98 vdd gnd cell_6t
Xbit_r99_c114 bl_114 br_114 wl_99 vdd gnd cell_6t
Xbit_r100_c114 bl_114 br_114 wl_100 vdd gnd cell_6t
Xbit_r101_c114 bl_114 br_114 wl_101 vdd gnd cell_6t
Xbit_r102_c114 bl_114 br_114 wl_102 vdd gnd cell_6t
Xbit_r103_c114 bl_114 br_114 wl_103 vdd gnd cell_6t
Xbit_r104_c114 bl_114 br_114 wl_104 vdd gnd cell_6t
Xbit_r105_c114 bl_114 br_114 wl_105 vdd gnd cell_6t
Xbit_r106_c114 bl_114 br_114 wl_106 vdd gnd cell_6t
Xbit_r107_c114 bl_114 br_114 wl_107 vdd gnd cell_6t
Xbit_r108_c114 bl_114 br_114 wl_108 vdd gnd cell_6t
Xbit_r109_c114 bl_114 br_114 wl_109 vdd gnd cell_6t
Xbit_r110_c114 bl_114 br_114 wl_110 vdd gnd cell_6t
Xbit_r111_c114 bl_114 br_114 wl_111 vdd gnd cell_6t
Xbit_r112_c114 bl_114 br_114 wl_112 vdd gnd cell_6t
Xbit_r113_c114 bl_114 br_114 wl_113 vdd gnd cell_6t
Xbit_r114_c114 bl_114 br_114 wl_114 vdd gnd cell_6t
Xbit_r115_c114 bl_114 br_114 wl_115 vdd gnd cell_6t
Xbit_r116_c114 bl_114 br_114 wl_116 vdd gnd cell_6t
Xbit_r117_c114 bl_114 br_114 wl_117 vdd gnd cell_6t
Xbit_r118_c114 bl_114 br_114 wl_118 vdd gnd cell_6t
Xbit_r119_c114 bl_114 br_114 wl_119 vdd gnd cell_6t
Xbit_r120_c114 bl_114 br_114 wl_120 vdd gnd cell_6t
Xbit_r121_c114 bl_114 br_114 wl_121 vdd gnd cell_6t
Xbit_r122_c114 bl_114 br_114 wl_122 vdd gnd cell_6t
Xbit_r123_c114 bl_114 br_114 wl_123 vdd gnd cell_6t
Xbit_r124_c114 bl_114 br_114 wl_124 vdd gnd cell_6t
Xbit_r125_c114 bl_114 br_114 wl_125 vdd gnd cell_6t
Xbit_r126_c114 bl_114 br_114 wl_126 vdd gnd cell_6t
Xbit_r127_c114 bl_114 br_114 wl_127 vdd gnd cell_6t
Xbit_r128_c114 bl_114 br_114 wl_128 vdd gnd cell_6t
Xbit_r129_c114 bl_114 br_114 wl_129 vdd gnd cell_6t
Xbit_r130_c114 bl_114 br_114 wl_130 vdd gnd cell_6t
Xbit_r131_c114 bl_114 br_114 wl_131 vdd gnd cell_6t
Xbit_r132_c114 bl_114 br_114 wl_132 vdd gnd cell_6t
Xbit_r133_c114 bl_114 br_114 wl_133 vdd gnd cell_6t
Xbit_r134_c114 bl_114 br_114 wl_134 vdd gnd cell_6t
Xbit_r135_c114 bl_114 br_114 wl_135 vdd gnd cell_6t
Xbit_r136_c114 bl_114 br_114 wl_136 vdd gnd cell_6t
Xbit_r137_c114 bl_114 br_114 wl_137 vdd gnd cell_6t
Xbit_r138_c114 bl_114 br_114 wl_138 vdd gnd cell_6t
Xbit_r139_c114 bl_114 br_114 wl_139 vdd gnd cell_6t
Xbit_r140_c114 bl_114 br_114 wl_140 vdd gnd cell_6t
Xbit_r141_c114 bl_114 br_114 wl_141 vdd gnd cell_6t
Xbit_r142_c114 bl_114 br_114 wl_142 vdd gnd cell_6t
Xbit_r143_c114 bl_114 br_114 wl_143 vdd gnd cell_6t
Xbit_r144_c114 bl_114 br_114 wl_144 vdd gnd cell_6t
Xbit_r145_c114 bl_114 br_114 wl_145 vdd gnd cell_6t
Xbit_r146_c114 bl_114 br_114 wl_146 vdd gnd cell_6t
Xbit_r147_c114 bl_114 br_114 wl_147 vdd gnd cell_6t
Xbit_r148_c114 bl_114 br_114 wl_148 vdd gnd cell_6t
Xbit_r149_c114 bl_114 br_114 wl_149 vdd gnd cell_6t
Xbit_r150_c114 bl_114 br_114 wl_150 vdd gnd cell_6t
Xbit_r151_c114 bl_114 br_114 wl_151 vdd gnd cell_6t
Xbit_r152_c114 bl_114 br_114 wl_152 vdd gnd cell_6t
Xbit_r153_c114 bl_114 br_114 wl_153 vdd gnd cell_6t
Xbit_r154_c114 bl_114 br_114 wl_154 vdd gnd cell_6t
Xbit_r155_c114 bl_114 br_114 wl_155 vdd gnd cell_6t
Xbit_r156_c114 bl_114 br_114 wl_156 vdd gnd cell_6t
Xbit_r157_c114 bl_114 br_114 wl_157 vdd gnd cell_6t
Xbit_r158_c114 bl_114 br_114 wl_158 vdd gnd cell_6t
Xbit_r159_c114 bl_114 br_114 wl_159 vdd gnd cell_6t
Xbit_r160_c114 bl_114 br_114 wl_160 vdd gnd cell_6t
Xbit_r161_c114 bl_114 br_114 wl_161 vdd gnd cell_6t
Xbit_r162_c114 bl_114 br_114 wl_162 vdd gnd cell_6t
Xbit_r163_c114 bl_114 br_114 wl_163 vdd gnd cell_6t
Xbit_r164_c114 bl_114 br_114 wl_164 vdd gnd cell_6t
Xbit_r165_c114 bl_114 br_114 wl_165 vdd gnd cell_6t
Xbit_r166_c114 bl_114 br_114 wl_166 vdd gnd cell_6t
Xbit_r167_c114 bl_114 br_114 wl_167 vdd gnd cell_6t
Xbit_r168_c114 bl_114 br_114 wl_168 vdd gnd cell_6t
Xbit_r169_c114 bl_114 br_114 wl_169 vdd gnd cell_6t
Xbit_r170_c114 bl_114 br_114 wl_170 vdd gnd cell_6t
Xbit_r171_c114 bl_114 br_114 wl_171 vdd gnd cell_6t
Xbit_r172_c114 bl_114 br_114 wl_172 vdd gnd cell_6t
Xbit_r173_c114 bl_114 br_114 wl_173 vdd gnd cell_6t
Xbit_r174_c114 bl_114 br_114 wl_174 vdd gnd cell_6t
Xbit_r175_c114 bl_114 br_114 wl_175 vdd gnd cell_6t
Xbit_r176_c114 bl_114 br_114 wl_176 vdd gnd cell_6t
Xbit_r177_c114 bl_114 br_114 wl_177 vdd gnd cell_6t
Xbit_r178_c114 bl_114 br_114 wl_178 vdd gnd cell_6t
Xbit_r179_c114 bl_114 br_114 wl_179 vdd gnd cell_6t
Xbit_r180_c114 bl_114 br_114 wl_180 vdd gnd cell_6t
Xbit_r181_c114 bl_114 br_114 wl_181 vdd gnd cell_6t
Xbit_r182_c114 bl_114 br_114 wl_182 vdd gnd cell_6t
Xbit_r183_c114 bl_114 br_114 wl_183 vdd gnd cell_6t
Xbit_r184_c114 bl_114 br_114 wl_184 vdd gnd cell_6t
Xbit_r185_c114 bl_114 br_114 wl_185 vdd gnd cell_6t
Xbit_r186_c114 bl_114 br_114 wl_186 vdd gnd cell_6t
Xbit_r187_c114 bl_114 br_114 wl_187 vdd gnd cell_6t
Xbit_r188_c114 bl_114 br_114 wl_188 vdd gnd cell_6t
Xbit_r189_c114 bl_114 br_114 wl_189 vdd gnd cell_6t
Xbit_r190_c114 bl_114 br_114 wl_190 vdd gnd cell_6t
Xbit_r191_c114 bl_114 br_114 wl_191 vdd gnd cell_6t
Xbit_r192_c114 bl_114 br_114 wl_192 vdd gnd cell_6t
Xbit_r193_c114 bl_114 br_114 wl_193 vdd gnd cell_6t
Xbit_r194_c114 bl_114 br_114 wl_194 vdd gnd cell_6t
Xbit_r195_c114 bl_114 br_114 wl_195 vdd gnd cell_6t
Xbit_r196_c114 bl_114 br_114 wl_196 vdd gnd cell_6t
Xbit_r197_c114 bl_114 br_114 wl_197 vdd gnd cell_6t
Xbit_r198_c114 bl_114 br_114 wl_198 vdd gnd cell_6t
Xbit_r199_c114 bl_114 br_114 wl_199 vdd gnd cell_6t
Xbit_r200_c114 bl_114 br_114 wl_200 vdd gnd cell_6t
Xbit_r201_c114 bl_114 br_114 wl_201 vdd gnd cell_6t
Xbit_r202_c114 bl_114 br_114 wl_202 vdd gnd cell_6t
Xbit_r203_c114 bl_114 br_114 wl_203 vdd gnd cell_6t
Xbit_r204_c114 bl_114 br_114 wl_204 vdd gnd cell_6t
Xbit_r205_c114 bl_114 br_114 wl_205 vdd gnd cell_6t
Xbit_r206_c114 bl_114 br_114 wl_206 vdd gnd cell_6t
Xbit_r207_c114 bl_114 br_114 wl_207 vdd gnd cell_6t
Xbit_r208_c114 bl_114 br_114 wl_208 vdd gnd cell_6t
Xbit_r209_c114 bl_114 br_114 wl_209 vdd gnd cell_6t
Xbit_r210_c114 bl_114 br_114 wl_210 vdd gnd cell_6t
Xbit_r211_c114 bl_114 br_114 wl_211 vdd gnd cell_6t
Xbit_r212_c114 bl_114 br_114 wl_212 vdd gnd cell_6t
Xbit_r213_c114 bl_114 br_114 wl_213 vdd gnd cell_6t
Xbit_r214_c114 bl_114 br_114 wl_214 vdd gnd cell_6t
Xbit_r215_c114 bl_114 br_114 wl_215 vdd gnd cell_6t
Xbit_r216_c114 bl_114 br_114 wl_216 vdd gnd cell_6t
Xbit_r217_c114 bl_114 br_114 wl_217 vdd gnd cell_6t
Xbit_r218_c114 bl_114 br_114 wl_218 vdd gnd cell_6t
Xbit_r219_c114 bl_114 br_114 wl_219 vdd gnd cell_6t
Xbit_r220_c114 bl_114 br_114 wl_220 vdd gnd cell_6t
Xbit_r221_c114 bl_114 br_114 wl_221 vdd gnd cell_6t
Xbit_r222_c114 bl_114 br_114 wl_222 vdd gnd cell_6t
Xbit_r223_c114 bl_114 br_114 wl_223 vdd gnd cell_6t
Xbit_r224_c114 bl_114 br_114 wl_224 vdd gnd cell_6t
Xbit_r225_c114 bl_114 br_114 wl_225 vdd gnd cell_6t
Xbit_r226_c114 bl_114 br_114 wl_226 vdd gnd cell_6t
Xbit_r227_c114 bl_114 br_114 wl_227 vdd gnd cell_6t
Xbit_r228_c114 bl_114 br_114 wl_228 vdd gnd cell_6t
Xbit_r229_c114 bl_114 br_114 wl_229 vdd gnd cell_6t
Xbit_r230_c114 bl_114 br_114 wl_230 vdd gnd cell_6t
Xbit_r231_c114 bl_114 br_114 wl_231 vdd gnd cell_6t
Xbit_r232_c114 bl_114 br_114 wl_232 vdd gnd cell_6t
Xbit_r233_c114 bl_114 br_114 wl_233 vdd gnd cell_6t
Xbit_r234_c114 bl_114 br_114 wl_234 vdd gnd cell_6t
Xbit_r235_c114 bl_114 br_114 wl_235 vdd gnd cell_6t
Xbit_r236_c114 bl_114 br_114 wl_236 vdd gnd cell_6t
Xbit_r237_c114 bl_114 br_114 wl_237 vdd gnd cell_6t
Xbit_r238_c114 bl_114 br_114 wl_238 vdd gnd cell_6t
Xbit_r239_c114 bl_114 br_114 wl_239 vdd gnd cell_6t
Xbit_r240_c114 bl_114 br_114 wl_240 vdd gnd cell_6t
Xbit_r241_c114 bl_114 br_114 wl_241 vdd gnd cell_6t
Xbit_r242_c114 bl_114 br_114 wl_242 vdd gnd cell_6t
Xbit_r243_c114 bl_114 br_114 wl_243 vdd gnd cell_6t
Xbit_r244_c114 bl_114 br_114 wl_244 vdd gnd cell_6t
Xbit_r245_c114 bl_114 br_114 wl_245 vdd gnd cell_6t
Xbit_r246_c114 bl_114 br_114 wl_246 vdd gnd cell_6t
Xbit_r247_c114 bl_114 br_114 wl_247 vdd gnd cell_6t
Xbit_r248_c114 bl_114 br_114 wl_248 vdd gnd cell_6t
Xbit_r249_c114 bl_114 br_114 wl_249 vdd gnd cell_6t
Xbit_r250_c114 bl_114 br_114 wl_250 vdd gnd cell_6t
Xbit_r251_c114 bl_114 br_114 wl_251 vdd gnd cell_6t
Xbit_r252_c114 bl_114 br_114 wl_252 vdd gnd cell_6t
Xbit_r253_c114 bl_114 br_114 wl_253 vdd gnd cell_6t
Xbit_r254_c114 bl_114 br_114 wl_254 vdd gnd cell_6t
Xbit_r255_c114 bl_114 br_114 wl_255 vdd gnd cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd cell_6t
Xbit_r1_c115 bl_115 br_115 wl_1 vdd gnd cell_6t
Xbit_r2_c115 bl_115 br_115 wl_2 vdd gnd cell_6t
Xbit_r3_c115 bl_115 br_115 wl_3 vdd gnd cell_6t
Xbit_r4_c115 bl_115 br_115 wl_4 vdd gnd cell_6t
Xbit_r5_c115 bl_115 br_115 wl_5 vdd gnd cell_6t
Xbit_r6_c115 bl_115 br_115 wl_6 vdd gnd cell_6t
Xbit_r7_c115 bl_115 br_115 wl_7 vdd gnd cell_6t
Xbit_r8_c115 bl_115 br_115 wl_8 vdd gnd cell_6t
Xbit_r9_c115 bl_115 br_115 wl_9 vdd gnd cell_6t
Xbit_r10_c115 bl_115 br_115 wl_10 vdd gnd cell_6t
Xbit_r11_c115 bl_115 br_115 wl_11 vdd gnd cell_6t
Xbit_r12_c115 bl_115 br_115 wl_12 vdd gnd cell_6t
Xbit_r13_c115 bl_115 br_115 wl_13 vdd gnd cell_6t
Xbit_r14_c115 bl_115 br_115 wl_14 vdd gnd cell_6t
Xbit_r15_c115 bl_115 br_115 wl_15 vdd gnd cell_6t
Xbit_r16_c115 bl_115 br_115 wl_16 vdd gnd cell_6t
Xbit_r17_c115 bl_115 br_115 wl_17 vdd gnd cell_6t
Xbit_r18_c115 bl_115 br_115 wl_18 vdd gnd cell_6t
Xbit_r19_c115 bl_115 br_115 wl_19 vdd gnd cell_6t
Xbit_r20_c115 bl_115 br_115 wl_20 vdd gnd cell_6t
Xbit_r21_c115 bl_115 br_115 wl_21 vdd gnd cell_6t
Xbit_r22_c115 bl_115 br_115 wl_22 vdd gnd cell_6t
Xbit_r23_c115 bl_115 br_115 wl_23 vdd gnd cell_6t
Xbit_r24_c115 bl_115 br_115 wl_24 vdd gnd cell_6t
Xbit_r25_c115 bl_115 br_115 wl_25 vdd gnd cell_6t
Xbit_r26_c115 bl_115 br_115 wl_26 vdd gnd cell_6t
Xbit_r27_c115 bl_115 br_115 wl_27 vdd gnd cell_6t
Xbit_r28_c115 bl_115 br_115 wl_28 vdd gnd cell_6t
Xbit_r29_c115 bl_115 br_115 wl_29 vdd gnd cell_6t
Xbit_r30_c115 bl_115 br_115 wl_30 vdd gnd cell_6t
Xbit_r31_c115 bl_115 br_115 wl_31 vdd gnd cell_6t
Xbit_r32_c115 bl_115 br_115 wl_32 vdd gnd cell_6t
Xbit_r33_c115 bl_115 br_115 wl_33 vdd gnd cell_6t
Xbit_r34_c115 bl_115 br_115 wl_34 vdd gnd cell_6t
Xbit_r35_c115 bl_115 br_115 wl_35 vdd gnd cell_6t
Xbit_r36_c115 bl_115 br_115 wl_36 vdd gnd cell_6t
Xbit_r37_c115 bl_115 br_115 wl_37 vdd gnd cell_6t
Xbit_r38_c115 bl_115 br_115 wl_38 vdd gnd cell_6t
Xbit_r39_c115 bl_115 br_115 wl_39 vdd gnd cell_6t
Xbit_r40_c115 bl_115 br_115 wl_40 vdd gnd cell_6t
Xbit_r41_c115 bl_115 br_115 wl_41 vdd gnd cell_6t
Xbit_r42_c115 bl_115 br_115 wl_42 vdd gnd cell_6t
Xbit_r43_c115 bl_115 br_115 wl_43 vdd gnd cell_6t
Xbit_r44_c115 bl_115 br_115 wl_44 vdd gnd cell_6t
Xbit_r45_c115 bl_115 br_115 wl_45 vdd gnd cell_6t
Xbit_r46_c115 bl_115 br_115 wl_46 vdd gnd cell_6t
Xbit_r47_c115 bl_115 br_115 wl_47 vdd gnd cell_6t
Xbit_r48_c115 bl_115 br_115 wl_48 vdd gnd cell_6t
Xbit_r49_c115 bl_115 br_115 wl_49 vdd gnd cell_6t
Xbit_r50_c115 bl_115 br_115 wl_50 vdd gnd cell_6t
Xbit_r51_c115 bl_115 br_115 wl_51 vdd gnd cell_6t
Xbit_r52_c115 bl_115 br_115 wl_52 vdd gnd cell_6t
Xbit_r53_c115 bl_115 br_115 wl_53 vdd gnd cell_6t
Xbit_r54_c115 bl_115 br_115 wl_54 vdd gnd cell_6t
Xbit_r55_c115 bl_115 br_115 wl_55 vdd gnd cell_6t
Xbit_r56_c115 bl_115 br_115 wl_56 vdd gnd cell_6t
Xbit_r57_c115 bl_115 br_115 wl_57 vdd gnd cell_6t
Xbit_r58_c115 bl_115 br_115 wl_58 vdd gnd cell_6t
Xbit_r59_c115 bl_115 br_115 wl_59 vdd gnd cell_6t
Xbit_r60_c115 bl_115 br_115 wl_60 vdd gnd cell_6t
Xbit_r61_c115 bl_115 br_115 wl_61 vdd gnd cell_6t
Xbit_r62_c115 bl_115 br_115 wl_62 vdd gnd cell_6t
Xbit_r63_c115 bl_115 br_115 wl_63 vdd gnd cell_6t
Xbit_r64_c115 bl_115 br_115 wl_64 vdd gnd cell_6t
Xbit_r65_c115 bl_115 br_115 wl_65 vdd gnd cell_6t
Xbit_r66_c115 bl_115 br_115 wl_66 vdd gnd cell_6t
Xbit_r67_c115 bl_115 br_115 wl_67 vdd gnd cell_6t
Xbit_r68_c115 bl_115 br_115 wl_68 vdd gnd cell_6t
Xbit_r69_c115 bl_115 br_115 wl_69 vdd gnd cell_6t
Xbit_r70_c115 bl_115 br_115 wl_70 vdd gnd cell_6t
Xbit_r71_c115 bl_115 br_115 wl_71 vdd gnd cell_6t
Xbit_r72_c115 bl_115 br_115 wl_72 vdd gnd cell_6t
Xbit_r73_c115 bl_115 br_115 wl_73 vdd gnd cell_6t
Xbit_r74_c115 bl_115 br_115 wl_74 vdd gnd cell_6t
Xbit_r75_c115 bl_115 br_115 wl_75 vdd gnd cell_6t
Xbit_r76_c115 bl_115 br_115 wl_76 vdd gnd cell_6t
Xbit_r77_c115 bl_115 br_115 wl_77 vdd gnd cell_6t
Xbit_r78_c115 bl_115 br_115 wl_78 vdd gnd cell_6t
Xbit_r79_c115 bl_115 br_115 wl_79 vdd gnd cell_6t
Xbit_r80_c115 bl_115 br_115 wl_80 vdd gnd cell_6t
Xbit_r81_c115 bl_115 br_115 wl_81 vdd gnd cell_6t
Xbit_r82_c115 bl_115 br_115 wl_82 vdd gnd cell_6t
Xbit_r83_c115 bl_115 br_115 wl_83 vdd gnd cell_6t
Xbit_r84_c115 bl_115 br_115 wl_84 vdd gnd cell_6t
Xbit_r85_c115 bl_115 br_115 wl_85 vdd gnd cell_6t
Xbit_r86_c115 bl_115 br_115 wl_86 vdd gnd cell_6t
Xbit_r87_c115 bl_115 br_115 wl_87 vdd gnd cell_6t
Xbit_r88_c115 bl_115 br_115 wl_88 vdd gnd cell_6t
Xbit_r89_c115 bl_115 br_115 wl_89 vdd gnd cell_6t
Xbit_r90_c115 bl_115 br_115 wl_90 vdd gnd cell_6t
Xbit_r91_c115 bl_115 br_115 wl_91 vdd gnd cell_6t
Xbit_r92_c115 bl_115 br_115 wl_92 vdd gnd cell_6t
Xbit_r93_c115 bl_115 br_115 wl_93 vdd gnd cell_6t
Xbit_r94_c115 bl_115 br_115 wl_94 vdd gnd cell_6t
Xbit_r95_c115 bl_115 br_115 wl_95 vdd gnd cell_6t
Xbit_r96_c115 bl_115 br_115 wl_96 vdd gnd cell_6t
Xbit_r97_c115 bl_115 br_115 wl_97 vdd gnd cell_6t
Xbit_r98_c115 bl_115 br_115 wl_98 vdd gnd cell_6t
Xbit_r99_c115 bl_115 br_115 wl_99 vdd gnd cell_6t
Xbit_r100_c115 bl_115 br_115 wl_100 vdd gnd cell_6t
Xbit_r101_c115 bl_115 br_115 wl_101 vdd gnd cell_6t
Xbit_r102_c115 bl_115 br_115 wl_102 vdd gnd cell_6t
Xbit_r103_c115 bl_115 br_115 wl_103 vdd gnd cell_6t
Xbit_r104_c115 bl_115 br_115 wl_104 vdd gnd cell_6t
Xbit_r105_c115 bl_115 br_115 wl_105 vdd gnd cell_6t
Xbit_r106_c115 bl_115 br_115 wl_106 vdd gnd cell_6t
Xbit_r107_c115 bl_115 br_115 wl_107 vdd gnd cell_6t
Xbit_r108_c115 bl_115 br_115 wl_108 vdd gnd cell_6t
Xbit_r109_c115 bl_115 br_115 wl_109 vdd gnd cell_6t
Xbit_r110_c115 bl_115 br_115 wl_110 vdd gnd cell_6t
Xbit_r111_c115 bl_115 br_115 wl_111 vdd gnd cell_6t
Xbit_r112_c115 bl_115 br_115 wl_112 vdd gnd cell_6t
Xbit_r113_c115 bl_115 br_115 wl_113 vdd gnd cell_6t
Xbit_r114_c115 bl_115 br_115 wl_114 vdd gnd cell_6t
Xbit_r115_c115 bl_115 br_115 wl_115 vdd gnd cell_6t
Xbit_r116_c115 bl_115 br_115 wl_116 vdd gnd cell_6t
Xbit_r117_c115 bl_115 br_115 wl_117 vdd gnd cell_6t
Xbit_r118_c115 bl_115 br_115 wl_118 vdd gnd cell_6t
Xbit_r119_c115 bl_115 br_115 wl_119 vdd gnd cell_6t
Xbit_r120_c115 bl_115 br_115 wl_120 vdd gnd cell_6t
Xbit_r121_c115 bl_115 br_115 wl_121 vdd gnd cell_6t
Xbit_r122_c115 bl_115 br_115 wl_122 vdd gnd cell_6t
Xbit_r123_c115 bl_115 br_115 wl_123 vdd gnd cell_6t
Xbit_r124_c115 bl_115 br_115 wl_124 vdd gnd cell_6t
Xbit_r125_c115 bl_115 br_115 wl_125 vdd gnd cell_6t
Xbit_r126_c115 bl_115 br_115 wl_126 vdd gnd cell_6t
Xbit_r127_c115 bl_115 br_115 wl_127 vdd gnd cell_6t
Xbit_r128_c115 bl_115 br_115 wl_128 vdd gnd cell_6t
Xbit_r129_c115 bl_115 br_115 wl_129 vdd gnd cell_6t
Xbit_r130_c115 bl_115 br_115 wl_130 vdd gnd cell_6t
Xbit_r131_c115 bl_115 br_115 wl_131 vdd gnd cell_6t
Xbit_r132_c115 bl_115 br_115 wl_132 vdd gnd cell_6t
Xbit_r133_c115 bl_115 br_115 wl_133 vdd gnd cell_6t
Xbit_r134_c115 bl_115 br_115 wl_134 vdd gnd cell_6t
Xbit_r135_c115 bl_115 br_115 wl_135 vdd gnd cell_6t
Xbit_r136_c115 bl_115 br_115 wl_136 vdd gnd cell_6t
Xbit_r137_c115 bl_115 br_115 wl_137 vdd gnd cell_6t
Xbit_r138_c115 bl_115 br_115 wl_138 vdd gnd cell_6t
Xbit_r139_c115 bl_115 br_115 wl_139 vdd gnd cell_6t
Xbit_r140_c115 bl_115 br_115 wl_140 vdd gnd cell_6t
Xbit_r141_c115 bl_115 br_115 wl_141 vdd gnd cell_6t
Xbit_r142_c115 bl_115 br_115 wl_142 vdd gnd cell_6t
Xbit_r143_c115 bl_115 br_115 wl_143 vdd gnd cell_6t
Xbit_r144_c115 bl_115 br_115 wl_144 vdd gnd cell_6t
Xbit_r145_c115 bl_115 br_115 wl_145 vdd gnd cell_6t
Xbit_r146_c115 bl_115 br_115 wl_146 vdd gnd cell_6t
Xbit_r147_c115 bl_115 br_115 wl_147 vdd gnd cell_6t
Xbit_r148_c115 bl_115 br_115 wl_148 vdd gnd cell_6t
Xbit_r149_c115 bl_115 br_115 wl_149 vdd gnd cell_6t
Xbit_r150_c115 bl_115 br_115 wl_150 vdd gnd cell_6t
Xbit_r151_c115 bl_115 br_115 wl_151 vdd gnd cell_6t
Xbit_r152_c115 bl_115 br_115 wl_152 vdd gnd cell_6t
Xbit_r153_c115 bl_115 br_115 wl_153 vdd gnd cell_6t
Xbit_r154_c115 bl_115 br_115 wl_154 vdd gnd cell_6t
Xbit_r155_c115 bl_115 br_115 wl_155 vdd gnd cell_6t
Xbit_r156_c115 bl_115 br_115 wl_156 vdd gnd cell_6t
Xbit_r157_c115 bl_115 br_115 wl_157 vdd gnd cell_6t
Xbit_r158_c115 bl_115 br_115 wl_158 vdd gnd cell_6t
Xbit_r159_c115 bl_115 br_115 wl_159 vdd gnd cell_6t
Xbit_r160_c115 bl_115 br_115 wl_160 vdd gnd cell_6t
Xbit_r161_c115 bl_115 br_115 wl_161 vdd gnd cell_6t
Xbit_r162_c115 bl_115 br_115 wl_162 vdd gnd cell_6t
Xbit_r163_c115 bl_115 br_115 wl_163 vdd gnd cell_6t
Xbit_r164_c115 bl_115 br_115 wl_164 vdd gnd cell_6t
Xbit_r165_c115 bl_115 br_115 wl_165 vdd gnd cell_6t
Xbit_r166_c115 bl_115 br_115 wl_166 vdd gnd cell_6t
Xbit_r167_c115 bl_115 br_115 wl_167 vdd gnd cell_6t
Xbit_r168_c115 bl_115 br_115 wl_168 vdd gnd cell_6t
Xbit_r169_c115 bl_115 br_115 wl_169 vdd gnd cell_6t
Xbit_r170_c115 bl_115 br_115 wl_170 vdd gnd cell_6t
Xbit_r171_c115 bl_115 br_115 wl_171 vdd gnd cell_6t
Xbit_r172_c115 bl_115 br_115 wl_172 vdd gnd cell_6t
Xbit_r173_c115 bl_115 br_115 wl_173 vdd gnd cell_6t
Xbit_r174_c115 bl_115 br_115 wl_174 vdd gnd cell_6t
Xbit_r175_c115 bl_115 br_115 wl_175 vdd gnd cell_6t
Xbit_r176_c115 bl_115 br_115 wl_176 vdd gnd cell_6t
Xbit_r177_c115 bl_115 br_115 wl_177 vdd gnd cell_6t
Xbit_r178_c115 bl_115 br_115 wl_178 vdd gnd cell_6t
Xbit_r179_c115 bl_115 br_115 wl_179 vdd gnd cell_6t
Xbit_r180_c115 bl_115 br_115 wl_180 vdd gnd cell_6t
Xbit_r181_c115 bl_115 br_115 wl_181 vdd gnd cell_6t
Xbit_r182_c115 bl_115 br_115 wl_182 vdd gnd cell_6t
Xbit_r183_c115 bl_115 br_115 wl_183 vdd gnd cell_6t
Xbit_r184_c115 bl_115 br_115 wl_184 vdd gnd cell_6t
Xbit_r185_c115 bl_115 br_115 wl_185 vdd gnd cell_6t
Xbit_r186_c115 bl_115 br_115 wl_186 vdd gnd cell_6t
Xbit_r187_c115 bl_115 br_115 wl_187 vdd gnd cell_6t
Xbit_r188_c115 bl_115 br_115 wl_188 vdd gnd cell_6t
Xbit_r189_c115 bl_115 br_115 wl_189 vdd gnd cell_6t
Xbit_r190_c115 bl_115 br_115 wl_190 vdd gnd cell_6t
Xbit_r191_c115 bl_115 br_115 wl_191 vdd gnd cell_6t
Xbit_r192_c115 bl_115 br_115 wl_192 vdd gnd cell_6t
Xbit_r193_c115 bl_115 br_115 wl_193 vdd gnd cell_6t
Xbit_r194_c115 bl_115 br_115 wl_194 vdd gnd cell_6t
Xbit_r195_c115 bl_115 br_115 wl_195 vdd gnd cell_6t
Xbit_r196_c115 bl_115 br_115 wl_196 vdd gnd cell_6t
Xbit_r197_c115 bl_115 br_115 wl_197 vdd gnd cell_6t
Xbit_r198_c115 bl_115 br_115 wl_198 vdd gnd cell_6t
Xbit_r199_c115 bl_115 br_115 wl_199 vdd gnd cell_6t
Xbit_r200_c115 bl_115 br_115 wl_200 vdd gnd cell_6t
Xbit_r201_c115 bl_115 br_115 wl_201 vdd gnd cell_6t
Xbit_r202_c115 bl_115 br_115 wl_202 vdd gnd cell_6t
Xbit_r203_c115 bl_115 br_115 wl_203 vdd gnd cell_6t
Xbit_r204_c115 bl_115 br_115 wl_204 vdd gnd cell_6t
Xbit_r205_c115 bl_115 br_115 wl_205 vdd gnd cell_6t
Xbit_r206_c115 bl_115 br_115 wl_206 vdd gnd cell_6t
Xbit_r207_c115 bl_115 br_115 wl_207 vdd gnd cell_6t
Xbit_r208_c115 bl_115 br_115 wl_208 vdd gnd cell_6t
Xbit_r209_c115 bl_115 br_115 wl_209 vdd gnd cell_6t
Xbit_r210_c115 bl_115 br_115 wl_210 vdd gnd cell_6t
Xbit_r211_c115 bl_115 br_115 wl_211 vdd gnd cell_6t
Xbit_r212_c115 bl_115 br_115 wl_212 vdd gnd cell_6t
Xbit_r213_c115 bl_115 br_115 wl_213 vdd gnd cell_6t
Xbit_r214_c115 bl_115 br_115 wl_214 vdd gnd cell_6t
Xbit_r215_c115 bl_115 br_115 wl_215 vdd gnd cell_6t
Xbit_r216_c115 bl_115 br_115 wl_216 vdd gnd cell_6t
Xbit_r217_c115 bl_115 br_115 wl_217 vdd gnd cell_6t
Xbit_r218_c115 bl_115 br_115 wl_218 vdd gnd cell_6t
Xbit_r219_c115 bl_115 br_115 wl_219 vdd gnd cell_6t
Xbit_r220_c115 bl_115 br_115 wl_220 vdd gnd cell_6t
Xbit_r221_c115 bl_115 br_115 wl_221 vdd gnd cell_6t
Xbit_r222_c115 bl_115 br_115 wl_222 vdd gnd cell_6t
Xbit_r223_c115 bl_115 br_115 wl_223 vdd gnd cell_6t
Xbit_r224_c115 bl_115 br_115 wl_224 vdd gnd cell_6t
Xbit_r225_c115 bl_115 br_115 wl_225 vdd gnd cell_6t
Xbit_r226_c115 bl_115 br_115 wl_226 vdd gnd cell_6t
Xbit_r227_c115 bl_115 br_115 wl_227 vdd gnd cell_6t
Xbit_r228_c115 bl_115 br_115 wl_228 vdd gnd cell_6t
Xbit_r229_c115 bl_115 br_115 wl_229 vdd gnd cell_6t
Xbit_r230_c115 bl_115 br_115 wl_230 vdd gnd cell_6t
Xbit_r231_c115 bl_115 br_115 wl_231 vdd gnd cell_6t
Xbit_r232_c115 bl_115 br_115 wl_232 vdd gnd cell_6t
Xbit_r233_c115 bl_115 br_115 wl_233 vdd gnd cell_6t
Xbit_r234_c115 bl_115 br_115 wl_234 vdd gnd cell_6t
Xbit_r235_c115 bl_115 br_115 wl_235 vdd gnd cell_6t
Xbit_r236_c115 bl_115 br_115 wl_236 vdd gnd cell_6t
Xbit_r237_c115 bl_115 br_115 wl_237 vdd gnd cell_6t
Xbit_r238_c115 bl_115 br_115 wl_238 vdd gnd cell_6t
Xbit_r239_c115 bl_115 br_115 wl_239 vdd gnd cell_6t
Xbit_r240_c115 bl_115 br_115 wl_240 vdd gnd cell_6t
Xbit_r241_c115 bl_115 br_115 wl_241 vdd gnd cell_6t
Xbit_r242_c115 bl_115 br_115 wl_242 vdd gnd cell_6t
Xbit_r243_c115 bl_115 br_115 wl_243 vdd gnd cell_6t
Xbit_r244_c115 bl_115 br_115 wl_244 vdd gnd cell_6t
Xbit_r245_c115 bl_115 br_115 wl_245 vdd gnd cell_6t
Xbit_r246_c115 bl_115 br_115 wl_246 vdd gnd cell_6t
Xbit_r247_c115 bl_115 br_115 wl_247 vdd gnd cell_6t
Xbit_r248_c115 bl_115 br_115 wl_248 vdd gnd cell_6t
Xbit_r249_c115 bl_115 br_115 wl_249 vdd gnd cell_6t
Xbit_r250_c115 bl_115 br_115 wl_250 vdd gnd cell_6t
Xbit_r251_c115 bl_115 br_115 wl_251 vdd gnd cell_6t
Xbit_r252_c115 bl_115 br_115 wl_252 vdd gnd cell_6t
Xbit_r253_c115 bl_115 br_115 wl_253 vdd gnd cell_6t
Xbit_r254_c115 bl_115 br_115 wl_254 vdd gnd cell_6t
Xbit_r255_c115 bl_115 br_115 wl_255 vdd gnd cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd cell_6t
Xbit_r1_c116 bl_116 br_116 wl_1 vdd gnd cell_6t
Xbit_r2_c116 bl_116 br_116 wl_2 vdd gnd cell_6t
Xbit_r3_c116 bl_116 br_116 wl_3 vdd gnd cell_6t
Xbit_r4_c116 bl_116 br_116 wl_4 vdd gnd cell_6t
Xbit_r5_c116 bl_116 br_116 wl_5 vdd gnd cell_6t
Xbit_r6_c116 bl_116 br_116 wl_6 vdd gnd cell_6t
Xbit_r7_c116 bl_116 br_116 wl_7 vdd gnd cell_6t
Xbit_r8_c116 bl_116 br_116 wl_8 vdd gnd cell_6t
Xbit_r9_c116 bl_116 br_116 wl_9 vdd gnd cell_6t
Xbit_r10_c116 bl_116 br_116 wl_10 vdd gnd cell_6t
Xbit_r11_c116 bl_116 br_116 wl_11 vdd gnd cell_6t
Xbit_r12_c116 bl_116 br_116 wl_12 vdd gnd cell_6t
Xbit_r13_c116 bl_116 br_116 wl_13 vdd gnd cell_6t
Xbit_r14_c116 bl_116 br_116 wl_14 vdd gnd cell_6t
Xbit_r15_c116 bl_116 br_116 wl_15 vdd gnd cell_6t
Xbit_r16_c116 bl_116 br_116 wl_16 vdd gnd cell_6t
Xbit_r17_c116 bl_116 br_116 wl_17 vdd gnd cell_6t
Xbit_r18_c116 bl_116 br_116 wl_18 vdd gnd cell_6t
Xbit_r19_c116 bl_116 br_116 wl_19 vdd gnd cell_6t
Xbit_r20_c116 bl_116 br_116 wl_20 vdd gnd cell_6t
Xbit_r21_c116 bl_116 br_116 wl_21 vdd gnd cell_6t
Xbit_r22_c116 bl_116 br_116 wl_22 vdd gnd cell_6t
Xbit_r23_c116 bl_116 br_116 wl_23 vdd gnd cell_6t
Xbit_r24_c116 bl_116 br_116 wl_24 vdd gnd cell_6t
Xbit_r25_c116 bl_116 br_116 wl_25 vdd gnd cell_6t
Xbit_r26_c116 bl_116 br_116 wl_26 vdd gnd cell_6t
Xbit_r27_c116 bl_116 br_116 wl_27 vdd gnd cell_6t
Xbit_r28_c116 bl_116 br_116 wl_28 vdd gnd cell_6t
Xbit_r29_c116 bl_116 br_116 wl_29 vdd gnd cell_6t
Xbit_r30_c116 bl_116 br_116 wl_30 vdd gnd cell_6t
Xbit_r31_c116 bl_116 br_116 wl_31 vdd gnd cell_6t
Xbit_r32_c116 bl_116 br_116 wl_32 vdd gnd cell_6t
Xbit_r33_c116 bl_116 br_116 wl_33 vdd gnd cell_6t
Xbit_r34_c116 bl_116 br_116 wl_34 vdd gnd cell_6t
Xbit_r35_c116 bl_116 br_116 wl_35 vdd gnd cell_6t
Xbit_r36_c116 bl_116 br_116 wl_36 vdd gnd cell_6t
Xbit_r37_c116 bl_116 br_116 wl_37 vdd gnd cell_6t
Xbit_r38_c116 bl_116 br_116 wl_38 vdd gnd cell_6t
Xbit_r39_c116 bl_116 br_116 wl_39 vdd gnd cell_6t
Xbit_r40_c116 bl_116 br_116 wl_40 vdd gnd cell_6t
Xbit_r41_c116 bl_116 br_116 wl_41 vdd gnd cell_6t
Xbit_r42_c116 bl_116 br_116 wl_42 vdd gnd cell_6t
Xbit_r43_c116 bl_116 br_116 wl_43 vdd gnd cell_6t
Xbit_r44_c116 bl_116 br_116 wl_44 vdd gnd cell_6t
Xbit_r45_c116 bl_116 br_116 wl_45 vdd gnd cell_6t
Xbit_r46_c116 bl_116 br_116 wl_46 vdd gnd cell_6t
Xbit_r47_c116 bl_116 br_116 wl_47 vdd gnd cell_6t
Xbit_r48_c116 bl_116 br_116 wl_48 vdd gnd cell_6t
Xbit_r49_c116 bl_116 br_116 wl_49 vdd gnd cell_6t
Xbit_r50_c116 bl_116 br_116 wl_50 vdd gnd cell_6t
Xbit_r51_c116 bl_116 br_116 wl_51 vdd gnd cell_6t
Xbit_r52_c116 bl_116 br_116 wl_52 vdd gnd cell_6t
Xbit_r53_c116 bl_116 br_116 wl_53 vdd gnd cell_6t
Xbit_r54_c116 bl_116 br_116 wl_54 vdd gnd cell_6t
Xbit_r55_c116 bl_116 br_116 wl_55 vdd gnd cell_6t
Xbit_r56_c116 bl_116 br_116 wl_56 vdd gnd cell_6t
Xbit_r57_c116 bl_116 br_116 wl_57 vdd gnd cell_6t
Xbit_r58_c116 bl_116 br_116 wl_58 vdd gnd cell_6t
Xbit_r59_c116 bl_116 br_116 wl_59 vdd gnd cell_6t
Xbit_r60_c116 bl_116 br_116 wl_60 vdd gnd cell_6t
Xbit_r61_c116 bl_116 br_116 wl_61 vdd gnd cell_6t
Xbit_r62_c116 bl_116 br_116 wl_62 vdd gnd cell_6t
Xbit_r63_c116 bl_116 br_116 wl_63 vdd gnd cell_6t
Xbit_r64_c116 bl_116 br_116 wl_64 vdd gnd cell_6t
Xbit_r65_c116 bl_116 br_116 wl_65 vdd gnd cell_6t
Xbit_r66_c116 bl_116 br_116 wl_66 vdd gnd cell_6t
Xbit_r67_c116 bl_116 br_116 wl_67 vdd gnd cell_6t
Xbit_r68_c116 bl_116 br_116 wl_68 vdd gnd cell_6t
Xbit_r69_c116 bl_116 br_116 wl_69 vdd gnd cell_6t
Xbit_r70_c116 bl_116 br_116 wl_70 vdd gnd cell_6t
Xbit_r71_c116 bl_116 br_116 wl_71 vdd gnd cell_6t
Xbit_r72_c116 bl_116 br_116 wl_72 vdd gnd cell_6t
Xbit_r73_c116 bl_116 br_116 wl_73 vdd gnd cell_6t
Xbit_r74_c116 bl_116 br_116 wl_74 vdd gnd cell_6t
Xbit_r75_c116 bl_116 br_116 wl_75 vdd gnd cell_6t
Xbit_r76_c116 bl_116 br_116 wl_76 vdd gnd cell_6t
Xbit_r77_c116 bl_116 br_116 wl_77 vdd gnd cell_6t
Xbit_r78_c116 bl_116 br_116 wl_78 vdd gnd cell_6t
Xbit_r79_c116 bl_116 br_116 wl_79 vdd gnd cell_6t
Xbit_r80_c116 bl_116 br_116 wl_80 vdd gnd cell_6t
Xbit_r81_c116 bl_116 br_116 wl_81 vdd gnd cell_6t
Xbit_r82_c116 bl_116 br_116 wl_82 vdd gnd cell_6t
Xbit_r83_c116 bl_116 br_116 wl_83 vdd gnd cell_6t
Xbit_r84_c116 bl_116 br_116 wl_84 vdd gnd cell_6t
Xbit_r85_c116 bl_116 br_116 wl_85 vdd gnd cell_6t
Xbit_r86_c116 bl_116 br_116 wl_86 vdd gnd cell_6t
Xbit_r87_c116 bl_116 br_116 wl_87 vdd gnd cell_6t
Xbit_r88_c116 bl_116 br_116 wl_88 vdd gnd cell_6t
Xbit_r89_c116 bl_116 br_116 wl_89 vdd gnd cell_6t
Xbit_r90_c116 bl_116 br_116 wl_90 vdd gnd cell_6t
Xbit_r91_c116 bl_116 br_116 wl_91 vdd gnd cell_6t
Xbit_r92_c116 bl_116 br_116 wl_92 vdd gnd cell_6t
Xbit_r93_c116 bl_116 br_116 wl_93 vdd gnd cell_6t
Xbit_r94_c116 bl_116 br_116 wl_94 vdd gnd cell_6t
Xbit_r95_c116 bl_116 br_116 wl_95 vdd gnd cell_6t
Xbit_r96_c116 bl_116 br_116 wl_96 vdd gnd cell_6t
Xbit_r97_c116 bl_116 br_116 wl_97 vdd gnd cell_6t
Xbit_r98_c116 bl_116 br_116 wl_98 vdd gnd cell_6t
Xbit_r99_c116 bl_116 br_116 wl_99 vdd gnd cell_6t
Xbit_r100_c116 bl_116 br_116 wl_100 vdd gnd cell_6t
Xbit_r101_c116 bl_116 br_116 wl_101 vdd gnd cell_6t
Xbit_r102_c116 bl_116 br_116 wl_102 vdd gnd cell_6t
Xbit_r103_c116 bl_116 br_116 wl_103 vdd gnd cell_6t
Xbit_r104_c116 bl_116 br_116 wl_104 vdd gnd cell_6t
Xbit_r105_c116 bl_116 br_116 wl_105 vdd gnd cell_6t
Xbit_r106_c116 bl_116 br_116 wl_106 vdd gnd cell_6t
Xbit_r107_c116 bl_116 br_116 wl_107 vdd gnd cell_6t
Xbit_r108_c116 bl_116 br_116 wl_108 vdd gnd cell_6t
Xbit_r109_c116 bl_116 br_116 wl_109 vdd gnd cell_6t
Xbit_r110_c116 bl_116 br_116 wl_110 vdd gnd cell_6t
Xbit_r111_c116 bl_116 br_116 wl_111 vdd gnd cell_6t
Xbit_r112_c116 bl_116 br_116 wl_112 vdd gnd cell_6t
Xbit_r113_c116 bl_116 br_116 wl_113 vdd gnd cell_6t
Xbit_r114_c116 bl_116 br_116 wl_114 vdd gnd cell_6t
Xbit_r115_c116 bl_116 br_116 wl_115 vdd gnd cell_6t
Xbit_r116_c116 bl_116 br_116 wl_116 vdd gnd cell_6t
Xbit_r117_c116 bl_116 br_116 wl_117 vdd gnd cell_6t
Xbit_r118_c116 bl_116 br_116 wl_118 vdd gnd cell_6t
Xbit_r119_c116 bl_116 br_116 wl_119 vdd gnd cell_6t
Xbit_r120_c116 bl_116 br_116 wl_120 vdd gnd cell_6t
Xbit_r121_c116 bl_116 br_116 wl_121 vdd gnd cell_6t
Xbit_r122_c116 bl_116 br_116 wl_122 vdd gnd cell_6t
Xbit_r123_c116 bl_116 br_116 wl_123 vdd gnd cell_6t
Xbit_r124_c116 bl_116 br_116 wl_124 vdd gnd cell_6t
Xbit_r125_c116 bl_116 br_116 wl_125 vdd gnd cell_6t
Xbit_r126_c116 bl_116 br_116 wl_126 vdd gnd cell_6t
Xbit_r127_c116 bl_116 br_116 wl_127 vdd gnd cell_6t
Xbit_r128_c116 bl_116 br_116 wl_128 vdd gnd cell_6t
Xbit_r129_c116 bl_116 br_116 wl_129 vdd gnd cell_6t
Xbit_r130_c116 bl_116 br_116 wl_130 vdd gnd cell_6t
Xbit_r131_c116 bl_116 br_116 wl_131 vdd gnd cell_6t
Xbit_r132_c116 bl_116 br_116 wl_132 vdd gnd cell_6t
Xbit_r133_c116 bl_116 br_116 wl_133 vdd gnd cell_6t
Xbit_r134_c116 bl_116 br_116 wl_134 vdd gnd cell_6t
Xbit_r135_c116 bl_116 br_116 wl_135 vdd gnd cell_6t
Xbit_r136_c116 bl_116 br_116 wl_136 vdd gnd cell_6t
Xbit_r137_c116 bl_116 br_116 wl_137 vdd gnd cell_6t
Xbit_r138_c116 bl_116 br_116 wl_138 vdd gnd cell_6t
Xbit_r139_c116 bl_116 br_116 wl_139 vdd gnd cell_6t
Xbit_r140_c116 bl_116 br_116 wl_140 vdd gnd cell_6t
Xbit_r141_c116 bl_116 br_116 wl_141 vdd gnd cell_6t
Xbit_r142_c116 bl_116 br_116 wl_142 vdd gnd cell_6t
Xbit_r143_c116 bl_116 br_116 wl_143 vdd gnd cell_6t
Xbit_r144_c116 bl_116 br_116 wl_144 vdd gnd cell_6t
Xbit_r145_c116 bl_116 br_116 wl_145 vdd gnd cell_6t
Xbit_r146_c116 bl_116 br_116 wl_146 vdd gnd cell_6t
Xbit_r147_c116 bl_116 br_116 wl_147 vdd gnd cell_6t
Xbit_r148_c116 bl_116 br_116 wl_148 vdd gnd cell_6t
Xbit_r149_c116 bl_116 br_116 wl_149 vdd gnd cell_6t
Xbit_r150_c116 bl_116 br_116 wl_150 vdd gnd cell_6t
Xbit_r151_c116 bl_116 br_116 wl_151 vdd gnd cell_6t
Xbit_r152_c116 bl_116 br_116 wl_152 vdd gnd cell_6t
Xbit_r153_c116 bl_116 br_116 wl_153 vdd gnd cell_6t
Xbit_r154_c116 bl_116 br_116 wl_154 vdd gnd cell_6t
Xbit_r155_c116 bl_116 br_116 wl_155 vdd gnd cell_6t
Xbit_r156_c116 bl_116 br_116 wl_156 vdd gnd cell_6t
Xbit_r157_c116 bl_116 br_116 wl_157 vdd gnd cell_6t
Xbit_r158_c116 bl_116 br_116 wl_158 vdd gnd cell_6t
Xbit_r159_c116 bl_116 br_116 wl_159 vdd gnd cell_6t
Xbit_r160_c116 bl_116 br_116 wl_160 vdd gnd cell_6t
Xbit_r161_c116 bl_116 br_116 wl_161 vdd gnd cell_6t
Xbit_r162_c116 bl_116 br_116 wl_162 vdd gnd cell_6t
Xbit_r163_c116 bl_116 br_116 wl_163 vdd gnd cell_6t
Xbit_r164_c116 bl_116 br_116 wl_164 vdd gnd cell_6t
Xbit_r165_c116 bl_116 br_116 wl_165 vdd gnd cell_6t
Xbit_r166_c116 bl_116 br_116 wl_166 vdd gnd cell_6t
Xbit_r167_c116 bl_116 br_116 wl_167 vdd gnd cell_6t
Xbit_r168_c116 bl_116 br_116 wl_168 vdd gnd cell_6t
Xbit_r169_c116 bl_116 br_116 wl_169 vdd gnd cell_6t
Xbit_r170_c116 bl_116 br_116 wl_170 vdd gnd cell_6t
Xbit_r171_c116 bl_116 br_116 wl_171 vdd gnd cell_6t
Xbit_r172_c116 bl_116 br_116 wl_172 vdd gnd cell_6t
Xbit_r173_c116 bl_116 br_116 wl_173 vdd gnd cell_6t
Xbit_r174_c116 bl_116 br_116 wl_174 vdd gnd cell_6t
Xbit_r175_c116 bl_116 br_116 wl_175 vdd gnd cell_6t
Xbit_r176_c116 bl_116 br_116 wl_176 vdd gnd cell_6t
Xbit_r177_c116 bl_116 br_116 wl_177 vdd gnd cell_6t
Xbit_r178_c116 bl_116 br_116 wl_178 vdd gnd cell_6t
Xbit_r179_c116 bl_116 br_116 wl_179 vdd gnd cell_6t
Xbit_r180_c116 bl_116 br_116 wl_180 vdd gnd cell_6t
Xbit_r181_c116 bl_116 br_116 wl_181 vdd gnd cell_6t
Xbit_r182_c116 bl_116 br_116 wl_182 vdd gnd cell_6t
Xbit_r183_c116 bl_116 br_116 wl_183 vdd gnd cell_6t
Xbit_r184_c116 bl_116 br_116 wl_184 vdd gnd cell_6t
Xbit_r185_c116 bl_116 br_116 wl_185 vdd gnd cell_6t
Xbit_r186_c116 bl_116 br_116 wl_186 vdd gnd cell_6t
Xbit_r187_c116 bl_116 br_116 wl_187 vdd gnd cell_6t
Xbit_r188_c116 bl_116 br_116 wl_188 vdd gnd cell_6t
Xbit_r189_c116 bl_116 br_116 wl_189 vdd gnd cell_6t
Xbit_r190_c116 bl_116 br_116 wl_190 vdd gnd cell_6t
Xbit_r191_c116 bl_116 br_116 wl_191 vdd gnd cell_6t
Xbit_r192_c116 bl_116 br_116 wl_192 vdd gnd cell_6t
Xbit_r193_c116 bl_116 br_116 wl_193 vdd gnd cell_6t
Xbit_r194_c116 bl_116 br_116 wl_194 vdd gnd cell_6t
Xbit_r195_c116 bl_116 br_116 wl_195 vdd gnd cell_6t
Xbit_r196_c116 bl_116 br_116 wl_196 vdd gnd cell_6t
Xbit_r197_c116 bl_116 br_116 wl_197 vdd gnd cell_6t
Xbit_r198_c116 bl_116 br_116 wl_198 vdd gnd cell_6t
Xbit_r199_c116 bl_116 br_116 wl_199 vdd gnd cell_6t
Xbit_r200_c116 bl_116 br_116 wl_200 vdd gnd cell_6t
Xbit_r201_c116 bl_116 br_116 wl_201 vdd gnd cell_6t
Xbit_r202_c116 bl_116 br_116 wl_202 vdd gnd cell_6t
Xbit_r203_c116 bl_116 br_116 wl_203 vdd gnd cell_6t
Xbit_r204_c116 bl_116 br_116 wl_204 vdd gnd cell_6t
Xbit_r205_c116 bl_116 br_116 wl_205 vdd gnd cell_6t
Xbit_r206_c116 bl_116 br_116 wl_206 vdd gnd cell_6t
Xbit_r207_c116 bl_116 br_116 wl_207 vdd gnd cell_6t
Xbit_r208_c116 bl_116 br_116 wl_208 vdd gnd cell_6t
Xbit_r209_c116 bl_116 br_116 wl_209 vdd gnd cell_6t
Xbit_r210_c116 bl_116 br_116 wl_210 vdd gnd cell_6t
Xbit_r211_c116 bl_116 br_116 wl_211 vdd gnd cell_6t
Xbit_r212_c116 bl_116 br_116 wl_212 vdd gnd cell_6t
Xbit_r213_c116 bl_116 br_116 wl_213 vdd gnd cell_6t
Xbit_r214_c116 bl_116 br_116 wl_214 vdd gnd cell_6t
Xbit_r215_c116 bl_116 br_116 wl_215 vdd gnd cell_6t
Xbit_r216_c116 bl_116 br_116 wl_216 vdd gnd cell_6t
Xbit_r217_c116 bl_116 br_116 wl_217 vdd gnd cell_6t
Xbit_r218_c116 bl_116 br_116 wl_218 vdd gnd cell_6t
Xbit_r219_c116 bl_116 br_116 wl_219 vdd gnd cell_6t
Xbit_r220_c116 bl_116 br_116 wl_220 vdd gnd cell_6t
Xbit_r221_c116 bl_116 br_116 wl_221 vdd gnd cell_6t
Xbit_r222_c116 bl_116 br_116 wl_222 vdd gnd cell_6t
Xbit_r223_c116 bl_116 br_116 wl_223 vdd gnd cell_6t
Xbit_r224_c116 bl_116 br_116 wl_224 vdd gnd cell_6t
Xbit_r225_c116 bl_116 br_116 wl_225 vdd gnd cell_6t
Xbit_r226_c116 bl_116 br_116 wl_226 vdd gnd cell_6t
Xbit_r227_c116 bl_116 br_116 wl_227 vdd gnd cell_6t
Xbit_r228_c116 bl_116 br_116 wl_228 vdd gnd cell_6t
Xbit_r229_c116 bl_116 br_116 wl_229 vdd gnd cell_6t
Xbit_r230_c116 bl_116 br_116 wl_230 vdd gnd cell_6t
Xbit_r231_c116 bl_116 br_116 wl_231 vdd gnd cell_6t
Xbit_r232_c116 bl_116 br_116 wl_232 vdd gnd cell_6t
Xbit_r233_c116 bl_116 br_116 wl_233 vdd gnd cell_6t
Xbit_r234_c116 bl_116 br_116 wl_234 vdd gnd cell_6t
Xbit_r235_c116 bl_116 br_116 wl_235 vdd gnd cell_6t
Xbit_r236_c116 bl_116 br_116 wl_236 vdd gnd cell_6t
Xbit_r237_c116 bl_116 br_116 wl_237 vdd gnd cell_6t
Xbit_r238_c116 bl_116 br_116 wl_238 vdd gnd cell_6t
Xbit_r239_c116 bl_116 br_116 wl_239 vdd gnd cell_6t
Xbit_r240_c116 bl_116 br_116 wl_240 vdd gnd cell_6t
Xbit_r241_c116 bl_116 br_116 wl_241 vdd gnd cell_6t
Xbit_r242_c116 bl_116 br_116 wl_242 vdd gnd cell_6t
Xbit_r243_c116 bl_116 br_116 wl_243 vdd gnd cell_6t
Xbit_r244_c116 bl_116 br_116 wl_244 vdd gnd cell_6t
Xbit_r245_c116 bl_116 br_116 wl_245 vdd gnd cell_6t
Xbit_r246_c116 bl_116 br_116 wl_246 vdd gnd cell_6t
Xbit_r247_c116 bl_116 br_116 wl_247 vdd gnd cell_6t
Xbit_r248_c116 bl_116 br_116 wl_248 vdd gnd cell_6t
Xbit_r249_c116 bl_116 br_116 wl_249 vdd gnd cell_6t
Xbit_r250_c116 bl_116 br_116 wl_250 vdd gnd cell_6t
Xbit_r251_c116 bl_116 br_116 wl_251 vdd gnd cell_6t
Xbit_r252_c116 bl_116 br_116 wl_252 vdd gnd cell_6t
Xbit_r253_c116 bl_116 br_116 wl_253 vdd gnd cell_6t
Xbit_r254_c116 bl_116 br_116 wl_254 vdd gnd cell_6t
Xbit_r255_c116 bl_116 br_116 wl_255 vdd gnd cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd cell_6t
Xbit_r1_c117 bl_117 br_117 wl_1 vdd gnd cell_6t
Xbit_r2_c117 bl_117 br_117 wl_2 vdd gnd cell_6t
Xbit_r3_c117 bl_117 br_117 wl_3 vdd gnd cell_6t
Xbit_r4_c117 bl_117 br_117 wl_4 vdd gnd cell_6t
Xbit_r5_c117 bl_117 br_117 wl_5 vdd gnd cell_6t
Xbit_r6_c117 bl_117 br_117 wl_6 vdd gnd cell_6t
Xbit_r7_c117 bl_117 br_117 wl_7 vdd gnd cell_6t
Xbit_r8_c117 bl_117 br_117 wl_8 vdd gnd cell_6t
Xbit_r9_c117 bl_117 br_117 wl_9 vdd gnd cell_6t
Xbit_r10_c117 bl_117 br_117 wl_10 vdd gnd cell_6t
Xbit_r11_c117 bl_117 br_117 wl_11 vdd gnd cell_6t
Xbit_r12_c117 bl_117 br_117 wl_12 vdd gnd cell_6t
Xbit_r13_c117 bl_117 br_117 wl_13 vdd gnd cell_6t
Xbit_r14_c117 bl_117 br_117 wl_14 vdd gnd cell_6t
Xbit_r15_c117 bl_117 br_117 wl_15 vdd gnd cell_6t
Xbit_r16_c117 bl_117 br_117 wl_16 vdd gnd cell_6t
Xbit_r17_c117 bl_117 br_117 wl_17 vdd gnd cell_6t
Xbit_r18_c117 bl_117 br_117 wl_18 vdd gnd cell_6t
Xbit_r19_c117 bl_117 br_117 wl_19 vdd gnd cell_6t
Xbit_r20_c117 bl_117 br_117 wl_20 vdd gnd cell_6t
Xbit_r21_c117 bl_117 br_117 wl_21 vdd gnd cell_6t
Xbit_r22_c117 bl_117 br_117 wl_22 vdd gnd cell_6t
Xbit_r23_c117 bl_117 br_117 wl_23 vdd gnd cell_6t
Xbit_r24_c117 bl_117 br_117 wl_24 vdd gnd cell_6t
Xbit_r25_c117 bl_117 br_117 wl_25 vdd gnd cell_6t
Xbit_r26_c117 bl_117 br_117 wl_26 vdd gnd cell_6t
Xbit_r27_c117 bl_117 br_117 wl_27 vdd gnd cell_6t
Xbit_r28_c117 bl_117 br_117 wl_28 vdd gnd cell_6t
Xbit_r29_c117 bl_117 br_117 wl_29 vdd gnd cell_6t
Xbit_r30_c117 bl_117 br_117 wl_30 vdd gnd cell_6t
Xbit_r31_c117 bl_117 br_117 wl_31 vdd gnd cell_6t
Xbit_r32_c117 bl_117 br_117 wl_32 vdd gnd cell_6t
Xbit_r33_c117 bl_117 br_117 wl_33 vdd gnd cell_6t
Xbit_r34_c117 bl_117 br_117 wl_34 vdd gnd cell_6t
Xbit_r35_c117 bl_117 br_117 wl_35 vdd gnd cell_6t
Xbit_r36_c117 bl_117 br_117 wl_36 vdd gnd cell_6t
Xbit_r37_c117 bl_117 br_117 wl_37 vdd gnd cell_6t
Xbit_r38_c117 bl_117 br_117 wl_38 vdd gnd cell_6t
Xbit_r39_c117 bl_117 br_117 wl_39 vdd gnd cell_6t
Xbit_r40_c117 bl_117 br_117 wl_40 vdd gnd cell_6t
Xbit_r41_c117 bl_117 br_117 wl_41 vdd gnd cell_6t
Xbit_r42_c117 bl_117 br_117 wl_42 vdd gnd cell_6t
Xbit_r43_c117 bl_117 br_117 wl_43 vdd gnd cell_6t
Xbit_r44_c117 bl_117 br_117 wl_44 vdd gnd cell_6t
Xbit_r45_c117 bl_117 br_117 wl_45 vdd gnd cell_6t
Xbit_r46_c117 bl_117 br_117 wl_46 vdd gnd cell_6t
Xbit_r47_c117 bl_117 br_117 wl_47 vdd gnd cell_6t
Xbit_r48_c117 bl_117 br_117 wl_48 vdd gnd cell_6t
Xbit_r49_c117 bl_117 br_117 wl_49 vdd gnd cell_6t
Xbit_r50_c117 bl_117 br_117 wl_50 vdd gnd cell_6t
Xbit_r51_c117 bl_117 br_117 wl_51 vdd gnd cell_6t
Xbit_r52_c117 bl_117 br_117 wl_52 vdd gnd cell_6t
Xbit_r53_c117 bl_117 br_117 wl_53 vdd gnd cell_6t
Xbit_r54_c117 bl_117 br_117 wl_54 vdd gnd cell_6t
Xbit_r55_c117 bl_117 br_117 wl_55 vdd gnd cell_6t
Xbit_r56_c117 bl_117 br_117 wl_56 vdd gnd cell_6t
Xbit_r57_c117 bl_117 br_117 wl_57 vdd gnd cell_6t
Xbit_r58_c117 bl_117 br_117 wl_58 vdd gnd cell_6t
Xbit_r59_c117 bl_117 br_117 wl_59 vdd gnd cell_6t
Xbit_r60_c117 bl_117 br_117 wl_60 vdd gnd cell_6t
Xbit_r61_c117 bl_117 br_117 wl_61 vdd gnd cell_6t
Xbit_r62_c117 bl_117 br_117 wl_62 vdd gnd cell_6t
Xbit_r63_c117 bl_117 br_117 wl_63 vdd gnd cell_6t
Xbit_r64_c117 bl_117 br_117 wl_64 vdd gnd cell_6t
Xbit_r65_c117 bl_117 br_117 wl_65 vdd gnd cell_6t
Xbit_r66_c117 bl_117 br_117 wl_66 vdd gnd cell_6t
Xbit_r67_c117 bl_117 br_117 wl_67 vdd gnd cell_6t
Xbit_r68_c117 bl_117 br_117 wl_68 vdd gnd cell_6t
Xbit_r69_c117 bl_117 br_117 wl_69 vdd gnd cell_6t
Xbit_r70_c117 bl_117 br_117 wl_70 vdd gnd cell_6t
Xbit_r71_c117 bl_117 br_117 wl_71 vdd gnd cell_6t
Xbit_r72_c117 bl_117 br_117 wl_72 vdd gnd cell_6t
Xbit_r73_c117 bl_117 br_117 wl_73 vdd gnd cell_6t
Xbit_r74_c117 bl_117 br_117 wl_74 vdd gnd cell_6t
Xbit_r75_c117 bl_117 br_117 wl_75 vdd gnd cell_6t
Xbit_r76_c117 bl_117 br_117 wl_76 vdd gnd cell_6t
Xbit_r77_c117 bl_117 br_117 wl_77 vdd gnd cell_6t
Xbit_r78_c117 bl_117 br_117 wl_78 vdd gnd cell_6t
Xbit_r79_c117 bl_117 br_117 wl_79 vdd gnd cell_6t
Xbit_r80_c117 bl_117 br_117 wl_80 vdd gnd cell_6t
Xbit_r81_c117 bl_117 br_117 wl_81 vdd gnd cell_6t
Xbit_r82_c117 bl_117 br_117 wl_82 vdd gnd cell_6t
Xbit_r83_c117 bl_117 br_117 wl_83 vdd gnd cell_6t
Xbit_r84_c117 bl_117 br_117 wl_84 vdd gnd cell_6t
Xbit_r85_c117 bl_117 br_117 wl_85 vdd gnd cell_6t
Xbit_r86_c117 bl_117 br_117 wl_86 vdd gnd cell_6t
Xbit_r87_c117 bl_117 br_117 wl_87 vdd gnd cell_6t
Xbit_r88_c117 bl_117 br_117 wl_88 vdd gnd cell_6t
Xbit_r89_c117 bl_117 br_117 wl_89 vdd gnd cell_6t
Xbit_r90_c117 bl_117 br_117 wl_90 vdd gnd cell_6t
Xbit_r91_c117 bl_117 br_117 wl_91 vdd gnd cell_6t
Xbit_r92_c117 bl_117 br_117 wl_92 vdd gnd cell_6t
Xbit_r93_c117 bl_117 br_117 wl_93 vdd gnd cell_6t
Xbit_r94_c117 bl_117 br_117 wl_94 vdd gnd cell_6t
Xbit_r95_c117 bl_117 br_117 wl_95 vdd gnd cell_6t
Xbit_r96_c117 bl_117 br_117 wl_96 vdd gnd cell_6t
Xbit_r97_c117 bl_117 br_117 wl_97 vdd gnd cell_6t
Xbit_r98_c117 bl_117 br_117 wl_98 vdd gnd cell_6t
Xbit_r99_c117 bl_117 br_117 wl_99 vdd gnd cell_6t
Xbit_r100_c117 bl_117 br_117 wl_100 vdd gnd cell_6t
Xbit_r101_c117 bl_117 br_117 wl_101 vdd gnd cell_6t
Xbit_r102_c117 bl_117 br_117 wl_102 vdd gnd cell_6t
Xbit_r103_c117 bl_117 br_117 wl_103 vdd gnd cell_6t
Xbit_r104_c117 bl_117 br_117 wl_104 vdd gnd cell_6t
Xbit_r105_c117 bl_117 br_117 wl_105 vdd gnd cell_6t
Xbit_r106_c117 bl_117 br_117 wl_106 vdd gnd cell_6t
Xbit_r107_c117 bl_117 br_117 wl_107 vdd gnd cell_6t
Xbit_r108_c117 bl_117 br_117 wl_108 vdd gnd cell_6t
Xbit_r109_c117 bl_117 br_117 wl_109 vdd gnd cell_6t
Xbit_r110_c117 bl_117 br_117 wl_110 vdd gnd cell_6t
Xbit_r111_c117 bl_117 br_117 wl_111 vdd gnd cell_6t
Xbit_r112_c117 bl_117 br_117 wl_112 vdd gnd cell_6t
Xbit_r113_c117 bl_117 br_117 wl_113 vdd gnd cell_6t
Xbit_r114_c117 bl_117 br_117 wl_114 vdd gnd cell_6t
Xbit_r115_c117 bl_117 br_117 wl_115 vdd gnd cell_6t
Xbit_r116_c117 bl_117 br_117 wl_116 vdd gnd cell_6t
Xbit_r117_c117 bl_117 br_117 wl_117 vdd gnd cell_6t
Xbit_r118_c117 bl_117 br_117 wl_118 vdd gnd cell_6t
Xbit_r119_c117 bl_117 br_117 wl_119 vdd gnd cell_6t
Xbit_r120_c117 bl_117 br_117 wl_120 vdd gnd cell_6t
Xbit_r121_c117 bl_117 br_117 wl_121 vdd gnd cell_6t
Xbit_r122_c117 bl_117 br_117 wl_122 vdd gnd cell_6t
Xbit_r123_c117 bl_117 br_117 wl_123 vdd gnd cell_6t
Xbit_r124_c117 bl_117 br_117 wl_124 vdd gnd cell_6t
Xbit_r125_c117 bl_117 br_117 wl_125 vdd gnd cell_6t
Xbit_r126_c117 bl_117 br_117 wl_126 vdd gnd cell_6t
Xbit_r127_c117 bl_117 br_117 wl_127 vdd gnd cell_6t
Xbit_r128_c117 bl_117 br_117 wl_128 vdd gnd cell_6t
Xbit_r129_c117 bl_117 br_117 wl_129 vdd gnd cell_6t
Xbit_r130_c117 bl_117 br_117 wl_130 vdd gnd cell_6t
Xbit_r131_c117 bl_117 br_117 wl_131 vdd gnd cell_6t
Xbit_r132_c117 bl_117 br_117 wl_132 vdd gnd cell_6t
Xbit_r133_c117 bl_117 br_117 wl_133 vdd gnd cell_6t
Xbit_r134_c117 bl_117 br_117 wl_134 vdd gnd cell_6t
Xbit_r135_c117 bl_117 br_117 wl_135 vdd gnd cell_6t
Xbit_r136_c117 bl_117 br_117 wl_136 vdd gnd cell_6t
Xbit_r137_c117 bl_117 br_117 wl_137 vdd gnd cell_6t
Xbit_r138_c117 bl_117 br_117 wl_138 vdd gnd cell_6t
Xbit_r139_c117 bl_117 br_117 wl_139 vdd gnd cell_6t
Xbit_r140_c117 bl_117 br_117 wl_140 vdd gnd cell_6t
Xbit_r141_c117 bl_117 br_117 wl_141 vdd gnd cell_6t
Xbit_r142_c117 bl_117 br_117 wl_142 vdd gnd cell_6t
Xbit_r143_c117 bl_117 br_117 wl_143 vdd gnd cell_6t
Xbit_r144_c117 bl_117 br_117 wl_144 vdd gnd cell_6t
Xbit_r145_c117 bl_117 br_117 wl_145 vdd gnd cell_6t
Xbit_r146_c117 bl_117 br_117 wl_146 vdd gnd cell_6t
Xbit_r147_c117 bl_117 br_117 wl_147 vdd gnd cell_6t
Xbit_r148_c117 bl_117 br_117 wl_148 vdd gnd cell_6t
Xbit_r149_c117 bl_117 br_117 wl_149 vdd gnd cell_6t
Xbit_r150_c117 bl_117 br_117 wl_150 vdd gnd cell_6t
Xbit_r151_c117 bl_117 br_117 wl_151 vdd gnd cell_6t
Xbit_r152_c117 bl_117 br_117 wl_152 vdd gnd cell_6t
Xbit_r153_c117 bl_117 br_117 wl_153 vdd gnd cell_6t
Xbit_r154_c117 bl_117 br_117 wl_154 vdd gnd cell_6t
Xbit_r155_c117 bl_117 br_117 wl_155 vdd gnd cell_6t
Xbit_r156_c117 bl_117 br_117 wl_156 vdd gnd cell_6t
Xbit_r157_c117 bl_117 br_117 wl_157 vdd gnd cell_6t
Xbit_r158_c117 bl_117 br_117 wl_158 vdd gnd cell_6t
Xbit_r159_c117 bl_117 br_117 wl_159 vdd gnd cell_6t
Xbit_r160_c117 bl_117 br_117 wl_160 vdd gnd cell_6t
Xbit_r161_c117 bl_117 br_117 wl_161 vdd gnd cell_6t
Xbit_r162_c117 bl_117 br_117 wl_162 vdd gnd cell_6t
Xbit_r163_c117 bl_117 br_117 wl_163 vdd gnd cell_6t
Xbit_r164_c117 bl_117 br_117 wl_164 vdd gnd cell_6t
Xbit_r165_c117 bl_117 br_117 wl_165 vdd gnd cell_6t
Xbit_r166_c117 bl_117 br_117 wl_166 vdd gnd cell_6t
Xbit_r167_c117 bl_117 br_117 wl_167 vdd gnd cell_6t
Xbit_r168_c117 bl_117 br_117 wl_168 vdd gnd cell_6t
Xbit_r169_c117 bl_117 br_117 wl_169 vdd gnd cell_6t
Xbit_r170_c117 bl_117 br_117 wl_170 vdd gnd cell_6t
Xbit_r171_c117 bl_117 br_117 wl_171 vdd gnd cell_6t
Xbit_r172_c117 bl_117 br_117 wl_172 vdd gnd cell_6t
Xbit_r173_c117 bl_117 br_117 wl_173 vdd gnd cell_6t
Xbit_r174_c117 bl_117 br_117 wl_174 vdd gnd cell_6t
Xbit_r175_c117 bl_117 br_117 wl_175 vdd gnd cell_6t
Xbit_r176_c117 bl_117 br_117 wl_176 vdd gnd cell_6t
Xbit_r177_c117 bl_117 br_117 wl_177 vdd gnd cell_6t
Xbit_r178_c117 bl_117 br_117 wl_178 vdd gnd cell_6t
Xbit_r179_c117 bl_117 br_117 wl_179 vdd gnd cell_6t
Xbit_r180_c117 bl_117 br_117 wl_180 vdd gnd cell_6t
Xbit_r181_c117 bl_117 br_117 wl_181 vdd gnd cell_6t
Xbit_r182_c117 bl_117 br_117 wl_182 vdd gnd cell_6t
Xbit_r183_c117 bl_117 br_117 wl_183 vdd gnd cell_6t
Xbit_r184_c117 bl_117 br_117 wl_184 vdd gnd cell_6t
Xbit_r185_c117 bl_117 br_117 wl_185 vdd gnd cell_6t
Xbit_r186_c117 bl_117 br_117 wl_186 vdd gnd cell_6t
Xbit_r187_c117 bl_117 br_117 wl_187 vdd gnd cell_6t
Xbit_r188_c117 bl_117 br_117 wl_188 vdd gnd cell_6t
Xbit_r189_c117 bl_117 br_117 wl_189 vdd gnd cell_6t
Xbit_r190_c117 bl_117 br_117 wl_190 vdd gnd cell_6t
Xbit_r191_c117 bl_117 br_117 wl_191 vdd gnd cell_6t
Xbit_r192_c117 bl_117 br_117 wl_192 vdd gnd cell_6t
Xbit_r193_c117 bl_117 br_117 wl_193 vdd gnd cell_6t
Xbit_r194_c117 bl_117 br_117 wl_194 vdd gnd cell_6t
Xbit_r195_c117 bl_117 br_117 wl_195 vdd gnd cell_6t
Xbit_r196_c117 bl_117 br_117 wl_196 vdd gnd cell_6t
Xbit_r197_c117 bl_117 br_117 wl_197 vdd gnd cell_6t
Xbit_r198_c117 bl_117 br_117 wl_198 vdd gnd cell_6t
Xbit_r199_c117 bl_117 br_117 wl_199 vdd gnd cell_6t
Xbit_r200_c117 bl_117 br_117 wl_200 vdd gnd cell_6t
Xbit_r201_c117 bl_117 br_117 wl_201 vdd gnd cell_6t
Xbit_r202_c117 bl_117 br_117 wl_202 vdd gnd cell_6t
Xbit_r203_c117 bl_117 br_117 wl_203 vdd gnd cell_6t
Xbit_r204_c117 bl_117 br_117 wl_204 vdd gnd cell_6t
Xbit_r205_c117 bl_117 br_117 wl_205 vdd gnd cell_6t
Xbit_r206_c117 bl_117 br_117 wl_206 vdd gnd cell_6t
Xbit_r207_c117 bl_117 br_117 wl_207 vdd gnd cell_6t
Xbit_r208_c117 bl_117 br_117 wl_208 vdd gnd cell_6t
Xbit_r209_c117 bl_117 br_117 wl_209 vdd gnd cell_6t
Xbit_r210_c117 bl_117 br_117 wl_210 vdd gnd cell_6t
Xbit_r211_c117 bl_117 br_117 wl_211 vdd gnd cell_6t
Xbit_r212_c117 bl_117 br_117 wl_212 vdd gnd cell_6t
Xbit_r213_c117 bl_117 br_117 wl_213 vdd gnd cell_6t
Xbit_r214_c117 bl_117 br_117 wl_214 vdd gnd cell_6t
Xbit_r215_c117 bl_117 br_117 wl_215 vdd gnd cell_6t
Xbit_r216_c117 bl_117 br_117 wl_216 vdd gnd cell_6t
Xbit_r217_c117 bl_117 br_117 wl_217 vdd gnd cell_6t
Xbit_r218_c117 bl_117 br_117 wl_218 vdd gnd cell_6t
Xbit_r219_c117 bl_117 br_117 wl_219 vdd gnd cell_6t
Xbit_r220_c117 bl_117 br_117 wl_220 vdd gnd cell_6t
Xbit_r221_c117 bl_117 br_117 wl_221 vdd gnd cell_6t
Xbit_r222_c117 bl_117 br_117 wl_222 vdd gnd cell_6t
Xbit_r223_c117 bl_117 br_117 wl_223 vdd gnd cell_6t
Xbit_r224_c117 bl_117 br_117 wl_224 vdd gnd cell_6t
Xbit_r225_c117 bl_117 br_117 wl_225 vdd gnd cell_6t
Xbit_r226_c117 bl_117 br_117 wl_226 vdd gnd cell_6t
Xbit_r227_c117 bl_117 br_117 wl_227 vdd gnd cell_6t
Xbit_r228_c117 bl_117 br_117 wl_228 vdd gnd cell_6t
Xbit_r229_c117 bl_117 br_117 wl_229 vdd gnd cell_6t
Xbit_r230_c117 bl_117 br_117 wl_230 vdd gnd cell_6t
Xbit_r231_c117 bl_117 br_117 wl_231 vdd gnd cell_6t
Xbit_r232_c117 bl_117 br_117 wl_232 vdd gnd cell_6t
Xbit_r233_c117 bl_117 br_117 wl_233 vdd gnd cell_6t
Xbit_r234_c117 bl_117 br_117 wl_234 vdd gnd cell_6t
Xbit_r235_c117 bl_117 br_117 wl_235 vdd gnd cell_6t
Xbit_r236_c117 bl_117 br_117 wl_236 vdd gnd cell_6t
Xbit_r237_c117 bl_117 br_117 wl_237 vdd gnd cell_6t
Xbit_r238_c117 bl_117 br_117 wl_238 vdd gnd cell_6t
Xbit_r239_c117 bl_117 br_117 wl_239 vdd gnd cell_6t
Xbit_r240_c117 bl_117 br_117 wl_240 vdd gnd cell_6t
Xbit_r241_c117 bl_117 br_117 wl_241 vdd gnd cell_6t
Xbit_r242_c117 bl_117 br_117 wl_242 vdd gnd cell_6t
Xbit_r243_c117 bl_117 br_117 wl_243 vdd gnd cell_6t
Xbit_r244_c117 bl_117 br_117 wl_244 vdd gnd cell_6t
Xbit_r245_c117 bl_117 br_117 wl_245 vdd gnd cell_6t
Xbit_r246_c117 bl_117 br_117 wl_246 vdd gnd cell_6t
Xbit_r247_c117 bl_117 br_117 wl_247 vdd gnd cell_6t
Xbit_r248_c117 bl_117 br_117 wl_248 vdd gnd cell_6t
Xbit_r249_c117 bl_117 br_117 wl_249 vdd gnd cell_6t
Xbit_r250_c117 bl_117 br_117 wl_250 vdd gnd cell_6t
Xbit_r251_c117 bl_117 br_117 wl_251 vdd gnd cell_6t
Xbit_r252_c117 bl_117 br_117 wl_252 vdd gnd cell_6t
Xbit_r253_c117 bl_117 br_117 wl_253 vdd gnd cell_6t
Xbit_r254_c117 bl_117 br_117 wl_254 vdd gnd cell_6t
Xbit_r255_c117 bl_117 br_117 wl_255 vdd gnd cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd cell_6t
Xbit_r1_c118 bl_118 br_118 wl_1 vdd gnd cell_6t
Xbit_r2_c118 bl_118 br_118 wl_2 vdd gnd cell_6t
Xbit_r3_c118 bl_118 br_118 wl_3 vdd gnd cell_6t
Xbit_r4_c118 bl_118 br_118 wl_4 vdd gnd cell_6t
Xbit_r5_c118 bl_118 br_118 wl_5 vdd gnd cell_6t
Xbit_r6_c118 bl_118 br_118 wl_6 vdd gnd cell_6t
Xbit_r7_c118 bl_118 br_118 wl_7 vdd gnd cell_6t
Xbit_r8_c118 bl_118 br_118 wl_8 vdd gnd cell_6t
Xbit_r9_c118 bl_118 br_118 wl_9 vdd gnd cell_6t
Xbit_r10_c118 bl_118 br_118 wl_10 vdd gnd cell_6t
Xbit_r11_c118 bl_118 br_118 wl_11 vdd gnd cell_6t
Xbit_r12_c118 bl_118 br_118 wl_12 vdd gnd cell_6t
Xbit_r13_c118 bl_118 br_118 wl_13 vdd gnd cell_6t
Xbit_r14_c118 bl_118 br_118 wl_14 vdd gnd cell_6t
Xbit_r15_c118 bl_118 br_118 wl_15 vdd gnd cell_6t
Xbit_r16_c118 bl_118 br_118 wl_16 vdd gnd cell_6t
Xbit_r17_c118 bl_118 br_118 wl_17 vdd gnd cell_6t
Xbit_r18_c118 bl_118 br_118 wl_18 vdd gnd cell_6t
Xbit_r19_c118 bl_118 br_118 wl_19 vdd gnd cell_6t
Xbit_r20_c118 bl_118 br_118 wl_20 vdd gnd cell_6t
Xbit_r21_c118 bl_118 br_118 wl_21 vdd gnd cell_6t
Xbit_r22_c118 bl_118 br_118 wl_22 vdd gnd cell_6t
Xbit_r23_c118 bl_118 br_118 wl_23 vdd gnd cell_6t
Xbit_r24_c118 bl_118 br_118 wl_24 vdd gnd cell_6t
Xbit_r25_c118 bl_118 br_118 wl_25 vdd gnd cell_6t
Xbit_r26_c118 bl_118 br_118 wl_26 vdd gnd cell_6t
Xbit_r27_c118 bl_118 br_118 wl_27 vdd gnd cell_6t
Xbit_r28_c118 bl_118 br_118 wl_28 vdd gnd cell_6t
Xbit_r29_c118 bl_118 br_118 wl_29 vdd gnd cell_6t
Xbit_r30_c118 bl_118 br_118 wl_30 vdd gnd cell_6t
Xbit_r31_c118 bl_118 br_118 wl_31 vdd gnd cell_6t
Xbit_r32_c118 bl_118 br_118 wl_32 vdd gnd cell_6t
Xbit_r33_c118 bl_118 br_118 wl_33 vdd gnd cell_6t
Xbit_r34_c118 bl_118 br_118 wl_34 vdd gnd cell_6t
Xbit_r35_c118 bl_118 br_118 wl_35 vdd gnd cell_6t
Xbit_r36_c118 bl_118 br_118 wl_36 vdd gnd cell_6t
Xbit_r37_c118 bl_118 br_118 wl_37 vdd gnd cell_6t
Xbit_r38_c118 bl_118 br_118 wl_38 vdd gnd cell_6t
Xbit_r39_c118 bl_118 br_118 wl_39 vdd gnd cell_6t
Xbit_r40_c118 bl_118 br_118 wl_40 vdd gnd cell_6t
Xbit_r41_c118 bl_118 br_118 wl_41 vdd gnd cell_6t
Xbit_r42_c118 bl_118 br_118 wl_42 vdd gnd cell_6t
Xbit_r43_c118 bl_118 br_118 wl_43 vdd gnd cell_6t
Xbit_r44_c118 bl_118 br_118 wl_44 vdd gnd cell_6t
Xbit_r45_c118 bl_118 br_118 wl_45 vdd gnd cell_6t
Xbit_r46_c118 bl_118 br_118 wl_46 vdd gnd cell_6t
Xbit_r47_c118 bl_118 br_118 wl_47 vdd gnd cell_6t
Xbit_r48_c118 bl_118 br_118 wl_48 vdd gnd cell_6t
Xbit_r49_c118 bl_118 br_118 wl_49 vdd gnd cell_6t
Xbit_r50_c118 bl_118 br_118 wl_50 vdd gnd cell_6t
Xbit_r51_c118 bl_118 br_118 wl_51 vdd gnd cell_6t
Xbit_r52_c118 bl_118 br_118 wl_52 vdd gnd cell_6t
Xbit_r53_c118 bl_118 br_118 wl_53 vdd gnd cell_6t
Xbit_r54_c118 bl_118 br_118 wl_54 vdd gnd cell_6t
Xbit_r55_c118 bl_118 br_118 wl_55 vdd gnd cell_6t
Xbit_r56_c118 bl_118 br_118 wl_56 vdd gnd cell_6t
Xbit_r57_c118 bl_118 br_118 wl_57 vdd gnd cell_6t
Xbit_r58_c118 bl_118 br_118 wl_58 vdd gnd cell_6t
Xbit_r59_c118 bl_118 br_118 wl_59 vdd gnd cell_6t
Xbit_r60_c118 bl_118 br_118 wl_60 vdd gnd cell_6t
Xbit_r61_c118 bl_118 br_118 wl_61 vdd gnd cell_6t
Xbit_r62_c118 bl_118 br_118 wl_62 vdd gnd cell_6t
Xbit_r63_c118 bl_118 br_118 wl_63 vdd gnd cell_6t
Xbit_r64_c118 bl_118 br_118 wl_64 vdd gnd cell_6t
Xbit_r65_c118 bl_118 br_118 wl_65 vdd gnd cell_6t
Xbit_r66_c118 bl_118 br_118 wl_66 vdd gnd cell_6t
Xbit_r67_c118 bl_118 br_118 wl_67 vdd gnd cell_6t
Xbit_r68_c118 bl_118 br_118 wl_68 vdd gnd cell_6t
Xbit_r69_c118 bl_118 br_118 wl_69 vdd gnd cell_6t
Xbit_r70_c118 bl_118 br_118 wl_70 vdd gnd cell_6t
Xbit_r71_c118 bl_118 br_118 wl_71 vdd gnd cell_6t
Xbit_r72_c118 bl_118 br_118 wl_72 vdd gnd cell_6t
Xbit_r73_c118 bl_118 br_118 wl_73 vdd gnd cell_6t
Xbit_r74_c118 bl_118 br_118 wl_74 vdd gnd cell_6t
Xbit_r75_c118 bl_118 br_118 wl_75 vdd gnd cell_6t
Xbit_r76_c118 bl_118 br_118 wl_76 vdd gnd cell_6t
Xbit_r77_c118 bl_118 br_118 wl_77 vdd gnd cell_6t
Xbit_r78_c118 bl_118 br_118 wl_78 vdd gnd cell_6t
Xbit_r79_c118 bl_118 br_118 wl_79 vdd gnd cell_6t
Xbit_r80_c118 bl_118 br_118 wl_80 vdd gnd cell_6t
Xbit_r81_c118 bl_118 br_118 wl_81 vdd gnd cell_6t
Xbit_r82_c118 bl_118 br_118 wl_82 vdd gnd cell_6t
Xbit_r83_c118 bl_118 br_118 wl_83 vdd gnd cell_6t
Xbit_r84_c118 bl_118 br_118 wl_84 vdd gnd cell_6t
Xbit_r85_c118 bl_118 br_118 wl_85 vdd gnd cell_6t
Xbit_r86_c118 bl_118 br_118 wl_86 vdd gnd cell_6t
Xbit_r87_c118 bl_118 br_118 wl_87 vdd gnd cell_6t
Xbit_r88_c118 bl_118 br_118 wl_88 vdd gnd cell_6t
Xbit_r89_c118 bl_118 br_118 wl_89 vdd gnd cell_6t
Xbit_r90_c118 bl_118 br_118 wl_90 vdd gnd cell_6t
Xbit_r91_c118 bl_118 br_118 wl_91 vdd gnd cell_6t
Xbit_r92_c118 bl_118 br_118 wl_92 vdd gnd cell_6t
Xbit_r93_c118 bl_118 br_118 wl_93 vdd gnd cell_6t
Xbit_r94_c118 bl_118 br_118 wl_94 vdd gnd cell_6t
Xbit_r95_c118 bl_118 br_118 wl_95 vdd gnd cell_6t
Xbit_r96_c118 bl_118 br_118 wl_96 vdd gnd cell_6t
Xbit_r97_c118 bl_118 br_118 wl_97 vdd gnd cell_6t
Xbit_r98_c118 bl_118 br_118 wl_98 vdd gnd cell_6t
Xbit_r99_c118 bl_118 br_118 wl_99 vdd gnd cell_6t
Xbit_r100_c118 bl_118 br_118 wl_100 vdd gnd cell_6t
Xbit_r101_c118 bl_118 br_118 wl_101 vdd gnd cell_6t
Xbit_r102_c118 bl_118 br_118 wl_102 vdd gnd cell_6t
Xbit_r103_c118 bl_118 br_118 wl_103 vdd gnd cell_6t
Xbit_r104_c118 bl_118 br_118 wl_104 vdd gnd cell_6t
Xbit_r105_c118 bl_118 br_118 wl_105 vdd gnd cell_6t
Xbit_r106_c118 bl_118 br_118 wl_106 vdd gnd cell_6t
Xbit_r107_c118 bl_118 br_118 wl_107 vdd gnd cell_6t
Xbit_r108_c118 bl_118 br_118 wl_108 vdd gnd cell_6t
Xbit_r109_c118 bl_118 br_118 wl_109 vdd gnd cell_6t
Xbit_r110_c118 bl_118 br_118 wl_110 vdd gnd cell_6t
Xbit_r111_c118 bl_118 br_118 wl_111 vdd gnd cell_6t
Xbit_r112_c118 bl_118 br_118 wl_112 vdd gnd cell_6t
Xbit_r113_c118 bl_118 br_118 wl_113 vdd gnd cell_6t
Xbit_r114_c118 bl_118 br_118 wl_114 vdd gnd cell_6t
Xbit_r115_c118 bl_118 br_118 wl_115 vdd gnd cell_6t
Xbit_r116_c118 bl_118 br_118 wl_116 vdd gnd cell_6t
Xbit_r117_c118 bl_118 br_118 wl_117 vdd gnd cell_6t
Xbit_r118_c118 bl_118 br_118 wl_118 vdd gnd cell_6t
Xbit_r119_c118 bl_118 br_118 wl_119 vdd gnd cell_6t
Xbit_r120_c118 bl_118 br_118 wl_120 vdd gnd cell_6t
Xbit_r121_c118 bl_118 br_118 wl_121 vdd gnd cell_6t
Xbit_r122_c118 bl_118 br_118 wl_122 vdd gnd cell_6t
Xbit_r123_c118 bl_118 br_118 wl_123 vdd gnd cell_6t
Xbit_r124_c118 bl_118 br_118 wl_124 vdd gnd cell_6t
Xbit_r125_c118 bl_118 br_118 wl_125 vdd gnd cell_6t
Xbit_r126_c118 bl_118 br_118 wl_126 vdd gnd cell_6t
Xbit_r127_c118 bl_118 br_118 wl_127 vdd gnd cell_6t
Xbit_r128_c118 bl_118 br_118 wl_128 vdd gnd cell_6t
Xbit_r129_c118 bl_118 br_118 wl_129 vdd gnd cell_6t
Xbit_r130_c118 bl_118 br_118 wl_130 vdd gnd cell_6t
Xbit_r131_c118 bl_118 br_118 wl_131 vdd gnd cell_6t
Xbit_r132_c118 bl_118 br_118 wl_132 vdd gnd cell_6t
Xbit_r133_c118 bl_118 br_118 wl_133 vdd gnd cell_6t
Xbit_r134_c118 bl_118 br_118 wl_134 vdd gnd cell_6t
Xbit_r135_c118 bl_118 br_118 wl_135 vdd gnd cell_6t
Xbit_r136_c118 bl_118 br_118 wl_136 vdd gnd cell_6t
Xbit_r137_c118 bl_118 br_118 wl_137 vdd gnd cell_6t
Xbit_r138_c118 bl_118 br_118 wl_138 vdd gnd cell_6t
Xbit_r139_c118 bl_118 br_118 wl_139 vdd gnd cell_6t
Xbit_r140_c118 bl_118 br_118 wl_140 vdd gnd cell_6t
Xbit_r141_c118 bl_118 br_118 wl_141 vdd gnd cell_6t
Xbit_r142_c118 bl_118 br_118 wl_142 vdd gnd cell_6t
Xbit_r143_c118 bl_118 br_118 wl_143 vdd gnd cell_6t
Xbit_r144_c118 bl_118 br_118 wl_144 vdd gnd cell_6t
Xbit_r145_c118 bl_118 br_118 wl_145 vdd gnd cell_6t
Xbit_r146_c118 bl_118 br_118 wl_146 vdd gnd cell_6t
Xbit_r147_c118 bl_118 br_118 wl_147 vdd gnd cell_6t
Xbit_r148_c118 bl_118 br_118 wl_148 vdd gnd cell_6t
Xbit_r149_c118 bl_118 br_118 wl_149 vdd gnd cell_6t
Xbit_r150_c118 bl_118 br_118 wl_150 vdd gnd cell_6t
Xbit_r151_c118 bl_118 br_118 wl_151 vdd gnd cell_6t
Xbit_r152_c118 bl_118 br_118 wl_152 vdd gnd cell_6t
Xbit_r153_c118 bl_118 br_118 wl_153 vdd gnd cell_6t
Xbit_r154_c118 bl_118 br_118 wl_154 vdd gnd cell_6t
Xbit_r155_c118 bl_118 br_118 wl_155 vdd gnd cell_6t
Xbit_r156_c118 bl_118 br_118 wl_156 vdd gnd cell_6t
Xbit_r157_c118 bl_118 br_118 wl_157 vdd gnd cell_6t
Xbit_r158_c118 bl_118 br_118 wl_158 vdd gnd cell_6t
Xbit_r159_c118 bl_118 br_118 wl_159 vdd gnd cell_6t
Xbit_r160_c118 bl_118 br_118 wl_160 vdd gnd cell_6t
Xbit_r161_c118 bl_118 br_118 wl_161 vdd gnd cell_6t
Xbit_r162_c118 bl_118 br_118 wl_162 vdd gnd cell_6t
Xbit_r163_c118 bl_118 br_118 wl_163 vdd gnd cell_6t
Xbit_r164_c118 bl_118 br_118 wl_164 vdd gnd cell_6t
Xbit_r165_c118 bl_118 br_118 wl_165 vdd gnd cell_6t
Xbit_r166_c118 bl_118 br_118 wl_166 vdd gnd cell_6t
Xbit_r167_c118 bl_118 br_118 wl_167 vdd gnd cell_6t
Xbit_r168_c118 bl_118 br_118 wl_168 vdd gnd cell_6t
Xbit_r169_c118 bl_118 br_118 wl_169 vdd gnd cell_6t
Xbit_r170_c118 bl_118 br_118 wl_170 vdd gnd cell_6t
Xbit_r171_c118 bl_118 br_118 wl_171 vdd gnd cell_6t
Xbit_r172_c118 bl_118 br_118 wl_172 vdd gnd cell_6t
Xbit_r173_c118 bl_118 br_118 wl_173 vdd gnd cell_6t
Xbit_r174_c118 bl_118 br_118 wl_174 vdd gnd cell_6t
Xbit_r175_c118 bl_118 br_118 wl_175 vdd gnd cell_6t
Xbit_r176_c118 bl_118 br_118 wl_176 vdd gnd cell_6t
Xbit_r177_c118 bl_118 br_118 wl_177 vdd gnd cell_6t
Xbit_r178_c118 bl_118 br_118 wl_178 vdd gnd cell_6t
Xbit_r179_c118 bl_118 br_118 wl_179 vdd gnd cell_6t
Xbit_r180_c118 bl_118 br_118 wl_180 vdd gnd cell_6t
Xbit_r181_c118 bl_118 br_118 wl_181 vdd gnd cell_6t
Xbit_r182_c118 bl_118 br_118 wl_182 vdd gnd cell_6t
Xbit_r183_c118 bl_118 br_118 wl_183 vdd gnd cell_6t
Xbit_r184_c118 bl_118 br_118 wl_184 vdd gnd cell_6t
Xbit_r185_c118 bl_118 br_118 wl_185 vdd gnd cell_6t
Xbit_r186_c118 bl_118 br_118 wl_186 vdd gnd cell_6t
Xbit_r187_c118 bl_118 br_118 wl_187 vdd gnd cell_6t
Xbit_r188_c118 bl_118 br_118 wl_188 vdd gnd cell_6t
Xbit_r189_c118 bl_118 br_118 wl_189 vdd gnd cell_6t
Xbit_r190_c118 bl_118 br_118 wl_190 vdd gnd cell_6t
Xbit_r191_c118 bl_118 br_118 wl_191 vdd gnd cell_6t
Xbit_r192_c118 bl_118 br_118 wl_192 vdd gnd cell_6t
Xbit_r193_c118 bl_118 br_118 wl_193 vdd gnd cell_6t
Xbit_r194_c118 bl_118 br_118 wl_194 vdd gnd cell_6t
Xbit_r195_c118 bl_118 br_118 wl_195 vdd gnd cell_6t
Xbit_r196_c118 bl_118 br_118 wl_196 vdd gnd cell_6t
Xbit_r197_c118 bl_118 br_118 wl_197 vdd gnd cell_6t
Xbit_r198_c118 bl_118 br_118 wl_198 vdd gnd cell_6t
Xbit_r199_c118 bl_118 br_118 wl_199 vdd gnd cell_6t
Xbit_r200_c118 bl_118 br_118 wl_200 vdd gnd cell_6t
Xbit_r201_c118 bl_118 br_118 wl_201 vdd gnd cell_6t
Xbit_r202_c118 bl_118 br_118 wl_202 vdd gnd cell_6t
Xbit_r203_c118 bl_118 br_118 wl_203 vdd gnd cell_6t
Xbit_r204_c118 bl_118 br_118 wl_204 vdd gnd cell_6t
Xbit_r205_c118 bl_118 br_118 wl_205 vdd gnd cell_6t
Xbit_r206_c118 bl_118 br_118 wl_206 vdd gnd cell_6t
Xbit_r207_c118 bl_118 br_118 wl_207 vdd gnd cell_6t
Xbit_r208_c118 bl_118 br_118 wl_208 vdd gnd cell_6t
Xbit_r209_c118 bl_118 br_118 wl_209 vdd gnd cell_6t
Xbit_r210_c118 bl_118 br_118 wl_210 vdd gnd cell_6t
Xbit_r211_c118 bl_118 br_118 wl_211 vdd gnd cell_6t
Xbit_r212_c118 bl_118 br_118 wl_212 vdd gnd cell_6t
Xbit_r213_c118 bl_118 br_118 wl_213 vdd gnd cell_6t
Xbit_r214_c118 bl_118 br_118 wl_214 vdd gnd cell_6t
Xbit_r215_c118 bl_118 br_118 wl_215 vdd gnd cell_6t
Xbit_r216_c118 bl_118 br_118 wl_216 vdd gnd cell_6t
Xbit_r217_c118 bl_118 br_118 wl_217 vdd gnd cell_6t
Xbit_r218_c118 bl_118 br_118 wl_218 vdd gnd cell_6t
Xbit_r219_c118 bl_118 br_118 wl_219 vdd gnd cell_6t
Xbit_r220_c118 bl_118 br_118 wl_220 vdd gnd cell_6t
Xbit_r221_c118 bl_118 br_118 wl_221 vdd gnd cell_6t
Xbit_r222_c118 bl_118 br_118 wl_222 vdd gnd cell_6t
Xbit_r223_c118 bl_118 br_118 wl_223 vdd gnd cell_6t
Xbit_r224_c118 bl_118 br_118 wl_224 vdd gnd cell_6t
Xbit_r225_c118 bl_118 br_118 wl_225 vdd gnd cell_6t
Xbit_r226_c118 bl_118 br_118 wl_226 vdd gnd cell_6t
Xbit_r227_c118 bl_118 br_118 wl_227 vdd gnd cell_6t
Xbit_r228_c118 bl_118 br_118 wl_228 vdd gnd cell_6t
Xbit_r229_c118 bl_118 br_118 wl_229 vdd gnd cell_6t
Xbit_r230_c118 bl_118 br_118 wl_230 vdd gnd cell_6t
Xbit_r231_c118 bl_118 br_118 wl_231 vdd gnd cell_6t
Xbit_r232_c118 bl_118 br_118 wl_232 vdd gnd cell_6t
Xbit_r233_c118 bl_118 br_118 wl_233 vdd gnd cell_6t
Xbit_r234_c118 bl_118 br_118 wl_234 vdd gnd cell_6t
Xbit_r235_c118 bl_118 br_118 wl_235 vdd gnd cell_6t
Xbit_r236_c118 bl_118 br_118 wl_236 vdd gnd cell_6t
Xbit_r237_c118 bl_118 br_118 wl_237 vdd gnd cell_6t
Xbit_r238_c118 bl_118 br_118 wl_238 vdd gnd cell_6t
Xbit_r239_c118 bl_118 br_118 wl_239 vdd gnd cell_6t
Xbit_r240_c118 bl_118 br_118 wl_240 vdd gnd cell_6t
Xbit_r241_c118 bl_118 br_118 wl_241 vdd gnd cell_6t
Xbit_r242_c118 bl_118 br_118 wl_242 vdd gnd cell_6t
Xbit_r243_c118 bl_118 br_118 wl_243 vdd gnd cell_6t
Xbit_r244_c118 bl_118 br_118 wl_244 vdd gnd cell_6t
Xbit_r245_c118 bl_118 br_118 wl_245 vdd gnd cell_6t
Xbit_r246_c118 bl_118 br_118 wl_246 vdd gnd cell_6t
Xbit_r247_c118 bl_118 br_118 wl_247 vdd gnd cell_6t
Xbit_r248_c118 bl_118 br_118 wl_248 vdd gnd cell_6t
Xbit_r249_c118 bl_118 br_118 wl_249 vdd gnd cell_6t
Xbit_r250_c118 bl_118 br_118 wl_250 vdd gnd cell_6t
Xbit_r251_c118 bl_118 br_118 wl_251 vdd gnd cell_6t
Xbit_r252_c118 bl_118 br_118 wl_252 vdd gnd cell_6t
Xbit_r253_c118 bl_118 br_118 wl_253 vdd gnd cell_6t
Xbit_r254_c118 bl_118 br_118 wl_254 vdd gnd cell_6t
Xbit_r255_c118 bl_118 br_118 wl_255 vdd gnd cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd cell_6t
Xbit_r1_c119 bl_119 br_119 wl_1 vdd gnd cell_6t
Xbit_r2_c119 bl_119 br_119 wl_2 vdd gnd cell_6t
Xbit_r3_c119 bl_119 br_119 wl_3 vdd gnd cell_6t
Xbit_r4_c119 bl_119 br_119 wl_4 vdd gnd cell_6t
Xbit_r5_c119 bl_119 br_119 wl_5 vdd gnd cell_6t
Xbit_r6_c119 bl_119 br_119 wl_6 vdd gnd cell_6t
Xbit_r7_c119 bl_119 br_119 wl_7 vdd gnd cell_6t
Xbit_r8_c119 bl_119 br_119 wl_8 vdd gnd cell_6t
Xbit_r9_c119 bl_119 br_119 wl_9 vdd gnd cell_6t
Xbit_r10_c119 bl_119 br_119 wl_10 vdd gnd cell_6t
Xbit_r11_c119 bl_119 br_119 wl_11 vdd gnd cell_6t
Xbit_r12_c119 bl_119 br_119 wl_12 vdd gnd cell_6t
Xbit_r13_c119 bl_119 br_119 wl_13 vdd gnd cell_6t
Xbit_r14_c119 bl_119 br_119 wl_14 vdd gnd cell_6t
Xbit_r15_c119 bl_119 br_119 wl_15 vdd gnd cell_6t
Xbit_r16_c119 bl_119 br_119 wl_16 vdd gnd cell_6t
Xbit_r17_c119 bl_119 br_119 wl_17 vdd gnd cell_6t
Xbit_r18_c119 bl_119 br_119 wl_18 vdd gnd cell_6t
Xbit_r19_c119 bl_119 br_119 wl_19 vdd gnd cell_6t
Xbit_r20_c119 bl_119 br_119 wl_20 vdd gnd cell_6t
Xbit_r21_c119 bl_119 br_119 wl_21 vdd gnd cell_6t
Xbit_r22_c119 bl_119 br_119 wl_22 vdd gnd cell_6t
Xbit_r23_c119 bl_119 br_119 wl_23 vdd gnd cell_6t
Xbit_r24_c119 bl_119 br_119 wl_24 vdd gnd cell_6t
Xbit_r25_c119 bl_119 br_119 wl_25 vdd gnd cell_6t
Xbit_r26_c119 bl_119 br_119 wl_26 vdd gnd cell_6t
Xbit_r27_c119 bl_119 br_119 wl_27 vdd gnd cell_6t
Xbit_r28_c119 bl_119 br_119 wl_28 vdd gnd cell_6t
Xbit_r29_c119 bl_119 br_119 wl_29 vdd gnd cell_6t
Xbit_r30_c119 bl_119 br_119 wl_30 vdd gnd cell_6t
Xbit_r31_c119 bl_119 br_119 wl_31 vdd gnd cell_6t
Xbit_r32_c119 bl_119 br_119 wl_32 vdd gnd cell_6t
Xbit_r33_c119 bl_119 br_119 wl_33 vdd gnd cell_6t
Xbit_r34_c119 bl_119 br_119 wl_34 vdd gnd cell_6t
Xbit_r35_c119 bl_119 br_119 wl_35 vdd gnd cell_6t
Xbit_r36_c119 bl_119 br_119 wl_36 vdd gnd cell_6t
Xbit_r37_c119 bl_119 br_119 wl_37 vdd gnd cell_6t
Xbit_r38_c119 bl_119 br_119 wl_38 vdd gnd cell_6t
Xbit_r39_c119 bl_119 br_119 wl_39 vdd gnd cell_6t
Xbit_r40_c119 bl_119 br_119 wl_40 vdd gnd cell_6t
Xbit_r41_c119 bl_119 br_119 wl_41 vdd gnd cell_6t
Xbit_r42_c119 bl_119 br_119 wl_42 vdd gnd cell_6t
Xbit_r43_c119 bl_119 br_119 wl_43 vdd gnd cell_6t
Xbit_r44_c119 bl_119 br_119 wl_44 vdd gnd cell_6t
Xbit_r45_c119 bl_119 br_119 wl_45 vdd gnd cell_6t
Xbit_r46_c119 bl_119 br_119 wl_46 vdd gnd cell_6t
Xbit_r47_c119 bl_119 br_119 wl_47 vdd gnd cell_6t
Xbit_r48_c119 bl_119 br_119 wl_48 vdd gnd cell_6t
Xbit_r49_c119 bl_119 br_119 wl_49 vdd gnd cell_6t
Xbit_r50_c119 bl_119 br_119 wl_50 vdd gnd cell_6t
Xbit_r51_c119 bl_119 br_119 wl_51 vdd gnd cell_6t
Xbit_r52_c119 bl_119 br_119 wl_52 vdd gnd cell_6t
Xbit_r53_c119 bl_119 br_119 wl_53 vdd gnd cell_6t
Xbit_r54_c119 bl_119 br_119 wl_54 vdd gnd cell_6t
Xbit_r55_c119 bl_119 br_119 wl_55 vdd gnd cell_6t
Xbit_r56_c119 bl_119 br_119 wl_56 vdd gnd cell_6t
Xbit_r57_c119 bl_119 br_119 wl_57 vdd gnd cell_6t
Xbit_r58_c119 bl_119 br_119 wl_58 vdd gnd cell_6t
Xbit_r59_c119 bl_119 br_119 wl_59 vdd gnd cell_6t
Xbit_r60_c119 bl_119 br_119 wl_60 vdd gnd cell_6t
Xbit_r61_c119 bl_119 br_119 wl_61 vdd gnd cell_6t
Xbit_r62_c119 bl_119 br_119 wl_62 vdd gnd cell_6t
Xbit_r63_c119 bl_119 br_119 wl_63 vdd gnd cell_6t
Xbit_r64_c119 bl_119 br_119 wl_64 vdd gnd cell_6t
Xbit_r65_c119 bl_119 br_119 wl_65 vdd gnd cell_6t
Xbit_r66_c119 bl_119 br_119 wl_66 vdd gnd cell_6t
Xbit_r67_c119 bl_119 br_119 wl_67 vdd gnd cell_6t
Xbit_r68_c119 bl_119 br_119 wl_68 vdd gnd cell_6t
Xbit_r69_c119 bl_119 br_119 wl_69 vdd gnd cell_6t
Xbit_r70_c119 bl_119 br_119 wl_70 vdd gnd cell_6t
Xbit_r71_c119 bl_119 br_119 wl_71 vdd gnd cell_6t
Xbit_r72_c119 bl_119 br_119 wl_72 vdd gnd cell_6t
Xbit_r73_c119 bl_119 br_119 wl_73 vdd gnd cell_6t
Xbit_r74_c119 bl_119 br_119 wl_74 vdd gnd cell_6t
Xbit_r75_c119 bl_119 br_119 wl_75 vdd gnd cell_6t
Xbit_r76_c119 bl_119 br_119 wl_76 vdd gnd cell_6t
Xbit_r77_c119 bl_119 br_119 wl_77 vdd gnd cell_6t
Xbit_r78_c119 bl_119 br_119 wl_78 vdd gnd cell_6t
Xbit_r79_c119 bl_119 br_119 wl_79 vdd gnd cell_6t
Xbit_r80_c119 bl_119 br_119 wl_80 vdd gnd cell_6t
Xbit_r81_c119 bl_119 br_119 wl_81 vdd gnd cell_6t
Xbit_r82_c119 bl_119 br_119 wl_82 vdd gnd cell_6t
Xbit_r83_c119 bl_119 br_119 wl_83 vdd gnd cell_6t
Xbit_r84_c119 bl_119 br_119 wl_84 vdd gnd cell_6t
Xbit_r85_c119 bl_119 br_119 wl_85 vdd gnd cell_6t
Xbit_r86_c119 bl_119 br_119 wl_86 vdd gnd cell_6t
Xbit_r87_c119 bl_119 br_119 wl_87 vdd gnd cell_6t
Xbit_r88_c119 bl_119 br_119 wl_88 vdd gnd cell_6t
Xbit_r89_c119 bl_119 br_119 wl_89 vdd gnd cell_6t
Xbit_r90_c119 bl_119 br_119 wl_90 vdd gnd cell_6t
Xbit_r91_c119 bl_119 br_119 wl_91 vdd gnd cell_6t
Xbit_r92_c119 bl_119 br_119 wl_92 vdd gnd cell_6t
Xbit_r93_c119 bl_119 br_119 wl_93 vdd gnd cell_6t
Xbit_r94_c119 bl_119 br_119 wl_94 vdd gnd cell_6t
Xbit_r95_c119 bl_119 br_119 wl_95 vdd gnd cell_6t
Xbit_r96_c119 bl_119 br_119 wl_96 vdd gnd cell_6t
Xbit_r97_c119 bl_119 br_119 wl_97 vdd gnd cell_6t
Xbit_r98_c119 bl_119 br_119 wl_98 vdd gnd cell_6t
Xbit_r99_c119 bl_119 br_119 wl_99 vdd gnd cell_6t
Xbit_r100_c119 bl_119 br_119 wl_100 vdd gnd cell_6t
Xbit_r101_c119 bl_119 br_119 wl_101 vdd gnd cell_6t
Xbit_r102_c119 bl_119 br_119 wl_102 vdd gnd cell_6t
Xbit_r103_c119 bl_119 br_119 wl_103 vdd gnd cell_6t
Xbit_r104_c119 bl_119 br_119 wl_104 vdd gnd cell_6t
Xbit_r105_c119 bl_119 br_119 wl_105 vdd gnd cell_6t
Xbit_r106_c119 bl_119 br_119 wl_106 vdd gnd cell_6t
Xbit_r107_c119 bl_119 br_119 wl_107 vdd gnd cell_6t
Xbit_r108_c119 bl_119 br_119 wl_108 vdd gnd cell_6t
Xbit_r109_c119 bl_119 br_119 wl_109 vdd gnd cell_6t
Xbit_r110_c119 bl_119 br_119 wl_110 vdd gnd cell_6t
Xbit_r111_c119 bl_119 br_119 wl_111 vdd gnd cell_6t
Xbit_r112_c119 bl_119 br_119 wl_112 vdd gnd cell_6t
Xbit_r113_c119 bl_119 br_119 wl_113 vdd gnd cell_6t
Xbit_r114_c119 bl_119 br_119 wl_114 vdd gnd cell_6t
Xbit_r115_c119 bl_119 br_119 wl_115 vdd gnd cell_6t
Xbit_r116_c119 bl_119 br_119 wl_116 vdd gnd cell_6t
Xbit_r117_c119 bl_119 br_119 wl_117 vdd gnd cell_6t
Xbit_r118_c119 bl_119 br_119 wl_118 vdd gnd cell_6t
Xbit_r119_c119 bl_119 br_119 wl_119 vdd gnd cell_6t
Xbit_r120_c119 bl_119 br_119 wl_120 vdd gnd cell_6t
Xbit_r121_c119 bl_119 br_119 wl_121 vdd gnd cell_6t
Xbit_r122_c119 bl_119 br_119 wl_122 vdd gnd cell_6t
Xbit_r123_c119 bl_119 br_119 wl_123 vdd gnd cell_6t
Xbit_r124_c119 bl_119 br_119 wl_124 vdd gnd cell_6t
Xbit_r125_c119 bl_119 br_119 wl_125 vdd gnd cell_6t
Xbit_r126_c119 bl_119 br_119 wl_126 vdd gnd cell_6t
Xbit_r127_c119 bl_119 br_119 wl_127 vdd gnd cell_6t
Xbit_r128_c119 bl_119 br_119 wl_128 vdd gnd cell_6t
Xbit_r129_c119 bl_119 br_119 wl_129 vdd gnd cell_6t
Xbit_r130_c119 bl_119 br_119 wl_130 vdd gnd cell_6t
Xbit_r131_c119 bl_119 br_119 wl_131 vdd gnd cell_6t
Xbit_r132_c119 bl_119 br_119 wl_132 vdd gnd cell_6t
Xbit_r133_c119 bl_119 br_119 wl_133 vdd gnd cell_6t
Xbit_r134_c119 bl_119 br_119 wl_134 vdd gnd cell_6t
Xbit_r135_c119 bl_119 br_119 wl_135 vdd gnd cell_6t
Xbit_r136_c119 bl_119 br_119 wl_136 vdd gnd cell_6t
Xbit_r137_c119 bl_119 br_119 wl_137 vdd gnd cell_6t
Xbit_r138_c119 bl_119 br_119 wl_138 vdd gnd cell_6t
Xbit_r139_c119 bl_119 br_119 wl_139 vdd gnd cell_6t
Xbit_r140_c119 bl_119 br_119 wl_140 vdd gnd cell_6t
Xbit_r141_c119 bl_119 br_119 wl_141 vdd gnd cell_6t
Xbit_r142_c119 bl_119 br_119 wl_142 vdd gnd cell_6t
Xbit_r143_c119 bl_119 br_119 wl_143 vdd gnd cell_6t
Xbit_r144_c119 bl_119 br_119 wl_144 vdd gnd cell_6t
Xbit_r145_c119 bl_119 br_119 wl_145 vdd gnd cell_6t
Xbit_r146_c119 bl_119 br_119 wl_146 vdd gnd cell_6t
Xbit_r147_c119 bl_119 br_119 wl_147 vdd gnd cell_6t
Xbit_r148_c119 bl_119 br_119 wl_148 vdd gnd cell_6t
Xbit_r149_c119 bl_119 br_119 wl_149 vdd gnd cell_6t
Xbit_r150_c119 bl_119 br_119 wl_150 vdd gnd cell_6t
Xbit_r151_c119 bl_119 br_119 wl_151 vdd gnd cell_6t
Xbit_r152_c119 bl_119 br_119 wl_152 vdd gnd cell_6t
Xbit_r153_c119 bl_119 br_119 wl_153 vdd gnd cell_6t
Xbit_r154_c119 bl_119 br_119 wl_154 vdd gnd cell_6t
Xbit_r155_c119 bl_119 br_119 wl_155 vdd gnd cell_6t
Xbit_r156_c119 bl_119 br_119 wl_156 vdd gnd cell_6t
Xbit_r157_c119 bl_119 br_119 wl_157 vdd gnd cell_6t
Xbit_r158_c119 bl_119 br_119 wl_158 vdd gnd cell_6t
Xbit_r159_c119 bl_119 br_119 wl_159 vdd gnd cell_6t
Xbit_r160_c119 bl_119 br_119 wl_160 vdd gnd cell_6t
Xbit_r161_c119 bl_119 br_119 wl_161 vdd gnd cell_6t
Xbit_r162_c119 bl_119 br_119 wl_162 vdd gnd cell_6t
Xbit_r163_c119 bl_119 br_119 wl_163 vdd gnd cell_6t
Xbit_r164_c119 bl_119 br_119 wl_164 vdd gnd cell_6t
Xbit_r165_c119 bl_119 br_119 wl_165 vdd gnd cell_6t
Xbit_r166_c119 bl_119 br_119 wl_166 vdd gnd cell_6t
Xbit_r167_c119 bl_119 br_119 wl_167 vdd gnd cell_6t
Xbit_r168_c119 bl_119 br_119 wl_168 vdd gnd cell_6t
Xbit_r169_c119 bl_119 br_119 wl_169 vdd gnd cell_6t
Xbit_r170_c119 bl_119 br_119 wl_170 vdd gnd cell_6t
Xbit_r171_c119 bl_119 br_119 wl_171 vdd gnd cell_6t
Xbit_r172_c119 bl_119 br_119 wl_172 vdd gnd cell_6t
Xbit_r173_c119 bl_119 br_119 wl_173 vdd gnd cell_6t
Xbit_r174_c119 bl_119 br_119 wl_174 vdd gnd cell_6t
Xbit_r175_c119 bl_119 br_119 wl_175 vdd gnd cell_6t
Xbit_r176_c119 bl_119 br_119 wl_176 vdd gnd cell_6t
Xbit_r177_c119 bl_119 br_119 wl_177 vdd gnd cell_6t
Xbit_r178_c119 bl_119 br_119 wl_178 vdd gnd cell_6t
Xbit_r179_c119 bl_119 br_119 wl_179 vdd gnd cell_6t
Xbit_r180_c119 bl_119 br_119 wl_180 vdd gnd cell_6t
Xbit_r181_c119 bl_119 br_119 wl_181 vdd gnd cell_6t
Xbit_r182_c119 bl_119 br_119 wl_182 vdd gnd cell_6t
Xbit_r183_c119 bl_119 br_119 wl_183 vdd gnd cell_6t
Xbit_r184_c119 bl_119 br_119 wl_184 vdd gnd cell_6t
Xbit_r185_c119 bl_119 br_119 wl_185 vdd gnd cell_6t
Xbit_r186_c119 bl_119 br_119 wl_186 vdd gnd cell_6t
Xbit_r187_c119 bl_119 br_119 wl_187 vdd gnd cell_6t
Xbit_r188_c119 bl_119 br_119 wl_188 vdd gnd cell_6t
Xbit_r189_c119 bl_119 br_119 wl_189 vdd gnd cell_6t
Xbit_r190_c119 bl_119 br_119 wl_190 vdd gnd cell_6t
Xbit_r191_c119 bl_119 br_119 wl_191 vdd gnd cell_6t
Xbit_r192_c119 bl_119 br_119 wl_192 vdd gnd cell_6t
Xbit_r193_c119 bl_119 br_119 wl_193 vdd gnd cell_6t
Xbit_r194_c119 bl_119 br_119 wl_194 vdd gnd cell_6t
Xbit_r195_c119 bl_119 br_119 wl_195 vdd gnd cell_6t
Xbit_r196_c119 bl_119 br_119 wl_196 vdd gnd cell_6t
Xbit_r197_c119 bl_119 br_119 wl_197 vdd gnd cell_6t
Xbit_r198_c119 bl_119 br_119 wl_198 vdd gnd cell_6t
Xbit_r199_c119 bl_119 br_119 wl_199 vdd gnd cell_6t
Xbit_r200_c119 bl_119 br_119 wl_200 vdd gnd cell_6t
Xbit_r201_c119 bl_119 br_119 wl_201 vdd gnd cell_6t
Xbit_r202_c119 bl_119 br_119 wl_202 vdd gnd cell_6t
Xbit_r203_c119 bl_119 br_119 wl_203 vdd gnd cell_6t
Xbit_r204_c119 bl_119 br_119 wl_204 vdd gnd cell_6t
Xbit_r205_c119 bl_119 br_119 wl_205 vdd gnd cell_6t
Xbit_r206_c119 bl_119 br_119 wl_206 vdd gnd cell_6t
Xbit_r207_c119 bl_119 br_119 wl_207 vdd gnd cell_6t
Xbit_r208_c119 bl_119 br_119 wl_208 vdd gnd cell_6t
Xbit_r209_c119 bl_119 br_119 wl_209 vdd gnd cell_6t
Xbit_r210_c119 bl_119 br_119 wl_210 vdd gnd cell_6t
Xbit_r211_c119 bl_119 br_119 wl_211 vdd gnd cell_6t
Xbit_r212_c119 bl_119 br_119 wl_212 vdd gnd cell_6t
Xbit_r213_c119 bl_119 br_119 wl_213 vdd gnd cell_6t
Xbit_r214_c119 bl_119 br_119 wl_214 vdd gnd cell_6t
Xbit_r215_c119 bl_119 br_119 wl_215 vdd gnd cell_6t
Xbit_r216_c119 bl_119 br_119 wl_216 vdd gnd cell_6t
Xbit_r217_c119 bl_119 br_119 wl_217 vdd gnd cell_6t
Xbit_r218_c119 bl_119 br_119 wl_218 vdd gnd cell_6t
Xbit_r219_c119 bl_119 br_119 wl_219 vdd gnd cell_6t
Xbit_r220_c119 bl_119 br_119 wl_220 vdd gnd cell_6t
Xbit_r221_c119 bl_119 br_119 wl_221 vdd gnd cell_6t
Xbit_r222_c119 bl_119 br_119 wl_222 vdd gnd cell_6t
Xbit_r223_c119 bl_119 br_119 wl_223 vdd gnd cell_6t
Xbit_r224_c119 bl_119 br_119 wl_224 vdd gnd cell_6t
Xbit_r225_c119 bl_119 br_119 wl_225 vdd gnd cell_6t
Xbit_r226_c119 bl_119 br_119 wl_226 vdd gnd cell_6t
Xbit_r227_c119 bl_119 br_119 wl_227 vdd gnd cell_6t
Xbit_r228_c119 bl_119 br_119 wl_228 vdd gnd cell_6t
Xbit_r229_c119 bl_119 br_119 wl_229 vdd gnd cell_6t
Xbit_r230_c119 bl_119 br_119 wl_230 vdd gnd cell_6t
Xbit_r231_c119 bl_119 br_119 wl_231 vdd gnd cell_6t
Xbit_r232_c119 bl_119 br_119 wl_232 vdd gnd cell_6t
Xbit_r233_c119 bl_119 br_119 wl_233 vdd gnd cell_6t
Xbit_r234_c119 bl_119 br_119 wl_234 vdd gnd cell_6t
Xbit_r235_c119 bl_119 br_119 wl_235 vdd gnd cell_6t
Xbit_r236_c119 bl_119 br_119 wl_236 vdd gnd cell_6t
Xbit_r237_c119 bl_119 br_119 wl_237 vdd gnd cell_6t
Xbit_r238_c119 bl_119 br_119 wl_238 vdd gnd cell_6t
Xbit_r239_c119 bl_119 br_119 wl_239 vdd gnd cell_6t
Xbit_r240_c119 bl_119 br_119 wl_240 vdd gnd cell_6t
Xbit_r241_c119 bl_119 br_119 wl_241 vdd gnd cell_6t
Xbit_r242_c119 bl_119 br_119 wl_242 vdd gnd cell_6t
Xbit_r243_c119 bl_119 br_119 wl_243 vdd gnd cell_6t
Xbit_r244_c119 bl_119 br_119 wl_244 vdd gnd cell_6t
Xbit_r245_c119 bl_119 br_119 wl_245 vdd gnd cell_6t
Xbit_r246_c119 bl_119 br_119 wl_246 vdd gnd cell_6t
Xbit_r247_c119 bl_119 br_119 wl_247 vdd gnd cell_6t
Xbit_r248_c119 bl_119 br_119 wl_248 vdd gnd cell_6t
Xbit_r249_c119 bl_119 br_119 wl_249 vdd gnd cell_6t
Xbit_r250_c119 bl_119 br_119 wl_250 vdd gnd cell_6t
Xbit_r251_c119 bl_119 br_119 wl_251 vdd gnd cell_6t
Xbit_r252_c119 bl_119 br_119 wl_252 vdd gnd cell_6t
Xbit_r253_c119 bl_119 br_119 wl_253 vdd gnd cell_6t
Xbit_r254_c119 bl_119 br_119 wl_254 vdd gnd cell_6t
Xbit_r255_c119 bl_119 br_119 wl_255 vdd gnd cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd cell_6t
Xbit_r1_c120 bl_120 br_120 wl_1 vdd gnd cell_6t
Xbit_r2_c120 bl_120 br_120 wl_2 vdd gnd cell_6t
Xbit_r3_c120 bl_120 br_120 wl_3 vdd gnd cell_6t
Xbit_r4_c120 bl_120 br_120 wl_4 vdd gnd cell_6t
Xbit_r5_c120 bl_120 br_120 wl_5 vdd gnd cell_6t
Xbit_r6_c120 bl_120 br_120 wl_6 vdd gnd cell_6t
Xbit_r7_c120 bl_120 br_120 wl_7 vdd gnd cell_6t
Xbit_r8_c120 bl_120 br_120 wl_8 vdd gnd cell_6t
Xbit_r9_c120 bl_120 br_120 wl_9 vdd gnd cell_6t
Xbit_r10_c120 bl_120 br_120 wl_10 vdd gnd cell_6t
Xbit_r11_c120 bl_120 br_120 wl_11 vdd gnd cell_6t
Xbit_r12_c120 bl_120 br_120 wl_12 vdd gnd cell_6t
Xbit_r13_c120 bl_120 br_120 wl_13 vdd gnd cell_6t
Xbit_r14_c120 bl_120 br_120 wl_14 vdd gnd cell_6t
Xbit_r15_c120 bl_120 br_120 wl_15 vdd gnd cell_6t
Xbit_r16_c120 bl_120 br_120 wl_16 vdd gnd cell_6t
Xbit_r17_c120 bl_120 br_120 wl_17 vdd gnd cell_6t
Xbit_r18_c120 bl_120 br_120 wl_18 vdd gnd cell_6t
Xbit_r19_c120 bl_120 br_120 wl_19 vdd gnd cell_6t
Xbit_r20_c120 bl_120 br_120 wl_20 vdd gnd cell_6t
Xbit_r21_c120 bl_120 br_120 wl_21 vdd gnd cell_6t
Xbit_r22_c120 bl_120 br_120 wl_22 vdd gnd cell_6t
Xbit_r23_c120 bl_120 br_120 wl_23 vdd gnd cell_6t
Xbit_r24_c120 bl_120 br_120 wl_24 vdd gnd cell_6t
Xbit_r25_c120 bl_120 br_120 wl_25 vdd gnd cell_6t
Xbit_r26_c120 bl_120 br_120 wl_26 vdd gnd cell_6t
Xbit_r27_c120 bl_120 br_120 wl_27 vdd gnd cell_6t
Xbit_r28_c120 bl_120 br_120 wl_28 vdd gnd cell_6t
Xbit_r29_c120 bl_120 br_120 wl_29 vdd gnd cell_6t
Xbit_r30_c120 bl_120 br_120 wl_30 vdd gnd cell_6t
Xbit_r31_c120 bl_120 br_120 wl_31 vdd gnd cell_6t
Xbit_r32_c120 bl_120 br_120 wl_32 vdd gnd cell_6t
Xbit_r33_c120 bl_120 br_120 wl_33 vdd gnd cell_6t
Xbit_r34_c120 bl_120 br_120 wl_34 vdd gnd cell_6t
Xbit_r35_c120 bl_120 br_120 wl_35 vdd gnd cell_6t
Xbit_r36_c120 bl_120 br_120 wl_36 vdd gnd cell_6t
Xbit_r37_c120 bl_120 br_120 wl_37 vdd gnd cell_6t
Xbit_r38_c120 bl_120 br_120 wl_38 vdd gnd cell_6t
Xbit_r39_c120 bl_120 br_120 wl_39 vdd gnd cell_6t
Xbit_r40_c120 bl_120 br_120 wl_40 vdd gnd cell_6t
Xbit_r41_c120 bl_120 br_120 wl_41 vdd gnd cell_6t
Xbit_r42_c120 bl_120 br_120 wl_42 vdd gnd cell_6t
Xbit_r43_c120 bl_120 br_120 wl_43 vdd gnd cell_6t
Xbit_r44_c120 bl_120 br_120 wl_44 vdd gnd cell_6t
Xbit_r45_c120 bl_120 br_120 wl_45 vdd gnd cell_6t
Xbit_r46_c120 bl_120 br_120 wl_46 vdd gnd cell_6t
Xbit_r47_c120 bl_120 br_120 wl_47 vdd gnd cell_6t
Xbit_r48_c120 bl_120 br_120 wl_48 vdd gnd cell_6t
Xbit_r49_c120 bl_120 br_120 wl_49 vdd gnd cell_6t
Xbit_r50_c120 bl_120 br_120 wl_50 vdd gnd cell_6t
Xbit_r51_c120 bl_120 br_120 wl_51 vdd gnd cell_6t
Xbit_r52_c120 bl_120 br_120 wl_52 vdd gnd cell_6t
Xbit_r53_c120 bl_120 br_120 wl_53 vdd gnd cell_6t
Xbit_r54_c120 bl_120 br_120 wl_54 vdd gnd cell_6t
Xbit_r55_c120 bl_120 br_120 wl_55 vdd gnd cell_6t
Xbit_r56_c120 bl_120 br_120 wl_56 vdd gnd cell_6t
Xbit_r57_c120 bl_120 br_120 wl_57 vdd gnd cell_6t
Xbit_r58_c120 bl_120 br_120 wl_58 vdd gnd cell_6t
Xbit_r59_c120 bl_120 br_120 wl_59 vdd gnd cell_6t
Xbit_r60_c120 bl_120 br_120 wl_60 vdd gnd cell_6t
Xbit_r61_c120 bl_120 br_120 wl_61 vdd gnd cell_6t
Xbit_r62_c120 bl_120 br_120 wl_62 vdd gnd cell_6t
Xbit_r63_c120 bl_120 br_120 wl_63 vdd gnd cell_6t
Xbit_r64_c120 bl_120 br_120 wl_64 vdd gnd cell_6t
Xbit_r65_c120 bl_120 br_120 wl_65 vdd gnd cell_6t
Xbit_r66_c120 bl_120 br_120 wl_66 vdd gnd cell_6t
Xbit_r67_c120 bl_120 br_120 wl_67 vdd gnd cell_6t
Xbit_r68_c120 bl_120 br_120 wl_68 vdd gnd cell_6t
Xbit_r69_c120 bl_120 br_120 wl_69 vdd gnd cell_6t
Xbit_r70_c120 bl_120 br_120 wl_70 vdd gnd cell_6t
Xbit_r71_c120 bl_120 br_120 wl_71 vdd gnd cell_6t
Xbit_r72_c120 bl_120 br_120 wl_72 vdd gnd cell_6t
Xbit_r73_c120 bl_120 br_120 wl_73 vdd gnd cell_6t
Xbit_r74_c120 bl_120 br_120 wl_74 vdd gnd cell_6t
Xbit_r75_c120 bl_120 br_120 wl_75 vdd gnd cell_6t
Xbit_r76_c120 bl_120 br_120 wl_76 vdd gnd cell_6t
Xbit_r77_c120 bl_120 br_120 wl_77 vdd gnd cell_6t
Xbit_r78_c120 bl_120 br_120 wl_78 vdd gnd cell_6t
Xbit_r79_c120 bl_120 br_120 wl_79 vdd gnd cell_6t
Xbit_r80_c120 bl_120 br_120 wl_80 vdd gnd cell_6t
Xbit_r81_c120 bl_120 br_120 wl_81 vdd gnd cell_6t
Xbit_r82_c120 bl_120 br_120 wl_82 vdd gnd cell_6t
Xbit_r83_c120 bl_120 br_120 wl_83 vdd gnd cell_6t
Xbit_r84_c120 bl_120 br_120 wl_84 vdd gnd cell_6t
Xbit_r85_c120 bl_120 br_120 wl_85 vdd gnd cell_6t
Xbit_r86_c120 bl_120 br_120 wl_86 vdd gnd cell_6t
Xbit_r87_c120 bl_120 br_120 wl_87 vdd gnd cell_6t
Xbit_r88_c120 bl_120 br_120 wl_88 vdd gnd cell_6t
Xbit_r89_c120 bl_120 br_120 wl_89 vdd gnd cell_6t
Xbit_r90_c120 bl_120 br_120 wl_90 vdd gnd cell_6t
Xbit_r91_c120 bl_120 br_120 wl_91 vdd gnd cell_6t
Xbit_r92_c120 bl_120 br_120 wl_92 vdd gnd cell_6t
Xbit_r93_c120 bl_120 br_120 wl_93 vdd gnd cell_6t
Xbit_r94_c120 bl_120 br_120 wl_94 vdd gnd cell_6t
Xbit_r95_c120 bl_120 br_120 wl_95 vdd gnd cell_6t
Xbit_r96_c120 bl_120 br_120 wl_96 vdd gnd cell_6t
Xbit_r97_c120 bl_120 br_120 wl_97 vdd gnd cell_6t
Xbit_r98_c120 bl_120 br_120 wl_98 vdd gnd cell_6t
Xbit_r99_c120 bl_120 br_120 wl_99 vdd gnd cell_6t
Xbit_r100_c120 bl_120 br_120 wl_100 vdd gnd cell_6t
Xbit_r101_c120 bl_120 br_120 wl_101 vdd gnd cell_6t
Xbit_r102_c120 bl_120 br_120 wl_102 vdd gnd cell_6t
Xbit_r103_c120 bl_120 br_120 wl_103 vdd gnd cell_6t
Xbit_r104_c120 bl_120 br_120 wl_104 vdd gnd cell_6t
Xbit_r105_c120 bl_120 br_120 wl_105 vdd gnd cell_6t
Xbit_r106_c120 bl_120 br_120 wl_106 vdd gnd cell_6t
Xbit_r107_c120 bl_120 br_120 wl_107 vdd gnd cell_6t
Xbit_r108_c120 bl_120 br_120 wl_108 vdd gnd cell_6t
Xbit_r109_c120 bl_120 br_120 wl_109 vdd gnd cell_6t
Xbit_r110_c120 bl_120 br_120 wl_110 vdd gnd cell_6t
Xbit_r111_c120 bl_120 br_120 wl_111 vdd gnd cell_6t
Xbit_r112_c120 bl_120 br_120 wl_112 vdd gnd cell_6t
Xbit_r113_c120 bl_120 br_120 wl_113 vdd gnd cell_6t
Xbit_r114_c120 bl_120 br_120 wl_114 vdd gnd cell_6t
Xbit_r115_c120 bl_120 br_120 wl_115 vdd gnd cell_6t
Xbit_r116_c120 bl_120 br_120 wl_116 vdd gnd cell_6t
Xbit_r117_c120 bl_120 br_120 wl_117 vdd gnd cell_6t
Xbit_r118_c120 bl_120 br_120 wl_118 vdd gnd cell_6t
Xbit_r119_c120 bl_120 br_120 wl_119 vdd gnd cell_6t
Xbit_r120_c120 bl_120 br_120 wl_120 vdd gnd cell_6t
Xbit_r121_c120 bl_120 br_120 wl_121 vdd gnd cell_6t
Xbit_r122_c120 bl_120 br_120 wl_122 vdd gnd cell_6t
Xbit_r123_c120 bl_120 br_120 wl_123 vdd gnd cell_6t
Xbit_r124_c120 bl_120 br_120 wl_124 vdd gnd cell_6t
Xbit_r125_c120 bl_120 br_120 wl_125 vdd gnd cell_6t
Xbit_r126_c120 bl_120 br_120 wl_126 vdd gnd cell_6t
Xbit_r127_c120 bl_120 br_120 wl_127 vdd gnd cell_6t
Xbit_r128_c120 bl_120 br_120 wl_128 vdd gnd cell_6t
Xbit_r129_c120 bl_120 br_120 wl_129 vdd gnd cell_6t
Xbit_r130_c120 bl_120 br_120 wl_130 vdd gnd cell_6t
Xbit_r131_c120 bl_120 br_120 wl_131 vdd gnd cell_6t
Xbit_r132_c120 bl_120 br_120 wl_132 vdd gnd cell_6t
Xbit_r133_c120 bl_120 br_120 wl_133 vdd gnd cell_6t
Xbit_r134_c120 bl_120 br_120 wl_134 vdd gnd cell_6t
Xbit_r135_c120 bl_120 br_120 wl_135 vdd gnd cell_6t
Xbit_r136_c120 bl_120 br_120 wl_136 vdd gnd cell_6t
Xbit_r137_c120 bl_120 br_120 wl_137 vdd gnd cell_6t
Xbit_r138_c120 bl_120 br_120 wl_138 vdd gnd cell_6t
Xbit_r139_c120 bl_120 br_120 wl_139 vdd gnd cell_6t
Xbit_r140_c120 bl_120 br_120 wl_140 vdd gnd cell_6t
Xbit_r141_c120 bl_120 br_120 wl_141 vdd gnd cell_6t
Xbit_r142_c120 bl_120 br_120 wl_142 vdd gnd cell_6t
Xbit_r143_c120 bl_120 br_120 wl_143 vdd gnd cell_6t
Xbit_r144_c120 bl_120 br_120 wl_144 vdd gnd cell_6t
Xbit_r145_c120 bl_120 br_120 wl_145 vdd gnd cell_6t
Xbit_r146_c120 bl_120 br_120 wl_146 vdd gnd cell_6t
Xbit_r147_c120 bl_120 br_120 wl_147 vdd gnd cell_6t
Xbit_r148_c120 bl_120 br_120 wl_148 vdd gnd cell_6t
Xbit_r149_c120 bl_120 br_120 wl_149 vdd gnd cell_6t
Xbit_r150_c120 bl_120 br_120 wl_150 vdd gnd cell_6t
Xbit_r151_c120 bl_120 br_120 wl_151 vdd gnd cell_6t
Xbit_r152_c120 bl_120 br_120 wl_152 vdd gnd cell_6t
Xbit_r153_c120 bl_120 br_120 wl_153 vdd gnd cell_6t
Xbit_r154_c120 bl_120 br_120 wl_154 vdd gnd cell_6t
Xbit_r155_c120 bl_120 br_120 wl_155 vdd gnd cell_6t
Xbit_r156_c120 bl_120 br_120 wl_156 vdd gnd cell_6t
Xbit_r157_c120 bl_120 br_120 wl_157 vdd gnd cell_6t
Xbit_r158_c120 bl_120 br_120 wl_158 vdd gnd cell_6t
Xbit_r159_c120 bl_120 br_120 wl_159 vdd gnd cell_6t
Xbit_r160_c120 bl_120 br_120 wl_160 vdd gnd cell_6t
Xbit_r161_c120 bl_120 br_120 wl_161 vdd gnd cell_6t
Xbit_r162_c120 bl_120 br_120 wl_162 vdd gnd cell_6t
Xbit_r163_c120 bl_120 br_120 wl_163 vdd gnd cell_6t
Xbit_r164_c120 bl_120 br_120 wl_164 vdd gnd cell_6t
Xbit_r165_c120 bl_120 br_120 wl_165 vdd gnd cell_6t
Xbit_r166_c120 bl_120 br_120 wl_166 vdd gnd cell_6t
Xbit_r167_c120 bl_120 br_120 wl_167 vdd gnd cell_6t
Xbit_r168_c120 bl_120 br_120 wl_168 vdd gnd cell_6t
Xbit_r169_c120 bl_120 br_120 wl_169 vdd gnd cell_6t
Xbit_r170_c120 bl_120 br_120 wl_170 vdd gnd cell_6t
Xbit_r171_c120 bl_120 br_120 wl_171 vdd gnd cell_6t
Xbit_r172_c120 bl_120 br_120 wl_172 vdd gnd cell_6t
Xbit_r173_c120 bl_120 br_120 wl_173 vdd gnd cell_6t
Xbit_r174_c120 bl_120 br_120 wl_174 vdd gnd cell_6t
Xbit_r175_c120 bl_120 br_120 wl_175 vdd gnd cell_6t
Xbit_r176_c120 bl_120 br_120 wl_176 vdd gnd cell_6t
Xbit_r177_c120 bl_120 br_120 wl_177 vdd gnd cell_6t
Xbit_r178_c120 bl_120 br_120 wl_178 vdd gnd cell_6t
Xbit_r179_c120 bl_120 br_120 wl_179 vdd gnd cell_6t
Xbit_r180_c120 bl_120 br_120 wl_180 vdd gnd cell_6t
Xbit_r181_c120 bl_120 br_120 wl_181 vdd gnd cell_6t
Xbit_r182_c120 bl_120 br_120 wl_182 vdd gnd cell_6t
Xbit_r183_c120 bl_120 br_120 wl_183 vdd gnd cell_6t
Xbit_r184_c120 bl_120 br_120 wl_184 vdd gnd cell_6t
Xbit_r185_c120 bl_120 br_120 wl_185 vdd gnd cell_6t
Xbit_r186_c120 bl_120 br_120 wl_186 vdd gnd cell_6t
Xbit_r187_c120 bl_120 br_120 wl_187 vdd gnd cell_6t
Xbit_r188_c120 bl_120 br_120 wl_188 vdd gnd cell_6t
Xbit_r189_c120 bl_120 br_120 wl_189 vdd gnd cell_6t
Xbit_r190_c120 bl_120 br_120 wl_190 vdd gnd cell_6t
Xbit_r191_c120 bl_120 br_120 wl_191 vdd gnd cell_6t
Xbit_r192_c120 bl_120 br_120 wl_192 vdd gnd cell_6t
Xbit_r193_c120 bl_120 br_120 wl_193 vdd gnd cell_6t
Xbit_r194_c120 bl_120 br_120 wl_194 vdd gnd cell_6t
Xbit_r195_c120 bl_120 br_120 wl_195 vdd gnd cell_6t
Xbit_r196_c120 bl_120 br_120 wl_196 vdd gnd cell_6t
Xbit_r197_c120 bl_120 br_120 wl_197 vdd gnd cell_6t
Xbit_r198_c120 bl_120 br_120 wl_198 vdd gnd cell_6t
Xbit_r199_c120 bl_120 br_120 wl_199 vdd gnd cell_6t
Xbit_r200_c120 bl_120 br_120 wl_200 vdd gnd cell_6t
Xbit_r201_c120 bl_120 br_120 wl_201 vdd gnd cell_6t
Xbit_r202_c120 bl_120 br_120 wl_202 vdd gnd cell_6t
Xbit_r203_c120 bl_120 br_120 wl_203 vdd gnd cell_6t
Xbit_r204_c120 bl_120 br_120 wl_204 vdd gnd cell_6t
Xbit_r205_c120 bl_120 br_120 wl_205 vdd gnd cell_6t
Xbit_r206_c120 bl_120 br_120 wl_206 vdd gnd cell_6t
Xbit_r207_c120 bl_120 br_120 wl_207 vdd gnd cell_6t
Xbit_r208_c120 bl_120 br_120 wl_208 vdd gnd cell_6t
Xbit_r209_c120 bl_120 br_120 wl_209 vdd gnd cell_6t
Xbit_r210_c120 bl_120 br_120 wl_210 vdd gnd cell_6t
Xbit_r211_c120 bl_120 br_120 wl_211 vdd gnd cell_6t
Xbit_r212_c120 bl_120 br_120 wl_212 vdd gnd cell_6t
Xbit_r213_c120 bl_120 br_120 wl_213 vdd gnd cell_6t
Xbit_r214_c120 bl_120 br_120 wl_214 vdd gnd cell_6t
Xbit_r215_c120 bl_120 br_120 wl_215 vdd gnd cell_6t
Xbit_r216_c120 bl_120 br_120 wl_216 vdd gnd cell_6t
Xbit_r217_c120 bl_120 br_120 wl_217 vdd gnd cell_6t
Xbit_r218_c120 bl_120 br_120 wl_218 vdd gnd cell_6t
Xbit_r219_c120 bl_120 br_120 wl_219 vdd gnd cell_6t
Xbit_r220_c120 bl_120 br_120 wl_220 vdd gnd cell_6t
Xbit_r221_c120 bl_120 br_120 wl_221 vdd gnd cell_6t
Xbit_r222_c120 bl_120 br_120 wl_222 vdd gnd cell_6t
Xbit_r223_c120 bl_120 br_120 wl_223 vdd gnd cell_6t
Xbit_r224_c120 bl_120 br_120 wl_224 vdd gnd cell_6t
Xbit_r225_c120 bl_120 br_120 wl_225 vdd gnd cell_6t
Xbit_r226_c120 bl_120 br_120 wl_226 vdd gnd cell_6t
Xbit_r227_c120 bl_120 br_120 wl_227 vdd gnd cell_6t
Xbit_r228_c120 bl_120 br_120 wl_228 vdd gnd cell_6t
Xbit_r229_c120 bl_120 br_120 wl_229 vdd gnd cell_6t
Xbit_r230_c120 bl_120 br_120 wl_230 vdd gnd cell_6t
Xbit_r231_c120 bl_120 br_120 wl_231 vdd gnd cell_6t
Xbit_r232_c120 bl_120 br_120 wl_232 vdd gnd cell_6t
Xbit_r233_c120 bl_120 br_120 wl_233 vdd gnd cell_6t
Xbit_r234_c120 bl_120 br_120 wl_234 vdd gnd cell_6t
Xbit_r235_c120 bl_120 br_120 wl_235 vdd gnd cell_6t
Xbit_r236_c120 bl_120 br_120 wl_236 vdd gnd cell_6t
Xbit_r237_c120 bl_120 br_120 wl_237 vdd gnd cell_6t
Xbit_r238_c120 bl_120 br_120 wl_238 vdd gnd cell_6t
Xbit_r239_c120 bl_120 br_120 wl_239 vdd gnd cell_6t
Xbit_r240_c120 bl_120 br_120 wl_240 vdd gnd cell_6t
Xbit_r241_c120 bl_120 br_120 wl_241 vdd gnd cell_6t
Xbit_r242_c120 bl_120 br_120 wl_242 vdd gnd cell_6t
Xbit_r243_c120 bl_120 br_120 wl_243 vdd gnd cell_6t
Xbit_r244_c120 bl_120 br_120 wl_244 vdd gnd cell_6t
Xbit_r245_c120 bl_120 br_120 wl_245 vdd gnd cell_6t
Xbit_r246_c120 bl_120 br_120 wl_246 vdd gnd cell_6t
Xbit_r247_c120 bl_120 br_120 wl_247 vdd gnd cell_6t
Xbit_r248_c120 bl_120 br_120 wl_248 vdd gnd cell_6t
Xbit_r249_c120 bl_120 br_120 wl_249 vdd gnd cell_6t
Xbit_r250_c120 bl_120 br_120 wl_250 vdd gnd cell_6t
Xbit_r251_c120 bl_120 br_120 wl_251 vdd gnd cell_6t
Xbit_r252_c120 bl_120 br_120 wl_252 vdd gnd cell_6t
Xbit_r253_c120 bl_120 br_120 wl_253 vdd gnd cell_6t
Xbit_r254_c120 bl_120 br_120 wl_254 vdd gnd cell_6t
Xbit_r255_c120 bl_120 br_120 wl_255 vdd gnd cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd cell_6t
Xbit_r1_c121 bl_121 br_121 wl_1 vdd gnd cell_6t
Xbit_r2_c121 bl_121 br_121 wl_2 vdd gnd cell_6t
Xbit_r3_c121 bl_121 br_121 wl_3 vdd gnd cell_6t
Xbit_r4_c121 bl_121 br_121 wl_4 vdd gnd cell_6t
Xbit_r5_c121 bl_121 br_121 wl_5 vdd gnd cell_6t
Xbit_r6_c121 bl_121 br_121 wl_6 vdd gnd cell_6t
Xbit_r7_c121 bl_121 br_121 wl_7 vdd gnd cell_6t
Xbit_r8_c121 bl_121 br_121 wl_8 vdd gnd cell_6t
Xbit_r9_c121 bl_121 br_121 wl_9 vdd gnd cell_6t
Xbit_r10_c121 bl_121 br_121 wl_10 vdd gnd cell_6t
Xbit_r11_c121 bl_121 br_121 wl_11 vdd gnd cell_6t
Xbit_r12_c121 bl_121 br_121 wl_12 vdd gnd cell_6t
Xbit_r13_c121 bl_121 br_121 wl_13 vdd gnd cell_6t
Xbit_r14_c121 bl_121 br_121 wl_14 vdd gnd cell_6t
Xbit_r15_c121 bl_121 br_121 wl_15 vdd gnd cell_6t
Xbit_r16_c121 bl_121 br_121 wl_16 vdd gnd cell_6t
Xbit_r17_c121 bl_121 br_121 wl_17 vdd gnd cell_6t
Xbit_r18_c121 bl_121 br_121 wl_18 vdd gnd cell_6t
Xbit_r19_c121 bl_121 br_121 wl_19 vdd gnd cell_6t
Xbit_r20_c121 bl_121 br_121 wl_20 vdd gnd cell_6t
Xbit_r21_c121 bl_121 br_121 wl_21 vdd gnd cell_6t
Xbit_r22_c121 bl_121 br_121 wl_22 vdd gnd cell_6t
Xbit_r23_c121 bl_121 br_121 wl_23 vdd gnd cell_6t
Xbit_r24_c121 bl_121 br_121 wl_24 vdd gnd cell_6t
Xbit_r25_c121 bl_121 br_121 wl_25 vdd gnd cell_6t
Xbit_r26_c121 bl_121 br_121 wl_26 vdd gnd cell_6t
Xbit_r27_c121 bl_121 br_121 wl_27 vdd gnd cell_6t
Xbit_r28_c121 bl_121 br_121 wl_28 vdd gnd cell_6t
Xbit_r29_c121 bl_121 br_121 wl_29 vdd gnd cell_6t
Xbit_r30_c121 bl_121 br_121 wl_30 vdd gnd cell_6t
Xbit_r31_c121 bl_121 br_121 wl_31 vdd gnd cell_6t
Xbit_r32_c121 bl_121 br_121 wl_32 vdd gnd cell_6t
Xbit_r33_c121 bl_121 br_121 wl_33 vdd gnd cell_6t
Xbit_r34_c121 bl_121 br_121 wl_34 vdd gnd cell_6t
Xbit_r35_c121 bl_121 br_121 wl_35 vdd gnd cell_6t
Xbit_r36_c121 bl_121 br_121 wl_36 vdd gnd cell_6t
Xbit_r37_c121 bl_121 br_121 wl_37 vdd gnd cell_6t
Xbit_r38_c121 bl_121 br_121 wl_38 vdd gnd cell_6t
Xbit_r39_c121 bl_121 br_121 wl_39 vdd gnd cell_6t
Xbit_r40_c121 bl_121 br_121 wl_40 vdd gnd cell_6t
Xbit_r41_c121 bl_121 br_121 wl_41 vdd gnd cell_6t
Xbit_r42_c121 bl_121 br_121 wl_42 vdd gnd cell_6t
Xbit_r43_c121 bl_121 br_121 wl_43 vdd gnd cell_6t
Xbit_r44_c121 bl_121 br_121 wl_44 vdd gnd cell_6t
Xbit_r45_c121 bl_121 br_121 wl_45 vdd gnd cell_6t
Xbit_r46_c121 bl_121 br_121 wl_46 vdd gnd cell_6t
Xbit_r47_c121 bl_121 br_121 wl_47 vdd gnd cell_6t
Xbit_r48_c121 bl_121 br_121 wl_48 vdd gnd cell_6t
Xbit_r49_c121 bl_121 br_121 wl_49 vdd gnd cell_6t
Xbit_r50_c121 bl_121 br_121 wl_50 vdd gnd cell_6t
Xbit_r51_c121 bl_121 br_121 wl_51 vdd gnd cell_6t
Xbit_r52_c121 bl_121 br_121 wl_52 vdd gnd cell_6t
Xbit_r53_c121 bl_121 br_121 wl_53 vdd gnd cell_6t
Xbit_r54_c121 bl_121 br_121 wl_54 vdd gnd cell_6t
Xbit_r55_c121 bl_121 br_121 wl_55 vdd gnd cell_6t
Xbit_r56_c121 bl_121 br_121 wl_56 vdd gnd cell_6t
Xbit_r57_c121 bl_121 br_121 wl_57 vdd gnd cell_6t
Xbit_r58_c121 bl_121 br_121 wl_58 vdd gnd cell_6t
Xbit_r59_c121 bl_121 br_121 wl_59 vdd gnd cell_6t
Xbit_r60_c121 bl_121 br_121 wl_60 vdd gnd cell_6t
Xbit_r61_c121 bl_121 br_121 wl_61 vdd gnd cell_6t
Xbit_r62_c121 bl_121 br_121 wl_62 vdd gnd cell_6t
Xbit_r63_c121 bl_121 br_121 wl_63 vdd gnd cell_6t
Xbit_r64_c121 bl_121 br_121 wl_64 vdd gnd cell_6t
Xbit_r65_c121 bl_121 br_121 wl_65 vdd gnd cell_6t
Xbit_r66_c121 bl_121 br_121 wl_66 vdd gnd cell_6t
Xbit_r67_c121 bl_121 br_121 wl_67 vdd gnd cell_6t
Xbit_r68_c121 bl_121 br_121 wl_68 vdd gnd cell_6t
Xbit_r69_c121 bl_121 br_121 wl_69 vdd gnd cell_6t
Xbit_r70_c121 bl_121 br_121 wl_70 vdd gnd cell_6t
Xbit_r71_c121 bl_121 br_121 wl_71 vdd gnd cell_6t
Xbit_r72_c121 bl_121 br_121 wl_72 vdd gnd cell_6t
Xbit_r73_c121 bl_121 br_121 wl_73 vdd gnd cell_6t
Xbit_r74_c121 bl_121 br_121 wl_74 vdd gnd cell_6t
Xbit_r75_c121 bl_121 br_121 wl_75 vdd gnd cell_6t
Xbit_r76_c121 bl_121 br_121 wl_76 vdd gnd cell_6t
Xbit_r77_c121 bl_121 br_121 wl_77 vdd gnd cell_6t
Xbit_r78_c121 bl_121 br_121 wl_78 vdd gnd cell_6t
Xbit_r79_c121 bl_121 br_121 wl_79 vdd gnd cell_6t
Xbit_r80_c121 bl_121 br_121 wl_80 vdd gnd cell_6t
Xbit_r81_c121 bl_121 br_121 wl_81 vdd gnd cell_6t
Xbit_r82_c121 bl_121 br_121 wl_82 vdd gnd cell_6t
Xbit_r83_c121 bl_121 br_121 wl_83 vdd gnd cell_6t
Xbit_r84_c121 bl_121 br_121 wl_84 vdd gnd cell_6t
Xbit_r85_c121 bl_121 br_121 wl_85 vdd gnd cell_6t
Xbit_r86_c121 bl_121 br_121 wl_86 vdd gnd cell_6t
Xbit_r87_c121 bl_121 br_121 wl_87 vdd gnd cell_6t
Xbit_r88_c121 bl_121 br_121 wl_88 vdd gnd cell_6t
Xbit_r89_c121 bl_121 br_121 wl_89 vdd gnd cell_6t
Xbit_r90_c121 bl_121 br_121 wl_90 vdd gnd cell_6t
Xbit_r91_c121 bl_121 br_121 wl_91 vdd gnd cell_6t
Xbit_r92_c121 bl_121 br_121 wl_92 vdd gnd cell_6t
Xbit_r93_c121 bl_121 br_121 wl_93 vdd gnd cell_6t
Xbit_r94_c121 bl_121 br_121 wl_94 vdd gnd cell_6t
Xbit_r95_c121 bl_121 br_121 wl_95 vdd gnd cell_6t
Xbit_r96_c121 bl_121 br_121 wl_96 vdd gnd cell_6t
Xbit_r97_c121 bl_121 br_121 wl_97 vdd gnd cell_6t
Xbit_r98_c121 bl_121 br_121 wl_98 vdd gnd cell_6t
Xbit_r99_c121 bl_121 br_121 wl_99 vdd gnd cell_6t
Xbit_r100_c121 bl_121 br_121 wl_100 vdd gnd cell_6t
Xbit_r101_c121 bl_121 br_121 wl_101 vdd gnd cell_6t
Xbit_r102_c121 bl_121 br_121 wl_102 vdd gnd cell_6t
Xbit_r103_c121 bl_121 br_121 wl_103 vdd gnd cell_6t
Xbit_r104_c121 bl_121 br_121 wl_104 vdd gnd cell_6t
Xbit_r105_c121 bl_121 br_121 wl_105 vdd gnd cell_6t
Xbit_r106_c121 bl_121 br_121 wl_106 vdd gnd cell_6t
Xbit_r107_c121 bl_121 br_121 wl_107 vdd gnd cell_6t
Xbit_r108_c121 bl_121 br_121 wl_108 vdd gnd cell_6t
Xbit_r109_c121 bl_121 br_121 wl_109 vdd gnd cell_6t
Xbit_r110_c121 bl_121 br_121 wl_110 vdd gnd cell_6t
Xbit_r111_c121 bl_121 br_121 wl_111 vdd gnd cell_6t
Xbit_r112_c121 bl_121 br_121 wl_112 vdd gnd cell_6t
Xbit_r113_c121 bl_121 br_121 wl_113 vdd gnd cell_6t
Xbit_r114_c121 bl_121 br_121 wl_114 vdd gnd cell_6t
Xbit_r115_c121 bl_121 br_121 wl_115 vdd gnd cell_6t
Xbit_r116_c121 bl_121 br_121 wl_116 vdd gnd cell_6t
Xbit_r117_c121 bl_121 br_121 wl_117 vdd gnd cell_6t
Xbit_r118_c121 bl_121 br_121 wl_118 vdd gnd cell_6t
Xbit_r119_c121 bl_121 br_121 wl_119 vdd gnd cell_6t
Xbit_r120_c121 bl_121 br_121 wl_120 vdd gnd cell_6t
Xbit_r121_c121 bl_121 br_121 wl_121 vdd gnd cell_6t
Xbit_r122_c121 bl_121 br_121 wl_122 vdd gnd cell_6t
Xbit_r123_c121 bl_121 br_121 wl_123 vdd gnd cell_6t
Xbit_r124_c121 bl_121 br_121 wl_124 vdd gnd cell_6t
Xbit_r125_c121 bl_121 br_121 wl_125 vdd gnd cell_6t
Xbit_r126_c121 bl_121 br_121 wl_126 vdd gnd cell_6t
Xbit_r127_c121 bl_121 br_121 wl_127 vdd gnd cell_6t
Xbit_r128_c121 bl_121 br_121 wl_128 vdd gnd cell_6t
Xbit_r129_c121 bl_121 br_121 wl_129 vdd gnd cell_6t
Xbit_r130_c121 bl_121 br_121 wl_130 vdd gnd cell_6t
Xbit_r131_c121 bl_121 br_121 wl_131 vdd gnd cell_6t
Xbit_r132_c121 bl_121 br_121 wl_132 vdd gnd cell_6t
Xbit_r133_c121 bl_121 br_121 wl_133 vdd gnd cell_6t
Xbit_r134_c121 bl_121 br_121 wl_134 vdd gnd cell_6t
Xbit_r135_c121 bl_121 br_121 wl_135 vdd gnd cell_6t
Xbit_r136_c121 bl_121 br_121 wl_136 vdd gnd cell_6t
Xbit_r137_c121 bl_121 br_121 wl_137 vdd gnd cell_6t
Xbit_r138_c121 bl_121 br_121 wl_138 vdd gnd cell_6t
Xbit_r139_c121 bl_121 br_121 wl_139 vdd gnd cell_6t
Xbit_r140_c121 bl_121 br_121 wl_140 vdd gnd cell_6t
Xbit_r141_c121 bl_121 br_121 wl_141 vdd gnd cell_6t
Xbit_r142_c121 bl_121 br_121 wl_142 vdd gnd cell_6t
Xbit_r143_c121 bl_121 br_121 wl_143 vdd gnd cell_6t
Xbit_r144_c121 bl_121 br_121 wl_144 vdd gnd cell_6t
Xbit_r145_c121 bl_121 br_121 wl_145 vdd gnd cell_6t
Xbit_r146_c121 bl_121 br_121 wl_146 vdd gnd cell_6t
Xbit_r147_c121 bl_121 br_121 wl_147 vdd gnd cell_6t
Xbit_r148_c121 bl_121 br_121 wl_148 vdd gnd cell_6t
Xbit_r149_c121 bl_121 br_121 wl_149 vdd gnd cell_6t
Xbit_r150_c121 bl_121 br_121 wl_150 vdd gnd cell_6t
Xbit_r151_c121 bl_121 br_121 wl_151 vdd gnd cell_6t
Xbit_r152_c121 bl_121 br_121 wl_152 vdd gnd cell_6t
Xbit_r153_c121 bl_121 br_121 wl_153 vdd gnd cell_6t
Xbit_r154_c121 bl_121 br_121 wl_154 vdd gnd cell_6t
Xbit_r155_c121 bl_121 br_121 wl_155 vdd gnd cell_6t
Xbit_r156_c121 bl_121 br_121 wl_156 vdd gnd cell_6t
Xbit_r157_c121 bl_121 br_121 wl_157 vdd gnd cell_6t
Xbit_r158_c121 bl_121 br_121 wl_158 vdd gnd cell_6t
Xbit_r159_c121 bl_121 br_121 wl_159 vdd gnd cell_6t
Xbit_r160_c121 bl_121 br_121 wl_160 vdd gnd cell_6t
Xbit_r161_c121 bl_121 br_121 wl_161 vdd gnd cell_6t
Xbit_r162_c121 bl_121 br_121 wl_162 vdd gnd cell_6t
Xbit_r163_c121 bl_121 br_121 wl_163 vdd gnd cell_6t
Xbit_r164_c121 bl_121 br_121 wl_164 vdd gnd cell_6t
Xbit_r165_c121 bl_121 br_121 wl_165 vdd gnd cell_6t
Xbit_r166_c121 bl_121 br_121 wl_166 vdd gnd cell_6t
Xbit_r167_c121 bl_121 br_121 wl_167 vdd gnd cell_6t
Xbit_r168_c121 bl_121 br_121 wl_168 vdd gnd cell_6t
Xbit_r169_c121 bl_121 br_121 wl_169 vdd gnd cell_6t
Xbit_r170_c121 bl_121 br_121 wl_170 vdd gnd cell_6t
Xbit_r171_c121 bl_121 br_121 wl_171 vdd gnd cell_6t
Xbit_r172_c121 bl_121 br_121 wl_172 vdd gnd cell_6t
Xbit_r173_c121 bl_121 br_121 wl_173 vdd gnd cell_6t
Xbit_r174_c121 bl_121 br_121 wl_174 vdd gnd cell_6t
Xbit_r175_c121 bl_121 br_121 wl_175 vdd gnd cell_6t
Xbit_r176_c121 bl_121 br_121 wl_176 vdd gnd cell_6t
Xbit_r177_c121 bl_121 br_121 wl_177 vdd gnd cell_6t
Xbit_r178_c121 bl_121 br_121 wl_178 vdd gnd cell_6t
Xbit_r179_c121 bl_121 br_121 wl_179 vdd gnd cell_6t
Xbit_r180_c121 bl_121 br_121 wl_180 vdd gnd cell_6t
Xbit_r181_c121 bl_121 br_121 wl_181 vdd gnd cell_6t
Xbit_r182_c121 bl_121 br_121 wl_182 vdd gnd cell_6t
Xbit_r183_c121 bl_121 br_121 wl_183 vdd gnd cell_6t
Xbit_r184_c121 bl_121 br_121 wl_184 vdd gnd cell_6t
Xbit_r185_c121 bl_121 br_121 wl_185 vdd gnd cell_6t
Xbit_r186_c121 bl_121 br_121 wl_186 vdd gnd cell_6t
Xbit_r187_c121 bl_121 br_121 wl_187 vdd gnd cell_6t
Xbit_r188_c121 bl_121 br_121 wl_188 vdd gnd cell_6t
Xbit_r189_c121 bl_121 br_121 wl_189 vdd gnd cell_6t
Xbit_r190_c121 bl_121 br_121 wl_190 vdd gnd cell_6t
Xbit_r191_c121 bl_121 br_121 wl_191 vdd gnd cell_6t
Xbit_r192_c121 bl_121 br_121 wl_192 vdd gnd cell_6t
Xbit_r193_c121 bl_121 br_121 wl_193 vdd gnd cell_6t
Xbit_r194_c121 bl_121 br_121 wl_194 vdd gnd cell_6t
Xbit_r195_c121 bl_121 br_121 wl_195 vdd gnd cell_6t
Xbit_r196_c121 bl_121 br_121 wl_196 vdd gnd cell_6t
Xbit_r197_c121 bl_121 br_121 wl_197 vdd gnd cell_6t
Xbit_r198_c121 bl_121 br_121 wl_198 vdd gnd cell_6t
Xbit_r199_c121 bl_121 br_121 wl_199 vdd gnd cell_6t
Xbit_r200_c121 bl_121 br_121 wl_200 vdd gnd cell_6t
Xbit_r201_c121 bl_121 br_121 wl_201 vdd gnd cell_6t
Xbit_r202_c121 bl_121 br_121 wl_202 vdd gnd cell_6t
Xbit_r203_c121 bl_121 br_121 wl_203 vdd gnd cell_6t
Xbit_r204_c121 bl_121 br_121 wl_204 vdd gnd cell_6t
Xbit_r205_c121 bl_121 br_121 wl_205 vdd gnd cell_6t
Xbit_r206_c121 bl_121 br_121 wl_206 vdd gnd cell_6t
Xbit_r207_c121 bl_121 br_121 wl_207 vdd gnd cell_6t
Xbit_r208_c121 bl_121 br_121 wl_208 vdd gnd cell_6t
Xbit_r209_c121 bl_121 br_121 wl_209 vdd gnd cell_6t
Xbit_r210_c121 bl_121 br_121 wl_210 vdd gnd cell_6t
Xbit_r211_c121 bl_121 br_121 wl_211 vdd gnd cell_6t
Xbit_r212_c121 bl_121 br_121 wl_212 vdd gnd cell_6t
Xbit_r213_c121 bl_121 br_121 wl_213 vdd gnd cell_6t
Xbit_r214_c121 bl_121 br_121 wl_214 vdd gnd cell_6t
Xbit_r215_c121 bl_121 br_121 wl_215 vdd gnd cell_6t
Xbit_r216_c121 bl_121 br_121 wl_216 vdd gnd cell_6t
Xbit_r217_c121 bl_121 br_121 wl_217 vdd gnd cell_6t
Xbit_r218_c121 bl_121 br_121 wl_218 vdd gnd cell_6t
Xbit_r219_c121 bl_121 br_121 wl_219 vdd gnd cell_6t
Xbit_r220_c121 bl_121 br_121 wl_220 vdd gnd cell_6t
Xbit_r221_c121 bl_121 br_121 wl_221 vdd gnd cell_6t
Xbit_r222_c121 bl_121 br_121 wl_222 vdd gnd cell_6t
Xbit_r223_c121 bl_121 br_121 wl_223 vdd gnd cell_6t
Xbit_r224_c121 bl_121 br_121 wl_224 vdd gnd cell_6t
Xbit_r225_c121 bl_121 br_121 wl_225 vdd gnd cell_6t
Xbit_r226_c121 bl_121 br_121 wl_226 vdd gnd cell_6t
Xbit_r227_c121 bl_121 br_121 wl_227 vdd gnd cell_6t
Xbit_r228_c121 bl_121 br_121 wl_228 vdd gnd cell_6t
Xbit_r229_c121 bl_121 br_121 wl_229 vdd gnd cell_6t
Xbit_r230_c121 bl_121 br_121 wl_230 vdd gnd cell_6t
Xbit_r231_c121 bl_121 br_121 wl_231 vdd gnd cell_6t
Xbit_r232_c121 bl_121 br_121 wl_232 vdd gnd cell_6t
Xbit_r233_c121 bl_121 br_121 wl_233 vdd gnd cell_6t
Xbit_r234_c121 bl_121 br_121 wl_234 vdd gnd cell_6t
Xbit_r235_c121 bl_121 br_121 wl_235 vdd gnd cell_6t
Xbit_r236_c121 bl_121 br_121 wl_236 vdd gnd cell_6t
Xbit_r237_c121 bl_121 br_121 wl_237 vdd gnd cell_6t
Xbit_r238_c121 bl_121 br_121 wl_238 vdd gnd cell_6t
Xbit_r239_c121 bl_121 br_121 wl_239 vdd gnd cell_6t
Xbit_r240_c121 bl_121 br_121 wl_240 vdd gnd cell_6t
Xbit_r241_c121 bl_121 br_121 wl_241 vdd gnd cell_6t
Xbit_r242_c121 bl_121 br_121 wl_242 vdd gnd cell_6t
Xbit_r243_c121 bl_121 br_121 wl_243 vdd gnd cell_6t
Xbit_r244_c121 bl_121 br_121 wl_244 vdd gnd cell_6t
Xbit_r245_c121 bl_121 br_121 wl_245 vdd gnd cell_6t
Xbit_r246_c121 bl_121 br_121 wl_246 vdd gnd cell_6t
Xbit_r247_c121 bl_121 br_121 wl_247 vdd gnd cell_6t
Xbit_r248_c121 bl_121 br_121 wl_248 vdd gnd cell_6t
Xbit_r249_c121 bl_121 br_121 wl_249 vdd gnd cell_6t
Xbit_r250_c121 bl_121 br_121 wl_250 vdd gnd cell_6t
Xbit_r251_c121 bl_121 br_121 wl_251 vdd gnd cell_6t
Xbit_r252_c121 bl_121 br_121 wl_252 vdd gnd cell_6t
Xbit_r253_c121 bl_121 br_121 wl_253 vdd gnd cell_6t
Xbit_r254_c121 bl_121 br_121 wl_254 vdd gnd cell_6t
Xbit_r255_c121 bl_121 br_121 wl_255 vdd gnd cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd cell_6t
Xbit_r1_c122 bl_122 br_122 wl_1 vdd gnd cell_6t
Xbit_r2_c122 bl_122 br_122 wl_2 vdd gnd cell_6t
Xbit_r3_c122 bl_122 br_122 wl_3 vdd gnd cell_6t
Xbit_r4_c122 bl_122 br_122 wl_4 vdd gnd cell_6t
Xbit_r5_c122 bl_122 br_122 wl_5 vdd gnd cell_6t
Xbit_r6_c122 bl_122 br_122 wl_6 vdd gnd cell_6t
Xbit_r7_c122 bl_122 br_122 wl_7 vdd gnd cell_6t
Xbit_r8_c122 bl_122 br_122 wl_8 vdd gnd cell_6t
Xbit_r9_c122 bl_122 br_122 wl_9 vdd gnd cell_6t
Xbit_r10_c122 bl_122 br_122 wl_10 vdd gnd cell_6t
Xbit_r11_c122 bl_122 br_122 wl_11 vdd gnd cell_6t
Xbit_r12_c122 bl_122 br_122 wl_12 vdd gnd cell_6t
Xbit_r13_c122 bl_122 br_122 wl_13 vdd gnd cell_6t
Xbit_r14_c122 bl_122 br_122 wl_14 vdd gnd cell_6t
Xbit_r15_c122 bl_122 br_122 wl_15 vdd gnd cell_6t
Xbit_r16_c122 bl_122 br_122 wl_16 vdd gnd cell_6t
Xbit_r17_c122 bl_122 br_122 wl_17 vdd gnd cell_6t
Xbit_r18_c122 bl_122 br_122 wl_18 vdd gnd cell_6t
Xbit_r19_c122 bl_122 br_122 wl_19 vdd gnd cell_6t
Xbit_r20_c122 bl_122 br_122 wl_20 vdd gnd cell_6t
Xbit_r21_c122 bl_122 br_122 wl_21 vdd gnd cell_6t
Xbit_r22_c122 bl_122 br_122 wl_22 vdd gnd cell_6t
Xbit_r23_c122 bl_122 br_122 wl_23 vdd gnd cell_6t
Xbit_r24_c122 bl_122 br_122 wl_24 vdd gnd cell_6t
Xbit_r25_c122 bl_122 br_122 wl_25 vdd gnd cell_6t
Xbit_r26_c122 bl_122 br_122 wl_26 vdd gnd cell_6t
Xbit_r27_c122 bl_122 br_122 wl_27 vdd gnd cell_6t
Xbit_r28_c122 bl_122 br_122 wl_28 vdd gnd cell_6t
Xbit_r29_c122 bl_122 br_122 wl_29 vdd gnd cell_6t
Xbit_r30_c122 bl_122 br_122 wl_30 vdd gnd cell_6t
Xbit_r31_c122 bl_122 br_122 wl_31 vdd gnd cell_6t
Xbit_r32_c122 bl_122 br_122 wl_32 vdd gnd cell_6t
Xbit_r33_c122 bl_122 br_122 wl_33 vdd gnd cell_6t
Xbit_r34_c122 bl_122 br_122 wl_34 vdd gnd cell_6t
Xbit_r35_c122 bl_122 br_122 wl_35 vdd gnd cell_6t
Xbit_r36_c122 bl_122 br_122 wl_36 vdd gnd cell_6t
Xbit_r37_c122 bl_122 br_122 wl_37 vdd gnd cell_6t
Xbit_r38_c122 bl_122 br_122 wl_38 vdd gnd cell_6t
Xbit_r39_c122 bl_122 br_122 wl_39 vdd gnd cell_6t
Xbit_r40_c122 bl_122 br_122 wl_40 vdd gnd cell_6t
Xbit_r41_c122 bl_122 br_122 wl_41 vdd gnd cell_6t
Xbit_r42_c122 bl_122 br_122 wl_42 vdd gnd cell_6t
Xbit_r43_c122 bl_122 br_122 wl_43 vdd gnd cell_6t
Xbit_r44_c122 bl_122 br_122 wl_44 vdd gnd cell_6t
Xbit_r45_c122 bl_122 br_122 wl_45 vdd gnd cell_6t
Xbit_r46_c122 bl_122 br_122 wl_46 vdd gnd cell_6t
Xbit_r47_c122 bl_122 br_122 wl_47 vdd gnd cell_6t
Xbit_r48_c122 bl_122 br_122 wl_48 vdd gnd cell_6t
Xbit_r49_c122 bl_122 br_122 wl_49 vdd gnd cell_6t
Xbit_r50_c122 bl_122 br_122 wl_50 vdd gnd cell_6t
Xbit_r51_c122 bl_122 br_122 wl_51 vdd gnd cell_6t
Xbit_r52_c122 bl_122 br_122 wl_52 vdd gnd cell_6t
Xbit_r53_c122 bl_122 br_122 wl_53 vdd gnd cell_6t
Xbit_r54_c122 bl_122 br_122 wl_54 vdd gnd cell_6t
Xbit_r55_c122 bl_122 br_122 wl_55 vdd gnd cell_6t
Xbit_r56_c122 bl_122 br_122 wl_56 vdd gnd cell_6t
Xbit_r57_c122 bl_122 br_122 wl_57 vdd gnd cell_6t
Xbit_r58_c122 bl_122 br_122 wl_58 vdd gnd cell_6t
Xbit_r59_c122 bl_122 br_122 wl_59 vdd gnd cell_6t
Xbit_r60_c122 bl_122 br_122 wl_60 vdd gnd cell_6t
Xbit_r61_c122 bl_122 br_122 wl_61 vdd gnd cell_6t
Xbit_r62_c122 bl_122 br_122 wl_62 vdd gnd cell_6t
Xbit_r63_c122 bl_122 br_122 wl_63 vdd gnd cell_6t
Xbit_r64_c122 bl_122 br_122 wl_64 vdd gnd cell_6t
Xbit_r65_c122 bl_122 br_122 wl_65 vdd gnd cell_6t
Xbit_r66_c122 bl_122 br_122 wl_66 vdd gnd cell_6t
Xbit_r67_c122 bl_122 br_122 wl_67 vdd gnd cell_6t
Xbit_r68_c122 bl_122 br_122 wl_68 vdd gnd cell_6t
Xbit_r69_c122 bl_122 br_122 wl_69 vdd gnd cell_6t
Xbit_r70_c122 bl_122 br_122 wl_70 vdd gnd cell_6t
Xbit_r71_c122 bl_122 br_122 wl_71 vdd gnd cell_6t
Xbit_r72_c122 bl_122 br_122 wl_72 vdd gnd cell_6t
Xbit_r73_c122 bl_122 br_122 wl_73 vdd gnd cell_6t
Xbit_r74_c122 bl_122 br_122 wl_74 vdd gnd cell_6t
Xbit_r75_c122 bl_122 br_122 wl_75 vdd gnd cell_6t
Xbit_r76_c122 bl_122 br_122 wl_76 vdd gnd cell_6t
Xbit_r77_c122 bl_122 br_122 wl_77 vdd gnd cell_6t
Xbit_r78_c122 bl_122 br_122 wl_78 vdd gnd cell_6t
Xbit_r79_c122 bl_122 br_122 wl_79 vdd gnd cell_6t
Xbit_r80_c122 bl_122 br_122 wl_80 vdd gnd cell_6t
Xbit_r81_c122 bl_122 br_122 wl_81 vdd gnd cell_6t
Xbit_r82_c122 bl_122 br_122 wl_82 vdd gnd cell_6t
Xbit_r83_c122 bl_122 br_122 wl_83 vdd gnd cell_6t
Xbit_r84_c122 bl_122 br_122 wl_84 vdd gnd cell_6t
Xbit_r85_c122 bl_122 br_122 wl_85 vdd gnd cell_6t
Xbit_r86_c122 bl_122 br_122 wl_86 vdd gnd cell_6t
Xbit_r87_c122 bl_122 br_122 wl_87 vdd gnd cell_6t
Xbit_r88_c122 bl_122 br_122 wl_88 vdd gnd cell_6t
Xbit_r89_c122 bl_122 br_122 wl_89 vdd gnd cell_6t
Xbit_r90_c122 bl_122 br_122 wl_90 vdd gnd cell_6t
Xbit_r91_c122 bl_122 br_122 wl_91 vdd gnd cell_6t
Xbit_r92_c122 bl_122 br_122 wl_92 vdd gnd cell_6t
Xbit_r93_c122 bl_122 br_122 wl_93 vdd gnd cell_6t
Xbit_r94_c122 bl_122 br_122 wl_94 vdd gnd cell_6t
Xbit_r95_c122 bl_122 br_122 wl_95 vdd gnd cell_6t
Xbit_r96_c122 bl_122 br_122 wl_96 vdd gnd cell_6t
Xbit_r97_c122 bl_122 br_122 wl_97 vdd gnd cell_6t
Xbit_r98_c122 bl_122 br_122 wl_98 vdd gnd cell_6t
Xbit_r99_c122 bl_122 br_122 wl_99 vdd gnd cell_6t
Xbit_r100_c122 bl_122 br_122 wl_100 vdd gnd cell_6t
Xbit_r101_c122 bl_122 br_122 wl_101 vdd gnd cell_6t
Xbit_r102_c122 bl_122 br_122 wl_102 vdd gnd cell_6t
Xbit_r103_c122 bl_122 br_122 wl_103 vdd gnd cell_6t
Xbit_r104_c122 bl_122 br_122 wl_104 vdd gnd cell_6t
Xbit_r105_c122 bl_122 br_122 wl_105 vdd gnd cell_6t
Xbit_r106_c122 bl_122 br_122 wl_106 vdd gnd cell_6t
Xbit_r107_c122 bl_122 br_122 wl_107 vdd gnd cell_6t
Xbit_r108_c122 bl_122 br_122 wl_108 vdd gnd cell_6t
Xbit_r109_c122 bl_122 br_122 wl_109 vdd gnd cell_6t
Xbit_r110_c122 bl_122 br_122 wl_110 vdd gnd cell_6t
Xbit_r111_c122 bl_122 br_122 wl_111 vdd gnd cell_6t
Xbit_r112_c122 bl_122 br_122 wl_112 vdd gnd cell_6t
Xbit_r113_c122 bl_122 br_122 wl_113 vdd gnd cell_6t
Xbit_r114_c122 bl_122 br_122 wl_114 vdd gnd cell_6t
Xbit_r115_c122 bl_122 br_122 wl_115 vdd gnd cell_6t
Xbit_r116_c122 bl_122 br_122 wl_116 vdd gnd cell_6t
Xbit_r117_c122 bl_122 br_122 wl_117 vdd gnd cell_6t
Xbit_r118_c122 bl_122 br_122 wl_118 vdd gnd cell_6t
Xbit_r119_c122 bl_122 br_122 wl_119 vdd gnd cell_6t
Xbit_r120_c122 bl_122 br_122 wl_120 vdd gnd cell_6t
Xbit_r121_c122 bl_122 br_122 wl_121 vdd gnd cell_6t
Xbit_r122_c122 bl_122 br_122 wl_122 vdd gnd cell_6t
Xbit_r123_c122 bl_122 br_122 wl_123 vdd gnd cell_6t
Xbit_r124_c122 bl_122 br_122 wl_124 vdd gnd cell_6t
Xbit_r125_c122 bl_122 br_122 wl_125 vdd gnd cell_6t
Xbit_r126_c122 bl_122 br_122 wl_126 vdd gnd cell_6t
Xbit_r127_c122 bl_122 br_122 wl_127 vdd gnd cell_6t
Xbit_r128_c122 bl_122 br_122 wl_128 vdd gnd cell_6t
Xbit_r129_c122 bl_122 br_122 wl_129 vdd gnd cell_6t
Xbit_r130_c122 bl_122 br_122 wl_130 vdd gnd cell_6t
Xbit_r131_c122 bl_122 br_122 wl_131 vdd gnd cell_6t
Xbit_r132_c122 bl_122 br_122 wl_132 vdd gnd cell_6t
Xbit_r133_c122 bl_122 br_122 wl_133 vdd gnd cell_6t
Xbit_r134_c122 bl_122 br_122 wl_134 vdd gnd cell_6t
Xbit_r135_c122 bl_122 br_122 wl_135 vdd gnd cell_6t
Xbit_r136_c122 bl_122 br_122 wl_136 vdd gnd cell_6t
Xbit_r137_c122 bl_122 br_122 wl_137 vdd gnd cell_6t
Xbit_r138_c122 bl_122 br_122 wl_138 vdd gnd cell_6t
Xbit_r139_c122 bl_122 br_122 wl_139 vdd gnd cell_6t
Xbit_r140_c122 bl_122 br_122 wl_140 vdd gnd cell_6t
Xbit_r141_c122 bl_122 br_122 wl_141 vdd gnd cell_6t
Xbit_r142_c122 bl_122 br_122 wl_142 vdd gnd cell_6t
Xbit_r143_c122 bl_122 br_122 wl_143 vdd gnd cell_6t
Xbit_r144_c122 bl_122 br_122 wl_144 vdd gnd cell_6t
Xbit_r145_c122 bl_122 br_122 wl_145 vdd gnd cell_6t
Xbit_r146_c122 bl_122 br_122 wl_146 vdd gnd cell_6t
Xbit_r147_c122 bl_122 br_122 wl_147 vdd gnd cell_6t
Xbit_r148_c122 bl_122 br_122 wl_148 vdd gnd cell_6t
Xbit_r149_c122 bl_122 br_122 wl_149 vdd gnd cell_6t
Xbit_r150_c122 bl_122 br_122 wl_150 vdd gnd cell_6t
Xbit_r151_c122 bl_122 br_122 wl_151 vdd gnd cell_6t
Xbit_r152_c122 bl_122 br_122 wl_152 vdd gnd cell_6t
Xbit_r153_c122 bl_122 br_122 wl_153 vdd gnd cell_6t
Xbit_r154_c122 bl_122 br_122 wl_154 vdd gnd cell_6t
Xbit_r155_c122 bl_122 br_122 wl_155 vdd gnd cell_6t
Xbit_r156_c122 bl_122 br_122 wl_156 vdd gnd cell_6t
Xbit_r157_c122 bl_122 br_122 wl_157 vdd gnd cell_6t
Xbit_r158_c122 bl_122 br_122 wl_158 vdd gnd cell_6t
Xbit_r159_c122 bl_122 br_122 wl_159 vdd gnd cell_6t
Xbit_r160_c122 bl_122 br_122 wl_160 vdd gnd cell_6t
Xbit_r161_c122 bl_122 br_122 wl_161 vdd gnd cell_6t
Xbit_r162_c122 bl_122 br_122 wl_162 vdd gnd cell_6t
Xbit_r163_c122 bl_122 br_122 wl_163 vdd gnd cell_6t
Xbit_r164_c122 bl_122 br_122 wl_164 vdd gnd cell_6t
Xbit_r165_c122 bl_122 br_122 wl_165 vdd gnd cell_6t
Xbit_r166_c122 bl_122 br_122 wl_166 vdd gnd cell_6t
Xbit_r167_c122 bl_122 br_122 wl_167 vdd gnd cell_6t
Xbit_r168_c122 bl_122 br_122 wl_168 vdd gnd cell_6t
Xbit_r169_c122 bl_122 br_122 wl_169 vdd gnd cell_6t
Xbit_r170_c122 bl_122 br_122 wl_170 vdd gnd cell_6t
Xbit_r171_c122 bl_122 br_122 wl_171 vdd gnd cell_6t
Xbit_r172_c122 bl_122 br_122 wl_172 vdd gnd cell_6t
Xbit_r173_c122 bl_122 br_122 wl_173 vdd gnd cell_6t
Xbit_r174_c122 bl_122 br_122 wl_174 vdd gnd cell_6t
Xbit_r175_c122 bl_122 br_122 wl_175 vdd gnd cell_6t
Xbit_r176_c122 bl_122 br_122 wl_176 vdd gnd cell_6t
Xbit_r177_c122 bl_122 br_122 wl_177 vdd gnd cell_6t
Xbit_r178_c122 bl_122 br_122 wl_178 vdd gnd cell_6t
Xbit_r179_c122 bl_122 br_122 wl_179 vdd gnd cell_6t
Xbit_r180_c122 bl_122 br_122 wl_180 vdd gnd cell_6t
Xbit_r181_c122 bl_122 br_122 wl_181 vdd gnd cell_6t
Xbit_r182_c122 bl_122 br_122 wl_182 vdd gnd cell_6t
Xbit_r183_c122 bl_122 br_122 wl_183 vdd gnd cell_6t
Xbit_r184_c122 bl_122 br_122 wl_184 vdd gnd cell_6t
Xbit_r185_c122 bl_122 br_122 wl_185 vdd gnd cell_6t
Xbit_r186_c122 bl_122 br_122 wl_186 vdd gnd cell_6t
Xbit_r187_c122 bl_122 br_122 wl_187 vdd gnd cell_6t
Xbit_r188_c122 bl_122 br_122 wl_188 vdd gnd cell_6t
Xbit_r189_c122 bl_122 br_122 wl_189 vdd gnd cell_6t
Xbit_r190_c122 bl_122 br_122 wl_190 vdd gnd cell_6t
Xbit_r191_c122 bl_122 br_122 wl_191 vdd gnd cell_6t
Xbit_r192_c122 bl_122 br_122 wl_192 vdd gnd cell_6t
Xbit_r193_c122 bl_122 br_122 wl_193 vdd gnd cell_6t
Xbit_r194_c122 bl_122 br_122 wl_194 vdd gnd cell_6t
Xbit_r195_c122 bl_122 br_122 wl_195 vdd gnd cell_6t
Xbit_r196_c122 bl_122 br_122 wl_196 vdd gnd cell_6t
Xbit_r197_c122 bl_122 br_122 wl_197 vdd gnd cell_6t
Xbit_r198_c122 bl_122 br_122 wl_198 vdd gnd cell_6t
Xbit_r199_c122 bl_122 br_122 wl_199 vdd gnd cell_6t
Xbit_r200_c122 bl_122 br_122 wl_200 vdd gnd cell_6t
Xbit_r201_c122 bl_122 br_122 wl_201 vdd gnd cell_6t
Xbit_r202_c122 bl_122 br_122 wl_202 vdd gnd cell_6t
Xbit_r203_c122 bl_122 br_122 wl_203 vdd gnd cell_6t
Xbit_r204_c122 bl_122 br_122 wl_204 vdd gnd cell_6t
Xbit_r205_c122 bl_122 br_122 wl_205 vdd gnd cell_6t
Xbit_r206_c122 bl_122 br_122 wl_206 vdd gnd cell_6t
Xbit_r207_c122 bl_122 br_122 wl_207 vdd gnd cell_6t
Xbit_r208_c122 bl_122 br_122 wl_208 vdd gnd cell_6t
Xbit_r209_c122 bl_122 br_122 wl_209 vdd gnd cell_6t
Xbit_r210_c122 bl_122 br_122 wl_210 vdd gnd cell_6t
Xbit_r211_c122 bl_122 br_122 wl_211 vdd gnd cell_6t
Xbit_r212_c122 bl_122 br_122 wl_212 vdd gnd cell_6t
Xbit_r213_c122 bl_122 br_122 wl_213 vdd gnd cell_6t
Xbit_r214_c122 bl_122 br_122 wl_214 vdd gnd cell_6t
Xbit_r215_c122 bl_122 br_122 wl_215 vdd gnd cell_6t
Xbit_r216_c122 bl_122 br_122 wl_216 vdd gnd cell_6t
Xbit_r217_c122 bl_122 br_122 wl_217 vdd gnd cell_6t
Xbit_r218_c122 bl_122 br_122 wl_218 vdd gnd cell_6t
Xbit_r219_c122 bl_122 br_122 wl_219 vdd gnd cell_6t
Xbit_r220_c122 bl_122 br_122 wl_220 vdd gnd cell_6t
Xbit_r221_c122 bl_122 br_122 wl_221 vdd gnd cell_6t
Xbit_r222_c122 bl_122 br_122 wl_222 vdd gnd cell_6t
Xbit_r223_c122 bl_122 br_122 wl_223 vdd gnd cell_6t
Xbit_r224_c122 bl_122 br_122 wl_224 vdd gnd cell_6t
Xbit_r225_c122 bl_122 br_122 wl_225 vdd gnd cell_6t
Xbit_r226_c122 bl_122 br_122 wl_226 vdd gnd cell_6t
Xbit_r227_c122 bl_122 br_122 wl_227 vdd gnd cell_6t
Xbit_r228_c122 bl_122 br_122 wl_228 vdd gnd cell_6t
Xbit_r229_c122 bl_122 br_122 wl_229 vdd gnd cell_6t
Xbit_r230_c122 bl_122 br_122 wl_230 vdd gnd cell_6t
Xbit_r231_c122 bl_122 br_122 wl_231 vdd gnd cell_6t
Xbit_r232_c122 bl_122 br_122 wl_232 vdd gnd cell_6t
Xbit_r233_c122 bl_122 br_122 wl_233 vdd gnd cell_6t
Xbit_r234_c122 bl_122 br_122 wl_234 vdd gnd cell_6t
Xbit_r235_c122 bl_122 br_122 wl_235 vdd gnd cell_6t
Xbit_r236_c122 bl_122 br_122 wl_236 vdd gnd cell_6t
Xbit_r237_c122 bl_122 br_122 wl_237 vdd gnd cell_6t
Xbit_r238_c122 bl_122 br_122 wl_238 vdd gnd cell_6t
Xbit_r239_c122 bl_122 br_122 wl_239 vdd gnd cell_6t
Xbit_r240_c122 bl_122 br_122 wl_240 vdd gnd cell_6t
Xbit_r241_c122 bl_122 br_122 wl_241 vdd gnd cell_6t
Xbit_r242_c122 bl_122 br_122 wl_242 vdd gnd cell_6t
Xbit_r243_c122 bl_122 br_122 wl_243 vdd gnd cell_6t
Xbit_r244_c122 bl_122 br_122 wl_244 vdd gnd cell_6t
Xbit_r245_c122 bl_122 br_122 wl_245 vdd gnd cell_6t
Xbit_r246_c122 bl_122 br_122 wl_246 vdd gnd cell_6t
Xbit_r247_c122 bl_122 br_122 wl_247 vdd gnd cell_6t
Xbit_r248_c122 bl_122 br_122 wl_248 vdd gnd cell_6t
Xbit_r249_c122 bl_122 br_122 wl_249 vdd gnd cell_6t
Xbit_r250_c122 bl_122 br_122 wl_250 vdd gnd cell_6t
Xbit_r251_c122 bl_122 br_122 wl_251 vdd gnd cell_6t
Xbit_r252_c122 bl_122 br_122 wl_252 vdd gnd cell_6t
Xbit_r253_c122 bl_122 br_122 wl_253 vdd gnd cell_6t
Xbit_r254_c122 bl_122 br_122 wl_254 vdd gnd cell_6t
Xbit_r255_c122 bl_122 br_122 wl_255 vdd gnd cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd cell_6t
Xbit_r1_c123 bl_123 br_123 wl_1 vdd gnd cell_6t
Xbit_r2_c123 bl_123 br_123 wl_2 vdd gnd cell_6t
Xbit_r3_c123 bl_123 br_123 wl_3 vdd gnd cell_6t
Xbit_r4_c123 bl_123 br_123 wl_4 vdd gnd cell_6t
Xbit_r5_c123 bl_123 br_123 wl_5 vdd gnd cell_6t
Xbit_r6_c123 bl_123 br_123 wl_6 vdd gnd cell_6t
Xbit_r7_c123 bl_123 br_123 wl_7 vdd gnd cell_6t
Xbit_r8_c123 bl_123 br_123 wl_8 vdd gnd cell_6t
Xbit_r9_c123 bl_123 br_123 wl_9 vdd gnd cell_6t
Xbit_r10_c123 bl_123 br_123 wl_10 vdd gnd cell_6t
Xbit_r11_c123 bl_123 br_123 wl_11 vdd gnd cell_6t
Xbit_r12_c123 bl_123 br_123 wl_12 vdd gnd cell_6t
Xbit_r13_c123 bl_123 br_123 wl_13 vdd gnd cell_6t
Xbit_r14_c123 bl_123 br_123 wl_14 vdd gnd cell_6t
Xbit_r15_c123 bl_123 br_123 wl_15 vdd gnd cell_6t
Xbit_r16_c123 bl_123 br_123 wl_16 vdd gnd cell_6t
Xbit_r17_c123 bl_123 br_123 wl_17 vdd gnd cell_6t
Xbit_r18_c123 bl_123 br_123 wl_18 vdd gnd cell_6t
Xbit_r19_c123 bl_123 br_123 wl_19 vdd gnd cell_6t
Xbit_r20_c123 bl_123 br_123 wl_20 vdd gnd cell_6t
Xbit_r21_c123 bl_123 br_123 wl_21 vdd gnd cell_6t
Xbit_r22_c123 bl_123 br_123 wl_22 vdd gnd cell_6t
Xbit_r23_c123 bl_123 br_123 wl_23 vdd gnd cell_6t
Xbit_r24_c123 bl_123 br_123 wl_24 vdd gnd cell_6t
Xbit_r25_c123 bl_123 br_123 wl_25 vdd gnd cell_6t
Xbit_r26_c123 bl_123 br_123 wl_26 vdd gnd cell_6t
Xbit_r27_c123 bl_123 br_123 wl_27 vdd gnd cell_6t
Xbit_r28_c123 bl_123 br_123 wl_28 vdd gnd cell_6t
Xbit_r29_c123 bl_123 br_123 wl_29 vdd gnd cell_6t
Xbit_r30_c123 bl_123 br_123 wl_30 vdd gnd cell_6t
Xbit_r31_c123 bl_123 br_123 wl_31 vdd gnd cell_6t
Xbit_r32_c123 bl_123 br_123 wl_32 vdd gnd cell_6t
Xbit_r33_c123 bl_123 br_123 wl_33 vdd gnd cell_6t
Xbit_r34_c123 bl_123 br_123 wl_34 vdd gnd cell_6t
Xbit_r35_c123 bl_123 br_123 wl_35 vdd gnd cell_6t
Xbit_r36_c123 bl_123 br_123 wl_36 vdd gnd cell_6t
Xbit_r37_c123 bl_123 br_123 wl_37 vdd gnd cell_6t
Xbit_r38_c123 bl_123 br_123 wl_38 vdd gnd cell_6t
Xbit_r39_c123 bl_123 br_123 wl_39 vdd gnd cell_6t
Xbit_r40_c123 bl_123 br_123 wl_40 vdd gnd cell_6t
Xbit_r41_c123 bl_123 br_123 wl_41 vdd gnd cell_6t
Xbit_r42_c123 bl_123 br_123 wl_42 vdd gnd cell_6t
Xbit_r43_c123 bl_123 br_123 wl_43 vdd gnd cell_6t
Xbit_r44_c123 bl_123 br_123 wl_44 vdd gnd cell_6t
Xbit_r45_c123 bl_123 br_123 wl_45 vdd gnd cell_6t
Xbit_r46_c123 bl_123 br_123 wl_46 vdd gnd cell_6t
Xbit_r47_c123 bl_123 br_123 wl_47 vdd gnd cell_6t
Xbit_r48_c123 bl_123 br_123 wl_48 vdd gnd cell_6t
Xbit_r49_c123 bl_123 br_123 wl_49 vdd gnd cell_6t
Xbit_r50_c123 bl_123 br_123 wl_50 vdd gnd cell_6t
Xbit_r51_c123 bl_123 br_123 wl_51 vdd gnd cell_6t
Xbit_r52_c123 bl_123 br_123 wl_52 vdd gnd cell_6t
Xbit_r53_c123 bl_123 br_123 wl_53 vdd gnd cell_6t
Xbit_r54_c123 bl_123 br_123 wl_54 vdd gnd cell_6t
Xbit_r55_c123 bl_123 br_123 wl_55 vdd gnd cell_6t
Xbit_r56_c123 bl_123 br_123 wl_56 vdd gnd cell_6t
Xbit_r57_c123 bl_123 br_123 wl_57 vdd gnd cell_6t
Xbit_r58_c123 bl_123 br_123 wl_58 vdd gnd cell_6t
Xbit_r59_c123 bl_123 br_123 wl_59 vdd gnd cell_6t
Xbit_r60_c123 bl_123 br_123 wl_60 vdd gnd cell_6t
Xbit_r61_c123 bl_123 br_123 wl_61 vdd gnd cell_6t
Xbit_r62_c123 bl_123 br_123 wl_62 vdd gnd cell_6t
Xbit_r63_c123 bl_123 br_123 wl_63 vdd gnd cell_6t
Xbit_r64_c123 bl_123 br_123 wl_64 vdd gnd cell_6t
Xbit_r65_c123 bl_123 br_123 wl_65 vdd gnd cell_6t
Xbit_r66_c123 bl_123 br_123 wl_66 vdd gnd cell_6t
Xbit_r67_c123 bl_123 br_123 wl_67 vdd gnd cell_6t
Xbit_r68_c123 bl_123 br_123 wl_68 vdd gnd cell_6t
Xbit_r69_c123 bl_123 br_123 wl_69 vdd gnd cell_6t
Xbit_r70_c123 bl_123 br_123 wl_70 vdd gnd cell_6t
Xbit_r71_c123 bl_123 br_123 wl_71 vdd gnd cell_6t
Xbit_r72_c123 bl_123 br_123 wl_72 vdd gnd cell_6t
Xbit_r73_c123 bl_123 br_123 wl_73 vdd gnd cell_6t
Xbit_r74_c123 bl_123 br_123 wl_74 vdd gnd cell_6t
Xbit_r75_c123 bl_123 br_123 wl_75 vdd gnd cell_6t
Xbit_r76_c123 bl_123 br_123 wl_76 vdd gnd cell_6t
Xbit_r77_c123 bl_123 br_123 wl_77 vdd gnd cell_6t
Xbit_r78_c123 bl_123 br_123 wl_78 vdd gnd cell_6t
Xbit_r79_c123 bl_123 br_123 wl_79 vdd gnd cell_6t
Xbit_r80_c123 bl_123 br_123 wl_80 vdd gnd cell_6t
Xbit_r81_c123 bl_123 br_123 wl_81 vdd gnd cell_6t
Xbit_r82_c123 bl_123 br_123 wl_82 vdd gnd cell_6t
Xbit_r83_c123 bl_123 br_123 wl_83 vdd gnd cell_6t
Xbit_r84_c123 bl_123 br_123 wl_84 vdd gnd cell_6t
Xbit_r85_c123 bl_123 br_123 wl_85 vdd gnd cell_6t
Xbit_r86_c123 bl_123 br_123 wl_86 vdd gnd cell_6t
Xbit_r87_c123 bl_123 br_123 wl_87 vdd gnd cell_6t
Xbit_r88_c123 bl_123 br_123 wl_88 vdd gnd cell_6t
Xbit_r89_c123 bl_123 br_123 wl_89 vdd gnd cell_6t
Xbit_r90_c123 bl_123 br_123 wl_90 vdd gnd cell_6t
Xbit_r91_c123 bl_123 br_123 wl_91 vdd gnd cell_6t
Xbit_r92_c123 bl_123 br_123 wl_92 vdd gnd cell_6t
Xbit_r93_c123 bl_123 br_123 wl_93 vdd gnd cell_6t
Xbit_r94_c123 bl_123 br_123 wl_94 vdd gnd cell_6t
Xbit_r95_c123 bl_123 br_123 wl_95 vdd gnd cell_6t
Xbit_r96_c123 bl_123 br_123 wl_96 vdd gnd cell_6t
Xbit_r97_c123 bl_123 br_123 wl_97 vdd gnd cell_6t
Xbit_r98_c123 bl_123 br_123 wl_98 vdd gnd cell_6t
Xbit_r99_c123 bl_123 br_123 wl_99 vdd gnd cell_6t
Xbit_r100_c123 bl_123 br_123 wl_100 vdd gnd cell_6t
Xbit_r101_c123 bl_123 br_123 wl_101 vdd gnd cell_6t
Xbit_r102_c123 bl_123 br_123 wl_102 vdd gnd cell_6t
Xbit_r103_c123 bl_123 br_123 wl_103 vdd gnd cell_6t
Xbit_r104_c123 bl_123 br_123 wl_104 vdd gnd cell_6t
Xbit_r105_c123 bl_123 br_123 wl_105 vdd gnd cell_6t
Xbit_r106_c123 bl_123 br_123 wl_106 vdd gnd cell_6t
Xbit_r107_c123 bl_123 br_123 wl_107 vdd gnd cell_6t
Xbit_r108_c123 bl_123 br_123 wl_108 vdd gnd cell_6t
Xbit_r109_c123 bl_123 br_123 wl_109 vdd gnd cell_6t
Xbit_r110_c123 bl_123 br_123 wl_110 vdd gnd cell_6t
Xbit_r111_c123 bl_123 br_123 wl_111 vdd gnd cell_6t
Xbit_r112_c123 bl_123 br_123 wl_112 vdd gnd cell_6t
Xbit_r113_c123 bl_123 br_123 wl_113 vdd gnd cell_6t
Xbit_r114_c123 bl_123 br_123 wl_114 vdd gnd cell_6t
Xbit_r115_c123 bl_123 br_123 wl_115 vdd gnd cell_6t
Xbit_r116_c123 bl_123 br_123 wl_116 vdd gnd cell_6t
Xbit_r117_c123 bl_123 br_123 wl_117 vdd gnd cell_6t
Xbit_r118_c123 bl_123 br_123 wl_118 vdd gnd cell_6t
Xbit_r119_c123 bl_123 br_123 wl_119 vdd gnd cell_6t
Xbit_r120_c123 bl_123 br_123 wl_120 vdd gnd cell_6t
Xbit_r121_c123 bl_123 br_123 wl_121 vdd gnd cell_6t
Xbit_r122_c123 bl_123 br_123 wl_122 vdd gnd cell_6t
Xbit_r123_c123 bl_123 br_123 wl_123 vdd gnd cell_6t
Xbit_r124_c123 bl_123 br_123 wl_124 vdd gnd cell_6t
Xbit_r125_c123 bl_123 br_123 wl_125 vdd gnd cell_6t
Xbit_r126_c123 bl_123 br_123 wl_126 vdd gnd cell_6t
Xbit_r127_c123 bl_123 br_123 wl_127 vdd gnd cell_6t
Xbit_r128_c123 bl_123 br_123 wl_128 vdd gnd cell_6t
Xbit_r129_c123 bl_123 br_123 wl_129 vdd gnd cell_6t
Xbit_r130_c123 bl_123 br_123 wl_130 vdd gnd cell_6t
Xbit_r131_c123 bl_123 br_123 wl_131 vdd gnd cell_6t
Xbit_r132_c123 bl_123 br_123 wl_132 vdd gnd cell_6t
Xbit_r133_c123 bl_123 br_123 wl_133 vdd gnd cell_6t
Xbit_r134_c123 bl_123 br_123 wl_134 vdd gnd cell_6t
Xbit_r135_c123 bl_123 br_123 wl_135 vdd gnd cell_6t
Xbit_r136_c123 bl_123 br_123 wl_136 vdd gnd cell_6t
Xbit_r137_c123 bl_123 br_123 wl_137 vdd gnd cell_6t
Xbit_r138_c123 bl_123 br_123 wl_138 vdd gnd cell_6t
Xbit_r139_c123 bl_123 br_123 wl_139 vdd gnd cell_6t
Xbit_r140_c123 bl_123 br_123 wl_140 vdd gnd cell_6t
Xbit_r141_c123 bl_123 br_123 wl_141 vdd gnd cell_6t
Xbit_r142_c123 bl_123 br_123 wl_142 vdd gnd cell_6t
Xbit_r143_c123 bl_123 br_123 wl_143 vdd gnd cell_6t
Xbit_r144_c123 bl_123 br_123 wl_144 vdd gnd cell_6t
Xbit_r145_c123 bl_123 br_123 wl_145 vdd gnd cell_6t
Xbit_r146_c123 bl_123 br_123 wl_146 vdd gnd cell_6t
Xbit_r147_c123 bl_123 br_123 wl_147 vdd gnd cell_6t
Xbit_r148_c123 bl_123 br_123 wl_148 vdd gnd cell_6t
Xbit_r149_c123 bl_123 br_123 wl_149 vdd gnd cell_6t
Xbit_r150_c123 bl_123 br_123 wl_150 vdd gnd cell_6t
Xbit_r151_c123 bl_123 br_123 wl_151 vdd gnd cell_6t
Xbit_r152_c123 bl_123 br_123 wl_152 vdd gnd cell_6t
Xbit_r153_c123 bl_123 br_123 wl_153 vdd gnd cell_6t
Xbit_r154_c123 bl_123 br_123 wl_154 vdd gnd cell_6t
Xbit_r155_c123 bl_123 br_123 wl_155 vdd gnd cell_6t
Xbit_r156_c123 bl_123 br_123 wl_156 vdd gnd cell_6t
Xbit_r157_c123 bl_123 br_123 wl_157 vdd gnd cell_6t
Xbit_r158_c123 bl_123 br_123 wl_158 vdd gnd cell_6t
Xbit_r159_c123 bl_123 br_123 wl_159 vdd gnd cell_6t
Xbit_r160_c123 bl_123 br_123 wl_160 vdd gnd cell_6t
Xbit_r161_c123 bl_123 br_123 wl_161 vdd gnd cell_6t
Xbit_r162_c123 bl_123 br_123 wl_162 vdd gnd cell_6t
Xbit_r163_c123 bl_123 br_123 wl_163 vdd gnd cell_6t
Xbit_r164_c123 bl_123 br_123 wl_164 vdd gnd cell_6t
Xbit_r165_c123 bl_123 br_123 wl_165 vdd gnd cell_6t
Xbit_r166_c123 bl_123 br_123 wl_166 vdd gnd cell_6t
Xbit_r167_c123 bl_123 br_123 wl_167 vdd gnd cell_6t
Xbit_r168_c123 bl_123 br_123 wl_168 vdd gnd cell_6t
Xbit_r169_c123 bl_123 br_123 wl_169 vdd gnd cell_6t
Xbit_r170_c123 bl_123 br_123 wl_170 vdd gnd cell_6t
Xbit_r171_c123 bl_123 br_123 wl_171 vdd gnd cell_6t
Xbit_r172_c123 bl_123 br_123 wl_172 vdd gnd cell_6t
Xbit_r173_c123 bl_123 br_123 wl_173 vdd gnd cell_6t
Xbit_r174_c123 bl_123 br_123 wl_174 vdd gnd cell_6t
Xbit_r175_c123 bl_123 br_123 wl_175 vdd gnd cell_6t
Xbit_r176_c123 bl_123 br_123 wl_176 vdd gnd cell_6t
Xbit_r177_c123 bl_123 br_123 wl_177 vdd gnd cell_6t
Xbit_r178_c123 bl_123 br_123 wl_178 vdd gnd cell_6t
Xbit_r179_c123 bl_123 br_123 wl_179 vdd gnd cell_6t
Xbit_r180_c123 bl_123 br_123 wl_180 vdd gnd cell_6t
Xbit_r181_c123 bl_123 br_123 wl_181 vdd gnd cell_6t
Xbit_r182_c123 bl_123 br_123 wl_182 vdd gnd cell_6t
Xbit_r183_c123 bl_123 br_123 wl_183 vdd gnd cell_6t
Xbit_r184_c123 bl_123 br_123 wl_184 vdd gnd cell_6t
Xbit_r185_c123 bl_123 br_123 wl_185 vdd gnd cell_6t
Xbit_r186_c123 bl_123 br_123 wl_186 vdd gnd cell_6t
Xbit_r187_c123 bl_123 br_123 wl_187 vdd gnd cell_6t
Xbit_r188_c123 bl_123 br_123 wl_188 vdd gnd cell_6t
Xbit_r189_c123 bl_123 br_123 wl_189 vdd gnd cell_6t
Xbit_r190_c123 bl_123 br_123 wl_190 vdd gnd cell_6t
Xbit_r191_c123 bl_123 br_123 wl_191 vdd gnd cell_6t
Xbit_r192_c123 bl_123 br_123 wl_192 vdd gnd cell_6t
Xbit_r193_c123 bl_123 br_123 wl_193 vdd gnd cell_6t
Xbit_r194_c123 bl_123 br_123 wl_194 vdd gnd cell_6t
Xbit_r195_c123 bl_123 br_123 wl_195 vdd gnd cell_6t
Xbit_r196_c123 bl_123 br_123 wl_196 vdd gnd cell_6t
Xbit_r197_c123 bl_123 br_123 wl_197 vdd gnd cell_6t
Xbit_r198_c123 bl_123 br_123 wl_198 vdd gnd cell_6t
Xbit_r199_c123 bl_123 br_123 wl_199 vdd gnd cell_6t
Xbit_r200_c123 bl_123 br_123 wl_200 vdd gnd cell_6t
Xbit_r201_c123 bl_123 br_123 wl_201 vdd gnd cell_6t
Xbit_r202_c123 bl_123 br_123 wl_202 vdd gnd cell_6t
Xbit_r203_c123 bl_123 br_123 wl_203 vdd gnd cell_6t
Xbit_r204_c123 bl_123 br_123 wl_204 vdd gnd cell_6t
Xbit_r205_c123 bl_123 br_123 wl_205 vdd gnd cell_6t
Xbit_r206_c123 bl_123 br_123 wl_206 vdd gnd cell_6t
Xbit_r207_c123 bl_123 br_123 wl_207 vdd gnd cell_6t
Xbit_r208_c123 bl_123 br_123 wl_208 vdd gnd cell_6t
Xbit_r209_c123 bl_123 br_123 wl_209 vdd gnd cell_6t
Xbit_r210_c123 bl_123 br_123 wl_210 vdd gnd cell_6t
Xbit_r211_c123 bl_123 br_123 wl_211 vdd gnd cell_6t
Xbit_r212_c123 bl_123 br_123 wl_212 vdd gnd cell_6t
Xbit_r213_c123 bl_123 br_123 wl_213 vdd gnd cell_6t
Xbit_r214_c123 bl_123 br_123 wl_214 vdd gnd cell_6t
Xbit_r215_c123 bl_123 br_123 wl_215 vdd gnd cell_6t
Xbit_r216_c123 bl_123 br_123 wl_216 vdd gnd cell_6t
Xbit_r217_c123 bl_123 br_123 wl_217 vdd gnd cell_6t
Xbit_r218_c123 bl_123 br_123 wl_218 vdd gnd cell_6t
Xbit_r219_c123 bl_123 br_123 wl_219 vdd gnd cell_6t
Xbit_r220_c123 bl_123 br_123 wl_220 vdd gnd cell_6t
Xbit_r221_c123 bl_123 br_123 wl_221 vdd gnd cell_6t
Xbit_r222_c123 bl_123 br_123 wl_222 vdd gnd cell_6t
Xbit_r223_c123 bl_123 br_123 wl_223 vdd gnd cell_6t
Xbit_r224_c123 bl_123 br_123 wl_224 vdd gnd cell_6t
Xbit_r225_c123 bl_123 br_123 wl_225 vdd gnd cell_6t
Xbit_r226_c123 bl_123 br_123 wl_226 vdd gnd cell_6t
Xbit_r227_c123 bl_123 br_123 wl_227 vdd gnd cell_6t
Xbit_r228_c123 bl_123 br_123 wl_228 vdd gnd cell_6t
Xbit_r229_c123 bl_123 br_123 wl_229 vdd gnd cell_6t
Xbit_r230_c123 bl_123 br_123 wl_230 vdd gnd cell_6t
Xbit_r231_c123 bl_123 br_123 wl_231 vdd gnd cell_6t
Xbit_r232_c123 bl_123 br_123 wl_232 vdd gnd cell_6t
Xbit_r233_c123 bl_123 br_123 wl_233 vdd gnd cell_6t
Xbit_r234_c123 bl_123 br_123 wl_234 vdd gnd cell_6t
Xbit_r235_c123 bl_123 br_123 wl_235 vdd gnd cell_6t
Xbit_r236_c123 bl_123 br_123 wl_236 vdd gnd cell_6t
Xbit_r237_c123 bl_123 br_123 wl_237 vdd gnd cell_6t
Xbit_r238_c123 bl_123 br_123 wl_238 vdd gnd cell_6t
Xbit_r239_c123 bl_123 br_123 wl_239 vdd gnd cell_6t
Xbit_r240_c123 bl_123 br_123 wl_240 vdd gnd cell_6t
Xbit_r241_c123 bl_123 br_123 wl_241 vdd gnd cell_6t
Xbit_r242_c123 bl_123 br_123 wl_242 vdd gnd cell_6t
Xbit_r243_c123 bl_123 br_123 wl_243 vdd gnd cell_6t
Xbit_r244_c123 bl_123 br_123 wl_244 vdd gnd cell_6t
Xbit_r245_c123 bl_123 br_123 wl_245 vdd gnd cell_6t
Xbit_r246_c123 bl_123 br_123 wl_246 vdd gnd cell_6t
Xbit_r247_c123 bl_123 br_123 wl_247 vdd gnd cell_6t
Xbit_r248_c123 bl_123 br_123 wl_248 vdd gnd cell_6t
Xbit_r249_c123 bl_123 br_123 wl_249 vdd gnd cell_6t
Xbit_r250_c123 bl_123 br_123 wl_250 vdd gnd cell_6t
Xbit_r251_c123 bl_123 br_123 wl_251 vdd gnd cell_6t
Xbit_r252_c123 bl_123 br_123 wl_252 vdd gnd cell_6t
Xbit_r253_c123 bl_123 br_123 wl_253 vdd gnd cell_6t
Xbit_r254_c123 bl_123 br_123 wl_254 vdd gnd cell_6t
Xbit_r255_c123 bl_123 br_123 wl_255 vdd gnd cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd cell_6t
Xbit_r1_c124 bl_124 br_124 wl_1 vdd gnd cell_6t
Xbit_r2_c124 bl_124 br_124 wl_2 vdd gnd cell_6t
Xbit_r3_c124 bl_124 br_124 wl_3 vdd gnd cell_6t
Xbit_r4_c124 bl_124 br_124 wl_4 vdd gnd cell_6t
Xbit_r5_c124 bl_124 br_124 wl_5 vdd gnd cell_6t
Xbit_r6_c124 bl_124 br_124 wl_6 vdd gnd cell_6t
Xbit_r7_c124 bl_124 br_124 wl_7 vdd gnd cell_6t
Xbit_r8_c124 bl_124 br_124 wl_8 vdd gnd cell_6t
Xbit_r9_c124 bl_124 br_124 wl_9 vdd gnd cell_6t
Xbit_r10_c124 bl_124 br_124 wl_10 vdd gnd cell_6t
Xbit_r11_c124 bl_124 br_124 wl_11 vdd gnd cell_6t
Xbit_r12_c124 bl_124 br_124 wl_12 vdd gnd cell_6t
Xbit_r13_c124 bl_124 br_124 wl_13 vdd gnd cell_6t
Xbit_r14_c124 bl_124 br_124 wl_14 vdd gnd cell_6t
Xbit_r15_c124 bl_124 br_124 wl_15 vdd gnd cell_6t
Xbit_r16_c124 bl_124 br_124 wl_16 vdd gnd cell_6t
Xbit_r17_c124 bl_124 br_124 wl_17 vdd gnd cell_6t
Xbit_r18_c124 bl_124 br_124 wl_18 vdd gnd cell_6t
Xbit_r19_c124 bl_124 br_124 wl_19 vdd gnd cell_6t
Xbit_r20_c124 bl_124 br_124 wl_20 vdd gnd cell_6t
Xbit_r21_c124 bl_124 br_124 wl_21 vdd gnd cell_6t
Xbit_r22_c124 bl_124 br_124 wl_22 vdd gnd cell_6t
Xbit_r23_c124 bl_124 br_124 wl_23 vdd gnd cell_6t
Xbit_r24_c124 bl_124 br_124 wl_24 vdd gnd cell_6t
Xbit_r25_c124 bl_124 br_124 wl_25 vdd gnd cell_6t
Xbit_r26_c124 bl_124 br_124 wl_26 vdd gnd cell_6t
Xbit_r27_c124 bl_124 br_124 wl_27 vdd gnd cell_6t
Xbit_r28_c124 bl_124 br_124 wl_28 vdd gnd cell_6t
Xbit_r29_c124 bl_124 br_124 wl_29 vdd gnd cell_6t
Xbit_r30_c124 bl_124 br_124 wl_30 vdd gnd cell_6t
Xbit_r31_c124 bl_124 br_124 wl_31 vdd gnd cell_6t
Xbit_r32_c124 bl_124 br_124 wl_32 vdd gnd cell_6t
Xbit_r33_c124 bl_124 br_124 wl_33 vdd gnd cell_6t
Xbit_r34_c124 bl_124 br_124 wl_34 vdd gnd cell_6t
Xbit_r35_c124 bl_124 br_124 wl_35 vdd gnd cell_6t
Xbit_r36_c124 bl_124 br_124 wl_36 vdd gnd cell_6t
Xbit_r37_c124 bl_124 br_124 wl_37 vdd gnd cell_6t
Xbit_r38_c124 bl_124 br_124 wl_38 vdd gnd cell_6t
Xbit_r39_c124 bl_124 br_124 wl_39 vdd gnd cell_6t
Xbit_r40_c124 bl_124 br_124 wl_40 vdd gnd cell_6t
Xbit_r41_c124 bl_124 br_124 wl_41 vdd gnd cell_6t
Xbit_r42_c124 bl_124 br_124 wl_42 vdd gnd cell_6t
Xbit_r43_c124 bl_124 br_124 wl_43 vdd gnd cell_6t
Xbit_r44_c124 bl_124 br_124 wl_44 vdd gnd cell_6t
Xbit_r45_c124 bl_124 br_124 wl_45 vdd gnd cell_6t
Xbit_r46_c124 bl_124 br_124 wl_46 vdd gnd cell_6t
Xbit_r47_c124 bl_124 br_124 wl_47 vdd gnd cell_6t
Xbit_r48_c124 bl_124 br_124 wl_48 vdd gnd cell_6t
Xbit_r49_c124 bl_124 br_124 wl_49 vdd gnd cell_6t
Xbit_r50_c124 bl_124 br_124 wl_50 vdd gnd cell_6t
Xbit_r51_c124 bl_124 br_124 wl_51 vdd gnd cell_6t
Xbit_r52_c124 bl_124 br_124 wl_52 vdd gnd cell_6t
Xbit_r53_c124 bl_124 br_124 wl_53 vdd gnd cell_6t
Xbit_r54_c124 bl_124 br_124 wl_54 vdd gnd cell_6t
Xbit_r55_c124 bl_124 br_124 wl_55 vdd gnd cell_6t
Xbit_r56_c124 bl_124 br_124 wl_56 vdd gnd cell_6t
Xbit_r57_c124 bl_124 br_124 wl_57 vdd gnd cell_6t
Xbit_r58_c124 bl_124 br_124 wl_58 vdd gnd cell_6t
Xbit_r59_c124 bl_124 br_124 wl_59 vdd gnd cell_6t
Xbit_r60_c124 bl_124 br_124 wl_60 vdd gnd cell_6t
Xbit_r61_c124 bl_124 br_124 wl_61 vdd gnd cell_6t
Xbit_r62_c124 bl_124 br_124 wl_62 vdd gnd cell_6t
Xbit_r63_c124 bl_124 br_124 wl_63 vdd gnd cell_6t
Xbit_r64_c124 bl_124 br_124 wl_64 vdd gnd cell_6t
Xbit_r65_c124 bl_124 br_124 wl_65 vdd gnd cell_6t
Xbit_r66_c124 bl_124 br_124 wl_66 vdd gnd cell_6t
Xbit_r67_c124 bl_124 br_124 wl_67 vdd gnd cell_6t
Xbit_r68_c124 bl_124 br_124 wl_68 vdd gnd cell_6t
Xbit_r69_c124 bl_124 br_124 wl_69 vdd gnd cell_6t
Xbit_r70_c124 bl_124 br_124 wl_70 vdd gnd cell_6t
Xbit_r71_c124 bl_124 br_124 wl_71 vdd gnd cell_6t
Xbit_r72_c124 bl_124 br_124 wl_72 vdd gnd cell_6t
Xbit_r73_c124 bl_124 br_124 wl_73 vdd gnd cell_6t
Xbit_r74_c124 bl_124 br_124 wl_74 vdd gnd cell_6t
Xbit_r75_c124 bl_124 br_124 wl_75 vdd gnd cell_6t
Xbit_r76_c124 bl_124 br_124 wl_76 vdd gnd cell_6t
Xbit_r77_c124 bl_124 br_124 wl_77 vdd gnd cell_6t
Xbit_r78_c124 bl_124 br_124 wl_78 vdd gnd cell_6t
Xbit_r79_c124 bl_124 br_124 wl_79 vdd gnd cell_6t
Xbit_r80_c124 bl_124 br_124 wl_80 vdd gnd cell_6t
Xbit_r81_c124 bl_124 br_124 wl_81 vdd gnd cell_6t
Xbit_r82_c124 bl_124 br_124 wl_82 vdd gnd cell_6t
Xbit_r83_c124 bl_124 br_124 wl_83 vdd gnd cell_6t
Xbit_r84_c124 bl_124 br_124 wl_84 vdd gnd cell_6t
Xbit_r85_c124 bl_124 br_124 wl_85 vdd gnd cell_6t
Xbit_r86_c124 bl_124 br_124 wl_86 vdd gnd cell_6t
Xbit_r87_c124 bl_124 br_124 wl_87 vdd gnd cell_6t
Xbit_r88_c124 bl_124 br_124 wl_88 vdd gnd cell_6t
Xbit_r89_c124 bl_124 br_124 wl_89 vdd gnd cell_6t
Xbit_r90_c124 bl_124 br_124 wl_90 vdd gnd cell_6t
Xbit_r91_c124 bl_124 br_124 wl_91 vdd gnd cell_6t
Xbit_r92_c124 bl_124 br_124 wl_92 vdd gnd cell_6t
Xbit_r93_c124 bl_124 br_124 wl_93 vdd gnd cell_6t
Xbit_r94_c124 bl_124 br_124 wl_94 vdd gnd cell_6t
Xbit_r95_c124 bl_124 br_124 wl_95 vdd gnd cell_6t
Xbit_r96_c124 bl_124 br_124 wl_96 vdd gnd cell_6t
Xbit_r97_c124 bl_124 br_124 wl_97 vdd gnd cell_6t
Xbit_r98_c124 bl_124 br_124 wl_98 vdd gnd cell_6t
Xbit_r99_c124 bl_124 br_124 wl_99 vdd gnd cell_6t
Xbit_r100_c124 bl_124 br_124 wl_100 vdd gnd cell_6t
Xbit_r101_c124 bl_124 br_124 wl_101 vdd gnd cell_6t
Xbit_r102_c124 bl_124 br_124 wl_102 vdd gnd cell_6t
Xbit_r103_c124 bl_124 br_124 wl_103 vdd gnd cell_6t
Xbit_r104_c124 bl_124 br_124 wl_104 vdd gnd cell_6t
Xbit_r105_c124 bl_124 br_124 wl_105 vdd gnd cell_6t
Xbit_r106_c124 bl_124 br_124 wl_106 vdd gnd cell_6t
Xbit_r107_c124 bl_124 br_124 wl_107 vdd gnd cell_6t
Xbit_r108_c124 bl_124 br_124 wl_108 vdd gnd cell_6t
Xbit_r109_c124 bl_124 br_124 wl_109 vdd gnd cell_6t
Xbit_r110_c124 bl_124 br_124 wl_110 vdd gnd cell_6t
Xbit_r111_c124 bl_124 br_124 wl_111 vdd gnd cell_6t
Xbit_r112_c124 bl_124 br_124 wl_112 vdd gnd cell_6t
Xbit_r113_c124 bl_124 br_124 wl_113 vdd gnd cell_6t
Xbit_r114_c124 bl_124 br_124 wl_114 vdd gnd cell_6t
Xbit_r115_c124 bl_124 br_124 wl_115 vdd gnd cell_6t
Xbit_r116_c124 bl_124 br_124 wl_116 vdd gnd cell_6t
Xbit_r117_c124 bl_124 br_124 wl_117 vdd gnd cell_6t
Xbit_r118_c124 bl_124 br_124 wl_118 vdd gnd cell_6t
Xbit_r119_c124 bl_124 br_124 wl_119 vdd gnd cell_6t
Xbit_r120_c124 bl_124 br_124 wl_120 vdd gnd cell_6t
Xbit_r121_c124 bl_124 br_124 wl_121 vdd gnd cell_6t
Xbit_r122_c124 bl_124 br_124 wl_122 vdd gnd cell_6t
Xbit_r123_c124 bl_124 br_124 wl_123 vdd gnd cell_6t
Xbit_r124_c124 bl_124 br_124 wl_124 vdd gnd cell_6t
Xbit_r125_c124 bl_124 br_124 wl_125 vdd gnd cell_6t
Xbit_r126_c124 bl_124 br_124 wl_126 vdd gnd cell_6t
Xbit_r127_c124 bl_124 br_124 wl_127 vdd gnd cell_6t
Xbit_r128_c124 bl_124 br_124 wl_128 vdd gnd cell_6t
Xbit_r129_c124 bl_124 br_124 wl_129 vdd gnd cell_6t
Xbit_r130_c124 bl_124 br_124 wl_130 vdd gnd cell_6t
Xbit_r131_c124 bl_124 br_124 wl_131 vdd gnd cell_6t
Xbit_r132_c124 bl_124 br_124 wl_132 vdd gnd cell_6t
Xbit_r133_c124 bl_124 br_124 wl_133 vdd gnd cell_6t
Xbit_r134_c124 bl_124 br_124 wl_134 vdd gnd cell_6t
Xbit_r135_c124 bl_124 br_124 wl_135 vdd gnd cell_6t
Xbit_r136_c124 bl_124 br_124 wl_136 vdd gnd cell_6t
Xbit_r137_c124 bl_124 br_124 wl_137 vdd gnd cell_6t
Xbit_r138_c124 bl_124 br_124 wl_138 vdd gnd cell_6t
Xbit_r139_c124 bl_124 br_124 wl_139 vdd gnd cell_6t
Xbit_r140_c124 bl_124 br_124 wl_140 vdd gnd cell_6t
Xbit_r141_c124 bl_124 br_124 wl_141 vdd gnd cell_6t
Xbit_r142_c124 bl_124 br_124 wl_142 vdd gnd cell_6t
Xbit_r143_c124 bl_124 br_124 wl_143 vdd gnd cell_6t
Xbit_r144_c124 bl_124 br_124 wl_144 vdd gnd cell_6t
Xbit_r145_c124 bl_124 br_124 wl_145 vdd gnd cell_6t
Xbit_r146_c124 bl_124 br_124 wl_146 vdd gnd cell_6t
Xbit_r147_c124 bl_124 br_124 wl_147 vdd gnd cell_6t
Xbit_r148_c124 bl_124 br_124 wl_148 vdd gnd cell_6t
Xbit_r149_c124 bl_124 br_124 wl_149 vdd gnd cell_6t
Xbit_r150_c124 bl_124 br_124 wl_150 vdd gnd cell_6t
Xbit_r151_c124 bl_124 br_124 wl_151 vdd gnd cell_6t
Xbit_r152_c124 bl_124 br_124 wl_152 vdd gnd cell_6t
Xbit_r153_c124 bl_124 br_124 wl_153 vdd gnd cell_6t
Xbit_r154_c124 bl_124 br_124 wl_154 vdd gnd cell_6t
Xbit_r155_c124 bl_124 br_124 wl_155 vdd gnd cell_6t
Xbit_r156_c124 bl_124 br_124 wl_156 vdd gnd cell_6t
Xbit_r157_c124 bl_124 br_124 wl_157 vdd gnd cell_6t
Xbit_r158_c124 bl_124 br_124 wl_158 vdd gnd cell_6t
Xbit_r159_c124 bl_124 br_124 wl_159 vdd gnd cell_6t
Xbit_r160_c124 bl_124 br_124 wl_160 vdd gnd cell_6t
Xbit_r161_c124 bl_124 br_124 wl_161 vdd gnd cell_6t
Xbit_r162_c124 bl_124 br_124 wl_162 vdd gnd cell_6t
Xbit_r163_c124 bl_124 br_124 wl_163 vdd gnd cell_6t
Xbit_r164_c124 bl_124 br_124 wl_164 vdd gnd cell_6t
Xbit_r165_c124 bl_124 br_124 wl_165 vdd gnd cell_6t
Xbit_r166_c124 bl_124 br_124 wl_166 vdd gnd cell_6t
Xbit_r167_c124 bl_124 br_124 wl_167 vdd gnd cell_6t
Xbit_r168_c124 bl_124 br_124 wl_168 vdd gnd cell_6t
Xbit_r169_c124 bl_124 br_124 wl_169 vdd gnd cell_6t
Xbit_r170_c124 bl_124 br_124 wl_170 vdd gnd cell_6t
Xbit_r171_c124 bl_124 br_124 wl_171 vdd gnd cell_6t
Xbit_r172_c124 bl_124 br_124 wl_172 vdd gnd cell_6t
Xbit_r173_c124 bl_124 br_124 wl_173 vdd gnd cell_6t
Xbit_r174_c124 bl_124 br_124 wl_174 vdd gnd cell_6t
Xbit_r175_c124 bl_124 br_124 wl_175 vdd gnd cell_6t
Xbit_r176_c124 bl_124 br_124 wl_176 vdd gnd cell_6t
Xbit_r177_c124 bl_124 br_124 wl_177 vdd gnd cell_6t
Xbit_r178_c124 bl_124 br_124 wl_178 vdd gnd cell_6t
Xbit_r179_c124 bl_124 br_124 wl_179 vdd gnd cell_6t
Xbit_r180_c124 bl_124 br_124 wl_180 vdd gnd cell_6t
Xbit_r181_c124 bl_124 br_124 wl_181 vdd gnd cell_6t
Xbit_r182_c124 bl_124 br_124 wl_182 vdd gnd cell_6t
Xbit_r183_c124 bl_124 br_124 wl_183 vdd gnd cell_6t
Xbit_r184_c124 bl_124 br_124 wl_184 vdd gnd cell_6t
Xbit_r185_c124 bl_124 br_124 wl_185 vdd gnd cell_6t
Xbit_r186_c124 bl_124 br_124 wl_186 vdd gnd cell_6t
Xbit_r187_c124 bl_124 br_124 wl_187 vdd gnd cell_6t
Xbit_r188_c124 bl_124 br_124 wl_188 vdd gnd cell_6t
Xbit_r189_c124 bl_124 br_124 wl_189 vdd gnd cell_6t
Xbit_r190_c124 bl_124 br_124 wl_190 vdd gnd cell_6t
Xbit_r191_c124 bl_124 br_124 wl_191 vdd gnd cell_6t
Xbit_r192_c124 bl_124 br_124 wl_192 vdd gnd cell_6t
Xbit_r193_c124 bl_124 br_124 wl_193 vdd gnd cell_6t
Xbit_r194_c124 bl_124 br_124 wl_194 vdd gnd cell_6t
Xbit_r195_c124 bl_124 br_124 wl_195 vdd gnd cell_6t
Xbit_r196_c124 bl_124 br_124 wl_196 vdd gnd cell_6t
Xbit_r197_c124 bl_124 br_124 wl_197 vdd gnd cell_6t
Xbit_r198_c124 bl_124 br_124 wl_198 vdd gnd cell_6t
Xbit_r199_c124 bl_124 br_124 wl_199 vdd gnd cell_6t
Xbit_r200_c124 bl_124 br_124 wl_200 vdd gnd cell_6t
Xbit_r201_c124 bl_124 br_124 wl_201 vdd gnd cell_6t
Xbit_r202_c124 bl_124 br_124 wl_202 vdd gnd cell_6t
Xbit_r203_c124 bl_124 br_124 wl_203 vdd gnd cell_6t
Xbit_r204_c124 bl_124 br_124 wl_204 vdd gnd cell_6t
Xbit_r205_c124 bl_124 br_124 wl_205 vdd gnd cell_6t
Xbit_r206_c124 bl_124 br_124 wl_206 vdd gnd cell_6t
Xbit_r207_c124 bl_124 br_124 wl_207 vdd gnd cell_6t
Xbit_r208_c124 bl_124 br_124 wl_208 vdd gnd cell_6t
Xbit_r209_c124 bl_124 br_124 wl_209 vdd gnd cell_6t
Xbit_r210_c124 bl_124 br_124 wl_210 vdd gnd cell_6t
Xbit_r211_c124 bl_124 br_124 wl_211 vdd gnd cell_6t
Xbit_r212_c124 bl_124 br_124 wl_212 vdd gnd cell_6t
Xbit_r213_c124 bl_124 br_124 wl_213 vdd gnd cell_6t
Xbit_r214_c124 bl_124 br_124 wl_214 vdd gnd cell_6t
Xbit_r215_c124 bl_124 br_124 wl_215 vdd gnd cell_6t
Xbit_r216_c124 bl_124 br_124 wl_216 vdd gnd cell_6t
Xbit_r217_c124 bl_124 br_124 wl_217 vdd gnd cell_6t
Xbit_r218_c124 bl_124 br_124 wl_218 vdd gnd cell_6t
Xbit_r219_c124 bl_124 br_124 wl_219 vdd gnd cell_6t
Xbit_r220_c124 bl_124 br_124 wl_220 vdd gnd cell_6t
Xbit_r221_c124 bl_124 br_124 wl_221 vdd gnd cell_6t
Xbit_r222_c124 bl_124 br_124 wl_222 vdd gnd cell_6t
Xbit_r223_c124 bl_124 br_124 wl_223 vdd gnd cell_6t
Xbit_r224_c124 bl_124 br_124 wl_224 vdd gnd cell_6t
Xbit_r225_c124 bl_124 br_124 wl_225 vdd gnd cell_6t
Xbit_r226_c124 bl_124 br_124 wl_226 vdd gnd cell_6t
Xbit_r227_c124 bl_124 br_124 wl_227 vdd gnd cell_6t
Xbit_r228_c124 bl_124 br_124 wl_228 vdd gnd cell_6t
Xbit_r229_c124 bl_124 br_124 wl_229 vdd gnd cell_6t
Xbit_r230_c124 bl_124 br_124 wl_230 vdd gnd cell_6t
Xbit_r231_c124 bl_124 br_124 wl_231 vdd gnd cell_6t
Xbit_r232_c124 bl_124 br_124 wl_232 vdd gnd cell_6t
Xbit_r233_c124 bl_124 br_124 wl_233 vdd gnd cell_6t
Xbit_r234_c124 bl_124 br_124 wl_234 vdd gnd cell_6t
Xbit_r235_c124 bl_124 br_124 wl_235 vdd gnd cell_6t
Xbit_r236_c124 bl_124 br_124 wl_236 vdd gnd cell_6t
Xbit_r237_c124 bl_124 br_124 wl_237 vdd gnd cell_6t
Xbit_r238_c124 bl_124 br_124 wl_238 vdd gnd cell_6t
Xbit_r239_c124 bl_124 br_124 wl_239 vdd gnd cell_6t
Xbit_r240_c124 bl_124 br_124 wl_240 vdd gnd cell_6t
Xbit_r241_c124 bl_124 br_124 wl_241 vdd gnd cell_6t
Xbit_r242_c124 bl_124 br_124 wl_242 vdd gnd cell_6t
Xbit_r243_c124 bl_124 br_124 wl_243 vdd gnd cell_6t
Xbit_r244_c124 bl_124 br_124 wl_244 vdd gnd cell_6t
Xbit_r245_c124 bl_124 br_124 wl_245 vdd gnd cell_6t
Xbit_r246_c124 bl_124 br_124 wl_246 vdd gnd cell_6t
Xbit_r247_c124 bl_124 br_124 wl_247 vdd gnd cell_6t
Xbit_r248_c124 bl_124 br_124 wl_248 vdd gnd cell_6t
Xbit_r249_c124 bl_124 br_124 wl_249 vdd gnd cell_6t
Xbit_r250_c124 bl_124 br_124 wl_250 vdd gnd cell_6t
Xbit_r251_c124 bl_124 br_124 wl_251 vdd gnd cell_6t
Xbit_r252_c124 bl_124 br_124 wl_252 vdd gnd cell_6t
Xbit_r253_c124 bl_124 br_124 wl_253 vdd gnd cell_6t
Xbit_r254_c124 bl_124 br_124 wl_254 vdd gnd cell_6t
Xbit_r255_c124 bl_124 br_124 wl_255 vdd gnd cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd cell_6t
Xbit_r1_c125 bl_125 br_125 wl_1 vdd gnd cell_6t
Xbit_r2_c125 bl_125 br_125 wl_2 vdd gnd cell_6t
Xbit_r3_c125 bl_125 br_125 wl_3 vdd gnd cell_6t
Xbit_r4_c125 bl_125 br_125 wl_4 vdd gnd cell_6t
Xbit_r5_c125 bl_125 br_125 wl_5 vdd gnd cell_6t
Xbit_r6_c125 bl_125 br_125 wl_6 vdd gnd cell_6t
Xbit_r7_c125 bl_125 br_125 wl_7 vdd gnd cell_6t
Xbit_r8_c125 bl_125 br_125 wl_8 vdd gnd cell_6t
Xbit_r9_c125 bl_125 br_125 wl_9 vdd gnd cell_6t
Xbit_r10_c125 bl_125 br_125 wl_10 vdd gnd cell_6t
Xbit_r11_c125 bl_125 br_125 wl_11 vdd gnd cell_6t
Xbit_r12_c125 bl_125 br_125 wl_12 vdd gnd cell_6t
Xbit_r13_c125 bl_125 br_125 wl_13 vdd gnd cell_6t
Xbit_r14_c125 bl_125 br_125 wl_14 vdd gnd cell_6t
Xbit_r15_c125 bl_125 br_125 wl_15 vdd gnd cell_6t
Xbit_r16_c125 bl_125 br_125 wl_16 vdd gnd cell_6t
Xbit_r17_c125 bl_125 br_125 wl_17 vdd gnd cell_6t
Xbit_r18_c125 bl_125 br_125 wl_18 vdd gnd cell_6t
Xbit_r19_c125 bl_125 br_125 wl_19 vdd gnd cell_6t
Xbit_r20_c125 bl_125 br_125 wl_20 vdd gnd cell_6t
Xbit_r21_c125 bl_125 br_125 wl_21 vdd gnd cell_6t
Xbit_r22_c125 bl_125 br_125 wl_22 vdd gnd cell_6t
Xbit_r23_c125 bl_125 br_125 wl_23 vdd gnd cell_6t
Xbit_r24_c125 bl_125 br_125 wl_24 vdd gnd cell_6t
Xbit_r25_c125 bl_125 br_125 wl_25 vdd gnd cell_6t
Xbit_r26_c125 bl_125 br_125 wl_26 vdd gnd cell_6t
Xbit_r27_c125 bl_125 br_125 wl_27 vdd gnd cell_6t
Xbit_r28_c125 bl_125 br_125 wl_28 vdd gnd cell_6t
Xbit_r29_c125 bl_125 br_125 wl_29 vdd gnd cell_6t
Xbit_r30_c125 bl_125 br_125 wl_30 vdd gnd cell_6t
Xbit_r31_c125 bl_125 br_125 wl_31 vdd gnd cell_6t
Xbit_r32_c125 bl_125 br_125 wl_32 vdd gnd cell_6t
Xbit_r33_c125 bl_125 br_125 wl_33 vdd gnd cell_6t
Xbit_r34_c125 bl_125 br_125 wl_34 vdd gnd cell_6t
Xbit_r35_c125 bl_125 br_125 wl_35 vdd gnd cell_6t
Xbit_r36_c125 bl_125 br_125 wl_36 vdd gnd cell_6t
Xbit_r37_c125 bl_125 br_125 wl_37 vdd gnd cell_6t
Xbit_r38_c125 bl_125 br_125 wl_38 vdd gnd cell_6t
Xbit_r39_c125 bl_125 br_125 wl_39 vdd gnd cell_6t
Xbit_r40_c125 bl_125 br_125 wl_40 vdd gnd cell_6t
Xbit_r41_c125 bl_125 br_125 wl_41 vdd gnd cell_6t
Xbit_r42_c125 bl_125 br_125 wl_42 vdd gnd cell_6t
Xbit_r43_c125 bl_125 br_125 wl_43 vdd gnd cell_6t
Xbit_r44_c125 bl_125 br_125 wl_44 vdd gnd cell_6t
Xbit_r45_c125 bl_125 br_125 wl_45 vdd gnd cell_6t
Xbit_r46_c125 bl_125 br_125 wl_46 vdd gnd cell_6t
Xbit_r47_c125 bl_125 br_125 wl_47 vdd gnd cell_6t
Xbit_r48_c125 bl_125 br_125 wl_48 vdd gnd cell_6t
Xbit_r49_c125 bl_125 br_125 wl_49 vdd gnd cell_6t
Xbit_r50_c125 bl_125 br_125 wl_50 vdd gnd cell_6t
Xbit_r51_c125 bl_125 br_125 wl_51 vdd gnd cell_6t
Xbit_r52_c125 bl_125 br_125 wl_52 vdd gnd cell_6t
Xbit_r53_c125 bl_125 br_125 wl_53 vdd gnd cell_6t
Xbit_r54_c125 bl_125 br_125 wl_54 vdd gnd cell_6t
Xbit_r55_c125 bl_125 br_125 wl_55 vdd gnd cell_6t
Xbit_r56_c125 bl_125 br_125 wl_56 vdd gnd cell_6t
Xbit_r57_c125 bl_125 br_125 wl_57 vdd gnd cell_6t
Xbit_r58_c125 bl_125 br_125 wl_58 vdd gnd cell_6t
Xbit_r59_c125 bl_125 br_125 wl_59 vdd gnd cell_6t
Xbit_r60_c125 bl_125 br_125 wl_60 vdd gnd cell_6t
Xbit_r61_c125 bl_125 br_125 wl_61 vdd gnd cell_6t
Xbit_r62_c125 bl_125 br_125 wl_62 vdd gnd cell_6t
Xbit_r63_c125 bl_125 br_125 wl_63 vdd gnd cell_6t
Xbit_r64_c125 bl_125 br_125 wl_64 vdd gnd cell_6t
Xbit_r65_c125 bl_125 br_125 wl_65 vdd gnd cell_6t
Xbit_r66_c125 bl_125 br_125 wl_66 vdd gnd cell_6t
Xbit_r67_c125 bl_125 br_125 wl_67 vdd gnd cell_6t
Xbit_r68_c125 bl_125 br_125 wl_68 vdd gnd cell_6t
Xbit_r69_c125 bl_125 br_125 wl_69 vdd gnd cell_6t
Xbit_r70_c125 bl_125 br_125 wl_70 vdd gnd cell_6t
Xbit_r71_c125 bl_125 br_125 wl_71 vdd gnd cell_6t
Xbit_r72_c125 bl_125 br_125 wl_72 vdd gnd cell_6t
Xbit_r73_c125 bl_125 br_125 wl_73 vdd gnd cell_6t
Xbit_r74_c125 bl_125 br_125 wl_74 vdd gnd cell_6t
Xbit_r75_c125 bl_125 br_125 wl_75 vdd gnd cell_6t
Xbit_r76_c125 bl_125 br_125 wl_76 vdd gnd cell_6t
Xbit_r77_c125 bl_125 br_125 wl_77 vdd gnd cell_6t
Xbit_r78_c125 bl_125 br_125 wl_78 vdd gnd cell_6t
Xbit_r79_c125 bl_125 br_125 wl_79 vdd gnd cell_6t
Xbit_r80_c125 bl_125 br_125 wl_80 vdd gnd cell_6t
Xbit_r81_c125 bl_125 br_125 wl_81 vdd gnd cell_6t
Xbit_r82_c125 bl_125 br_125 wl_82 vdd gnd cell_6t
Xbit_r83_c125 bl_125 br_125 wl_83 vdd gnd cell_6t
Xbit_r84_c125 bl_125 br_125 wl_84 vdd gnd cell_6t
Xbit_r85_c125 bl_125 br_125 wl_85 vdd gnd cell_6t
Xbit_r86_c125 bl_125 br_125 wl_86 vdd gnd cell_6t
Xbit_r87_c125 bl_125 br_125 wl_87 vdd gnd cell_6t
Xbit_r88_c125 bl_125 br_125 wl_88 vdd gnd cell_6t
Xbit_r89_c125 bl_125 br_125 wl_89 vdd gnd cell_6t
Xbit_r90_c125 bl_125 br_125 wl_90 vdd gnd cell_6t
Xbit_r91_c125 bl_125 br_125 wl_91 vdd gnd cell_6t
Xbit_r92_c125 bl_125 br_125 wl_92 vdd gnd cell_6t
Xbit_r93_c125 bl_125 br_125 wl_93 vdd gnd cell_6t
Xbit_r94_c125 bl_125 br_125 wl_94 vdd gnd cell_6t
Xbit_r95_c125 bl_125 br_125 wl_95 vdd gnd cell_6t
Xbit_r96_c125 bl_125 br_125 wl_96 vdd gnd cell_6t
Xbit_r97_c125 bl_125 br_125 wl_97 vdd gnd cell_6t
Xbit_r98_c125 bl_125 br_125 wl_98 vdd gnd cell_6t
Xbit_r99_c125 bl_125 br_125 wl_99 vdd gnd cell_6t
Xbit_r100_c125 bl_125 br_125 wl_100 vdd gnd cell_6t
Xbit_r101_c125 bl_125 br_125 wl_101 vdd gnd cell_6t
Xbit_r102_c125 bl_125 br_125 wl_102 vdd gnd cell_6t
Xbit_r103_c125 bl_125 br_125 wl_103 vdd gnd cell_6t
Xbit_r104_c125 bl_125 br_125 wl_104 vdd gnd cell_6t
Xbit_r105_c125 bl_125 br_125 wl_105 vdd gnd cell_6t
Xbit_r106_c125 bl_125 br_125 wl_106 vdd gnd cell_6t
Xbit_r107_c125 bl_125 br_125 wl_107 vdd gnd cell_6t
Xbit_r108_c125 bl_125 br_125 wl_108 vdd gnd cell_6t
Xbit_r109_c125 bl_125 br_125 wl_109 vdd gnd cell_6t
Xbit_r110_c125 bl_125 br_125 wl_110 vdd gnd cell_6t
Xbit_r111_c125 bl_125 br_125 wl_111 vdd gnd cell_6t
Xbit_r112_c125 bl_125 br_125 wl_112 vdd gnd cell_6t
Xbit_r113_c125 bl_125 br_125 wl_113 vdd gnd cell_6t
Xbit_r114_c125 bl_125 br_125 wl_114 vdd gnd cell_6t
Xbit_r115_c125 bl_125 br_125 wl_115 vdd gnd cell_6t
Xbit_r116_c125 bl_125 br_125 wl_116 vdd gnd cell_6t
Xbit_r117_c125 bl_125 br_125 wl_117 vdd gnd cell_6t
Xbit_r118_c125 bl_125 br_125 wl_118 vdd gnd cell_6t
Xbit_r119_c125 bl_125 br_125 wl_119 vdd gnd cell_6t
Xbit_r120_c125 bl_125 br_125 wl_120 vdd gnd cell_6t
Xbit_r121_c125 bl_125 br_125 wl_121 vdd gnd cell_6t
Xbit_r122_c125 bl_125 br_125 wl_122 vdd gnd cell_6t
Xbit_r123_c125 bl_125 br_125 wl_123 vdd gnd cell_6t
Xbit_r124_c125 bl_125 br_125 wl_124 vdd gnd cell_6t
Xbit_r125_c125 bl_125 br_125 wl_125 vdd gnd cell_6t
Xbit_r126_c125 bl_125 br_125 wl_126 vdd gnd cell_6t
Xbit_r127_c125 bl_125 br_125 wl_127 vdd gnd cell_6t
Xbit_r128_c125 bl_125 br_125 wl_128 vdd gnd cell_6t
Xbit_r129_c125 bl_125 br_125 wl_129 vdd gnd cell_6t
Xbit_r130_c125 bl_125 br_125 wl_130 vdd gnd cell_6t
Xbit_r131_c125 bl_125 br_125 wl_131 vdd gnd cell_6t
Xbit_r132_c125 bl_125 br_125 wl_132 vdd gnd cell_6t
Xbit_r133_c125 bl_125 br_125 wl_133 vdd gnd cell_6t
Xbit_r134_c125 bl_125 br_125 wl_134 vdd gnd cell_6t
Xbit_r135_c125 bl_125 br_125 wl_135 vdd gnd cell_6t
Xbit_r136_c125 bl_125 br_125 wl_136 vdd gnd cell_6t
Xbit_r137_c125 bl_125 br_125 wl_137 vdd gnd cell_6t
Xbit_r138_c125 bl_125 br_125 wl_138 vdd gnd cell_6t
Xbit_r139_c125 bl_125 br_125 wl_139 vdd gnd cell_6t
Xbit_r140_c125 bl_125 br_125 wl_140 vdd gnd cell_6t
Xbit_r141_c125 bl_125 br_125 wl_141 vdd gnd cell_6t
Xbit_r142_c125 bl_125 br_125 wl_142 vdd gnd cell_6t
Xbit_r143_c125 bl_125 br_125 wl_143 vdd gnd cell_6t
Xbit_r144_c125 bl_125 br_125 wl_144 vdd gnd cell_6t
Xbit_r145_c125 bl_125 br_125 wl_145 vdd gnd cell_6t
Xbit_r146_c125 bl_125 br_125 wl_146 vdd gnd cell_6t
Xbit_r147_c125 bl_125 br_125 wl_147 vdd gnd cell_6t
Xbit_r148_c125 bl_125 br_125 wl_148 vdd gnd cell_6t
Xbit_r149_c125 bl_125 br_125 wl_149 vdd gnd cell_6t
Xbit_r150_c125 bl_125 br_125 wl_150 vdd gnd cell_6t
Xbit_r151_c125 bl_125 br_125 wl_151 vdd gnd cell_6t
Xbit_r152_c125 bl_125 br_125 wl_152 vdd gnd cell_6t
Xbit_r153_c125 bl_125 br_125 wl_153 vdd gnd cell_6t
Xbit_r154_c125 bl_125 br_125 wl_154 vdd gnd cell_6t
Xbit_r155_c125 bl_125 br_125 wl_155 vdd gnd cell_6t
Xbit_r156_c125 bl_125 br_125 wl_156 vdd gnd cell_6t
Xbit_r157_c125 bl_125 br_125 wl_157 vdd gnd cell_6t
Xbit_r158_c125 bl_125 br_125 wl_158 vdd gnd cell_6t
Xbit_r159_c125 bl_125 br_125 wl_159 vdd gnd cell_6t
Xbit_r160_c125 bl_125 br_125 wl_160 vdd gnd cell_6t
Xbit_r161_c125 bl_125 br_125 wl_161 vdd gnd cell_6t
Xbit_r162_c125 bl_125 br_125 wl_162 vdd gnd cell_6t
Xbit_r163_c125 bl_125 br_125 wl_163 vdd gnd cell_6t
Xbit_r164_c125 bl_125 br_125 wl_164 vdd gnd cell_6t
Xbit_r165_c125 bl_125 br_125 wl_165 vdd gnd cell_6t
Xbit_r166_c125 bl_125 br_125 wl_166 vdd gnd cell_6t
Xbit_r167_c125 bl_125 br_125 wl_167 vdd gnd cell_6t
Xbit_r168_c125 bl_125 br_125 wl_168 vdd gnd cell_6t
Xbit_r169_c125 bl_125 br_125 wl_169 vdd gnd cell_6t
Xbit_r170_c125 bl_125 br_125 wl_170 vdd gnd cell_6t
Xbit_r171_c125 bl_125 br_125 wl_171 vdd gnd cell_6t
Xbit_r172_c125 bl_125 br_125 wl_172 vdd gnd cell_6t
Xbit_r173_c125 bl_125 br_125 wl_173 vdd gnd cell_6t
Xbit_r174_c125 bl_125 br_125 wl_174 vdd gnd cell_6t
Xbit_r175_c125 bl_125 br_125 wl_175 vdd gnd cell_6t
Xbit_r176_c125 bl_125 br_125 wl_176 vdd gnd cell_6t
Xbit_r177_c125 bl_125 br_125 wl_177 vdd gnd cell_6t
Xbit_r178_c125 bl_125 br_125 wl_178 vdd gnd cell_6t
Xbit_r179_c125 bl_125 br_125 wl_179 vdd gnd cell_6t
Xbit_r180_c125 bl_125 br_125 wl_180 vdd gnd cell_6t
Xbit_r181_c125 bl_125 br_125 wl_181 vdd gnd cell_6t
Xbit_r182_c125 bl_125 br_125 wl_182 vdd gnd cell_6t
Xbit_r183_c125 bl_125 br_125 wl_183 vdd gnd cell_6t
Xbit_r184_c125 bl_125 br_125 wl_184 vdd gnd cell_6t
Xbit_r185_c125 bl_125 br_125 wl_185 vdd gnd cell_6t
Xbit_r186_c125 bl_125 br_125 wl_186 vdd gnd cell_6t
Xbit_r187_c125 bl_125 br_125 wl_187 vdd gnd cell_6t
Xbit_r188_c125 bl_125 br_125 wl_188 vdd gnd cell_6t
Xbit_r189_c125 bl_125 br_125 wl_189 vdd gnd cell_6t
Xbit_r190_c125 bl_125 br_125 wl_190 vdd gnd cell_6t
Xbit_r191_c125 bl_125 br_125 wl_191 vdd gnd cell_6t
Xbit_r192_c125 bl_125 br_125 wl_192 vdd gnd cell_6t
Xbit_r193_c125 bl_125 br_125 wl_193 vdd gnd cell_6t
Xbit_r194_c125 bl_125 br_125 wl_194 vdd gnd cell_6t
Xbit_r195_c125 bl_125 br_125 wl_195 vdd gnd cell_6t
Xbit_r196_c125 bl_125 br_125 wl_196 vdd gnd cell_6t
Xbit_r197_c125 bl_125 br_125 wl_197 vdd gnd cell_6t
Xbit_r198_c125 bl_125 br_125 wl_198 vdd gnd cell_6t
Xbit_r199_c125 bl_125 br_125 wl_199 vdd gnd cell_6t
Xbit_r200_c125 bl_125 br_125 wl_200 vdd gnd cell_6t
Xbit_r201_c125 bl_125 br_125 wl_201 vdd gnd cell_6t
Xbit_r202_c125 bl_125 br_125 wl_202 vdd gnd cell_6t
Xbit_r203_c125 bl_125 br_125 wl_203 vdd gnd cell_6t
Xbit_r204_c125 bl_125 br_125 wl_204 vdd gnd cell_6t
Xbit_r205_c125 bl_125 br_125 wl_205 vdd gnd cell_6t
Xbit_r206_c125 bl_125 br_125 wl_206 vdd gnd cell_6t
Xbit_r207_c125 bl_125 br_125 wl_207 vdd gnd cell_6t
Xbit_r208_c125 bl_125 br_125 wl_208 vdd gnd cell_6t
Xbit_r209_c125 bl_125 br_125 wl_209 vdd gnd cell_6t
Xbit_r210_c125 bl_125 br_125 wl_210 vdd gnd cell_6t
Xbit_r211_c125 bl_125 br_125 wl_211 vdd gnd cell_6t
Xbit_r212_c125 bl_125 br_125 wl_212 vdd gnd cell_6t
Xbit_r213_c125 bl_125 br_125 wl_213 vdd gnd cell_6t
Xbit_r214_c125 bl_125 br_125 wl_214 vdd gnd cell_6t
Xbit_r215_c125 bl_125 br_125 wl_215 vdd gnd cell_6t
Xbit_r216_c125 bl_125 br_125 wl_216 vdd gnd cell_6t
Xbit_r217_c125 bl_125 br_125 wl_217 vdd gnd cell_6t
Xbit_r218_c125 bl_125 br_125 wl_218 vdd gnd cell_6t
Xbit_r219_c125 bl_125 br_125 wl_219 vdd gnd cell_6t
Xbit_r220_c125 bl_125 br_125 wl_220 vdd gnd cell_6t
Xbit_r221_c125 bl_125 br_125 wl_221 vdd gnd cell_6t
Xbit_r222_c125 bl_125 br_125 wl_222 vdd gnd cell_6t
Xbit_r223_c125 bl_125 br_125 wl_223 vdd gnd cell_6t
Xbit_r224_c125 bl_125 br_125 wl_224 vdd gnd cell_6t
Xbit_r225_c125 bl_125 br_125 wl_225 vdd gnd cell_6t
Xbit_r226_c125 bl_125 br_125 wl_226 vdd gnd cell_6t
Xbit_r227_c125 bl_125 br_125 wl_227 vdd gnd cell_6t
Xbit_r228_c125 bl_125 br_125 wl_228 vdd gnd cell_6t
Xbit_r229_c125 bl_125 br_125 wl_229 vdd gnd cell_6t
Xbit_r230_c125 bl_125 br_125 wl_230 vdd gnd cell_6t
Xbit_r231_c125 bl_125 br_125 wl_231 vdd gnd cell_6t
Xbit_r232_c125 bl_125 br_125 wl_232 vdd gnd cell_6t
Xbit_r233_c125 bl_125 br_125 wl_233 vdd gnd cell_6t
Xbit_r234_c125 bl_125 br_125 wl_234 vdd gnd cell_6t
Xbit_r235_c125 bl_125 br_125 wl_235 vdd gnd cell_6t
Xbit_r236_c125 bl_125 br_125 wl_236 vdd gnd cell_6t
Xbit_r237_c125 bl_125 br_125 wl_237 vdd gnd cell_6t
Xbit_r238_c125 bl_125 br_125 wl_238 vdd gnd cell_6t
Xbit_r239_c125 bl_125 br_125 wl_239 vdd gnd cell_6t
Xbit_r240_c125 bl_125 br_125 wl_240 vdd gnd cell_6t
Xbit_r241_c125 bl_125 br_125 wl_241 vdd gnd cell_6t
Xbit_r242_c125 bl_125 br_125 wl_242 vdd gnd cell_6t
Xbit_r243_c125 bl_125 br_125 wl_243 vdd gnd cell_6t
Xbit_r244_c125 bl_125 br_125 wl_244 vdd gnd cell_6t
Xbit_r245_c125 bl_125 br_125 wl_245 vdd gnd cell_6t
Xbit_r246_c125 bl_125 br_125 wl_246 vdd gnd cell_6t
Xbit_r247_c125 bl_125 br_125 wl_247 vdd gnd cell_6t
Xbit_r248_c125 bl_125 br_125 wl_248 vdd gnd cell_6t
Xbit_r249_c125 bl_125 br_125 wl_249 vdd gnd cell_6t
Xbit_r250_c125 bl_125 br_125 wl_250 vdd gnd cell_6t
Xbit_r251_c125 bl_125 br_125 wl_251 vdd gnd cell_6t
Xbit_r252_c125 bl_125 br_125 wl_252 vdd gnd cell_6t
Xbit_r253_c125 bl_125 br_125 wl_253 vdd gnd cell_6t
Xbit_r254_c125 bl_125 br_125 wl_254 vdd gnd cell_6t
Xbit_r255_c125 bl_125 br_125 wl_255 vdd gnd cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd cell_6t
Xbit_r1_c126 bl_126 br_126 wl_1 vdd gnd cell_6t
Xbit_r2_c126 bl_126 br_126 wl_2 vdd gnd cell_6t
Xbit_r3_c126 bl_126 br_126 wl_3 vdd gnd cell_6t
Xbit_r4_c126 bl_126 br_126 wl_4 vdd gnd cell_6t
Xbit_r5_c126 bl_126 br_126 wl_5 vdd gnd cell_6t
Xbit_r6_c126 bl_126 br_126 wl_6 vdd gnd cell_6t
Xbit_r7_c126 bl_126 br_126 wl_7 vdd gnd cell_6t
Xbit_r8_c126 bl_126 br_126 wl_8 vdd gnd cell_6t
Xbit_r9_c126 bl_126 br_126 wl_9 vdd gnd cell_6t
Xbit_r10_c126 bl_126 br_126 wl_10 vdd gnd cell_6t
Xbit_r11_c126 bl_126 br_126 wl_11 vdd gnd cell_6t
Xbit_r12_c126 bl_126 br_126 wl_12 vdd gnd cell_6t
Xbit_r13_c126 bl_126 br_126 wl_13 vdd gnd cell_6t
Xbit_r14_c126 bl_126 br_126 wl_14 vdd gnd cell_6t
Xbit_r15_c126 bl_126 br_126 wl_15 vdd gnd cell_6t
Xbit_r16_c126 bl_126 br_126 wl_16 vdd gnd cell_6t
Xbit_r17_c126 bl_126 br_126 wl_17 vdd gnd cell_6t
Xbit_r18_c126 bl_126 br_126 wl_18 vdd gnd cell_6t
Xbit_r19_c126 bl_126 br_126 wl_19 vdd gnd cell_6t
Xbit_r20_c126 bl_126 br_126 wl_20 vdd gnd cell_6t
Xbit_r21_c126 bl_126 br_126 wl_21 vdd gnd cell_6t
Xbit_r22_c126 bl_126 br_126 wl_22 vdd gnd cell_6t
Xbit_r23_c126 bl_126 br_126 wl_23 vdd gnd cell_6t
Xbit_r24_c126 bl_126 br_126 wl_24 vdd gnd cell_6t
Xbit_r25_c126 bl_126 br_126 wl_25 vdd gnd cell_6t
Xbit_r26_c126 bl_126 br_126 wl_26 vdd gnd cell_6t
Xbit_r27_c126 bl_126 br_126 wl_27 vdd gnd cell_6t
Xbit_r28_c126 bl_126 br_126 wl_28 vdd gnd cell_6t
Xbit_r29_c126 bl_126 br_126 wl_29 vdd gnd cell_6t
Xbit_r30_c126 bl_126 br_126 wl_30 vdd gnd cell_6t
Xbit_r31_c126 bl_126 br_126 wl_31 vdd gnd cell_6t
Xbit_r32_c126 bl_126 br_126 wl_32 vdd gnd cell_6t
Xbit_r33_c126 bl_126 br_126 wl_33 vdd gnd cell_6t
Xbit_r34_c126 bl_126 br_126 wl_34 vdd gnd cell_6t
Xbit_r35_c126 bl_126 br_126 wl_35 vdd gnd cell_6t
Xbit_r36_c126 bl_126 br_126 wl_36 vdd gnd cell_6t
Xbit_r37_c126 bl_126 br_126 wl_37 vdd gnd cell_6t
Xbit_r38_c126 bl_126 br_126 wl_38 vdd gnd cell_6t
Xbit_r39_c126 bl_126 br_126 wl_39 vdd gnd cell_6t
Xbit_r40_c126 bl_126 br_126 wl_40 vdd gnd cell_6t
Xbit_r41_c126 bl_126 br_126 wl_41 vdd gnd cell_6t
Xbit_r42_c126 bl_126 br_126 wl_42 vdd gnd cell_6t
Xbit_r43_c126 bl_126 br_126 wl_43 vdd gnd cell_6t
Xbit_r44_c126 bl_126 br_126 wl_44 vdd gnd cell_6t
Xbit_r45_c126 bl_126 br_126 wl_45 vdd gnd cell_6t
Xbit_r46_c126 bl_126 br_126 wl_46 vdd gnd cell_6t
Xbit_r47_c126 bl_126 br_126 wl_47 vdd gnd cell_6t
Xbit_r48_c126 bl_126 br_126 wl_48 vdd gnd cell_6t
Xbit_r49_c126 bl_126 br_126 wl_49 vdd gnd cell_6t
Xbit_r50_c126 bl_126 br_126 wl_50 vdd gnd cell_6t
Xbit_r51_c126 bl_126 br_126 wl_51 vdd gnd cell_6t
Xbit_r52_c126 bl_126 br_126 wl_52 vdd gnd cell_6t
Xbit_r53_c126 bl_126 br_126 wl_53 vdd gnd cell_6t
Xbit_r54_c126 bl_126 br_126 wl_54 vdd gnd cell_6t
Xbit_r55_c126 bl_126 br_126 wl_55 vdd gnd cell_6t
Xbit_r56_c126 bl_126 br_126 wl_56 vdd gnd cell_6t
Xbit_r57_c126 bl_126 br_126 wl_57 vdd gnd cell_6t
Xbit_r58_c126 bl_126 br_126 wl_58 vdd gnd cell_6t
Xbit_r59_c126 bl_126 br_126 wl_59 vdd gnd cell_6t
Xbit_r60_c126 bl_126 br_126 wl_60 vdd gnd cell_6t
Xbit_r61_c126 bl_126 br_126 wl_61 vdd gnd cell_6t
Xbit_r62_c126 bl_126 br_126 wl_62 vdd gnd cell_6t
Xbit_r63_c126 bl_126 br_126 wl_63 vdd gnd cell_6t
Xbit_r64_c126 bl_126 br_126 wl_64 vdd gnd cell_6t
Xbit_r65_c126 bl_126 br_126 wl_65 vdd gnd cell_6t
Xbit_r66_c126 bl_126 br_126 wl_66 vdd gnd cell_6t
Xbit_r67_c126 bl_126 br_126 wl_67 vdd gnd cell_6t
Xbit_r68_c126 bl_126 br_126 wl_68 vdd gnd cell_6t
Xbit_r69_c126 bl_126 br_126 wl_69 vdd gnd cell_6t
Xbit_r70_c126 bl_126 br_126 wl_70 vdd gnd cell_6t
Xbit_r71_c126 bl_126 br_126 wl_71 vdd gnd cell_6t
Xbit_r72_c126 bl_126 br_126 wl_72 vdd gnd cell_6t
Xbit_r73_c126 bl_126 br_126 wl_73 vdd gnd cell_6t
Xbit_r74_c126 bl_126 br_126 wl_74 vdd gnd cell_6t
Xbit_r75_c126 bl_126 br_126 wl_75 vdd gnd cell_6t
Xbit_r76_c126 bl_126 br_126 wl_76 vdd gnd cell_6t
Xbit_r77_c126 bl_126 br_126 wl_77 vdd gnd cell_6t
Xbit_r78_c126 bl_126 br_126 wl_78 vdd gnd cell_6t
Xbit_r79_c126 bl_126 br_126 wl_79 vdd gnd cell_6t
Xbit_r80_c126 bl_126 br_126 wl_80 vdd gnd cell_6t
Xbit_r81_c126 bl_126 br_126 wl_81 vdd gnd cell_6t
Xbit_r82_c126 bl_126 br_126 wl_82 vdd gnd cell_6t
Xbit_r83_c126 bl_126 br_126 wl_83 vdd gnd cell_6t
Xbit_r84_c126 bl_126 br_126 wl_84 vdd gnd cell_6t
Xbit_r85_c126 bl_126 br_126 wl_85 vdd gnd cell_6t
Xbit_r86_c126 bl_126 br_126 wl_86 vdd gnd cell_6t
Xbit_r87_c126 bl_126 br_126 wl_87 vdd gnd cell_6t
Xbit_r88_c126 bl_126 br_126 wl_88 vdd gnd cell_6t
Xbit_r89_c126 bl_126 br_126 wl_89 vdd gnd cell_6t
Xbit_r90_c126 bl_126 br_126 wl_90 vdd gnd cell_6t
Xbit_r91_c126 bl_126 br_126 wl_91 vdd gnd cell_6t
Xbit_r92_c126 bl_126 br_126 wl_92 vdd gnd cell_6t
Xbit_r93_c126 bl_126 br_126 wl_93 vdd gnd cell_6t
Xbit_r94_c126 bl_126 br_126 wl_94 vdd gnd cell_6t
Xbit_r95_c126 bl_126 br_126 wl_95 vdd gnd cell_6t
Xbit_r96_c126 bl_126 br_126 wl_96 vdd gnd cell_6t
Xbit_r97_c126 bl_126 br_126 wl_97 vdd gnd cell_6t
Xbit_r98_c126 bl_126 br_126 wl_98 vdd gnd cell_6t
Xbit_r99_c126 bl_126 br_126 wl_99 vdd gnd cell_6t
Xbit_r100_c126 bl_126 br_126 wl_100 vdd gnd cell_6t
Xbit_r101_c126 bl_126 br_126 wl_101 vdd gnd cell_6t
Xbit_r102_c126 bl_126 br_126 wl_102 vdd gnd cell_6t
Xbit_r103_c126 bl_126 br_126 wl_103 vdd gnd cell_6t
Xbit_r104_c126 bl_126 br_126 wl_104 vdd gnd cell_6t
Xbit_r105_c126 bl_126 br_126 wl_105 vdd gnd cell_6t
Xbit_r106_c126 bl_126 br_126 wl_106 vdd gnd cell_6t
Xbit_r107_c126 bl_126 br_126 wl_107 vdd gnd cell_6t
Xbit_r108_c126 bl_126 br_126 wl_108 vdd gnd cell_6t
Xbit_r109_c126 bl_126 br_126 wl_109 vdd gnd cell_6t
Xbit_r110_c126 bl_126 br_126 wl_110 vdd gnd cell_6t
Xbit_r111_c126 bl_126 br_126 wl_111 vdd gnd cell_6t
Xbit_r112_c126 bl_126 br_126 wl_112 vdd gnd cell_6t
Xbit_r113_c126 bl_126 br_126 wl_113 vdd gnd cell_6t
Xbit_r114_c126 bl_126 br_126 wl_114 vdd gnd cell_6t
Xbit_r115_c126 bl_126 br_126 wl_115 vdd gnd cell_6t
Xbit_r116_c126 bl_126 br_126 wl_116 vdd gnd cell_6t
Xbit_r117_c126 bl_126 br_126 wl_117 vdd gnd cell_6t
Xbit_r118_c126 bl_126 br_126 wl_118 vdd gnd cell_6t
Xbit_r119_c126 bl_126 br_126 wl_119 vdd gnd cell_6t
Xbit_r120_c126 bl_126 br_126 wl_120 vdd gnd cell_6t
Xbit_r121_c126 bl_126 br_126 wl_121 vdd gnd cell_6t
Xbit_r122_c126 bl_126 br_126 wl_122 vdd gnd cell_6t
Xbit_r123_c126 bl_126 br_126 wl_123 vdd gnd cell_6t
Xbit_r124_c126 bl_126 br_126 wl_124 vdd gnd cell_6t
Xbit_r125_c126 bl_126 br_126 wl_125 vdd gnd cell_6t
Xbit_r126_c126 bl_126 br_126 wl_126 vdd gnd cell_6t
Xbit_r127_c126 bl_126 br_126 wl_127 vdd gnd cell_6t
Xbit_r128_c126 bl_126 br_126 wl_128 vdd gnd cell_6t
Xbit_r129_c126 bl_126 br_126 wl_129 vdd gnd cell_6t
Xbit_r130_c126 bl_126 br_126 wl_130 vdd gnd cell_6t
Xbit_r131_c126 bl_126 br_126 wl_131 vdd gnd cell_6t
Xbit_r132_c126 bl_126 br_126 wl_132 vdd gnd cell_6t
Xbit_r133_c126 bl_126 br_126 wl_133 vdd gnd cell_6t
Xbit_r134_c126 bl_126 br_126 wl_134 vdd gnd cell_6t
Xbit_r135_c126 bl_126 br_126 wl_135 vdd gnd cell_6t
Xbit_r136_c126 bl_126 br_126 wl_136 vdd gnd cell_6t
Xbit_r137_c126 bl_126 br_126 wl_137 vdd gnd cell_6t
Xbit_r138_c126 bl_126 br_126 wl_138 vdd gnd cell_6t
Xbit_r139_c126 bl_126 br_126 wl_139 vdd gnd cell_6t
Xbit_r140_c126 bl_126 br_126 wl_140 vdd gnd cell_6t
Xbit_r141_c126 bl_126 br_126 wl_141 vdd gnd cell_6t
Xbit_r142_c126 bl_126 br_126 wl_142 vdd gnd cell_6t
Xbit_r143_c126 bl_126 br_126 wl_143 vdd gnd cell_6t
Xbit_r144_c126 bl_126 br_126 wl_144 vdd gnd cell_6t
Xbit_r145_c126 bl_126 br_126 wl_145 vdd gnd cell_6t
Xbit_r146_c126 bl_126 br_126 wl_146 vdd gnd cell_6t
Xbit_r147_c126 bl_126 br_126 wl_147 vdd gnd cell_6t
Xbit_r148_c126 bl_126 br_126 wl_148 vdd gnd cell_6t
Xbit_r149_c126 bl_126 br_126 wl_149 vdd gnd cell_6t
Xbit_r150_c126 bl_126 br_126 wl_150 vdd gnd cell_6t
Xbit_r151_c126 bl_126 br_126 wl_151 vdd gnd cell_6t
Xbit_r152_c126 bl_126 br_126 wl_152 vdd gnd cell_6t
Xbit_r153_c126 bl_126 br_126 wl_153 vdd gnd cell_6t
Xbit_r154_c126 bl_126 br_126 wl_154 vdd gnd cell_6t
Xbit_r155_c126 bl_126 br_126 wl_155 vdd gnd cell_6t
Xbit_r156_c126 bl_126 br_126 wl_156 vdd gnd cell_6t
Xbit_r157_c126 bl_126 br_126 wl_157 vdd gnd cell_6t
Xbit_r158_c126 bl_126 br_126 wl_158 vdd gnd cell_6t
Xbit_r159_c126 bl_126 br_126 wl_159 vdd gnd cell_6t
Xbit_r160_c126 bl_126 br_126 wl_160 vdd gnd cell_6t
Xbit_r161_c126 bl_126 br_126 wl_161 vdd gnd cell_6t
Xbit_r162_c126 bl_126 br_126 wl_162 vdd gnd cell_6t
Xbit_r163_c126 bl_126 br_126 wl_163 vdd gnd cell_6t
Xbit_r164_c126 bl_126 br_126 wl_164 vdd gnd cell_6t
Xbit_r165_c126 bl_126 br_126 wl_165 vdd gnd cell_6t
Xbit_r166_c126 bl_126 br_126 wl_166 vdd gnd cell_6t
Xbit_r167_c126 bl_126 br_126 wl_167 vdd gnd cell_6t
Xbit_r168_c126 bl_126 br_126 wl_168 vdd gnd cell_6t
Xbit_r169_c126 bl_126 br_126 wl_169 vdd gnd cell_6t
Xbit_r170_c126 bl_126 br_126 wl_170 vdd gnd cell_6t
Xbit_r171_c126 bl_126 br_126 wl_171 vdd gnd cell_6t
Xbit_r172_c126 bl_126 br_126 wl_172 vdd gnd cell_6t
Xbit_r173_c126 bl_126 br_126 wl_173 vdd gnd cell_6t
Xbit_r174_c126 bl_126 br_126 wl_174 vdd gnd cell_6t
Xbit_r175_c126 bl_126 br_126 wl_175 vdd gnd cell_6t
Xbit_r176_c126 bl_126 br_126 wl_176 vdd gnd cell_6t
Xbit_r177_c126 bl_126 br_126 wl_177 vdd gnd cell_6t
Xbit_r178_c126 bl_126 br_126 wl_178 vdd gnd cell_6t
Xbit_r179_c126 bl_126 br_126 wl_179 vdd gnd cell_6t
Xbit_r180_c126 bl_126 br_126 wl_180 vdd gnd cell_6t
Xbit_r181_c126 bl_126 br_126 wl_181 vdd gnd cell_6t
Xbit_r182_c126 bl_126 br_126 wl_182 vdd gnd cell_6t
Xbit_r183_c126 bl_126 br_126 wl_183 vdd gnd cell_6t
Xbit_r184_c126 bl_126 br_126 wl_184 vdd gnd cell_6t
Xbit_r185_c126 bl_126 br_126 wl_185 vdd gnd cell_6t
Xbit_r186_c126 bl_126 br_126 wl_186 vdd gnd cell_6t
Xbit_r187_c126 bl_126 br_126 wl_187 vdd gnd cell_6t
Xbit_r188_c126 bl_126 br_126 wl_188 vdd gnd cell_6t
Xbit_r189_c126 bl_126 br_126 wl_189 vdd gnd cell_6t
Xbit_r190_c126 bl_126 br_126 wl_190 vdd gnd cell_6t
Xbit_r191_c126 bl_126 br_126 wl_191 vdd gnd cell_6t
Xbit_r192_c126 bl_126 br_126 wl_192 vdd gnd cell_6t
Xbit_r193_c126 bl_126 br_126 wl_193 vdd gnd cell_6t
Xbit_r194_c126 bl_126 br_126 wl_194 vdd gnd cell_6t
Xbit_r195_c126 bl_126 br_126 wl_195 vdd gnd cell_6t
Xbit_r196_c126 bl_126 br_126 wl_196 vdd gnd cell_6t
Xbit_r197_c126 bl_126 br_126 wl_197 vdd gnd cell_6t
Xbit_r198_c126 bl_126 br_126 wl_198 vdd gnd cell_6t
Xbit_r199_c126 bl_126 br_126 wl_199 vdd gnd cell_6t
Xbit_r200_c126 bl_126 br_126 wl_200 vdd gnd cell_6t
Xbit_r201_c126 bl_126 br_126 wl_201 vdd gnd cell_6t
Xbit_r202_c126 bl_126 br_126 wl_202 vdd gnd cell_6t
Xbit_r203_c126 bl_126 br_126 wl_203 vdd gnd cell_6t
Xbit_r204_c126 bl_126 br_126 wl_204 vdd gnd cell_6t
Xbit_r205_c126 bl_126 br_126 wl_205 vdd gnd cell_6t
Xbit_r206_c126 bl_126 br_126 wl_206 vdd gnd cell_6t
Xbit_r207_c126 bl_126 br_126 wl_207 vdd gnd cell_6t
Xbit_r208_c126 bl_126 br_126 wl_208 vdd gnd cell_6t
Xbit_r209_c126 bl_126 br_126 wl_209 vdd gnd cell_6t
Xbit_r210_c126 bl_126 br_126 wl_210 vdd gnd cell_6t
Xbit_r211_c126 bl_126 br_126 wl_211 vdd gnd cell_6t
Xbit_r212_c126 bl_126 br_126 wl_212 vdd gnd cell_6t
Xbit_r213_c126 bl_126 br_126 wl_213 vdd gnd cell_6t
Xbit_r214_c126 bl_126 br_126 wl_214 vdd gnd cell_6t
Xbit_r215_c126 bl_126 br_126 wl_215 vdd gnd cell_6t
Xbit_r216_c126 bl_126 br_126 wl_216 vdd gnd cell_6t
Xbit_r217_c126 bl_126 br_126 wl_217 vdd gnd cell_6t
Xbit_r218_c126 bl_126 br_126 wl_218 vdd gnd cell_6t
Xbit_r219_c126 bl_126 br_126 wl_219 vdd gnd cell_6t
Xbit_r220_c126 bl_126 br_126 wl_220 vdd gnd cell_6t
Xbit_r221_c126 bl_126 br_126 wl_221 vdd gnd cell_6t
Xbit_r222_c126 bl_126 br_126 wl_222 vdd gnd cell_6t
Xbit_r223_c126 bl_126 br_126 wl_223 vdd gnd cell_6t
Xbit_r224_c126 bl_126 br_126 wl_224 vdd gnd cell_6t
Xbit_r225_c126 bl_126 br_126 wl_225 vdd gnd cell_6t
Xbit_r226_c126 bl_126 br_126 wl_226 vdd gnd cell_6t
Xbit_r227_c126 bl_126 br_126 wl_227 vdd gnd cell_6t
Xbit_r228_c126 bl_126 br_126 wl_228 vdd gnd cell_6t
Xbit_r229_c126 bl_126 br_126 wl_229 vdd gnd cell_6t
Xbit_r230_c126 bl_126 br_126 wl_230 vdd gnd cell_6t
Xbit_r231_c126 bl_126 br_126 wl_231 vdd gnd cell_6t
Xbit_r232_c126 bl_126 br_126 wl_232 vdd gnd cell_6t
Xbit_r233_c126 bl_126 br_126 wl_233 vdd gnd cell_6t
Xbit_r234_c126 bl_126 br_126 wl_234 vdd gnd cell_6t
Xbit_r235_c126 bl_126 br_126 wl_235 vdd gnd cell_6t
Xbit_r236_c126 bl_126 br_126 wl_236 vdd gnd cell_6t
Xbit_r237_c126 bl_126 br_126 wl_237 vdd gnd cell_6t
Xbit_r238_c126 bl_126 br_126 wl_238 vdd gnd cell_6t
Xbit_r239_c126 bl_126 br_126 wl_239 vdd gnd cell_6t
Xbit_r240_c126 bl_126 br_126 wl_240 vdd gnd cell_6t
Xbit_r241_c126 bl_126 br_126 wl_241 vdd gnd cell_6t
Xbit_r242_c126 bl_126 br_126 wl_242 vdd gnd cell_6t
Xbit_r243_c126 bl_126 br_126 wl_243 vdd gnd cell_6t
Xbit_r244_c126 bl_126 br_126 wl_244 vdd gnd cell_6t
Xbit_r245_c126 bl_126 br_126 wl_245 vdd gnd cell_6t
Xbit_r246_c126 bl_126 br_126 wl_246 vdd gnd cell_6t
Xbit_r247_c126 bl_126 br_126 wl_247 vdd gnd cell_6t
Xbit_r248_c126 bl_126 br_126 wl_248 vdd gnd cell_6t
Xbit_r249_c126 bl_126 br_126 wl_249 vdd gnd cell_6t
Xbit_r250_c126 bl_126 br_126 wl_250 vdd gnd cell_6t
Xbit_r251_c126 bl_126 br_126 wl_251 vdd gnd cell_6t
Xbit_r252_c126 bl_126 br_126 wl_252 vdd gnd cell_6t
Xbit_r253_c126 bl_126 br_126 wl_253 vdd gnd cell_6t
Xbit_r254_c126 bl_126 br_126 wl_254 vdd gnd cell_6t
Xbit_r255_c126 bl_126 br_126 wl_255 vdd gnd cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd cell_6t
Xbit_r1_c127 bl_127 br_127 wl_1 vdd gnd cell_6t
Xbit_r2_c127 bl_127 br_127 wl_2 vdd gnd cell_6t
Xbit_r3_c127 bl_127 br_127 wl_3 vdd gnd cell_6t
Xbit_r4_c127 bl_127 br_127 wl_4 vdd gnd cell_6t
Xbit_r5_c127 bl_127 br_127 wl_5 vdd gnd cell_6t
Xbit_r6_c127 bl_127 br_127 wl_6 vdd gnd cell_6t
Xbit_r7_c127 bl_127 br_127 wl_7 vdd gnd cell_6t
Xbit_r8_c127 bl_127 br_127 wl_8 vdd gnd cell_6t
Xbit_r9_c127 bl_127 br_127 wl_9 vdd gnd cell_6t
Xbit_r10_c127 bl_127 br_127 wl_10 vdd gnd cell_6t
Xbit_r11_c127 bl_127 br_127 wl_11 vdd gnd cell_6t
Xbit_r12_c127 bl_127 br_127 wl_12 vdd gnd cell_6t
Xbit_r13_c127 bl_127 br_127 wl_13 vdd gnd cell_6t
Xbit_r14_c127 bl_127 br_127 wl_14 vdd gnd cell_6t
Xbit_r15_c127 bl_127 br_127 wl_15 vdd gnd cell_6t
Xbit_r16_c127 bl_127 br_127 wl_16 vdd gnd cell_6t
Xbit_r17_c127 bl_127 br_127 wl_17 vdd gnd cell_6t
Xbit_r18_c127 bl_127 br_127 wl_18 vdd gnd cell_6t
Xbit_r19_c127 bl_127 br_127 wl_19 vdd gnd cell_6t
Xbit_r20_c127 bl_127 br_127 wl_20 vdd gnd cell_6t
Xbit_r21_c127 bl_127 br_127 wl_21 vdd gnd cell_6t
Xbit_r22_c127 bl_127 br_127 wl_22 vdd gnd cell_6t
Xbit_r23_c127 bl_127 br_127 wl_23 vdd gnd cell_6t
Xbit_r24_c127 bl_127 br_127 wl_24 vdd gnd cell_6t
Xbit_r25_c127 bl_127 br_127 wl_25 vdd gnd cell_6t
Xbit_r26_c127 bl_127 br_127 wl_26 vdd gnd cell_6t
Xbit_r27_c127 bl_127 br_127 wl_27 vdd gnd cell_6t
Xbit_r28_c127 bl_127 br_127 wl_28 vdd gnd cell_6t
Xbit_r29_c127 bl_127 br_127 wl_29 vdd gnd cell_6t
Xbit_r30_c127 bl_127 br_127 wl_30 vdd gnd cell_6t
Xbit_r31_c127 bl_127 br_127 wl_31 vdd gnd cell_6t
Xbit_r32_c127 bl_127 br_127 wl_32 vdd gnd cell_6t
Xbit_r33_c127 bl_127 br_127 wl_33 vdd gnd cell_6t
Xbit_r34_c127 bl_127 br_127 wl_34 vdd gnd cell_6t
Xbit_r35_c127 bl_127 br_127 wl_35 vdd gnd cell_6t
Xbit_r36_c127 bl_127 br_127 wl_36 vdd gnd cell_6t
Xbit_r37_c127 bl_127 br_127 wl_37 vdd gnd cell_6t
Xbit_r38_c127 bl_127 br_127 wl_38 vdd gnd cell_6t
Xbit_r39_c127 bl_127 br_127 wl_39 vdd gnd cell_6t
Xbit_r40_c127 bl_127 br_127 wl_40 vdd gnd cell_6t
Xbit_r41_c127 bl_127 br_127 wl_41 vdd gnd cell_6t
Xbit_r42_c127 bl_127 br_127 wl_42 vdd gnd cell_6t
Xbit_r43_c127 bl_127 br_127 wl_43 vdd gnd cell_6t
Xbit_r44_c127 bl_127 br_127 wl_44 vdd gnd cell_6t
Xbit_r45_c127 bl_127 br_127 wl_45 vdd gnd cell_6t
Xbit_r46_c127 bl_127 br_127 wl_46 vdd gnd cell_6t
Xbit_r47_c127 bl_127 br_127 wl_47 vdd gnd cell_6t
Xbit_r48_c127 bl_127 br_127 wl_48 vdd gnd cell_6t
Xbit_r49_c127 bl_127 br_127 wl_49 vdd gnd cell_6t
Xbit_r50_c127 bl_127 br_127 wl_50 vdd gnd cell_6t
Xbit_r51_c127 bl_127 br_127 wl_51 vdd gnd cell_6t
Xbit_r52_c127 bl_127 br_127 wl_52 vdd gnd cell_6t
Xbit_r53_c127 bl_127 br_127 wl_53 vdd gnd cell_6t
Xbit_r54_c127 bl_127 br_127 wl_54 vdd gnd cell_6t
Xbit_r55_c127 bl_127 br_127 wl_55 vdd gnd cell_6t
Xbit_r56_c127 bl_127 br_127 wl_56 vdd gnd cell_6t
Xbit_r57_c127 bl_127 br_127 wl_57 vdd gnd cell_6t
Xbit_r58_c127 bl_127 br_127 wl_58 vdd gnd cell_6t
Xbit_r59_c127 bl_127 br_127 wl_59 vdd gnd cell_6t
Xbit_r60_c127 bl_127 br_127 wl_60 vdd gnd cell_6t
Xbit_r61_c127 bl_127 br_127 wl_61 vdd gnd cell_6t
Xbit_r62_c127 bl_127 br_127 wl_62 vdd gnd cell_6t
Xbit_r63_c127 bl_127 br_127 wl_63 vdd gnd cell_6t
Xbit_r64_c127 bl_127 br_127 wl_64 vdd gnd cell_6t
Xbit_r65_c127 bl_127 br_127 wl_65 vdd gnd cell_6t
Xbit_r66_c127 bl_127 br_127 wl_66 vdd gnd cell_6t
Xbit_r67_c127 bl_127 br_127 wl_67 vdd gnd cell_6t
Xbit_r68_c127 bl_127 br_127 wl_68 vdd gnd cell_6t
Xbit_r69_c127 bl_127 br_127 wl_69 vdd gnd cell_6t
Xbit_r70_c127 bl_127 br_127 wl_70 vdd gnd cell_6t
Xbit_r71_c127 bl_127 br_127 wl_71 vdd gnd cell_6t
Xbit_r72_c127 bl_127 br_127 wl_72 vdd gnd cell_6t
Xbit_r73_c127 bl_127 br_127 wl_73 vdd gnd cell_6t
Xbit_r74_c127 bl_127 br_127 wl_74 vdd gnd cell_6t
Xbit_r75_c127 bl_127 br_127 wl_75 vdd gnd cell_6t
Xbit_r76_c127 bl_127 br_127 wl_76 vdd gnd cell_6t
Xbit_r77_c127 bl_127 br_127 wl_77 vdd gnd cell_6t
Xbit_r78_c127 bl_127 br_127 wl_78 vdd gnd cell_6t
Xbit_r79_c127 bl_127 br_127 wl_79 vdd gnd cell_6t
Xbit_r80_c127 bl_127 br_127 wl_80 vdd gnd cell_6t
Xbit_r81_c127 bl_127 br_127 wl_81 vdd gnd cell_6t
Xbit_r82_c127 bl_127 br_127 wl_82 vdd gnd cell_6t
Xbit_r83_c127 bl_127 br_127 wl_83 vdd gnd cell_6t
Xbit_r84_c127 bl_127 br_127 wl_84 vdd gnd cell_6t
Xbit_r85_c127 bl_127 br_127 wl_85 vdd gnd cell_6t
Xbit_r86_c127 bl_127 br_127 wl_86 vdd gnd cell_6t
Xbit_r87_c127 bl_127 br_127 wl_87 vdd gnd cell_6t
Xbit_r88_c127 bl_127 br_127 wl_88 vdd gnd cell_6t
Xbit_r89_c127 bl_127 br_127 wl_89 vdd gnd cell_6t
Xbit_r90_c127 bl_127 br_127 wl_90 vdd gnd cell_6t
Xbit_r91_c127 bl_127 br_127 wl_91 vdd gnd cell_6t
Xbit_r92_c127 bl_127 br_127 wl_92 vdd gnd cell_6t
Xbit_r93_c127 bl_127 br_127 wl_93 vdd gnd cell_6t
Xbit_r94_c127 bl_127 br_127 wl_94 vdd gnd cell_6t
Xbit_r95_c127 bl_127 br_127 wl_95 vdd gnd cell_6t
Xbit_r96_c127 bl_127 br_127 wl_96 vdd gnd cell_6t
Xbit_r97_c127 bl_127 br_127 wl_97 vdd gnd cell_6t
Xbit_r98_c127 bl_127 br_127 wl_98 vdd gnd cell_6t
Xbit_r99_c127 bl_127 br_127 wl_99 vdd gnd cell_6t
Xbit_r100_c127 bl_127 br_127 wl_100 vdd gnd cell_6t
Xbit_r101_c127 bl_127 br_127 wl_101 vdd gnd cell_6t
Xbit_r102_c127 bl_127 br_127 wl_102 vdd gnd cell_6t
Xbit_r103_c127 bl_127 br_127 wl_103 vdd gnd cell_6t
Xbit_r104_c127 bl_127 br_127 wl_104 vdd gnd cell_6t
Xbit_r105_c127 bl_127 br_127 wl_105 vdd gnd cell_6t
Xbit_r106_c127 bl_127 br_127 wl_106 vdd gnd cell_6t
Xbit_r107_c127 bl_127 br_127 wl_107 vdd gnd cell_6t
Xbit_r108_c127 bl_127 br_127 wl_108 vdd gnd cell_6t
Xbit_r109_c127 bl_127 br_127 wl_109 vdd gnd cell_6t
Xbit_r110_c127 bl_127 br_127 wl_110 vdd gnd cell_6t
Xbit_r111_c127 bl_127 br_127 wl_111 vdd gnd cell_6t
Xbit_r112_c127 bl_127 br_127 wl_112 vdd gnd cell_6t
Xbit_r113_c127 bl_127 br_127 wl_113 vdd gnd cell_6t
Xbit_r114_c127 bl_127 br_127 wl_114 vdd gnd cell_6t
Xbit_r115_c127 bl_127 br_127 wl_115 vdd gnd cell_6t
Xbit_r116_c127 bl_127 br_127 wl_116 vdd gnd cell_6t
Xbit_r117_c127 bl_127 br_127 wl_117 vdd gnd cell_6t
Xbit_r118_c127 bl_127 br_127 wl_118 vdd gnd cell_6t
Xbit_r119_c127 bl_127 br_127 wl_119 vdd gnd cell_6t
Xbit_r120_c127 bl_127 br_127 wl_120 vdd gnd cell_6t
Xbit_r121_c127 bl_127 br_127 wl_121 vdd gnd cell_6t
Xbit_r122_c127 bl_127 br_127 wl_122 vdd gnd cell_6t
Xbit_r123_c127 bl_127 br_127 wl_123 vdd gnd cell_6t
Xbit_r124_c127 bl_127 br_127 wl_124 vdd gnd cell_6t
Xbit_r125_c127 bl_127 br_127 wl_125 vdd gnd cell_6t
Xbit_r126_c127 bl_127 br_127 wl_126 vdd gnd cell_6t
Xbit_r127_c127 bl_127 br_127 wl_127 vdd gnd cell_6t
Xbit_r128_c127 bl_127 br_127 wl_128 vdd gnd cell_6t
Xbit_r129_c127 bl_127 br_127 wl_129 vdd gnd cell_6t
Xbit_r130_c127 bl_127 br_127 wl_130 vdd gnd cell_6t
Xbit_r131_c127 bl_127 br_127 wl_131 vdd gnd cell_6t
Xbit_r132_c127 bl_127 br_127 wl_132 vdd gnd cell_6t
Xbit_r133_c127 bl_127 br_127 wl_133 vdd gnd cell_6t
Xbit_r134_c127 bl_127 br_127 wl_134 vdd gnd cell_6t
Xbit_r135_c127 bl_127 br_127 wl_135 vdd gnd cell_6t
Xbit_r136_c127 bl_127 br_127 wl_136 vdd gnd cell_6t
Xbit_r137_c127 bl_127 br_127 wl_137 vdd gnd cell_6t
Xbit_r138_c127 bl_127 br_127 wl_138 vdd gnd cell_6t
Xbit_r139_c127 bl_127 br_127 wl_139 vdd gnd cell_6t
Xbit_r140_c127 bl_127 br_127 wl_140 vdd gnd cell_6t
Xbit_r141_c127 bl_127 br_127 wl_141 vdd gnd cell_6t
Xbit_r142_c127 bl_127 br_127 wl_142 vdd gnd cell_6t
Xbit_r143_c127 bl_127 br_127 wl_143 vdd gnd cell_6t
Xbit_r144_c127 bl_127 br_127 wl_144 vdd gnd cell_6t
Xbit_r145_c127 bl_127 br_127 wl_145 vdd gnd cell_6t
Xbit_r146_c127 bl_127 br_127 wl_146 vdd gnd cell_6t
Xbit_r147_c127 bl_127 br_127 wl_147 vdd gnd cell_6t
Xbit_r148_c127 bl_127 br_127 wl_148 vdd gnd cell_6t
Xbit_r149_c127 bl_127 br_127 wl_149 vdd gnd cell_6t
Xbit_r150_c127 bl_127 br_127 wl_150 vdd gnd cell_6t
Xbit_r151_c127 bl_127 br_127 wl_151 vdd gnd cell_6t
Xbit_r152_c127 bl_127 br_127 wl_152 vdd gnd cell_6t
Xbit_r153_c127 bl_127 br_127 wl_153 vdd gnd cell_6t
Xbit_r154_c127 bl_127 br_127 wl_154 vdd gnd cell_6t
Xbit_r155_c127 bl_127 br_127 wl_155 vdd gnd cell_6t
Xbit_r156_c127 bl_127 br_127 wl_156 vdd gnd cell_6t
Xbit_r157_c127 bl_127 br_127 wl_157 vdd gnd cell_6t
Xbit_r158_c127 bl_127 br_127 wl_158 vdd gnd cell_6t
Xbit_r159_c127 bl_127 br_127 wl_159 vdd gnd cell_6t
Xbit_r160_c127 bl_127 br_127 wl_160 vdd gnd cell_6t
Xbit_r161_c127 bl_127 br_127 wl_161 vdd gnd cell_6t
Xbit_r162_c127 bl_127 br_127 wl_162 vdd gnd cell_6t
Xbit_r163_c127 bl_127 br_127 wl_163 vdd gnd cell_6t
Xbit_r164_c127 bl_127 br_127 wl_164 vdd gnd cell_6t
Xbit_r165_c127 bl_127 br_127 wl_165 vdd gnd cell_6t
Xbit_r166_c127 bl_127 br_127 wl_166 vdd gnd cell_6t
Xbit_r167_c127 bl_127 br_127 wl_167 vdd gnd cell_6t
Xbit_r168_c127 bl_127 br_127 wl_168 vdd gnd cell_6t
Xbit_r169_c127 bl_127 br_127 wl_169 vdd gnd cell_6t
Xbit_r170_c127 bl_127 br_127 wl_170 vdd gnd cell_6t
Xbit_r171_c127 bl_127 br_127 wl_171 vdd gnd cell_6t
Xbit_r172_c127 bl_127 br_127 wl_172 vdd gnd cell_6t
Xbit_r173_c127 bl_127 br_127 wl_173 vdd gnd cell_6t
Xbit_r174_c127 bl_127 br_127 wl_174 vdd gnd cell_6t
Xbit_r175_c127 bl_127 br_127 wl_175 vdd gnd cell_6t
Xbit_r176_c127 bl_127 br_127 wl_176 vdd gnd cell_6t
Xbit_r177_c127 bl_127 br_127 wl_177 vdd gnd cell_6t
Xbit_r178_c127 bl_127 br_127 wl_178 vdd gnd cell_6t
Xbit_r179_c127 bl_127 br_127 wl_179 vdd gnd cell_6t
Xbit_r180_c127 bl_127 br_127 wl_180 vdd gnd cell_6t
Xbit_r181_c127 bl_127 br_127 wl_181 vdd gnd cell_6t
Xbit_r182_c127 bl_127 br_127 wl_182 vdd gnd cell_6t
Xbit_r183_c127 bl_127 br_127 wl_183 vdd gnd cell_6t
Xbit_r184_c127 bl_127 br_127 wl_184 vdd gnd cell_6t
Xbit_r185_c127 bl_127 br_127 wl_185 vdd gnd cell_6t
Xbit_r186_c127 bl_127 br_127 wl_186 vdd gnd cell_6t
Xbit_r187_c127 bl_127 br_127 wl_187 vdd gnd cell_6t
Xbit_r188_c127 bl_127 br_127 wl_188 vdd gnd cell_6t
Xbit_r189_c127 bl_127 br_127 wl_189 vdd gnd cell_6t
Xbit_r190_c127 bl_127 br_127 wl_190 vdd gnd cell_6t
Xbit_r191_c127 bl_127 br_127 wl_191 vdd gnd cell_6t
Xbit_r192_c127 bl_127 br_127 wl_192 vdd gnd cell_6t
Xbit_r193_c127 bl_127 br_127 wl_193 vdd gnd cell_6t
Xbit_r194_c127 bl_127 br_127 wl_194 vdd gnd cell_6t
Xbit_r195_c127 bl_127 br_127 wl_195 vdd gnd cell_6t
Xbit_r196_c127 bl_127 br_127 wl_196 vdd gnd cell_6t
Xbit_r197_c127 bl_127 br_127 wl_197 vdd gnd cell_6t
Xbit_r198_c127 bl_127 br_127 wl_198 vdd gnd cell_6t
Xbit_r199_c127 bl_127 br_127 wl_199 vdd gnd cell_6t
Xbit_r200_c127 bl_127 br_127 wl_200 vdd gnd cell_6t
Xbit_r201_c127 bl_127 br_127 wl_201 vdd gnd cell_6t
Xbit_r202_c127 bl_127 br_127 wl_202 vdd gnd cell_6t
Xbit_r203_c127 bl_127 br_127 wl_203 vdd gnd cell_6t
Xbit_r204_c127 bl_127 br_127 wl_204 vdd gnd cell_6t
Xbit_r205_c127 bl_127 br_127 wl_205 vdd gnd cell_6t
Xbit_r206_c127 bl_127 br_127 wl_206 vdd gnd cell_6t
Xbit_r207_c127 bl_127 br_127 wl_207 vdd gnd cell_6t
Xbit_r208_c127 bl_127 br_127 wl_208 vdd gnd cell_6t
Xbit_r209_c127 bl_127 br_127 wl_209 vdd gnd cell_6t
Xbit_r210_c127 bl_127 br_127 wl_210 vdd gnd cell_6t
Xbit_r211_c127 bl_127 br_127 wl_211 vdd gnd cell_6t
Xbit_r212_c127 bl_127 br_127 wl_212 vdd gnd cell_6t
Xbit_r213_c127 bl_127 br_127 wl_213 vdd gnd cell_6t
Xbit_r214_c127 bl_127 br_127 wl_214 vdd gnd cell_6t
Xbit_r215_c127 bl_127 br_127 wl_215 vdd gnd cell_6t
Xbit_r216_c127 bl_127 br_127 wl_216 vdd gnd cell_6t
Xbit_r217_c127 bl_127 br_127 wl_217 vdd gnd cell_6t
Xbit_r218_c127 bl_127 br_127 wl_218 vdd gnd cell_6t
Xbit_r219_c127 bl_127 br_127 wl_219 vdd gnd cell_6t
Xbit_r220_c127 bl_127 br_127 wl_220 vdd gnd cell_6t
Xbit_r221_c127 bl_127 br_127 wl_221 vdd gnd cell_6t
Xbit_r222_c127 bl_127 br_127 wl_222 vdd gnd cell_6t
Xbit_r223_c127 bl_127 br_127 wl_223 vdd gnd cell_6t
Xbit_r224_c127 bl_127 br_127 wl_224 vdd gnd cell_6t
Xbit_r225_c127 bl_127 br_127 wl_225 vdd gnd cell_6t
Xbit_r226_c127 bl_127 br_127 wl_226 vdd gnd cell_6t
Xbit_r227_c127 bl_127 br_127 wl_227 vdd gnd cell_6t
Xbit_r228_c127 bl_127 br_127 wl_228 vdd gnd cell_6t
Xbit_r229_c127 bl_127 br_127 wl_229 vdd gnd cell_6t
Xbit_r230_c127 bl_127 br_127 wl_230 vdd gnd cell_6t
Xbit_r231_c127 bl_127 br_127 wl_231 vdd gnd cell_6t
Xbit_r232_c127 bl_127 br_127 wl_232 vdd gnd cell_6t
Xbit_r233_c127 bl_127 br_127 wl_233 vdd gnd cell_6t
Xbit_r234_c127 bl_127 br_127 wl_234 vdd gnd cell_6t
Xbit_r235_c127 bl_127 br_127 wl_235 vdd gnd cell_6t
Xbit_r236_c127 bl_127 br_127 wl_236 vdd gnd cell_6t
Xbit_r237_c127 bl_127 br_127 wl_237 vdd gnd cell_6t
Xbit_r238_c127 bl_127 br_127 wl_238 vdd gnd cell_6t
Xbit_r239_c127 bl_127 br_127 wl_239 vdd gnd cell_6t
Xbit_r240_c127 bl_127 br_127 wl_240 vdd gnd cell_6t
Xbit_r241_c127 bl_127 br_127 wl_241 vdd gnd cell_6t
Xbit_r242_c127 bl_127 br_127 wl_242 vdd gnd cell_6t
Xbit_r243_c127 bl_127 br_127 wl_243 vdd gnd cell_6t
Xbit_r244_c127 bl_127 br_127 wl_244 vdd gnd cell_6t
Xbit_r245_c127 bl_127 br_127 wl_245 vdd gnd cell_6t
Xbit_r246_c127 bl_127 br_127 wl_246 vdd gnd cell_6t
Xbit_r247_c127 bl_127 br_127 wl_247 vdd gnd cell_6t
Xbit_r248_c127 bl_127 br_127 wl_248 vdd gnd cell_6t
Xbit_r249_c127 bl_127 br_127 wl_249 vdd gnd cell_6t
Xbit_r250_c127 bl_127 br_127 wl_250 vdd gnd cell_6t
Xbit_r251_c127 bl_127 br_127 wl_251 vdd gnd cell_6t
Xbit_r252_c127 bl_127 br_127 wl_252 vdd gnd cell_6t
Xbit_r253_c127 bl_127 br_127 wl_253 vdd gnd cell_6t
Xbit_r254_c127 bl_127 br_127 wl_254 vdd gnd cell_6t
Xbit_r255_c127 bl_127 br_127 wl_255 vdd gnd cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd cell_6t
Xbit_r1_c128 bl_128 br_128 wl_1 vdd gnd cell_6t
Xbit_r2_c128 bl_128 br_128 wl_2 vdd gnd cell_6t
Xbit_r3_c128 bl_128 br_128 wl_3 vdd gnd cell_6t
Xbit_r4_c128 bl_128 br_128 wl_4 vdd gnd cell_6t
Xbit_r5_c128 bl_128 br_128 wl_5 vdd gnd cell_6t
Xbit_r6_c128 bl_128 br_128 wl_6 vdd gnd cell_6t
Xbit_r7_c128 bl_128 br_128 wl_7 vdd gnd cell_6t
Xbit_r8_c128 bl_128 br_128 wl_8 vdd gnd cell_6t
Xbit_r9_c128 bl_128 br_128 wl_9 vdd gnd cell_6t
Xbit_r10_c128 bl_128 br_128 wl_10 vdd gnd cell_6t
Xbit_r11_c128 bl_128 br_128 wl_11 vdd gnd cell_6t
Xbit_r12_c128 bl_128 br_128 wl_12 vdd gnd cell_6t
Xbit_r13_c128 bl_128 br_128 wl_13 vdd gnd cell_6t
Xbit_r14_c128 bl_128 br_128 wl_14 vdd gnd cell_6t
Xbit_r15_c128 bl_128 br_128 wl_15 vdd gnd cell_6t
Xbit_r16_c128 bl_128 br_128 wl_16 vdd gnd cell_6t
Xbit_r17_c128 bl_128 br_128 wl_17 vdd gnd cell_6t
Xbit_r18_c128 bl_128 br_128 wl_18 vdd gnd cell_6t
Xbit_r19_c128 bl_128 br_128 wl_19 vdd gnd cell_6t
Xbit_r20_c128 bl_128 br_128 wl_20 vdd gnd cell_6t
Xbit_r21_c128 bl_128 br_128 wl_21 vdd gnd cell_6t
Xbit_r22_c128 bl_128 br_128 wl_22 vdd gnd cell_6t
Xbit_r23_c128 bl_128 br_128 wl_23 vdd gnd cell_6t
Xbit_r24_c128 bl_128 br_128 wl_24 vdd gnd cell_6t
Xbit_r25_c128 bl_128 br_128 wl_25 vdd gnd cell_6t
Xbit_r26_c128 bl_128 br_128 wl_26 vdd gnd cell_6t
Xbit_r27_c128 bl_128 br_128 wl_27 vdd gnd cell_6t
Xbit_r28_c128 bl_128 br_128 wl_28 vdd gnd cell_6t
Xbit_r29_c128 bl_128 br_128 wl_29 vdd gnd cell_6t
Xbit_r30_c128 bl_128 br_128 wl_30 vdd gnd cell_6t
Xbit_r31_c128 bl_128 br_128 wl_31 vdd gnd cell_6t
Xbit_r32_c128 bl_128 br_128 wl_32 vdd gnd cell_6t
Xbit_r33_c128 bl_128 br_128 wl_33 vdd gnd cell_6t
Xbit_r34_c128 bl_128 br_128 wl_34 vdd gnd cell_6t
Xbit_r35_c128 bl_128 br_128 wl_35 vdd gnd cell_6t
Xbit_r36_c128 bl_128 br_128 wl_36 vdd gnd cell_6t
Xbit_r37_c128 bl_128 br_128 wl_37 vdd gnd cell_6t
Xbit_r38_c128 bl_128 br_128 wl_38 vdd gnd cell_6t
Xbit_r39_c128 bl_128 br_128 wl_39 vdd gnd cell_6t
Xbit_r40_c128 bl_128 br_128 wl_40 vdd gnd cell_6t
Xbit_r41_c128 bl_128 br_128 wl_41 vdd gnd cell_6t
Xbit_r42_c128 bl_128 br_128 wl_42 vdd gnd cell_6t
Xbit_r43_c128 bl_128 br_128 wl_43 vdd gnd cell_6t
Xbit_r44_c128 bl_128 br_128 wl_44 vdd gnd cell_6t
Xbit_r45_c128 bl_128 br_128 wl_45 vdd gnd cell_6t
Xbit_r46_c128 bl_128 br_128 wl_46 vdd gnd cell_6t
Xbit_r47_c128 bl_128 br_128 wl_47 vdd gnd cell_6t
Xbit_r48_c128 bl_128 br_128 wl_48 vdd gnd cell_6t
Xbit_r49_c128 bl_128 br_128 wl_49 vdd gnd cell_6t
Xbit_r50_c128 bl_128 br_128 wl_50 vdd gnd cell_6t
Xbit_r51_c128 bl_128 br_128 wl_51 vdd gnd cell_6t
Xbit_r52_c128 bl_128 br_128 wl_52 vdd gnd cell_6t
Xbit_r53_c128 bl_128 br_128 wl_53 vdd gnd cell_6t
Xbit_r54_c128 bl_128 br_128 wl_54 vdd gnd cell_6t
Xbit_r55_c128 bl_128 br_128 wl_55 vdd gnd cell_6t
Xbit_r56_c128 bl_128 br_128 wl_56 vdd gnd cell_6t
Xbit_r57_c128 bl_128 br_128 wl_57 vdd gnd cell_6t
Xbit_r58_c128 bl_128 br_128 wl_58 vdd gnd cell_6t
Xbit_r59_c128 bl_128 br_128 wl_59 vdd gnd cell_6t
Xbit_r60_c128 bl_128 br_128 wl_60 vdd gnd cell_6t
Xbit_r61_c128 bl_128 br_128 wl_61 vdd gnd cell_6t
Xbit_r62_c128 bl_128 br_128 wl_62 vdd gnd cell_6t
Xbit_r63_c128 bl_128 br_128 wl_63 vdd gnd cell_6t
Xbit_r64_c128 bl_128 br_128 wl_64 vdd gnd cell_6t
Xbit_r65_c128 bl_128 br_128 wl_65 vdd gnd cell_6t
Xbit_r66_c128 bl_128 br_128 wl_66 vdd gnd cell_6t
Xbit_r67_c128 bl_128 br_128 wl_67 vdd gnd cell_6t
Xbit_r68_c128 bl_128 br_128 wl_68 vdd gnd cell_6t
Xbit_r69_c128 bl_128 br_128 wl_69 vdd gnd cell_6t
Xbit_r70_c128 bl_128 br_128 wl_70 vdd gnd cell_6t
Xbit_r71_c128 bl_128 br_128 wl_71 vdd gnd cell_6t
Xbit_r72_c128 bl_128 br_128 wl_72 vdd gnd cell_6t
Xbit_r73_c128 bl_128 br_128 wl_73 vdd gnd cell_6t
Xbit_r74_c128 bl_128 br_128 wl_74 vdd gnd cell_6t
Xbit_r75_c128 bl_128 br_128 wl_75 vdd gnd cell_6t
Xbit_r76_c128 bl_128 br_128 wl_76 vdd gnd cell_6t
Xbit_r77_c128 bl_128 br_128 wl_77 vdd gnd cell_6t
Xbit_r78_c128 bl_128 br_128 wl_78 vdd gnd cell_6t
Xbit_r79_c128 bl_128 br_128 wl_79 vdd gnd cell_6t
Xbit_r80_c128 bl_128 br_128 wl_80 vdd gnd cell_6t
Xbit_r81_c128 bl_128 br_128 wl_81 vdd gnd cell_6t
Xbit_r82_c128 bl_128 br_128 wl_82 vdd gnd cell_6t
Xbit_r83_c128 bl_128 br_128 wl_83 vdd gnd cell_6t
Xbit_r84_c128 bl_128 br_128 wl_84 vdd gnd cell_6t
Xbit_r85_c128 bl_128 br_128 wl_85 vdd gnd cell_6t
Xbit_r86_c128 bl_128 br_128 wl_86 vdd gnd cell_6t
Xbit_r87_c128 bl_128 br_128 wl_87 vdd gnd cell_6t
Xbit_r88_c128 bl_128 br_128 wl_88 vdd gnd cell_6t
Xbit_r89_c128 bl_128 br_128 wl_89 vdd gnd cell_6t
Xbit_r90_c128 bl_128 br_128 wl_90 vdd gnd cell_6t
Xbit_r91_c128 bl_128 br_128 wl_91 vdd gnd cell_6t
Xbit_r92_c128 bl_128 br_128 wl_92 vdd gnd cell_6t
Xbit_r93_c128 bl_128 br_128 wl_93 vdd gnd cell_6t
Xbit_r94_c128 bl_128 br_128 wl_94 vdd gnd cell_6t
Xbit_r95_c128 bl_128 br_128 wl_95 vdd gnd cell_6t
Xbit_r96_c128 bl_128 br_128 wl_96 vdd gnd cell_6t
Xbit_r97_c128 bl_128 br_128 wl_97 vdd gnd cell_6t
Xbit_r98_c128 bl_128 br_128 wl_98 vdd gnd cell_6t
Xbit_r99_c128 bl_128 br_128 wl_99 vdd gnd cell_6t
Xbit_r100_c128 bl_128 br_128 wl_100 vdd gnd cell_6t
Xbit_r101_c128 bl_128 br_128 wl_101 vdd gnd cell_6t
Xbit_r102_c128 bl_128 br_128 wl_102 vdd gnd cell_6t
Xbit_r103_c128 bl_128 br_128 wl_103 vdd gnd cell_6t
Xbit_r104_c128 bl_128 br_128 wl_104 vdd gnd cell_6t
Xbit_r105_c128 bl_128 br_128 wl_105 vdd gnd cell_6t
Xbit_r106_c128 bl_128 br_128 wl_106 vdd gnd cell_6t
Xbit_r107_c128 bl_128 br_128 wl_107 vdd gnd cell_6t
Xbit_r108_c128 bl_128 br_128 wl_108 vdd gnd cell_6t
Xbit_r109_c128 bl_128 br_128 wl_109 vdd gnd cell_6t
Xbit_r110_c128 bl_128 br_128 wl_110 vdd gnd cell_6t
Xbit_r111_c128 bl_128 br_128 wl_111 vdd gnd cell_6t
Xbit_r112_c128 bl_128 br_128 wl_112 vdd gnd cell_6t
Xbit_r113_c128 bl_128 br_128 wl_113 vdd gnd cell_6t
Xbit_r114_c128 bl_128 br_128 wl_114 vdd gnd cell_6t
Xbit_r115_c128 bl_128 br_128 wl_115 vdd gnd cell_6t
Xbit_r116_c128 bl_128 br_128 wl_116 vdd gnd cell_6t
Xbit_r117_c128 bl_128 br_128 wl_117 vdd gnd cell_6t
Xbit_r118_c128 bl_128 br_128 wl_118 vdd gnd cell_6t
Xbit_r119_c128 bl_128 br_128 wl_119 vdd gnd cell_6t
Xbit_r120_c128 bl_128 br_128 wl_120 vdd gnd cell_6t
Xbit_r121_c128 bl_128 br_128 wl_121 vdd gnd cell_6t
Xbit_r122_c128 bl_128 br_128 wl_122 vdd gnd cell_6t
Xbit_r123_c128 bl_128 br_128 wl_123 vdd gnd cell_6t
Xbit_r124_c128 bl_128 br_128 wl_124 vdd gnd cell_6t
Xbit_r125_c128 bl_128 br_128 wl_125 vdd gnd cell_6t
Xbit_r126_c128 bl_128 br_128 wl_126 vdd gnd cell_6t
Xbit_r127_c128 bl_128 br_128 wl_127 vdd gnd cell_6t
Xbit_r128_c128 bl_128 br_128 wl_128 vdd gnd cell_6t
Xbit_r129_c128 bl_128 br_128 wl_129 vdd gnd cell_6t
Xbit_r130_c128 bl_128 br_128 wl_130 vdd gnd cell_6t
Xbit_r131_c128 bl_128 br_128 wl_131 vdd gnd cell_6t
Xbit_r132_c128 bl_128 br_128 wl_132 vdd gnd cell_6t
Xbit_r133_c128 bl_128 br_128 wl_133 vdd gnd cell_6t
Xbit_r134_c128 bl_128 br_128 wl_134 vdd gnd cell_6t
Xbit_r135_c128 bl_128 br_128 wl_135 vdd gnd cell_6t
Xbit_r136_c128 bl_128 br_128 wl_136 vdd gnd cell_6t
Xbit_r137_c128 bl_128 br_128 wl_137 vdd gnd cell_6t
Xbit_r138_c128 bl_128 br_128 wl_138 vdd gnd cell_6t
Xbit_r139_c128 bl_128 br_128 wl_139 vdd gnd cell_6t
Xbit_r140_c128 bl_128 br_128 wl_140 vdd gnd cell_6t
Xbit_r141_c128 bl_128 br_128 wl_141 vdd gnd cell_6t
Xbit_r142_c128 bl_128 br_128 wl_142 vdd gnd cell_6t
Xbit_r143_c128 bl_128 br_128 wl_143 vdd gnd cell_6t
Xbit_r144_c128 bl_128 br_128 wl_144 vdd gnd cell_6t
Xbit_r145_c128 bl_128 br_128 wl_145 vdd gnd cell_6t
Xbit_r146_c128 bl_128 br_128 wl_146 vdd gnd cell_6t
Xbit_r147_c128 bl_128 br_128 wl_147 vdd gnd cell_6t
Xbit_r148_c128 bl_128 br_128 wl_148 vdd gnd cell_6t
Xbit_r149_c128 bl_128 br_128 wl_149 vdd gnd cell_6t
Xbit_r150_c128 bl_128 br_128 wl_150 vdd gnd cell_6t
Xbit_r151_c128 bl_128 br_128 wl_151 vdd gnd cell_6t
Xbit_r152_c128 bl_128 br_128 wl_152 vdd gnd cell_6t
Xbit_r153_c128 bl_128 br_128 wl_153 vdd gnd cell_6t
Xbit_r154_c128 bl_128 br_128 wl_154 vdd gnd cell_6t
Xbit_r155_c128 bl_128 br_128 wl_155 vdd gnd cell_6t
Xbit_r156_c128 bl_128 br_128 wl_156 vdd gnd cell_6t
Xbit_r157_c128 bl_128 br_128 wl_157 vdd gnd cell_6t
Xbit_r158_c128 bl_128 br_128 wl_158 vdd gnd cell_6t
Xbit_r159_c128 bl_128 br_128 wl_159 vdd gnd cell_6t
Xbit_r160_c128 bl_128 br_128 wl_160 vdd gnd cell_6t
Xbit_r161_c128 bl_128 br_128 wl_161 vdd gnd cell_6t
Xbit_r162_c128 bl_128 br_128 wl_162 vdd gnd cell_6t
Xbit_r163_c128 bl_128 br_128 wl_163 vdd gnd cell_6t
Xbit_r164_c128 bl_128 br_128 wl_164 vdd gnd cell_6t
Xbit_r165_c128 bl_128 br_128 wl_165 vdd gnd cell_6t
Xbit_r166_c128 bl_128 br_128 wl_166 vdd gnd cell_6t
Xbit_r167_c128 bl_128 br_128 wl_167 vdd gnd cell_6t
Xbit_r168_c128 bl_128 br_128 wl_168 vdd gnd cell_6t
Xbit_r169_c128 bl_128 br_128 wl_169 vdd gnd cell_6t
Xbit_r170_c128 bl_128 br_128 wl_170 vdd gnd cell_6t
Xbit_r171_c128 bl_128 br_128 wl_171 vdd gnd cell_6t
Xbit_r172_c128 bl_128 br_128 wl_172 vdd gnd cell_6t
Xbit_r173_c128 bl_128 br_128 wl_173 vdd gnd cell_6t
Xbit_r174_c128 bl_128 br_128 wl_174 vdd gnd cell_6t
Xbit_r175_c128 bl_128 br_128 wl_175 vdd gnd cell_6t
Xbit_r176_c128 bl_128 br_128 wl_176 vdd gnd cell_6t
Xbit_r177_c128 bl_128 br_128 wl_177 vdd gnd cell_6t
Xbit_r178_c128 bl_128 br_128 wl_178 vdd gnd cell_6t
Xbit_r179_c128 bl_128 br_128 wl_179 vdd gnd cell_6t
Xbit_r180_c128 bl_128 br_128 wl_180 vdd gnd cell_6t
Xbit_r181_c128 bl_128 br_128 wl_181 vdd gnd cell_6t
Xbit_r182_c128 bl_128 br_128 wl_182 vdd gnd cell_6t
Xbit_r183_c128 bl_128 br_128 wl_183 vdd gnd cell_6t
Xbit_r184_c128 bl_128 br_128 wl_184 vdd gnd cell_6t
Xbit_r185_c128 bl_128 br_128 wl_185 vdd gnd cell_6t
Xbit_r186_c128 bl_128 br_128 wl_186 vdd gnd cell_6t
Xbit_r187_c128 bl_128 br_128 wl_187 vdd gnd cell_6t
Xbit_r188_c128 bl_128 br_128 wl_188 vdd gnd cell_6t
Xbit_r189_c128 bl_128 br_128 wl_189 vdd gnd cell_6t
Xbit_r190_c128 bl_128 br_128 wl_190 vdd gnd cell_6t
Xbit_r191_c128 bl_128 br_128 wl_191 vdd gnd cell_6t
Xbit_r192_c128 bl_128 br_128 wl_192 vdd gnd cell_6t
Xbit_r193_c128 bl_128 br_128 wl_193 vdd gnd cell_6t
Xbit_r194_c128 bl_128 br_128 wl_194 vdd gnd cell_6t
Xbit_r195_c128 bl_128 br_128 wl_195 vdd gnd cell_6t
Xbit_r196_c128 bl_128 br_128 wl_196 vdd gnd cell_6t
Xbit_r197_c128 bl_128 br_128 wl_197 vdd gnd cell_6t
Xbit_r198_c128 bl_128 br_128 wl_198 vdd gnd cell_6t
Xbit_r199_c128 bl_128 br_128 wl_199 vdd gnd cell_6t
Xbit_r200_c128 bl_128 br_128 wl_200 vdd gnd cell_6t
Xbit_r201_c128 bl_128 br_128 wl_201 vdd gnd cell_6t
Xbit_r202_c128 bl_128 br_128 wl_202 vdd gnd cell_6t
Xbit_r203_c128 bl_128 br_128 wl_203 vdd gnd cell_6t
Xbit_r204_c128 bl_128 br_128 wl_204 vdd gnd cell_6t
Xbit_r205_c128 bl_128 br_128 wl_205 vdd gnd cell_6t
Xbit_r206_c128 bl_128 br_128 wl_206 vdd gnd cell_6t
Xbit_r207_c128 bl_128 br_128 wl_207 vdd gnd cell_6t
Xbit_r208_c128 bl_128 br_128 wl_208 vdd gnd cell_6t
Xbit_r209_c128 bl_128 br_128 wl_209 vdd gnd cell_6t
Xbit_r210_c128 bl_128 br_128 wl_210 vdd gnd cell_6t
Xbit_r211_c128 bl_128 br_128 wl_211 vdd gnd cell_6t
Xbit_r212_c128 bl_128 br_128 wl_212 vdd gnd cell_6t
Xbit_r213_c128 bl_128 br_128 wl_213 vdd gnd cell_6t
Xbit_r214_c128 bl_128 br_128 wl_214 vdd gnd cell_6t
Xbit_r215_c128 bl_128 br_128 wl_215 vdd gnd cell_6t
Xbit_r216_c128 bl_128 br_128 wl_216 vdd gnd cell_6t
Xbit_r217_c128 bl_128 br_128 wl_217 vdd gnd cell_6t
Xbit_r218_c128 bl_128 br_128 wl_218 vdd gnd cell_6t
Xbit_r219_c128 bl_128 br_128 wl_219 vdd gnd cell_6t
Xbit_r220_c128 bl_128 br_128 wl_220 vdd gnd cell_6t
Xbit_r221_c128 bl_128 br_128 wl_221 vdd gnd cell_6t
Xbit_r222_c128 bl_128 br_128 wl_222 vdd gnd cell_6t
Xbit_r223_c128 bl_128 br_128 wl_223 vdd gnd cell_6t
Xbit_r224_c128 bl_128 br_128 wl_224 vdd gnd cell_6t
Xbit_r225_c128 bl_128 br_128 wl_225 vdd gnd cell_6t
Xbit_r226_c128 bl_128 br_128 wl_226 vdd gnd cell_6t
Xbit_r227_c128 bl_128 br_128 wl_227 vdd gnd cell_6t
Xbit_r228_c128 bl_128 br_128 wl_228 vdd gnd cell_6t
Xbit_r229_c128 bl_128 br_128 wl_229 vdd gnd cell_6t
Xbit_r230_c128 bl_128 br_128 wl_230 vdd gnd cell_6t
Xbit_r231_c128 bl_128 br_128 wl_231 vdd gnd cell_6t
Xbit_r232_c128 bl_128 br_128 wl_232 vdd gnd cell_6t
Xbit_r233_c128 bl_128 br_128 wl_233 vdd gnd cell_6t
Xbit_r234_c128 bl_128 br_128 wl_234 vdd gnd cell_6t
Xbit_r235_c128 bl_128 br_128 wl_235 vdd gnd cell_6t
Xbit_r236_c128 bl_128 br_128 wl_236 vdd gnd cell_6t
Xbit_r237_c128 bl_128 br_128 wl_237 vdd gnd cell_6t
Xbit_r238_c128 bl_128 br_128 wl_238 vdd gnd cell_6t
Xbit_r239_c128 bl_128 br_128 wl_239 vdd gnd cell_6t
Xbit_r240_c128 bl_128 br_128 wl_240 vdd gnd cell_6t
Xbit_r241_c128 bl_128 br_128 wl_241 vdd gnd cell_6t
Xbit_r242_c128 bl_128 br_128 wl_242 vdd gnd cell_6t
Xbit_r243_c128 bl_128 br_128 wl_243 vdd gnd cell_6t
Xbit_r244_c128 bl_128 br_128 wl_244 vdd gnd cell_6t
Xbit_r245_c128 bl_128 br_128 wl_245 vdd gnd cell_6t
Xbit_r246_c128 bl_128 br_128 wl_246 vdd gnd cell_6t
Xbit_r247_c128 bl_128 br_128 wl_247 vdd gnd cell_6t
Xbit_r248_c128 bl_128 br_128 wl_248 vdd gnd cell_6t
Xbit_r249_c128 bl_128 br_128 wl_249 vdd gnd cell_6t
Xbit_r250_c128 bl_128 br_128 wl_250 vdd gnd cell_6t
Xbit_r251_c128 bl_128 br_128 wl_251 vdd gnd cell_6t
Xbit_r252_c128 bl_128 br_128 wl_252 vdd gnd cell_6t
Xbit_r253_c128 bl_128 br_128 wl_253 vdd gnd cell_6t
Xbit_r254_c128 bl_128 br_128 wl_254 vdd gnd cell_6t
Xbit_r255_c128 bl_128 br_128 wl_255 vdd gnd cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd cell_6t
Xbit_r1_c129 bl_129 br_129 wl_1 vdd gnd cell_6t
Xbit_r2_c129 bl_129 br_129 wl_2 vdd gnd cell_6t
Xbit_r3_c129 bl_129 br_129 wl_3 vdd gnd cell_6t
Xbit_r4_c129 bl_129 br_129 wl_4 vdd gnd cell_6t
Xbit_r5_c129 bl_129 br_129 wl_5 vdd gnd cell_6t
Xbit_r6_c129 bl_129 br_129 wl_6 vdd gnd cell_6t
Xbit_r7_c129 bl_129 br_129 wl_7 vdd gnd cell_6t
Xbit_r8_c129 bl_129 br_129 wl_8 vdd gnd cell_6t
Xbit_r9_c129 bl_129 br_129 wl_9 vdd gnd cell_6t
Xbit_r10_c129 bl_129 br_129 wl_10 vdd gnd cell_6t
Xbit_r11_c129 bl_129 br_129 wl_11 vdd gnd cell_6t
Xbit_r12_c129 bl_129 br_129 wl_12 vdd gnd cell_6t
Xbit_r13_c129 bl_129 br_129 wl_13 vdd gnd cell_6t
Xbit_r14_c129 bl_129 br_129 wl_14 vdd gnd cell_6t
Xbit_r15_c129 bl_129 br_129 wl_15 vdd gnd cell_6t
Xbit_r16_c129 bl_129 br_129 wl_16 vdd gnd cell_6t
Xbit_r17_c129 bl_129 br_129 wl_17 vdd gnd cell_6t
Xbit_r18_c129 bl_129 br_129 wl_18 vdd gnd cell_6t
Xbit_r19_c129 bl_129 br_129 wl_19 vdd gnd cell_6t
Xbit_r20_c129 bl_129 br_129 wl_20 vdd gnd cell_6t
Xbit_r21_c129 bl_129 br_129 wl_21 vdd gnd cell_6t
Xbit_r22_c129 bl_129 br_129 wl_22 vdd gnd cell_6t
Xbit_r23_c129 bl_129 br_129 wl_23 vdd gnd cell_6t
Xbit_r24_c129 bl_129 br_129 wl_24 vdd gnd cell_6t
Xbit_r25_c129 bl_129 br_129 wl_25 vdd gnd cell_6t
Xbit_r26_c129 bl_129 br_129 wl_26 vdd gnd cell_6t
Xbit_r27_c129 bl_129 br_129 wl_27 vdd gnd cell_6t
Xbit_r28_c129 bl_129 br_129 wl_28 vdd gnd cell_6t
Xbit_r29_c129 bl_129 br_129 wl_29 vdd gnd cell_6t
Xbit_r30_c129 bl_129 br_129 wl_30 vdd gnd cell_6t
Xbit_r31_c129 bl_129 br_129 wl_31 vdd gnd cell_6t
Xbit_r32_c129 bl_129 br_129 wl_32 vdd gnd cell_6t
Xbit_r33_c129 bl_129 br_129 wl_33 vdd gnd cell_6t
Xbit_r34_c129 bl_129 br_129 wl_34 vdd gnd cell_6t
Xbit_r35_c129 bl_129 br_129 wl_35 vdd gnd cell_6t
Xbit_r36_c129 bl_129 br_129 wl_36 vdd gnd cell_6t
Xbit_r37_c129 bl_129 br_129 wl_37 vdd gnd cell_6t
Xbit_r38_c129 bl_129 br_129 wl_38 vdd gnd cell_6t
Xbit_r39_c129 bl_129 br_129 wl_39 vdd gnd cell_6t
Xbit_r40_c129 bl_129 br_129 wl_40 vdd gnd cell_6t
Xbit_r41_c129 bl_129 br_129 wl_41 vdd gnd cell_6t
Xbit_r42_c129 bl_129 br_129 wl_42 vdd gnd cell_6t
Xbit_r43_c129 bl_129 br_129 wl_43 vdd gnd cell_6t
Xbit_r44_c129 bl_129 br_129 wl_44 vdd gnd cell_6t
Xbit_r45_c129 bl_129 br_129 wl_45 vdd gnd cell_6t
Xbit_r46_c129 bl_129 br_129 wl_46 vdd gnd cell_6t
Xbit_r47_c129 bl_129 br_129 wl_47 vdd gnd cell_6t
Xbit_r48_c129 bl_129 br_129 wl_48 vdd gnd cell_6t
Xbit_r49_c129 bl_129 br_129 wl_49 vdd gnd cell_6t
Xbit_r50_c129 bl_129 br_129 wl_50 vdd gnd cell_6t
Xbit_r51_c129 bl_129 br_129 wl_51 vdd gnd cell_6t
Xbit_r52_c129 bl_129 br_129 wl_52 vdd gnd cell_6t
Xbit_r53_c129 bl_129 br_129 wl_53 vdd gnd cell_6t
Xbit_r54_c129 bl_129 br_129 wl_54 vdd gnd cell_6t
Xbit_r55_c129 bl_129 br_129 wl_55 vdd gnd cell_6t
Xbit_r56_c129 bl_129 br_129 wl_56 vdd gnd cell_6t
Xbit_r57_c129 bl_129 br_129 wl_57 vdd gnd cell_6t
Xbit_r58_c129 bl_129 br_129 wl_58 vdd gnd cell_6t
Xbit_r59_c129 bl_129 br_129 wl_59 vdd gnd cell_6t
Xbit_r60_c129 bl_129 br_129 wl_60 vdd gnd cell_6t
Xbit_r61_c129 bl_129 br_129 wl_61 vdd gnd cell_6t
Xbit_r62_c129 bl_129 br_129 wl_62 vdd gnd cell_6t
Xbit_r63_c129 bl_129 br_129 wl_63 vdd gnd cell_6t
Xbit_r64_c129 bl_129 br_129 wl_64 vdd gnd cell_6t
Xbit_r65_c129 bl_129 br_129 wl_65 vdd gnd cell_6t
Xbit_r66_c129 bl_129 br_129 wl_66 vdd gnd cell_6t
Xbit_r67_c129 bl_129 br_129 wl_67 vdd gnd cell_6t
Xbit_r68_c129 bl_129 br_129 wl_68 vdd gnd cell_6t
Xbit_r69_c129 bl_129 br_129 wl_69 vdd gnd cell_6t
Xbit_r70_c129 bl_129 br_129 wl_70 vdd gnd cell_6t
Xbit_r71_c129 bl_129 br_129 wl_71 vdd gnd cell_6t
Xbit_r72_c129 bl_129 br_129 wl_72 vdd gnd cell_6t
Xbit_r73_c129 bl_129 br_129 wl_73 vdd gnd cell_6t
Xbit_r74_c129 bl_129 br_129 wl_74 vdd gnd cell_6t
Xbit_r75_c129 bl_129 br_129 wl_75 vdd gnd cell_6t
Xbit_r76_c129 bl_129 br_129 wl_76 vdd gnd cell_6t
Xbit_r77_c129 bl_129 br_129 wl_77 vdd gnd cell_6t
Xbit_r78_c129 bl_129 br_129 wl_78 vdd gnd cell_6t
Xbit_r79_c129 bl_129 br_129 wl_79 vdd gnd cell_6t
Xbit_r80_c129 bl_129 br_129 wl_80 vdd gnd cell_6t
Xbit_r81_c129 bl_129 br_129 wl_81 vdd gnd cell_6t
Xbit_r82_c129 bl_129 br_129 wl_82 vdd gnd cell_6t
Xbit_r83_c129 bl_129 br_129 wl_83 vdd gnd cell_6t
Xbit_r84_c129 bl_129 br_129 wl_84 vdd gnd cell_6t
Xbit_r85_c129 bl_129 br_129 wl_85 vdd gnd cell_6t
Xbit_r86_c129 bl_129 br_129 wl_86 vdd gnd cell_6t
Xbit_r87_c129 bl_129 br_129 wl_87 vdd gnd cell_6t
Xbit_r88_c129 bl_129 br_129 wl_88 vdd gnd cell_6t
Xbit_r89_c129 bl_129 br_129 wl_89 vdd gnd cell_6t
Xbit_r90_c129 bl_129 br_129 wl_90 vdd gnd cell_6t
Xbit_r91_c129 bl_129 br_129 wl_91 vdd gnd cell_6t
Xbit_r92_c129 bl_129 br_129 wl_92 vdd gnd cell_6t
Xbit_r93_c129 bl_129 br_129 wl_93 vdd gnd cell_6t
Xbit_r94_c129 bl_129 br_129 wl_94 vdd gnd cell_6t
Xbit_r95_c129 bl_129 br_129 wl_95 vdd gnd cell_6t
Xbit_r96_c129 bl_129 br_129 wl_96 vdd gnd cell_6t
Xbit_r97_c129 bl_129 br_129 wl_97 vdd gnd cell_6t
Xbit_r98_c129 bl_129 br_129 wl_98 vdd gnd cell_6t
Xbit_r99_c129 bl_129 br_129 wl_99 vdd gnd cell_6t
Xbit_r100_c129 bl_129 br_129 wl_100 vdd gnd cell_6t
Xbit_r101_c129 bl_129 br_129 wl_101 vdd gnd cell_6t
Xbit_r102_c129 bl_129 br_129 wl_102 vdd gnd cell_6t
Xbit_r103_c129 bl_129 br_129 wl_103 vdd gnd cell_6t
Xbit_r104_c129 bl_129 br_129 wl_104 vdd gnd cell_6t
Xbit_r105_c129 bl_129 br_129 wl_105 vdd gnd cell_6t
Xbit_r106_c129 bl_129 br_129 wl_106 vdd gnd cell_6t
Xbit_r107_c129 bl_129 br_129 wl_107 vdd gnd cell_6t
Xbit_r108_c129 bl_129 br_129 wl_108 vdd gnd cell_6t
Xbit_r109_c129 bl_129 br_129 wl_109 vdd gnd cell_6t
Xbit_r110_c129 bl_129 br_129 wl_110 vdd gnd cell_6t
Xbit_r111_c129 bl_129 br_129 wl_111 vdd gnd cell_6t
Xbit_r112_c129 bl_129 br_129 wl_112 vdd gnd cell_6t
Xbit_r113_c129 bl_129 br_129 wl_113 vdd gnd cell_6t
Xbit_r114_c129 bl_129 br_129 wl_114 vdd gnd cell_6t
Xbit_r115_c129 bl_129 br_129 wl_115 vdd gnd cell_6t
Xbit_r116_c129 bl_129 br_129 wl_116 vdd gnd cell_6t
Xbit_r117_c129 bl_129 br_129 wl_117 vdd gnd cell_6t
Xbit_r118_c129 bl_129 br_129 wl_118 vdd gnd cell_6t
Xbit_r119_c129 bl_129 br_129 wl_119 vdd gnd cell_6t
Xbit_r120_c129 bl_129 br_129 wl_120 vdd gnd cell_6t
Xbit_r121_c129 bl_129 br_129 wl_121 vdd gnd cell_6t
Xbit_r122_c129 bl_129 br_129 wl_122 vdd gnd cell_6t
Xbit_r123_c129 bl_129 br_129 wl_123 vdd gnd cell_6t
Xbit_r124_c129 bl_129 br_129 wl_124 vdd gnd cell_6t
Xbit_r125_c129 bl_129 br_129 wl_125 vdd gnd cell_6t
Xbit_r126_c129 bl_129 br_129 wl_126 vdd gnd cell_6t
Xbit_r127_c129 bl_129 br_129 wl_127 vdd gnd cell_6t
Xbit_r128_c129 bl_129 br_129 wl_128 vdd gnd cell_6t
Xbit_r129_c129 bl_129 br_129 wl_129 vdd gnd cell_6t
Xbit_r130_c129 bl_129 br_129 wl_130 vdd gnd cell_6t
Xbit_r131_c129 bl_129 br_129 wl_131 vdd gnd cell_6t
Xbit_r132_c129 bl_129 br_129 wl_132 vdd gnd cell_6t
Xbit_r133_c129 bl_129 br_129 wl_133 vdd gnd cell_6t
Xbit_r134_c129 bl_129 br_129 wl_134 vdd gnd cell_6t
Xbit_r135_c129 bl_129 br_129 wl_135 vdd gnd cell_6t
Xbit_r136_c129 bl_129 br_129 wl_136 vdd gnd cell_6t
Xbit_r137_c129 bl_129 br_129 wl_137 vdd gnd cell_6t
Xbit_r138_c129 bl_129 br_129 wl_138 vdd gnd cell_6t
Xbit_r139_c129 bl_129 br_129 wl_139 vdd gnd cell_6t
Xbit_r140_c129 bl_129 br_129 wl_140 vdd gnd cell_6t
Xbit_r141_c129 bl_129 br_129 wl_141 vdd gnd cell_6t
Xbit_r142_c129 bl_129 br_129 wl_142 vdd gnd cell_6t
Xbit_r143_c129 bl_129 br_129 wl_143 vdd gnd cell_6t
Xbit_r144_c129 bl_129 br_129 wl_144 vdd gnd cell_6t
Xbit_r145_c129 bl_129 br_129 wl_145 vdd gnd cell_6t
Xbit_r146_c129 bl_129 br_129 wl_146 vdd gnd cell_6t
Xbit_r147_c129 bl_129 br_129 wl_147 vdd gnd cell_6t
Xbit_r148_c129 bl_129 br_129 wl_148 vdd gnd cell_6t
Xbit_r149_c129 bl_129 br_129 wl_149 vdd gnd cell_6t
Xbit_r150_c129 bl_129 br_129 wl_150 vdd gnd cell_6t
Xbit_r151_c129 bl_129 br_129 wl_151 vdd gnd cell_6t
Xbit_r152_c129 bl_129 br_129 wl_152 vdd gnd cell_6t
Xbit_r153_c129 bl_129 br_129 wl_153 vdd gnd cell_6t
Xbit_r154_c129 bl_129 br_129 wl_154 vdd gnd cell_6t
Xbit_r155_c129 bl_129 br_129 wl_155 vdd gnd cell_6t
Xbit_r156_c129 bl_129 br_129 wl_156 vdd gnd cell_6t
Xbit_r157_c129 bl_129 br_129 wl_157 vdd gnd cell_6t
Xbit_r158_c129 bl_129 br_129 wl_158 vdd gnd cell_6t
Xbit_r159_c129 bl_129 br_129 wl_159 vdd gnd cell_6t
Xbit_r160_c129 bl_129 br_129 wl_160 vdd gnd cell_6t
Xbit_r161_c129 bl_129 br_129 wl_161 vdd gnd cell_6t
Xbit_r162_c129 bl_129 br_129 wl_162 vdd gnd cell_6t
Xbit_r163_c129 bl_129 br_129 wl_163 vdd gnd cell_6t
Xbit_r164_c129 bl_129 br_129 wl_164 vdd gnd cell_6t
Xbit_r165_c129 bl_129 br_129 wl_165 vdd gnd cell_6t
Xbit_r166_c129 bl_129 br_129 wl_166 vdd gnd cell_6t
Xbit_r167_c129 bl_129 br_129 wl_167 vdd gnd cell_6t
Xbit_r168_c129 bl_129 br_129 wl_168 vdd gnd cell_6t
Xbit_r169_c129 bl_129 br_129 wl_169 vdd gnd cell_6t
Xbit_r170_c129 bl_129 br_129 wl_170 vdd gnd cell_6t
Xbit_r171_c129 bl_129 br_129 wl_171 vdd gnd cell_6t
Xbit_r172_c129 bl_129 br_129 wl_172 vdd gnd cell_6t
Xbit_r173_c129 bl_129 br_129 wl_173 vdd gnd cell_6t
Xbit_r174_c129 bl_129 br_129 wl_174 vdd gnd cell_6t
Xbit_r175_c129 bl_129 br_129 wl_175 vdd gnd cell_6t
Xbit_r176_c129 bl_129 br_129 wl_176 vdd gnd cell_6t
Xbit_r177_c129 bl_129 br_129 wl_177 vdd gnd cell_6t
Xbit_r178_c129 bl_129 br_129 wl_178 vdd gnd cell_6t
Xbit_r179_c129 bl_129 br_129 wl_179 vdd gnd cell_6t
Xbit_r180_c129 bl_129 br_129 wl_180 vdd gnd cell_6t
Xbit_r181_c129 bl_129 br_129 wl_181 vdd gnd cell_6t
Xbit_r182_c129 bl_129 br_129 wl_182 vdd gnd cell_6t
Xbit_r183_c129 bl_129 br_129 wl_183 vdd gnd cell_6t
Xbit_r184_c129 bl_129 br_129 wl_184 vdd gnd cell_6t
Xbit_r185_c129 bl_129 br_129 wl_185 vdd gnd cell_6t
Xbit_r186_c129 bl_129 br_129 wl_186 vdd gnd cell_6t
Xbit_r187_c129 bl_129 br_129 wl_187 vdd gnd cell_6t
Xbit_r188_c129 bl_129 br_129 wl_188 vdd gnd cell_6t
Xbit_r189_c129 bl_129 br_129 wl_189 vdd gnd cell_6t
Xbit_r190_c129 bl_129 br_129 wl_190 vdd gnd cell_6t
Xbit_r191_c129 bl_129 br_129 wl_191 vdd gnd cell_6t
Xbit_r192_c129 bl_129 br_129 wl_192 vdd gnd cell_6t
Xbit_r193_c129 bl_129 br_129 wl_193 vdd gnd cell_6t
Xbit_r194_c129 bl_129 br_129 wl_194 vdd gnd cell_6t
Xbit_r195_c129 bl_129 br_129 wl_195 vdd gnd cell_6t
Xbit_r196_c129 bl_129 br_129 wl_196 vdd gnd cell_6t
Xbit_r197_c129 bl_129 br_129 wl_197 vdd gnd cell_6t
Xbit_r198_c129 bl_129 br_129 wl_198 vdd gnd cell_6t
Xbit_r199_c129 bl_129 br_129 wl_199 vdd gnd cell_6t
Xbit_r200_c129 bl_129 br_129 wl_200 vdd gnd cell_6t
Xbit_r201_c129 bl_129 br_129 wl_201 vdd gnd cell_6t
Xbit_r202_c129 bl_129 br_129 wl_202 vdd gnd cell_6t
Xbit_r203_c129 bl_129 br_129 wl_203 vdd gnd cell_6t
Xbit_r204_c129 bl_129 br_129 wl_204 vdd gnd cell_6t
Xbit_r205_c129 bl_129 br_129 wl_205 vdd gnd cell_6t
Xbit_r206_c129 bl_129 br_129 wl_206 vdd gnd cell_6t
Xbit_r207_c129 bl_129 br_129 wl_207 vdd gnd cell_6t
Xbit_r208_c129 bl_129 br_129 wl_208 vdd gnd cell_6t
Xbit_r209_c129 bl_129 br_129 wl_209 vdd gnd cell_6t
Xbit_r210_c129 bl_129 br_129 wl_210 vdd gnd cell_6t
Xbit_r211_c129 bl_129 br_129 wl_211 vdd gnd cell_6t
Xbit_r212_c129 bl_129 br_129 wl_212 vdd gnd cell_6t
Xbit_r213_c129 bl_129 br_129 wl_213 vdd gnd cell_6t
Xbit_r214_c129 bl_129 br_129 wl_214 vdd gnd cell_6t
Xbit_r215_c129 bl_129 br_129 wl_215 vdd gnd cell_6t
Xbit_r216_c129 bl_129 br_129 wl_216 vdd gnd cell_6t
Xbit_r217_c129 bl_129 br_129 wl_217 vdd gnd cell_6t
Xbit_r218_c129 bl_129 br_129 wl_218 vdd gnd cell_6t
Xbit_r219_c129 bl_129 br_129 wl_219 vdd gnd cell_6t
Xbit_r220_c129 bl_129 br_129 wl_220 vdd gnd cell_6t
Xbit_r221_c129 bl_129 br_129 wl_221 vdd gnd cell_6t
Xbit_r222_c129 bl_129 br_129 wl_222 vdd gnd cell_6t
Xbit_r223_c129 bl_129 br_129 wl_223 vdd gnd cell_6t
Xbit_r224_c129 bl_129 br_129 wl_224 vdd gnd cell_6t
Xbit_r225_c129 bl_129 br_129 wl_225 vdd gnd cell_6t
Xbit_r226_c129 bl_129 br_129 wl_226 vdd gnd cell_6t
Xbit_r227_c129 bl_129 br_129 wl_227 vdd gnd cell_6t
Xbit_r228_c129 bl_129 br_129 wl_228 vdd gnd cell_6t
Xbit_r229_c129 bl_129 br_129 wl_229 vdd gnd cell_6t
Xbit_r230_c129 bl_129 br_129 wl_230 vdd gnd cell_6t
Xbit_r231_c129 bl_129 br_129 wl_231 vdd gnd cell_6t
Xbit_r232_c129 bl_129 br_129 wl_232 vdd gnd cell_6t
Xbit_r233_c129 bl_129 br_129 wl_233 vdd gnd cell_6t
Xbit_r234_c129 bl_129 br_129 wl_234 vdd gnd cell_6t
Xbit_r235_c129 bl_129 br_129 wl_235 vdd gnd cell_6t
Xbit_r236_c129 bl_129 br_129 wl_236 vdd gnd cell_6t
Xbit_r237_c129 bl_129 br_129 wl_237 vdd gnd cell_6t
Xbit_r238_c129 bl_129 br_129 wl_238 vdd gnd cell_6t
Xbit_r239_c129 bl_129 br_129 wl_239 vdd gnd cell_6t
Xbit_r240_c129 bl_129 br_129 wl_240 vdd gnd cell_6t
Xbit_r241_c129 bl_129 br_129 wl_241 vdd gnd cell_6t
Xbit_r242_c129 bl_129 br_129 wl_242 vdd gnd cell_6t
Xbit_r243_c129 bl_129 br_129 wl_243 vdd gnd cell_6t
Xbit_r244_c129 bl_129 br_129 wl_244 vdd gnd cell_6t
Xbit_r245_c129 bl_129 br_129 wl_245 vdd gnd cell_6t
Xbit_r246_c129 bl_129 br_129 wl_246 vdd gnd cell_6t
Xbit_r247_c129 bl_129 br_129 wl_247 vdd gnd cell_6t
Xbit_r248_c129 bl_129 br_129 wl_248 vdd gnd cell_6t
Xbit_r249_c129 bl_129 br_129 wl_249 vdd gnd cell_6t
Xbit_r250_c129 bl_129 br_129 wl_250 vdd gnd cell_6t
Xbit_r251_c129 bl_129 br_129 wl_251 vdd gnd cell_6t
Xbit_r252_c129 bl_129 br_129 wl_252 vdd gnd cell_6t
Xbit_r253_c129 bl_129 br_129 wl_253 vdd gnd cell_6t
Xbit_r254_c129 bl_129 br_129 wl_254 vdd gnd cell_6t
Xbit_r255_c129 bl_129 br_129 wl_255 vdd gnd cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd cell_6t
Xbit_r1_c130 bl_130 br_130 wl_1 vdd gnd cell_6t
Xbit_r2_c130 bl_130 br_130 wl_2 vdd gnd cell_6t
Xbit_r3_c130 bl_130 br_130 wl_3 vdd gnd cell_6t
Xbit_r4_c130 bl_130 br_130 wl_4 vdd gnd cell_6t
Xbit_r5_c130 bl_130 br_130 wl_5 vdd gnd cell_6t
Xbit_r6_c130 bl_130 br_130 wl_6 vdd gnd cell_6t
Xbit_r7_c130 bl_130 br_130 wl_7 vdd gnd cell_6t
Xbit_r8_c130 bl_130 br_130 wl_8 vdd gnd cell_6t
Xbit_r9_c130 bl_130 br_130 wl_9 vdd gnd cell_6t
Xbit_r10_c130 bl_130 br_130 wl_10 vdd gnd cell_6t
Xbit_r11_c130 bl_130 br_130 wl_11 vdd gnd cell_6t
Xbit_r12_c130 bl_130 br_130 wl_12 vdd gnd cell_6t
Xbit_r13_c130 bl_130 br_130 wl_13 vdd gnd cell_6t
Xbit_r14_c130 bl_130 br_130 wl_14 vdd gnd cell_6t
Xbit_r15_c130 bl_130 br_130 wl_15 vdd gnd cell_6t
Xbit_r16_c130 bl_130 br_130 wl_16 vdd gnd cell_6t
Xbit_r17_c130 bl_130 br_130 wl_17 vdd gnd cell_6t
Xbit_r18_c130 bl_130 br_130 wl_18 vdd gnd cell_6t
Xbit_r19_c130 bl_130 br_130 wl_19 vdd gnd cell_6t
Xbit_r20_c130 bl_130 br_130 wl_20 vdd gnd cell_6t
Xbit_r21_c130 bl_130 br_130 wl_21 vdd gnd cell_6t
Xbit_r22_c130 bl_130 br_130 wl_22 vdd gnd cell_6t
Xbit_r23_c130 bl_130 br_130 wl_23 vdd gnd cell_6t
Xbit_r24_c130 bl_130 br_130 wl_24 vdd gnd cell_6t
Xbit_r25_c130 bl_130 br_130 wl_25 vdd gnd cell_6t
Xbit_r26_c130 bl_130 br_130 wl_26 vdd gnd cell_6t
Xbit_r27_c130 bl_130 br_130 wl_27 vdd gnd cell_6t
Xbit_r28_c130 bl_130 br_130 wl_28 vdd gnd cell_6t
Xbit_r29_c130 bl_130 br_130 wl_29 vdd gnd cell_6t
Xbit_r30_c130 bl_130 br_130 wl_30 vdd gnd cell_6t
Xbit_r31_c130 bl_130 br_130 wl_31 vdd gnd cell_6t
Xbit_r32_c130 bl_130 br_130 wl_32 vdd gnd cell_6t
Xbit_r33_c130 bl_130 br_130 wl_33 vdd gnd cell_6t
Xbit_r34_c130 bl_130 br_130 wl_34 vdd gnd cell_6t
Xbit_r35_c130 bl_130 br_130 wl_35 vdd gnd cell_6t
Xbit_r36_c130 bl_130 br_130 wl_36 vdd gnd cell_6t
Xbit_r37_c130 bl_130 br_130 wl_37 vdd gnd cell_6t
Xbit_r38_c130 bl_130 br_130 wl_38 vdd gnd cell_6t
Xbit_r39_c130 bl_130 br_130 wl_39 vdd gnd cell_6t
Xbit_r40_c130 bl_130 br_130 wl_40 vdd gnd cell_6t
Xbit_r41_c130 bl_130 br_130 wl_41 vdd gnd cell_6t
Xbit_r42_c130 bl_130 br_130 wl_42 vdd gnd cell_6t
Xbit_r43_c130 bl_130 br_130 wl_43 vdd gnd cell_6t
Xbit_r44_c130 bl_130 br_130 wl_44 vdd gnd cell_6t
Xbit_r45_c130 bl_130 br_130 wl_45 vdd gnd cell_6t
Xbit_r46_c130 bl_130 br_130 wl_46 vdd gnd cell_6t
Xbit_r47_c130 bl_130 br_130 wl_47 vdd gnd cell_6t
Xbit_r48_c130 bl_130 br_130 wl_48 vdd gnd cell_6t
Xbit_r49_c130 bl_130 br_130 wl_49 vdd gnd cell_6t
Xbit_r50_c130 bl_130 br_130 wl_50 vdd gnd cell_6t
Xbit_r51_c130 bl_130 br_130 wl_51 vdd gnd cell_6t
Xbit_r52_c130 bl_130 br_130 wl_52 vdd gnd cell_6t
Xbit_r53_c130 bl_130 br_130 wl_53 vdd gnd cell_6t
Xbit_r54_c130 bl_130 br_130 wl_54 vdd gnd cell_6t
Xbit_r55_c130 bl_130 br_130 wl_55 vdd gnd cell_6t
Xbit_r56_c130 bl_130 br_130 wl_56 vdd gnd cell_6t
Xbit_r57_c130 bl_130 br_130 wl_57 vdd gnd cell_6t
Xbit_r58_c130 bl_130 br_130 wl_58 vdd gnd cell_6t
Xbit_r59_c130 bl_130 br_130 wl_59 vdd gnd cell_6t
Xbit_r60_c130 bl_130 br_130 wl_60 vdd gnd cell_6t
Xbit_r61_c130 bl_130 br_130 wl_61 vdd gnd cell_6t
Xbit_r62_c130 bl_130 br_130 wl_62 vdd gnd cell_6t
Xbit_r63_c130 bl_130 br_130 wl_63 vdd gnd cell_6t
Xbit_r64_c130 bl_130 br_130 wl_64 vdd gnd cell_6t
Xbit_r65_c130 bl_130 br_130 wl_65 vdd gnd cell_6t
Xbit_r66_c130 bl_130 br_130 wl_66 vdd gnd cell_6t
Xbit_r67_c130 bl_130 br_130 wl_67 vdd gnd cell_6t
Xbit_r68_c130 bl_130 br_130 wl_68 vdd gnd cell_6t
Xbit_r69_c130 bl_130 br_130 wl_69 vdd gnd cell_6t
Xbit_r70_c130 bl_130 br_130 wl_70 vdd gnd cell_6t
Xbit_r71_c130 bl_130 br_130 wl_71 vdd gnd cell_6t
Xbit_r72_c130 bl_130 br_130 wl_72 vdd gnd cell_6t
Xbit_r73_c130 bl_130 br_130 wl_73 vdd gnd cell_6t
Xbit_r74_c130 bl_130 br_130 wl_74 vdd gnd cell_6t
Xbit_r75_c130 bl_130 br_130 wl_75 vdd gnd cell_6t
Xbit_r76_c130 bl_130 br_130 wl_76 vdd gnd cell_6t
Xbit_r77_c130 bl_130 br_130 wl_77 vdd gnd cell_6t
Xbit_r78_c130 bl_130 br_130 wl_78 vdd gnd cell_6t
Xbit_r79_c130 bl_130 br_130 wl_79 vdd gnd cell_6t
Xbit_r80_c130 bl_130 br_130 wl_80 vdd gnd cell_6t
Xbit_r81_c130 bl_130 br_130 wl_81 vdd gnd cell_6t
Xbit_r82_c130 bl_130 br_130 wl_82 vdd gnd cell_6t
Xbit_r83_c130 bl_130 br_130 wl_83 vdd gnd cell_6t
Xbit_r84_c130 bl_130 br_130 wl_84 vdd gnd cell_6t
Xbit_r85_c130 bl_130 br_130 wl_85 vdd gnd cell_6t
Xbit_r86_c130 bl_130 br_130 wl_86 vdd gnd cell_6t
Xbit_r87_c130 bl_130 br_130 wl_87 vdd gnd cell_6t
Xbit_r88_c130 bl_130 br_130 wl_88 vdd gnd cell_6t
Xbit_r89_c130 bl_130 br_130 wl_89 vdd gnd cell_6t
Xbit_r90_c130 bl_130 br_130 wl_90 vdd gnd cell_6t
Xbit_r91_c130 bl_130 br_130 wl_91 vdd gnd cell_6t
Xbit_r92_c130 bl_130 br_130 wl_92 vdd gnd cell_6t
Xbit_r93_c130 bl_130 br_130 wl_93 vdd gnd cell_6t
Xbit_r94_c130 bl_130 br_130 wl_94 vdd gnd cell_6t
Xbit_r95_c130 bl_130 br_130 wl_95 vdd gnd cell_6t
Xbit_r96_c130 bl_130 br_130 wl_96 vdd gnd cell_6t
Xbit_r97_c130 bl_130 br_130 wl_97 vdd gnd cell_6t
Xbit_r98_c130 bl_130 br_130 wl_98 vdd gnd cell_6t
Xbit_r99_c130 bl_130 br_130 wl_99 vdd gnd cell_6t
Xbit_r100_c130 bl_130 br_130 wl_100 vdd gnd cell_6t
Xbit_r101_c130 bl_130 br_130 wl_101 vdd gnd cell_6t
Xbit_r102_c130 bl_130 br_130 wl_102 vdd gnd cell_6t
Xbit_r103_c130 bl_130 br_130 wl_103 vdd gnd cell_6t
Xbit_r104_c130 bl_130 br_130 wl_104 vdd gnd cell_6t
Xbit_r105_c130 bl_130 br_130 wl_105 vdd gnd cell_6t
Xbit_r106_c130 bl_130 br_130 wl_106 vdd gnd cell_6t
Xbit_r107_c130 bl_130 br_130 wl_107 vdd gnd cell_6t
Xbit_r108_c130 bl_130 br_130 wl_108 vdd gnd cell_6t
Xbit_r109_c130 bl_130 br_130 wl_109 vdd gnd cell_6t
Xbit_r110_c130 bl_130 br_130 wl_110 vdd gnd cell_6t
Xbit_r111_c130 bl_130 br_130 wl_111 vdd gnd cell_6t
Xbit_r112_c130 bl_130 br_130 wl_112 vdd gnd cell_6t
Xbit_r113_c130 bl_130 br_130 wl_113 vdd gnd cell_6t
Xbit_r114_c130 bl_130 br_130 wl_114 vdd gnd cell_6t
Xbit_r115_c130 bl_130 br_130 wl_115 vdd gnd cell_6t
Xbit_r116_c130 bl_130 br_130 wl_116 vdd gnd cell_6t
Xbit_r117_c130 bl_130 br_130 wl_117 vdd gnd cell_6t
Xbit_r118_c130 bl_130 br_130 wl_118 vdd gnd cell_6t
Xbit_r119_c130 bl_130 br_130 wl_119 vdd gnd cell_6t
Xbit_r120_c130 bl_130 br_130 wl_120 vdd gnd cell_6t
Xbit_r121_c130 bl_130 br_130 wl_121 vdd gnd cell_6t
Xbit_r122_c130 bl_130 br_130 wl_122 vdd gnd cell_6t
Xbit_r123_c130 bl_130 br_130 wl_123 vdd gnd cell_6t
Xbit_r124_c130 bl_130 br_130 wl_124 vdd gnd cell_6t
Xbit_r125_c130 bl_130 br_130 wl_125 vdd gnd cell_6t
Xbit_r126_c130 bl_130 br_130 wl_126 vdd gnd cell_6t
Xbit_r127_c130 bl_130 br_130 wl_127 vdd gnd cell_6t
Xbit_r128_c130 bl_130 br_130 wl_128 vdd gnd cell_6t
Xbit_r129_c130 bl_130 br_130 wl_129 vdd gnd cell_6t
Xbit_r130_c130 bl_130 br_130 wl_130 vdd gnd cell_6t
Xbit_r131_c130 bl_130 br_130 wl_131 vdd gnd cell_6t
Xbit_r132_c130 bl_130 br_130 wl_132 vdd gnd cell_6t
Xbit_r133_c130 bl_130 br_130 wl_133 vdd gnd cell_6t
Xbit_r134_c130 bl_130 br_130 wl_134 vdd gnd cell_6t
Xbit_r135_c130 bl_130 br_130 wl_135 vdd gnd cell_6t
Xbit_r136_c130 bl_130 br_130 wl_136 vdd gnd cell_6t
Xbit_r137_c130 bl_130 br_130 wl_137 vdd gnd cell_6t
Xbit_r138_c130 bl_130 br_130 wl_138 vdd gnd cell_6t
Xbit_r139_c130 bl_130 br_130 wl_139 vdd gnd cell_6t
Xbit_r140_c130 bl_130 br_130 wl_140 vdd gnd cell_6t
Xbit_r141_c130 bl_130 br_130 wl_141 vdd gnd cell_6t
Xbit_r142_c130 bl_130 br_130 wl_142 vdd gnd cell_6t
Xbit_r143_c130 bl_130 br_130 wl_143 vdd gnd cell_6t
Xbit_r144_c130 bl_130 br_130 wl_144 vdd gnd cell_6t
Xbit_r145_c130 bl_130 br_130 wl_145 vdd gnd cell_6t
Xbit_r146_c130 bl_130 br_130 wl_146 vdd gnd cell_6t
Xbit_r147_c130 bl_130 br_130 wl_147 vdd gnd cell_6t
Xbit_r148_c130 bl_130 br_130 wl_148 vdd gnd cell_6t
Xbit_r149_c130 bl_130 br_130 wl_149 vdd gnd cell_6t
Xbit_r150_c130 bl_130 br_130 wl_150 vdd gnd cell_6t
Xbit_r151_c130 bl_130 br_130 wl_151 vdd gnd cell_6t
Xbit_r152_c130 bl_130 br_130 wl_152 vdd gnd cell_6t
Xbit_r153_c130 bl_130 br_130 wl_153 vdd gnd cell_6t
Xbit_r154_c130 bl_130 br_130 wl_154 vdd gnd cell_6t
Xbit_r155_c130 bl_130 br_130 wl_155 vdd gnd cell_6t
Xbit_r156_c130 bl_130 br_130 wl_156 vdd gnd cell_6t
Xbit_r157_c130 bl_130 br_130 wl_157 vdd gnd cell_6t
Xbit_r158_c130 bl_130 br_130 wl_158 vdd gnd cell_6t
Xbit_r159_c130 bl_130 br_130 wl_159 vdd gnd cell_6t
Xbit_r160_c130 bl_130 br_130 wl_160 vdd gnd cell_6t
Xbit_r161_c130 bl_130 br_130 wl_161 vdd gnd cell_6t
Xbit_r162_c130 bl_130 br_130 wl_162 vdd gnd cell_6t
Xbit_r163_c130 bl_130 br_130 wl_163 vdd gnd cell_6t
Xbit_r164_c130 bl_130 br_130 wl_164 vdd gnd cell_6t
Xbit_r165_c130 bl_130 br_130 wl_165 vdd gnd cell_6t
Xbit_r166_c130 bl_130 br_130 wl_166 vdd gnd cell_6t
Xbit_r167_c130 bl_130 br_130 wl_167 vdd gnd cell_6t
Xbit_r168_c130 bl_130 br_130 wl_168 vdd gnd cell_6t
Xbit_r169_c130 bl_130 br_130 wl_169 vdd gnd cell_6t
Xbit_r170_c130 bl_130 br_130 wl_170 vdd gnd cell_6t
Xbit_r171_c130 bl_130 br_130 wl_171 vdd gnd cell_6t
Xbit_r172_c130 bl_130 br_130 wl_172 vdd gnd cell_6t
Xbit_r173_c130 bl_130 br_130 wl_173 vdd gnd cell_6t
Xbit_r174_c130 bl_130 br_130 wl_174 vdd gnd cell_6t
Xbit_r175_c130 bl_130 br_130 wl_175 vdd gnd cell_6t
Xbit_r176_c130 bl_130 br_130 wl_176 vdd gnd cell_6t
Xbit_r177_c130 bl_130 br_130 wl_177 vdd gnd cell_6t
Xbit_r178_c130 bl_130 br_130 wl_178 vdd gnd cell_6t
Xbit_r179_c130 bl_130 br_130 wl_179 vdd gnd cell_6t
Xbit_r180_c130 bl_130 br_130 wl_180 vdd gnd cell_6t
Xbit_r181_c130 bl_130 br_130 wl_181 vdd gnd cell_6t
Xbit_r182_c130 bl_130 br_130 wl_182 vdd gnd cell_6t
Xbit_r183_c130 bl_130 br_130 wl_183 vdd gnd cell_6t
Xbit_r184_c130 bl_130 br_130 wl_184 vdd gnd cell_6t
Xbit_r185_c130 bl_130 br_130 wl_185 vdd gnd cell_6t
Xbit_r186_c130 bl_130 br_130 wl_186 vdd gnd cell_6t
Xbit_r187_c130 bl_130 br_130 wl_187 vdd gnd cell_6t
Xbit_r188_c130 bl_130 br_130 wl_188 vdd gnd cell_6t
Xbit_r189_c130 bl_130 br_130 wl_189 vdd gnd cell_6t
Xbit_r190_c130 bl_130 br_130 wl_190 vdd gnd cell_6t
Xbit_r191_c130 bl_130 br_130 wl_191 vdd gnd cell_6t
Xbit_r192_c130 bl_130 br_130 wl_192 vdd gnd cell_6t
Xbit_r193_c130 bl_130 br_130 wl_193 vdd gnd cell_6t
Xbit_r194_c130 bl_130 br_130 wl_194 vdd gnd cell_6t
Xbit_r195_c130 bl_130 br_130 wl_195 vdd gnd cell_6t
Xbit_r196_c130 bl_130 br_130 wl_196 vdd gnd cell_6t
Xbit_r197_c130 bl_130 br_130 wl_197 vdd gnd cell_6t
Xbit_r198_c130 bl_130 br_130 wl_198 vdd gnd cell_6t
Xbit_r199_c130 bl_130 br_130 wl_199 vdd gnd cell_6t
Xbit_r200_c130 bl_130 br_130 wl_200 vdd gnd cell_6t
Xbit_r201_c130 bl_130 br_130 wl_201 vdd gnd cell_6t
Xbit_r202_c130 bl_130 br_130 wl_202 vdd gnd cell_6t
Xbit_r203_c130 bl_130 br_130 wl_203 vdd gnd cell_6t
Xbit_r204_c130 bl_130 br_130 wl_204 vdd gnd cell_6t
Xbit_r205_c130 bl_130 br_130 wl_205 vdd gnd cell_6t
Xbit_r206_c130 bl_130 br_130 wl_206 vdd gnd cell_6t
Xbit_r207_c130 bl_130 br_130 wl_207 vdd gnd cell_6t
Xbit_r208_c130 bl_130 br_130 wl_208 vdd gnd cell_6t
Xbit_r209_c130 bl_130 br_130 wl_209 vdd gnd cell_6t
Xbit_r210_c130 bl_130 br_130 wl_210 vdd gnd cell_6t
Xbit_r211_c130 bl_130 br_130 wl_211 vdd gnd cell_6t
Xbit_r212_c130 bl_130 br_130 wl_212 vdd gnd cell_6t
Xbit_r213_c130 bl_130 br_130 wl_213 vdd gnd cell_6t
Xbit_r214_c130 bl_130 br_130 wl_214 vdd gnd cell_6t
Xbit_r215_c130 bl_130 br_130 wl_215 vdd gnd cell_6t
Xbit_r216_c130 bl_130 br_130 wl_216 vdd gnd cell_6t
Xbit_r217_c130 bl_130 br_130 wl_217 vdd gnd cell_6t
Xbit_r218_c130 bl_130 br_130 wl_218 vdd gnd cell_6t
Xbit_r219_c130 bl_130 br_130 wl_219 vdd gnd cell_6t
Xbit_r220_c130 bl_130 br_130 wl_220 vdd gnd cell_6t
Xbit_r221_c130 bl_130 br_130 wl_221 vdd gnd cell_6t
Xbit_r222_c130 bl_130 br_130 wl_222 vdd gnd cell_6t
Xbit_r223_c130 bl_130 br_130 wl_223 vdd gnd cell_6t
Xbit_r224_c130 bl_130 br_130 wl_224 vdd gnd cell_6t
Xbit_r225_c130 bl_130 br_130 wl_225 vdd gnd cell_6t
Xbit_r226_c130 bl_130 br_130 wl_226 vdd gnd cell_6t
Xbit_r227_c130 bl_130 br_130 wl_227 vdd gnd cell_6t
Xbit_r228_c130 bl_130 br_130 wl_228 vdd gnd cell_6t
Xbit_r229_c130 bl_130 br_130 wl_229 vdd gnd cell_6t
Xbit_r230_c130 bl_130 br_130 wl_230 vdd gnd cell_6t
Xbit_r231_c130 bl_130 br_130 wl_231 vdd gnd cell_6t
Xbit_r232_c130 bl_130 br_130 wl_232 vdd gnd cell_6t
Xbit_r233_c130 bl_130 br_130 wl_233 vdd gnd cell_6t
Xbit_r234_c130 bl_130 br_130 wl_234 vdd gnd cell_6t
Xbit_r235_c130 bl_130 br_130 wl_235 vdd gnd cell_6t
Xbit_r236_c130 bl_130 br_130 wl_236 vdd gnd cell_6t
Xbit_r237_c130 bl_130 br_130 wl_237 vdd gnd cell_6t
Xbit_r238_c130 bl_130 br_130 wl_238 vdd gnd cell_6t
Xbit_r239_c130 bl_130 br_130 wl_239 vdd gnd cell_6t
Xbit_r240_c130 bl_130 br_130 wl_240 vdd gnd cell_6t
Xbit_r241_c130 bl_130 br_130 wl_241 vdd gnd cell_6t
Xbit_r242_c130 bl_130 br_130 wl_242 vdd gnd cell_6t
Xbit_r243_c130 bl_130 br_130 wl_243 vdd gnd cell_6t
Xbit_r244_c130 bl_130 br_130 wl_244 vdd gnd cell_6t
Xbit_r245_c130 bl_130 br_130 wl_245 vdd gnd cell_6t
Xbit_r246_c130 bl_130 br_130 wl_246 vdd gnd cell_6t
Xbit_r247_c130 bl_130 br_130 wl_247 vdd gnd cell_6t
Xbit_r248_c130 bl_130 br_130 wl_248 vdd gnd cell_6t
Xbit_r249_c130 bl_130 br_130 wl_249 vdd gnd cell_6t
Xbit_r250_c130 bl_130 br_130 wl_250 vdd gnd cell_6t
Xbit_r251_c130 bl_130 br_130 wl_251 vdd gnd cell_6t
Xbit_r252_c130 bl_130 br_130 wl_252 vdd gnd cell_6t
Xbit_r253_c130 bl_130 br_130 wl_253 vdd gnd cell_6t
Xbit_r254_c130 bl_130 br_130 wl_254 vdd gnd cell_6t
Xbit_r255_c130 bl_130 br_130 wl_255 vdd gnd cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd cell_6t
Xbit_r1_c131 bl_131 br_131 wl_1 vdd gnd cell_6t
Xbit_r2_c131 bl_131 br_131 wl_2 vdd gnd cell_6t
Xbit_r3_c131 bl_131 br_131 wl_3 vdd gnd cell_6t
Xbit_r4_c131 bl_131 br_131 wl_4 vdd gnd cell_6t
Xbit_r5_c131 bl_131 br_131 wl_5 vdd gnd cell_6t
Xbit_r6_c131 bl_131 br_131 wl_6 vdd gnd cell_6t
Xbit_r7_c131 bl_131 br_131 wl_7 vdd gnd cell_6t
Xbit_r8_c131 bl_131 br_131 wl_8 vdd gnd cell_6t
Xbit_r9_c131 bl_131 br_131 wl_9 vdd gnd cell_6t
Xbit_r10_c131 bl_131 br_131 wl_10 vdd gnd cell_6t
Xbit_r11_c131 bl_131 br_131 wl_11 vdd gnd cell_6t
Xbit_r12_c131 bl_131 br_131 wl_12 vdd gnd cell_6t
Xbit_r13_c131 bl_131 br_131 wl_13 vdd gnd cell_6t
Xbit_r14_c131 bl_131 br_131 wl_14 vdd gnd cell_6t
Xbit_r15_c131 bl_131 br_131 wl_15 vdd gnd cell_6t
Xbit_r16_c131 bl_131 br_131 wl_16 vdd gnd cell_6t
Xbit_r17_c131 bl_131 br_131 wl_17 vdd gnd cell_6t
Xbit_r18_c131 bl_131 br_131 wl_18 vdd gnd cell_6t
Xbit_r19_c131 bl_131 br_131 wl_19 vdd gnd cell_6t
Xbit_r20_c131 bl_131 br_131 wl_20 vdd gnd cell_6t
Xbit_r21_c131 bl_131 br_131 wl_21 vdd gnd cell_6t
Xbit_r22_c131 bl_131 br_131 wl_22 vdd gnd cell_6t
Xbit_r23_c131 bl_131 br_131 wl_23 vdd gnd cell_6t
Xbit_r24_c131 bl_131 br_131 wl_24 vdd gnd cell_6t
Xbit_r25_c131 bl_131 br_131 wl_25 vdd gnd cell_6t
Xbit_r26_c131 bl_131 br_131 wl_26 vdd gnd cell_6t
Xbit_r27_c131 bl_131 br_131 wl_27 vdd gnd cell_6t
Xbit_r28_c131 bl_131 br_131 wl_28 vdd gnd cell_6t
Xbit_r29_c131 bl_131 br_131 wl_29 vdd gnd cell_6t
Xbit_r30_c131 bl_131 br_131 wl_30 vdd gnd cell_6t
Xbit_r31_c131 bl_131 br_131 wl_31 vdd gnd cell_6t
Xbit_r32_c131 bl_131 br_131 wl_32 vdd gnd cell_6t
Xbit_r33_c131 bl_131 br_131 wl_33 vdd gnd cell_6t
Xbit_r34_c131 bl_131 br_131 wl_34 vdd gnd cell_6t
Xbit_r35_c131 bl_131 br_131 wl_35 vdd gnd cell_6t
Xbit_r36_c131 bl_131 br_131 wl_36 vdd gnd cell_6t
Xbit_r37_c131 bl_131 br_131 wl_37 vdd gnd cell_6t
Xbit_r38_c131 bl_131 br_131 wl_38 vdd gnd cell_6t
Xbit_r39_c131 bl_131 br_131 wl_39 vdd gnd cell_6t
Xbit_r40_c131 bl_131 br_131 wl_40 vdd gnd cell_6t
Xbit_r41_c131 bl_131 br_131 wl_41 vdd gnd cell_6t
Xbit_r42_c131 bl_131 br_131 wl_42 vdd gnd cell_6t
Xbit_r43_c131 bl_131 br_131 wl_43 vdd gnd cell_6t
Xbit_r44_c131 bl_131 br_131 wl_44 vdd gnd cell_6t
Xbit_r45_c131 bl_131 br_131 wl_45 vdd gnd cell_6t
Xbit_r46_c131 bl_131 br_131 wl_46 vdd gnd cell_6t
Xbit_r47_c131 bl_131 br_131 wl_47 vdd gnd cell_6t
Xbit_r48_c131 bl_131 br_131 wl_48 vdd gnd cell_6t
Xbit_r49_c131 bl_131 br_131 wl_49 vdd gnd cell_6t
Xbit_r50_c131 bl_131 br_131 wl_50 vdd gnd cell_6t
Xbit_r51_c131 bl_131 br_131 wl_51 vdd gnd cell_6t
Xbit_r52_c131 bl_131 br_131 wl_52 vdd gnd cell_6t
Xbit_r53_c131 bl_131 br_131 wl_53 vdd gnd cell_6t
Xbit_r54_c131 bl_131 br_131 wl_54 vdd gnd cell_6t
Xbit_r55_c131 bl_131 br_131 wl_55 vdd gnd cell_6t
Xbit_r56_c131 bl_131 br_131 wl_56 vdd gnd cell_6t
Xbit_r57_c131 bl_131 br_131 wl_57 vdd gnd cell_6t
Xbit_r58_c131 bl_131 br_131 wl_58 vdd gnd cell_6t
Xbit_r59_c131 bl_131 br_131 wl_59 vdd gnd cell_6t
Xbit_r60_c131 bl_131 br_131 wl_60 vdd gnd cell_6t
Xbit_r61_c131 bl_131 br_131 wl_61 vdd gnd cell_6t
Xbit_r62_c131 bl_131 br_131 wl_62 vdd gnd cell_6t
Xbit_r63_c131 bl_131 br_131 wl_63 vdd gnd cell_6t
Xbit_r64_c131 bl_131 br_131 wl_64 vdd gnd cell_6t
Xbit_r65_c131 bl_131 br_131 wl_65 vdd gnd cell_6t
Xbit_r66_c131 bl_131 br_131 wl_66 vdd gnd cell_6t
Xbit_r67_c131 bl_131 br_131 wl_67 vdd gnd cell_6t
Xbit_r68_c131 bl_131 br_131 wl_68 vdd gnd cell_6t
Xbit_r69_c131 bl_131 br_131 wl_69 vdd gnd cell_6t
Xbit_r70_c131 bl_131 br_131 wl_70 vdd gnd cell_6t
Xbit_r71_c131 bl_131 br_131 wl_71 vdd gnd cell_6t
Xbit_r72_c131 bl_131 br_131 wl_72 vdd gnd cell_6t
Xbit_r73_c131 bl_131 br_131 wl_73 vdd gnd cell_6t
Xbit_r74_c131 bl_131 br_131 wl_74 vdd gnd cell_6t
Xbit_r75_c131 bl_131 br_131 wl_75 vdd gnd cell_6t
Xbit_r76_c131 bl_131 br_131 wl_76 vdd gnd cell_6t
Xbit_r77_c131 bl_131 br_131 wl_77 vdd gnd cell_6t
Xbit_r78_c131 bl_131 br_131 wl_78 vdd gnd cell_6t
Xbit_r79_c131 bl_131 br_131 wl_79 vdd gnd cell_6t
Xbit_r80_c131 bl_131 br_131 wl_80 vdd gnd cell_6t
Xbit_r81_c131 bl_131 br_131 wl_81 vdd gnd cell_6t
Xbit_r82_c131 bl_131 br_131 wl_82 vdd gnd cell_6t
Xbit_r83_c131 bl_131 br_131 wl_83 vdd gnd cell_6t
Xbit_r84_c131 bl_131 br_131 wl_84 vdd gnd cell_6t
Xbit_r85_c131 bl_131 br_131 wl_85 vdd gnd cell_6t
Xbit_r86_c131 bl_131 br_131 wl_86 vdd gnd cell_6t
Xbit_r87_c131 bl_131 br_131 wl_87 vdd gnd cell_6t
Xbit_r88_c131 bl_131 br_131 wl_88 vdd gnd cell_6t
Xbit_r89_c131 bl_131 br_131 wl_89 vdd gnd cell_6t
Xbit_r90_c131 bl_131 br_131 wl_90 vdd gnd cell_6t
Xbit_r91_c131 bl_131 br_131 wl_91 vdd gnd cell_6t
Xbit_r92_c131 bl_131 br_131 wl_92 vdd gnd cell_6t
Xbit_r93_c131 bl_131 br_131 wl_93 vdd gnd cell_6t
Xbit_r94_c131 bl_131 br_131 wl_94 vdd gnd cell_6t
Xbit_r95_c131 bl_131 br_131 wl_95 vdd gnd cell_6t
Xbit_r96_c131 bl_131 br_131 wl_96 vdd gnd cell_6t
Xbit_r97_c131 bl_131 br_131 wl_97 vdd gnd cell_6t
Xbit_r98_c131 bl_131 br_131 wl_98 vdd gnd cell_6t
Xbit_r99_c131 bl_131 br_131 wl_99 vdd gnd cell_6t
Xbit_r100_c131 bl_131 br_131 wl_100 vdd gnd cell_6t
Xbit_r101_c131 bl_131 br_131 wl_101 vdd gnd cell_6t
Xbit_r102_c131 bl_131 br_131 wl_102 vdd gnd cell_6t
Xbit_r103_c131 bl_131 br_131 wl_103 vdd gnd cell_6t
Xbit_r104_c131 bl_131 br_131 wl_104 vdd gnd cell_6t
Xbit_r105_c131 bl_131 br_131 wl_105 vdd gnd cell_6t
Xbit_r106_c131 bl_131 br_131 wl_106 vdd gnd cell_6t
Xbit_r107_c131 bl_131 br_131 wl_107 vdd gnd cell_6t
Xbit_r108_c131 bl_131 br_131 wl_108 vdd gnd cell_6t
Xbit_r109_c131 bl_131 br_131 wl_109 vdd gnd cell_6t
Xbit_r110_c131 bl_131 br_131 wl_110 vdd gnd cell_6t
Xbit_r111_c131 bl_131 br_131 wl_111 vdd gnd cell_6t
Xbit_r112_c131 bl_131 br_131 wl_112 vdd gnd cell_6t
Xbit_r113_c131 bl_131 br_131 wl_113 vdd gnd cell_6t
Xbit_r114_c131 bl_131 br_131 wl_114 vdd gnd cell_6t
Xbit_r115_c131 bl_131 br_131 wl_115 vdd gnd cell_6t
Xbit_r116_c131 bl_131 br_131 wl_116 vdd gnd cell_6t
Xbit_r117_c131 bl_131 br_131 wl_117 vdd gnd cell_6t
Xbit_r118_c131 bl_131 br_131 wl_118 vdd gnd cell_6t
Xbit_r119_c131 bl_131 br_131 wl_119 vdd gnd cell_6t
Xbit_r120_c131 bl_131 br_131 wl_120 vdd gnd cell_6t
Xbit_r121_c131 bl_131 br_131 wl_121 vdd gnd cell_6t
Xbit_r122_c131 bl_131 br_131 wl_122 vdd gnd cell_6t
Xbit_r123_c131 bl_131 br_131 wl_123 vdd gnd cell_6t
Xbit_r124_c131 bl_131 br_131 wl_124 vdd gnd cell_6t
Xbit_r125_c131 bl_131 br_131 wl_125 vdd gnd cell_6t
Xbit_r126_c131 bl_131 br_131 wl_126 vdd gnd cell_6t
Xbit_r127_c131 bl_131 br_131 wl_127 vdd gnd cell_6t
Xbit_r128_c131 bl_131 br_131 wl_128 vdd gnd cell_6t
Xbit_r129_c131 bl_131 br_131 wl_129 vdd gnd cell_6t
Xbit_r130_c131 bl_131 br_131 wl_130 vdd gnd cell_6t
Xbit_r131_c131 bl_131 br_131 wl_131 vdd gnd cell_6t
Xbit_r132_c131 bl_131 br_131 wl_132 vdd gnd cell_6t
Xbit_r133_c131 bl_131 br_131 wl_133 vdd gnd cell_6t
Xbit_r134_c131 bl_131 br_131 wl_134 vdd gnd cell_6t
Xbit_r135_c131 bl_131 br_131 wl_135 vdd gnd cell_6t
Xbit_r136_c131 bl_131 br_131 wl_136 vdd gnd cell_6t
Xbit_r137_c131 bl_131 br_131 wl_137 vdd gnd cell_6t
Xbit_r138_c131 bl_131 br_131 wl_138 vdd gnd cell_6t
Xbit_r139_c131 bl_131 br_131 wl_139 vdd gnd cell_6t
Xbit_r140_c131 bl_131 br_131 wl_140 vdd gnd cell_6t
Xbit_r141_c131 bl_131 br_131 wl_141 vdd gnd cell_6t
Xbit_r142_c131 bl_131 br_131 wl_142 vdd gnd cell_6t
Xbit_r143_c131 bl_131 br_131 wl_143 vdd gnd cell_6t
Xbit_r144_c131 bl_131 br_131 wl_144 vdd gnd cell_6t
Xbit_r145_c131 bl_131 br_131 wl_145 vdd gnd cell_6t
Xbit_r146_c131 bl_131 br_131 wl_146 vdd gnd cell_6t
Xbit_r147_c131 bl_131 br_131 wl_147 vdd gnd cell_6t
Xbit_r148_c131 bl_131 br_131 wl_148 vdd gnd cell_6t
Xbit_r149_c131 bl_131 br_131 wl_149 vdd gnd cell_6t
Xbit_r150_c131 bl_131 br_131 wl_150 vdd gnd cell_6t
Xbit_r151_c131 bl_131 br_131 wl_151 vdd gnd cell_6t
Xbit_r152_c131 bl_131 br_131 wl_152 vdd gnd cell_6t
Xbit_r153_c131 bl_131 br_131 wl_153 vdd gnd cell_6t
Xbit_r154_c131 bl_131 br_131 wl_154 vdd gnd cell_6t
Xbit_r155_c131 bl_131 br_131 wl_155 vdd gnd cell_6t
Xbit_r156_c131 bl_131 br_131 wl_156 vdd gnd cell_6t
Xbit_r157_c131 bl_131 br_131 wl_157 vdd gnd cell_6t
Xbit_r158_c131 bl_131 br_131 wl_158 vdd gnd cell_6t
Xbit_r159_c131 bl_131 br_131 wl_159 vdd gnd cell_6t
Xbit_r160_c131 bl_131 br_131 wl_160 vdd gnd cell_6t
Xbit_r161_c131 bl_131 br_131 wl_161 vdd gnd cell_6t
Xbit_r162_c131 bl_131 br_131 wl_162 vdd gnd cell_6t
Xbit_r163_c131 bl_131 br_131 wl_163 vdd gnd cell_6t
Xbit_r164_c131 bl_131 br_131 wl_164 vdd gnd cell_6t
Xbit_r165_c131 bl_131 br_131 wl_165 vdd gnd cell_6t
Xbit_r166_c131 bl_131 br_131 wl_166 vdd gnd cell_6t
Xbit_r167_c131 bl_131 br_131 wl_167 vdd gnd cell_6t
Xbit_r168_c131 bl_131 br_131 wl_168 vdd gnd cell_6t
Xbit_r169_c131 bl_131 br_131 wl_169 vdd gnd cell_6t
Xbit_r170_c131 bl_131 br_131 wl_170 vdd gnd cell_6t
Xbit_r171_c131 bl_131 br_131 wl_171 vdd gnd cell_6t
Xbit_r172_c131 bl_131 br_131 wl_172 vdd gnd cell_6t
Xbit_r173_c131 bl_131 br_131 wl_173 vdd gnd cell_6t
Xbit_r174_c131 bl_131 br_131 wl_174 vdd gnd cell_6t
Xbit_r175_c131 bl_131 br_131 wl_175 vdd gnd cell_6t
Xbit_r176_c131 bl_131 br_131 wl_176 vdd gnd cell_6t
Xbit_r177_c131 bl_131 br_131 wl_177 vdd gnd cell_6t
Xbit_r178_c131 bl_131 br_131 wl_178 vdd gnd cell_6t
Xbit_r179_c131 bl_131 br_131 wl_179 vdd gnd cell_6t
Xbit_r180_c131 bl_131 br_131 wl_180 vdd gnd cell_6t
Xbit_r181_c131 bl_131 br_131 wl_181 vdd gnd cell_6t
Xbit_r182_c131 bl_131 br_131 wl_182 vdd gnd cell_6t
Xbit_r183_c131 bl_131 br_131 wl_183 vdd gnd cell_6t
Xbit_r184_c131 bl_131 br_131 wl_184 vdd gnd cell_6t
Xbit_r185_c131 bl_131 br_131 wl_185 vdd gnd cell_6t
Xbit_r186_c131 bl_131 br_131 wl_186 vdd gnd cell_6t
Xbit_r187_c131 bl_131 br_131 wl_187 vdd gnd cell_6t
Xbit_r188_c131 bl_131 br_131 wl_188 vdd gnd cell_6t
Xbit_r189_c131 bl_131 br_131 wl_189 vdd gnd cell_6t
Xbit_r190_c131 bl_131 br_131 wl_190 vdd gnd cell_6t
Xbit_r191_c131 bl_131 br_131 wl_191 vdd gnd cell_6t
Xbit_r192_c131 bl_131 br_131 wl_192 vdd gnd cell_6t
Xbit_r193_c131 bl_131 br_131 wl_193 vdd gnd cell_6t
Xbit_r194_c131 bl_131 br_131 wl_194 vdd gnd cell_6t
Xbit_r195_c131 bl_131 br_131 wl_195 vdd gnd cell_6t
Xbit_r196_c131 bl_131 br_131 wl_196 vdd gnd cell_6t
Xbit_r197_c131 bl_131 br_131 wl_197 vdd gnd cell_6t
Xbit_r198_c131 bl_131 br_131 wl_198 vdd gnd cell_6t
Xbit_r199_c131 bl_131 br_131 wl_199 vdd gnd cell_6t
Xbit_r200_c131 bl_131 br_131 wl_200 vdd gnd cell_6t
Xbit_r201_c131 bl_131 br_131 wl_201 vdd gnd cell_6t
Xbit_r202_c131 bl_131 br_131 wl_202 vdd gnd cell_6t
Xbit_r203_c131 bl_131 br_131 wl_203 vdd gnd cell_6t
Xbit_r204_c131 bl_131 br_131 wl_204 vdd gnd cell_6t
Xbit_r205_c131 bl_131 br_131 wl_205 vdd gnd cell_6t
Xbit_r206_c131 bl_131 br_131 wl_206 vdd gnd cell_6t
Xbit_r207_c131 bl_131 br_131 wl_207 vdd gnd cell_6t
Xbit_r208_c131 bl_131 br_131 wl_208 vdd gnd cell_6t
Xbit_r209_c131 bl_131 br_131 wl_209 vdd gnd cell_6t
Xbit_r210_c131 bl_131 br_131 wl_210 vdd gnd cell_6t
Xbit_r211_c131 bl_131 br_131 wl_211 vdd gnd cell_6t
Xbit_r212_c131 bl_131 br_131 wl_212 vdd gnd cell_6t
Xbit_r213_c131 bl_131 br_131 wl_213 vdd gnd cell_6t
Xbit_r214_c131 bl_131 br_131 wl_214 vdd gnd cell_6t
Xbit_r215_c131 bl_131 br_131 wl_215 vdd gnd cell_6t
Xbit_r216_c131 bl_131 br_131 wl_216 vdd gnd cell_6t
Xbit_r217_c131 bl_131 br_131 wl_217 vdd gnd cell_6t
Xbit_r218_c131 bl_131 br_131 wl_218 vdd gnd cell_6t
Xbit_r219_c131 bl_131 br_131 wl_219 vdd gnd cell_6t
Xbit_r220_c131 bl_131 br_131 wl_220 vdd gnd cell_6t
Xbit_r221_c131 bl_131 br_131 wl_221 vdd gnd cell_6t
Xbit_r222_c131 bl_131 br_131 wl_222 vdd gnd cell_6t
Xbit_r223_c131 bl_131 br_131 wl_223 vdd gnd cell_6t
Xbit_r224_c131 bl_131 br_131 wl_224 vdd gnd cell_6t
Xbit_r225_c131 bl_131 br_131 wl_225 vdd gnd cell_6t
Xbit_r226_c131 bl_131 br_131 wl_226 vdd gnd cell_6t
Xbit_r227_c131 bl_131 br_131 wl_227 vdd gnd cell_6t
Xbit_r228_c131 bl_131 br_131 wl_228 vdd gnd cell_6t
Xbit_r229_c131 bl_131 br_131 wl_229 vdd gnd cell_6t
Xbit_r230_c131 bl_131 br_131 wl_230 vdd gnd cell_6t
Xbit_r231_c131 bl_131 br_131 wl_231 vdd gnd cell_6t
Xbit_r232_c131 bl_131 br_131 wl_232 vdd gnd cell_6t
Xbit_r233_c131 bl_131 br_131 wl_233 vdd gnd cell_6t
Xbit_r234_c131 bl_131 br_131 wl_234 vdd gnd cell_6t
Xbit_r235_c131 bl_131 br_131 wl_235 vdd gnd cell_6t
Xbit_r236_c131 bl_131 br_131 wl_236 vdd gnd cell_6t
Xbit_r237_c131 bl_131 br_131 wl_237 vdd gnd cell_6t
Xbit_r238_c131 bl_131 br_131 wl_238 vdd gnd cell_6t
Xbit_r239_c131 bl_131 br_131 wl_239 vdd gnd cell_6t
Xbit_r240_c131 bl_131 br_131 wl_240 vdd gnd cell_6t
Xbit_r241_c131 bl_131 br_131 wl_241 vdd gnd cell_6t
Xbit_r242_c131 bl_131 br_131 wl_242 vdd gnd cell_6t
Xbit_r243_c131 bl_131 br_131 wl_243 vdd gnd cell_6t
Xbit_r244_c131 bl_131 br_131 wl_244 vdd gnd cell_6t
Xbit_r245_c131 bl_131 br_131 wl_245 vdd gnd cell_6t
Xbit_r246_c131 bl_131 br_131 wl_246 vdd gnd cell_6t
Xbit_r247_c131 bl_131 br_131 wl_247 vdd gnd cell_6t
Xbit_r248_c131 bl_131 br_131 wl_248 vdd gnd cell_6t
Xbit_r249_c131 bl_131 br_131 wl_249 vdd gnd cell_6t
Xbit_r250_c131 bl_131 br_131 wl_250 vdd gnd cell_6t
Xbit_r251_c131 bl_131 br_131 wl_251 vdd gnd cell_6t
Xbit_r252_c131 bl_131 br_131 wl_252 vdd gnd cell_6t
Xbit_r253_c131 bl_131 br_131 wl_253 vdd gnd cell_6t
Xbit_r254_c131 bl_131 br_131 wl_254 vdd gnd cell_6t
Xbit_r255_c131 bl_131 br_131 wl_255 vdd gnd cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd cell_6t
Xbit_r1_c132 bl_132 br_132 wl_1 vdd gnd cell_6t
Xbit_r2_c132 bl_132 br_132 wl_2 vdd gnd cell_6t
Xbit_r3_c132 bl_132 br_132 wl_3 vdd gnd cell_6t
Xbit_r4_c132 bl_132 br_132 wl_4 vdd gnd cell_6t
Xbit_r5_c132 bl_132 br_132 wl_5 vdd gnd cell_6t
Xbit_r6_c132 bl_132 br_132 wl_6 vdd gnd cell_6t
Xbit_r7_c132 bl_132 br_132 wl_7 vdd gnd cell_6t
Xbit_r8_c132 bl_132 br_132 wl_8 vdd gnd cell_6t
Xbit_r9_c132 bl_132 br_132 wl_9 vdd gnd cell_6t
Xbit_r10_c132 bl_132 br_132 wl_10 vdd gnd cell_6t
Xbit_r11_c132 bl_132 br_132 wl_11 vdd gnd cell_6t
Xbit_r12_c132 bl_132 br_132 wl_12 vdd gnd cell_6t
Xbit_r13_c132 bl_132 br_132 wl_13 vdd gnd cell_6t
Xbit_r14_c132 bl_132 br_132 wl_14 vdd gnd cell_6t
Xbit_r15_c132 bl_132 br_132 wl_15 vdd gnd cell_6t
Xbit_r16_c132 bl_132 br_132 wl_16 vdd gnd cell_6t
Xbit_r17_c132 bl_132 br_132 wl_17 vdd gnd cell_6t
Xbit_r18_c132 bl_132 br_132 wl_18 vdd gnd cell_6t
Xbit_r19_c132 bl_132 br_132 wl_19 vdd gnd cell_6t
Xbit_r20_c132 bl_132 br_132 wl_20 vdd gnd cell_6t
Xbit_r21_c132 bl_132 br_132 wl_21 vdd gnd cell_6t
Xbit_r22_c132 bl_132 br_132 wl_22 vdd gnd cell_6t
Xbit_r23_c132 bl_132 br_132 wl_23 vdd gnd cell_6t
Xbit_r24_c132 bl_132 br_132 wl_24 vdd gnd cell_6t
Xbit_r25_c132 bl_132 br_132 wl_25 vdd gnd cell_6t
Xbit_r26_c132 bl_132 br_132 wl_26 vdd gnd cell_6t
Xbit_r27_c132 bl_132 br_132 wl_27 vdd gnd cell_6t
Xbit_r28_c132 bl_132 br_132 wl_28 vdd gnd cell_6t
Xbit_r29_c132 bl_132 br_132 wl_29 vdd gnd cell_6t
Xbit_r30_c132 bl_132 br_132 wl_30 vdd gnd cell_6t
Xbit_r31_c132 bl_132 br_132 wl_31 vdd gnd cell_6t
Xbit_r32_c132 bl_132 br_132 wl_32 vdd gnd cell_6t
Xbit_r33_c132 bl_132 br_132 wl_33 vdd gnd cell_6t
Xbit_r34_c132 bl_132 br_132 wl_34 vdd gnd cell_6t
Xbit_r35_c132 bl_132 br_132 wl_35 vdd gnd cell_6t
Xbit_r36_c132 bl_132 br_132 wl_36 vdd gnd cell_6t
Xbit_r37_c132 bl_132 br_132 wl_37 vdd gnd cell_6t
Xbit_r38_c132 bl_132 br_132 wl_38 vdd gnd cell_6t
Xbit_r39_c132 bl_132 br_132 wl_39 vdd gnd cell_6t
Xbit_r40_c132 bl_132 br_132 wl_40 vdd gnd cell_6t
Xbit_r41_c132 bl_132 br_132 wl_41 vdd gnd cell_6t
Xbit_r42_c132 bl_132 br_132 wl_42 vdd gnd cell_6t
Xbit_r43_c132 bl_132 br_132 wl_43 vdd gnd cell_6t
Xbit_r44_c132 bl_132 br_132 wl_44 vdd gnd cell_6t
Xbit_r45_c132 bl_132 br_132 wl_45 vdd gnd cell_6t
Xbit_r46_c132 bl_132 br_132 wl_46 vdd gnd cell_6t
Xbit_r47_c132 bl_132 br_132 wl_47 vdd gnd cell_6t
Xbit_r48_c132 bl_132 br_132 wl_48 vdd gnd cell_6t
Xbit_r49_c132 bl_132 br_132 wl_49 vdd gnd cell_6t
Xbit_r50_c132 bl_132 br_132 wl_50 vdd gnd cell_6t
Xbit_r51_c132 bl_132 br_132 wl_51 vdd gnd cell_6t
Xbit_r52_c132 bl_132 br_132 wl_52 vdd gnd cell_6t
Xbit_r53_c132 bl_132 br_132 wl_53 vdd gnd cell_6t
Xbit_r54_c132 bl_132 br_132 wl_54 vdd gnd cell_6t
Xbit_r55_c132 bl_132 br_132 wl_55 vdd gnd cell_6t
Xbit_r56_c132 bl_132 br_132 wl_56 vdd gnd cell_6t
Xbit_r57_c132 bl_132 br_132 wl_57 vdd gnd cell_6t
Xbit_r58_c132 bl_132 br_132 wl_58 vdd gnd cell_6t
Xbit_r59_c132 bl_132 br_132 wl_59 vdd gnd cell_6t
Xbit_r60_c132 bl_132 br_132 wl_60 vdd gnd cell_6t
Xbit_r61_c132 bl_132 br_132 wl_61 vdd gnd cell_6t
Xbit_r62_c132 bl_132 br_132 wl_62 vdd gnd cell_6t
Xbit_r63_c132 bl_132 br_132 wl_63 vdd gnd cell_6t
Xbit_r64_c132 bl_132 br_132 wl_64 vdd gnd cell_6t
Xbit_r65_c132 bl_132 br_132 wl_65 vdd gnd cell_6t
Xbit_r66_c132 bl_132 br_132 wl_66 vdd gnd cell_6t
Xbit_r67_c132 bl_132 br_132 wl_67 vdd gnd cell_6t
Xbit_r68_c132 bl_132 br_132 wl_68 vdd gnd cell_6t
Xbit_r69_c132 bl_132 br_132 wl_69 vdd gnd cell_6t
Xbit_r70_c132 bl_132 br_132 wl_70 vdd gnd cell_6t
Xbit_r71_c132 bl_132 br_132 wl_71 vdd gnd cell_6t
Xbit_r72_c132 bl_132 br_132 wl_72 vdd gnd cell_6t
Xbit_r73_c132 bl_132 br_132 wl_73 vdd gnd cell_6t
Xbit_r74_c132 bl_132 br_132 wl_74 vdd gnd cell_6t
Xbit_r75_c132 bl_132 br_132 wl_75 vdd gnd cell_6t
Xbit_r76_c132 bl_132 br_132 wl_76 vdd gnd cell_6t
Xbit_r77_c132 bl_132 br_132 wl_77 vdd gnd cell_6t
Xbit_r78_c132 bl_132 br_132 wl_78 vdd gnd cell_6t
Xbit_r79_c132 bl_132 br_132 wl_79 vdd gnd cell_6t
Xbit_r80_c132 bl_132 br_132 wl_80 vdd gnd cell_6t
Xbit_r81_c132 bl_132 br_132 wl_81 vdd gnd cell_6t
Xbit_r82_c132 bl_132 br_132 wl_82 vdd gnd cell_6t
Xbit_r83_c132 bl_132 br_132 wl_83 vdd gnd cell_6t
Xbit_r84_c132 bl_132 br_132 wl_84 vdd gnd cell_6t
Xbit_r85_c132 bl_132 br_132 wl_85 vdd gnd cell_6t
Xbit_r86_c132 bl_132 br_132 wl_86 vdd gnd cell_6t
Xbit_r87_c132 bl_132 br_132 wl_87 vdd gnd cell_6t
Xbit_r88_c132 bl_132 br_132 wl_88 vdd gnd cell_6t
Xbit_r89_c132 bl_132 br_132 wl_89 vdd gnd cell_6t
Xbit_r90_c132 bl_132 br_132 wl_90 vdd gnd cell_6t
Xbit_r91_c132 bl_132 br_132 wl_91 vdd gnd cell_6t
Xbit_r92_c132 bl_132 br_132 wl_92 vdd gnd cell_6t
Xbit_r93_c132 bl_132 br_132 wl_93 vdd gnd cell_6t
Xbit_r94_c132 bl_132 br_132 wl_94 vdd gnd cell_6t
Xbit_r95_c132 bl_132 br_132 wl_95 vdd gnd cell_6t
Xbit_r96_c132 bl_132 br_132 wl_96 vdd gnd cell_6t
Xbit_r97_c132 bl_132 br_132 wl_97 vdd gnd cell_6t
Xbit_r98_c132 bl_132 br_132 wl_98 vdd gnd cell_6t
Xbit_r99_c132 bl_132 br_132 wl_99 vdd gnd cell_6t
Xbit_r100_c132 bl_132 br_132 wl_100 vdd gnd cell_6t
Xbit_r101_c132 bl_132 br_132 wl_101 vdd gnd cell_6t
Xbit_r102_c132 bl_132 br_132 wl_102 vdd gnd cell_6t
Xbit_r103_c132 bl_132 br_132 wl_103 vdd gnd cell_6t
Xbit_r104_c132 bl_132 br_132 wl_104 vdd gnd cell_6t
Xbit_r105_c132 bl_132 br_132 wl_105 vdd gnd cell_6t
Xbit_r106_c132 bl_132 br_132 wl_106 vdd gnd cell_6t
Xbit_r107_c132 bl_132 br_132 wl_107 vdd gnd cell_6t
Xbit_r108_c132 bl_132 br_132 wl_108 vdd gnd cell_6t
Xbit_r109_c132 bl_132 br_132 wl_109 vdd gnd cell_6t
Xbit_r110_c132 bl_132 br_132 wl_110 vdd gnd cell_6t
Xbit_r111_c132 bl_132 br_132 wl_111 vdd gnd cell_6t
Xbit_r112_c132 bl_132 br_132 wl_112 vdd gnd cell_6t
Xbit_r113_c132 bl_132 br_132 wl_113 vdd gnd cell_6t
Xbit_r114_c132 bl_132 br_132 wl_114 vdd gnd cell_6t
Xbit_r115_c132 bl_132 br_132 wl_115 vdd gnd cell_6t
Xbit_r116_c132 bl_132 br_132 wl_116 vdd gnd cell_6t
Xbit_r117_c132 bl_132 br_132 wl_117 vdd gnd cell_6t
Xbit_r118_c132 bl_132 br_132 wl_118 vdd gnd cell_6t
Xbit_r119_c132 bl_132 br_132 wl_119 vdd gnd cell_6t
Xbit_r120_c132 bl_132 br_132 wl_120 vdd gnd cell_6t
Xbit_r121_c132 bl_132 br_132 wl_121 vdd gnd cell_6t
Xbit_r122_c132 bl_132 br_132 wl_122 vdd gnd cell_6t
Xbit_r123_c132 bl_132 br_132 wl_123 vdd gnd cell_6t
Xbit_r124_c132 bl_132 br_132 wl_124 vdd gnd cell_6t
Xbit_r125_c132 bl_132 br_132 wl_125 vdd gnd cell_6t
Xbit_r126_c132 bl_132 br_132 wl_126 vdd gnd cell_6t
Xbit_r127_c132 bl_132 br_132 wl_127 vdd gnd cell_6t
Xbit_r128_c132 bl_132 br_132 wl_128 vdd gnd cell_6t
Xbit_r129_c132 bl_132 br_132 wl_129 vdd gnd cell_6t
Xbit_r130_c132 bl_132 br_132 wl_130 vdd gnd cell_6t
Xbit_r131_c132 bl_132 br_132 wl_131 vdd gnd cell_6t
Xbit_r132_c132 bl_132 br_132 wl_132 vdd gnd cell_6t
Xbit_r133_c132 bl_132 br_132 wl_133 vdd gnd cell_6t
Xbit_r134_c132 bl_132 br_132 wl_134 vdd gnd cell_6t
Xbit_r135_c132 bl_132 br_132 wl_135 vdd gnd cell_6t
Xbit_r136_c132 bl_132 br_132 wl_136 vdd gnd cell_6t
Xbit_r137_c132 bl_132 br_132 wl_137 vdd gnd cell_6t
Xbit_r138_c132 bl_132 br_132 wl_138 vdd gnd cell_6t
Xbit_r139_c132 bl_132 br_132 wl_139 vdd gnd cell_6t
Xbit_r140_c132 bl_132 br_132 wl_140 vdd gnd cell_6t
Xbit_r141_c132 bl_132 br_132 wl_141 vdd gnd cell_6t
Xbit_r142_c132 bl_132 br_132 wl_142 vdd gnd cell_6t
Xbit_r143_c132 bl_132 br_132 wl_143 vdd gnd cell_6t
Xbit_r144_c132 bl_132 br_132 wl_144 vdd gnd cell_6t
Xbit_r145_c132 bl_132 br_132 wl_145 vdd gnd cell_6t
Xbit_r146_c132 bl_132 br_132 wl_146 vdd gnd cell_6t
Xbit_r147_c132 bl_132 br_132 wl_147 vdd gnd cell_6t
Xbit_r148_c132 bl_132 br_132 wl_148 vdd gnd cell_6t
Xbit_r149_c132 bl_132 br_132 wl_149 vdd gnd cell_6t
Xbit_r150_c132 bl_132 br_132 wl_150 vdd gnd cell_6t
Xbit_r151_c132 bl_132 br_132 wl_151 vdd gnd cell_6t
Xbit_r152_c132 bl_132 br_132 wl_152 vdd gnd cell_6t
Xbit_r153_c132 bl_132 br_132 wl_153 vdd gnd cell_6t
Xbit_r154_c132 bl_132 br_132 wl_154 vdd gnd cell_6t
Xbit_r155_c132 bl_132 br_132 wl_155 vdd gnd cell_6t
Xbit_r156_c132 bl_132 br_132 wl_156 vdd gnd cell_6t
Xbit_r157_c132 bl_132 br_132 wl_157 vdd gnd cell_6t
Xbit_r158_c132 bl_132 br_132 wl_158 vdd gnd cell_6t
Xbit_r159_c132 bl_132 br_132 wl_159 vdd gnd cell_6t
Xbit_r160_c132 bl_132 br_132 wl_160 vdd gnd cell_6t
Xbit_r161_c132 bl_132 br_132 wl_161 vdd gnd cell_6t
Xbit_r162_c132 bl_132 br_132 wl_162 vdd gnd cell_6t
Xbit_r163_c132 bl_132 br_132 wl_163 vdd gnd cell_6t
Xbit_r164_c132 bl_132 br_132 wl_164 vdd gnd cell_6t
Xbit_r165_c132 bl_132 br_132 wl_165 vdd gnd cell_6t
Xbit_r166_c132 bl_132 br_132 wl_166 vdd gnd cell_6t
Xbit_r167_c132 bl_132 br_132 wl_167 vdd gnd cell_6t
Xbit_r168_c132 bl_132 br_132 wl_168 vdd gnd cell_6t
Xbit_r169_c132 bl_132 br_132 wl_169 vdd gnd cell_6t
Xbit_r170_c132 bl_132 br_132 wl_170 vdd gnd cell_6t
Xbit_r171_c132 bl_132 br_132 wl_171 vdd gnd cell_6t
Xbit_r172_c132 bl_132 br_132 wl_172 vdd gnd cell_6t
Xbit_r173_c132 bl_132 br_132 wl_173 vdd gnd cell_6t
Xbit_r174_c132 bl_132 br_132 wl_174 vdd gnd cell_6t
Xbit_r175_c132 bl_132 br_132 wl_175 vdd gnd cell_6t
Xbit_r176_c132 bl_132 br_132 wl_176 vdd gnd cell_6t
Xbit_r177_c132 bl_132 br_132 wl_177 vdd gnd cell_6t
Xbit_r178_c132 bl_132 br_132 wl_178 vdd gnd cell_6t
Xbit_r179_c132 bl_132 br_132 wl_179 vdd gnd cell_6t
Xbit_r180_c132 bl_132 br_132 wl_180 vdd gnd cell_6t
Xbit_r181_c132 bl_132 br_132 wl_181 vdd gnd cell_6t
Xbit_r182_c132 bl_132 br_132 wl_182 vdd gnd cell_6t
Xbit_r183_c132 bl_132 br_132 wl_183 vdd gnd cell_6t
Xbit_r184_c132 bl_132 br_132 wl_184 vdd gnd cell_6t
Xbit_r185_c132 bl_132 br_132 wl_185 vdd gnd cell_6t
Xbit_r186_c132 bl_132 br_132 wl_186 vdd gnd cell_6t
Xbit_r187_c132 bl_132 br_132 wl_187 vdd gnd cell_6t
Xbit_r188_c132 bl_132 br_132 wl_188 vdd gnd cell_6t
Xbit_r189_c132 bl_132 br_132 wl_189 vdd gnd cell_6t
Xbit_r190_c132 bl_132 br_132 wl_190 vdd gnd cell_6t
Xbit_r191_c132 bl_132 br_132 wl_191 vdd gnd cell_6t
Xbit_r192_c132 bl_132 br_132 wl_192 vdd gnd cell_6t
Xbit_r193_c132 bl_132 br_132 wl_193 vdd gnd cell_6t
Xbit_r194_c132 bl_132 br_132 wl_194 vdd gnd cell_6t
Xbit_r195_c132 bl_132 br_132 wl_195 vdd gnd cell_6t
Xbit_r196_c132 bl_132 br_132 wl_196 vdd gnd cell_6t
Xbit_r197_c132 bl_132 br_132 wl_197 vdd gnd cell_6t
Xbit_r198_c132 bl_132 br_132 wl_198 vdd gnd cell_6t
Xbit_r199_c132 bl_132 br_132 wl_199 vdd gnd cell_6t
Xbit_r200_c132 bl_132 br_132 wl_200 vdd gnd cell_6t
Xbit_r201_c132 bl_132 br_132 wl_201 vdd gnd cell_6t
Xbit_r202_c132 bl_132 br_132 wl_202 vdd gnd cell_6t
Xbit_r203_c132 bl_132 br_132 wl_203 vdd gnd cell_6t
Xbit_r204_c132 bl_132 br_132 wl_204 vdd gnd cell_6t
Xbit_r205_c132 bl_132 br_132 wl_205 vdd gnd cell_6t
Xbit_r206_c132 bl_132 br_132 wl_206 vdd gnd cell_6t
Xbit_r207_c132 bl_132 br_132 wl_207 vdd gnd cell_6t
Xbit_r208_c132 bl_132 br_132 wl_208 vdd gnd cell_6t
Xbit_r209_c132 bl_132 br_132 wl_209 vdd gnd cell_6t
Xbit_r210_c132 bl_132 br_132 wl_210 vdd gnd cell_6t
Xbit_r211_c132 bl_132 br_132 wl_211 vdd gnd cell_6t
Xbit_r212_c132 bl_132 br_132 wl_212 vdd gnd cell_6t
Xbit_r213_c132 bl_132 br_132 wl_213 vdd gnd cell_6t
Xbit_r214_c132 bl_132 br_132 wl_214 vdd gnd cell_6t
Xbit_r215_c132 bl_132 br_132 wl_215 vdd gnd cell_6t
Xbit_r216_c132 bl_132 br_132 wl_216 vdd gnd cell_6t
Xbit_r217_c132 bl_132 br_132 wl_217 vdd gnd cell_6t
Xbit_r218_c132 bl_132 br_132 wl_218 vdd gnd cell_6t
Xbit_r219_c132 bl_132 br_132 wl_219 vdd gnd cell_6t
Xbit_r220_c132 bl_132 br_132 wl_220 vdd gnd cell_6t
Xbit_r221_c132 bl_132 br_132 wl_221 vdd gnd cell_6t
Xbit_r222_c132 bl_132 br_132 wl_222 vdd gnd cell_6t
Xbit_r223_c132 bl_132 br_132 wl_223 vdd gnd cell_6t
Xbit_r224_c132 bl_132 br_132 wl_224 vdd gnd cell_6t
Xbit_r225_c132 bl_132 br_132 wl_225 vdd gnd cell_6t
Xbit_r226_c132 bl_132 br_132 wl_226 vdd gnd cell_6t
Xbit_r227_c132 bl_132 br_132 wl_227 vdd gnd cell_6t
Xbit_r228_c132 bl_132 br_132 wl_228 vdd gnd cell_6t
Xbit_r229_c132 bl_132 br_132 wl_229 vdd gnd cell_6t
Xbit_r230_c132 bl_132 br_132 wl_230 vdd gnd cell_6t
Xbit_r231_c132 bl_132 br_132 wl_231 vdd gnd cell_6t
Xbit_r232_c132 bl_132 br_132 wl_232 vdd gnd cell_6t
Xbit_r233_c132 bl_132 br_132 wl_233 vdd gnd cell_6t
Xbit_r234_c132 bl_132 br_132 wl_234 vdd gnd cell_6t
Xbit_r235_c132 bl_132 br_132 wl_235 vdd gnd cell_6t
Xbit_r236_c132 bl_132 br_132 wl_236 vdd gnd cell_6t
Xbit_r237_c132 bl_132 br_132 wl_237 vdd gnd cell_6t
Xbit_r238_c132 bl_132 br_132 wl_238 vdd gnd cell_6t
Xbit_r239_c132 bl_132 br_132 wl_239 vdd gnd cell_6t
Xbit_r240_c132 bl_132 br_132 wl_240 vdd gnd cell_6t
Xbit_r241_c132 bl_132 br_132 wl_241 vdd gnd cell_6t
Xbit_r242_c132 bl_132 br_132 wl_242 vdd gnd cell_6t
Xbit_r243_c132 bl_132 br_132 wl_243 vdd gnd cell_6t
Xbit_r244_c132 bl_132 br_132 wl_244 vdd gnd cell_6t
Xbit_r245_c132 bl_132 br_132 wl_245 vdd gnd cell_6t
Xbit_r246_c132 bl_132 br_132 wl_246 vdd gnd cell_6t
Xbit_r247_c132 bl_132 br_132 wl_247 vdd gnd cell_6t
Xbit_r248_c132 bl_132 br_132 wl_248 vdd gnd cell_6t
Xbit_r249_c132 bl_132 br_132 wl_249 vdd gnd cell_6t
Xbit_r250_c132 bl_132 br_132 wl_250 vdd gnd cell_6t
Xbit_r251_c132 bl_132 br_132 wl_251 vdd gnd cell_6t
Xbit_r252_c132 bl_132 br_132 wl_252 vdd gnd cell_6t
Xbit_r253_c132 bl_132 br_132 wl_253 vdd gnd cell_6t
Xbit_r254_c132 bl_132 br_132 wl_254 vdd gnd cell_6t
Xbit_r255_c132 bl_132 br_132 wl_255 vdd gnd cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd cell_6t
Xbit_r1_c133 bl_133 br_133 wl_1 vdd gnd cell_6t
Xbit_r2_c133 bl_133 br_133 wl_2 vdd gnd cell_6t
Xbit_r3_c133 bl_133 br_133 wl_3 vdd gnd cell_6t
Xbit_r4_c133 bl_133 br_133 wl_4 vdd gnd cell_6t
Xbit_r5_c133 bl_133 br_133 wl_5 vdd gnd cell_6t
Xbit_r6_c133 bl_133 br_133 wl_6 vdd gnd cell_6t
Xbit_r7_c133 bl_133 br_133 wl_7 vdd gnd cell_6t
Xbit_r8_c133 bl_133 br_133 wl_8 vdd gnd cell_6t
Xbit_r9_c133 bl_133 br_133 wl_9 vdd gnd cell_6t
Xbit_r10_c133 bl_133 br_133 wl_10 vdd gnd cell_6t
Xbit_r11_c133 bl_133 br_133 wl_11 vdd gnd cell_6t
Xbit_r12_c133 bl_133 br_133 wl_12 vdd gnd cell_6t
Xbit_r13_c133 bl_133 br_133 wl_13 vdd gnd cell_6t
Xbit_r14_c133 bl_133 br_133 wl_14 vdd gnd cell_6t
Xbit_r15_c133 bl_133 br_133 wl_15 vdd gnd cell_6t
Xbit_r16_c133 bl_133 br_133 wl_16 vdd gnd cell_6t
Xbit_r17_c133 bl_133 br_133 wl_17 vdd gnd cell_6t
Xbit_r18_c133 bl_133 br_133 wl_18 vdd gnd cell_6t
Xbit_r19_c133 bl_133 br_133 wl_19 vdd gnd cell_6t
Xbit_r20_c133 bl_133 br_133 wl_20 vdd gnd cell_6t
Xbit_r21_c133 bl_133 br_133 wl_21 vdd gnd cell_6t
Xbit_r22_c133 bl_133 br_133 wl_22 vdd gnd cell_6t
Xbit_r23_c133 bl_133 br_133 wl_23 vdd gnd cell_6t
Xbit_r24_c133 bl_133 br_133 wl_24 vdd gnd cell_6t
Xbit_r25_c133 bl_133 br_133 wl_25 vdd gnd cell_6t
Xbit_r26_c133 bl_133 br_133 wl_26 vdd gnd cell_6t
Xbit_r27_c133 bl_133 br_133 wl_27 vdd gnd cell_6t
Xbit_r28_c133 bl_133 br_133 wl_28 vdd gnd cell_6t
Xbit_r29_c133 bl_133 br_133 wl_29 vdd gnd cell_6t
Xbit_r30_c133 bl_133 br_133 wl_30 vdd gnd cell_6t
Xbit_r31_c133 bl_133 br_133 wl_31 vdd gnd cell_6t
Xbit_r32_c133 bl_133 br_133 wl_32 vdd gnd cell_6t
Xbit_r33_c133 bl_133 br_133 wl_33 vdd gnd cell_6t
Xbit_r34_c133 bl_133 br_133 wl_34 vdd gnd cell_6t
Xbit_r35_c133 bl_133 br_133 wl_35 vdd gnd cell_6t
Xbit_r36_c133 bl_133 br_133 wl_36 vdd gnd cell_6t
Xbit_r37_c133 bl_133 br_133 wl_37 vdd gnd cell_6t
Xbit_r38_c133 bl_133 br_133 wl_38 vdd gnd cell_6t
Xbit_r39_c133 bl_133 br_133 wl_39 vdd gnd cell_6t
Xbit_r40_c133 bl_133 br_133 wl_40 vdd gnd cell_6t
Xbit_r41_c133 bl_133 br_133 wl_41 vdd gnd cell_6t
Xbit_r42_c133 bl_133 br_133 wl_42 vdd gnd cell_6t
Xbit_r43_c133 bl_133 br_133 wl_43 vdd gnd cell_6t
Xbit_r44_c133 bl_133 br_133 wl_44 vdd gnd cell_6t
Xbit_r45_c133 bl_133 br_133 wl_45 vdd gnd cell_6t
Xbit_r46_c133 bl_133 br_133 wl_46 vdd gnd cell_6t
Xbit_r47_c133 bl_133 br_133 wl_47 vdd gnd cell_6t
Xbit_r48_c133 bl_133 br_133 wl_48 vdd gnd cell_6t
Xbit_r49_c133 bl_133 br_133 wl_49 vdd gnd cell_6t
Xbit_r50_c133 bl_133 br_133 wl_50 vdd gnd cell_6t
Xbit_r51_c133 bl_133 br_133 wl_51 vdd gnd cell_6t
Xbit_r52_c133 bl_133 br_133 wl_52 vdd gnd cell_6t
Xbit_r53_c133 bl_133 br_133 wl_53 vdd gnd cell_6t
Xbit_r54_c133 bl_133 br_133 wl_54 vdd gnd cell_6t
Xbit_r55_c133 bl_133 br_133 wl_55 vdd gnd cell_6t
Xbit_r56_c133 bl_133 br_133 wl_56 vdd gnd cell_6t
Xbit_r57_c133 bl_133 br_133 wl_57 vdd gnd cell_6t
Xbit_r58_c133 bl_133 br_133 wl_58 vdd gnd cell_6t
Xbit_r59_c133 bl_133 br_133 wl_59 vdd gnd cell_6t
Xbit_r60_c133 bl_133 br_133 wl_60 vdd gnd cell_6t
Xbit_r61_c133 bl_133 br_133 wl_61 vdd gnd cell_6t
Xbit_r62_c133 bl_133 br_133 wl_62 vdd gnd cell_6t
Xbit_r63_c133 bl_133 br_133 wl_63 vdd gnd cell_6t
Xbit_r64_c133 bl_133 br_133 wl_64 vdd gnd cell_6t
Xbit_r65_c133 bl_133 br_133 wl_65 vdd gnd cell_6t
Xbit_r66_c133 bl_133 br_133 wl_66 vdd gnd cell_6t
Xbit_r67_c133 bl_133 br_133 wl_67 vdd gnd cell_6t
Xbit_r68_c133 bl_133 br_133 wl_68 vdd gnd cell_6t
Xbit_r69_c133 bl_133 br_133 wl_69 vdd gnd cell_6t
Xbit_r70_c133 bl_133 br_133 wl_70 vdd gnd cell_6t
Xbit_r71_c133 bl_133 br_133 wl_71 vdd gnd cell_6t
Xbit_r72_c133 bl_133 br_133 wl_72 vdd gnd cell_6t
Xbit_r73_c133 bl_133 br_133 wl_73 vdd gnd cell_6t
Xbit_r74_c133 bl_133 br_133 wl_74 vdd gnd cell_6t
Xbit_r75_c133 bl_133 br_133 wl_75 vdd gnd cell_6t
Xbit_r76_c133 bl_133 br_133 wl_76 vdd gnd cell_6t
Xbit_r77_c133 bl_133 br_133 wl_77 vdd gnd cell_6t
Xbit_r78_c133 bl_133 br_133 wl_78 vdd gnd cell_6t
Xbit_r79_c133 bl_133 br_133 wl_79 vdd gnd cell_6t
Xbit_r80_c133 bl_133 br_133 wl_80 vdd gnd cell_6t
Xbit_r81_c133 bl_133 br_133 wl_81 vdd gnd cell_6t
Xbit_r82_c133 bl_133 br_133 wl_82 vdd gnd cell_6t
Xbit_r83_c133 bl_133 br_133 wl_83 vdd gnd cell_6t
Xbit_r84_c133 bl_133 br_133 wl_84 vdd gnd cell_6t
Xbit_r85_c133 bl_133 br_133 wl_85 vdd gnd cell_6t
Xbit_r86_c133 bl_133 br_133 wl_86 vdd gnd cell_6t
Xbit_r87_c133 bl_133 br_133 wl_87 vdd gnd cell_6t
Xbit_r88_c133 bl_133 br_133 wl_88 vdd gnd cell_6t
Xbit_r89_c133 bl_133 br_133 wl_89 vdd gnd cell_6t
Xbit_r90_c133 bl_133 br_133 wl_90 vdd gnd cell_6t
Xbit_r91_c133 bl_133 br_133 wl_91 vdd gnd cell_6t
Xbit_r92_c133 bl_133 br_133 wl_92 vdd gnd cell_6t
Xbit_r93_c133 bl_133 br_133 wl_93 vdd gnd cell_6t
Xbit_r94_c133 bl_133 br_133 wl_94 vdd gnd cell_6t
Xbit_r95_c133 bl_133 br_133 wl_95 vdd gnd cell_6t
Xbit_r96_c133 bl_133 br_133 wl_96 vdd gnd cell_6t
Xbit_r97_c133 bl_133 br_133 wl_97 vdd gnd cell_6t
Xbit_r98_c133 bl_133 br_133 wl_98 vdd gnd cell_6t
Xbit_r99_c133 bl_133 br_133 wl_99 vdd gnd cell_6t
Xbit_r100_c133 bl_133 br_133 wl_100 vdd gnd cell_6t
Xbit_r101_c133 bl_133 br_133 wl_101 vdd gnd cell_6t
Xbit_r102_c133 bl_133 br_133 wl_102 vdd gnd cell_6t
Xbit_r103_c133 bl_133 br_133 wl_103 vdd gnd cell_6t
Xbit_r104_c133 bl_133 br_133 wl_104 vdd gnd cell_6t
Xbit_r105_c133 bl_133 br_133 wl_105 vdd gnd cell_6t
Xbit_r106_c133 bl_133 br_133 wl_106 vdd gnd cell_6t
Xbit_r107_c133 bl_133 br_133 wl_107 vdd gnd cell_6t
Xbit_r108_c133 bl_133 br_133 wl_108 vdd gnd cell_6t
Xbit_r109_c133 bl_133 br_133 wl_109 vdd gnd cell_6t
Xbit_r110_c133 bl_133 br_133 wl_110 vdd gnd cell_6t
Xbit_r111_c133 bl_133 br_133 wl_111 vdd gnd cell_6t
Xbit_r112_c133 bl_133 br_133 wl_112 vdd gnd cell_6t
Xbit_r113_c133 bl_133 br_133 wl_113 vdd gnd cell_6t
Xbit_r114_c133 bl_133 br_133 wl_114 vdd gnd cell_6t
Xbit_r115_c133 bl_133 br_133 wl_115 vdd gnd cell_6t
Xbit_r116_c133 bl_133 br_133 wl_116 vdd gnd cell_6t
Xbit_r117_c133 bl_133 br_133 wl_117 vdd gnd cell_6t
Xbit_r118_c133 bl_133 br_133 wl_118 vdd gnd cell_6t
Xbit_r119_c133 bl_133 br_133 wl_119 vdd gnd cell_6t
Xbit_r120_c133 bl_133 br_133 wl_120 vdd gnd cell_6t
Xbit_r121_c133 bl_133 br_133 wl_121 vdd gnd cell_6t
Xbit_r122_c133 bl_133 br_133 wl_122 vdd gnd cell_6t
Xbit_r123_c133 bl_133 br_133 wl_123 vdd gnd cell_6t
Xbit_r124_c133 bl_133 br_133 wl_124 vdd gnd cell_6t
Xbit_r125_c133 bl_133 br_133 wl_125 vdd gnd cell_6t
Xbit_r126_c133 bl_133 br_133 wl_126 vdd gnd cell_6t
Xbit_r127_c133 bl_133 br_133 wl_127 vdd gnd cell_6t
Xbit_r128_c133 bl_133 br_133 wl_128 vdd gnd cell_6t
Xbit_r129_c133 bl_133 br_133 wl_129 vdd gnd cell_6t
Xbit_r130_c133 bl_133 br_133 wl_130 vdd gnd cell_6t
Xbit_r131_c133 bl_133 br_133 wl_131 vdd gnd cell_6t
Xbit_r132_c133 bl_133 br_133 wl_132 vdd gnd cell_6t
Xbit_r133_c133 bl_133 br_133 wl_133 vdd gnd cell_6t
Xbit_r134_c133 bl_133 br_133 wl_134 vdd gnd cell_6t
Xbit_r135_c133 bl_133 br_133 wl_135 vdd gnd cell_6t
Xbit_r136_c133 bl_133 br_133 wl_136 vdd gnd cell_6t
Xbit_r137_c133 bl_133 br_133 wl_137 vdd gnd cell_6t
Xbit_r138_c133 bl_133 br_133 wl_138 vdd gnd cell_6t
Xbit_r139_c133 bl_133 br_133 wl_139 vdd gnd cell_6t
Xbit_r140_c133 bl_133 br_133 wl_140 vdd gnd cell_6t
Xbit_r141_c133 bl_133 br_133 wl_141 vdd gnd cell_6t
Xbit_r142_c133 bl_133 br_133 wl_142 vdd gnd cell_6t
Xbit_r143_c133 bl_133 br_133 wl_143 vdd gnd cell_6t
Xbit_r144_c133 bl_133 br_133 wl_144 vdd gnd cell_6t
Xbit_r145_c133 bl_133 br_133 wl_145 vdd gnd cell_6t
Xbit_r146_c133 bl_133 br_133 wl_146 vdd gnd cell_6t
Xbit_r147_c133 bl_133 br_133 wl_147 vdd gnd cell_6t
Xbit_r148_c133 bl_133 br_133 wl_148 vdd gnd cell_6t
Xbit_r149_c133 bl_133 br_133 wl_149 vdd gnd cell_6t
Xbit_r150_c133 bl_133 br_133 wl_150 vdd gnd cell_6t
Xbit_r151_c133 bl_133 br_133 wl_151 vdd gnd cell_6t
Xbit_r152_c133 bl_133 br_133 wl_152 vdd gnd cell_6t
Xbit_r153_c133 bl_133 br_133 wl_153 vdd gnd cell_6t
Xbit_r154_c133 bl_133 br_133 wl_154 vdd gnd cell_6t
Xbit_r155_c133 bl_133 br_133 wl_155 vdd gnd cell_6t
Xbit_r156_c133 bl_133 br_133 wl_156 vdd gnd cell_6t
Xbit_r157_c133 bl_133 br_133 wl_157 vdd gnd cell_6t
Xbit_r158_c133 bl_133 br_133 wl_158 vdd gnd cell_6t
Xbit_r159_c133 bl_133 br_133 wl_159 vdd gnd cell_6t
Xbit_r160_c133 bl_133 br_133 wl_160 vdd gnd cell_6t
Xbit_r161_c133 bl_133 br_133 wl_161 vdd gnd cell_6t
Xbit_r162_c133 bl_133 br_133 wl_162 vdd gnd cell_6t
Xbit_r163_c133 bl_133 br_133 wl_163 vdd gnd cell_6t
Xbit_r164_c133 bl_133 br_133 wl_164 vdd gnd cell_6t
Xbit_r165_c133 bl_133 br_133 wl_165 vdd gnd cell_6t
Xbit_r166_c133 bl_133 br_133 wl_166 vdd gnd cell_6t
Xbit_r167_c133 bl_133 br_133 wl_167 vdd gnd cell_6t
Xbit_r168_c133 bl_133 br_133 wl_168 vdd gnd cell_6t
Xbit_r169_c133 bl_133 br_133 wl_169 vdd gnd cell_6t
Xbit_r170_c133 bl_133 br_133 wl_170 vdd gnd cell_6t
Xbit_r171_c133 bl_133 br_133 wl_171 vdd gnd cell_6t
Xbit_r172_c133 bl_133 br_133 wl_172 vdd gnd cell_6t
Xbit_r173_c133 bl_133 br_133 wl_173 vdd gnd cell_6t
Xbit_r174_c133 bl_133 br_133 wl_174 vdd gnd cell_6t
Xbit_r175_c133 bl_133 br_133 wl_175 vdd gnd cell_6t
Xbit_r176_c133 bl_133 br_133 wl_176 vdd gnd cell_6t
Xbit_r177_c133 bl_133 br_133 wl_177 vdd gnd cell_6t
Xbit_r178_c133 bl_133 br_133 wl_178 vdd gnd cell_6t
Xbit_r179_c133 bl_133 br_133 wl_179 vdd gnd cell_6t
Xbit_r180_c133 bl_133 br_133 wl_180 vdd gnd cell_6t
Xbit_r181_c133 bl_133 br_133 wl_181 vdd gnd cell_6t
Xbit_r182_c133 bl_133 br_133 wl_182 vdd gnd cell_6t
Xbit_r183_c133 bl_133 br_133 wl_183 vdd gnd cell_6t
Xbit_r184_c133 bl_133 br_133 wl_184 vdd gnd cell_6t
Xbit_r185_c133 bl_133 br_133 wl_185 vdd gnd cell_6t
Xbit_r186_c133 bl_133 br_133 wl_186 vdd gnd cell_6t
Xbit_r187_c133 bl_133 br_133 wl_187 vdd gnd cell_6t
Xbit_r188_c133 bl_133 br_133 wl_188 vdd gnd cell_6t
Xbit_r189_c133 bl_133 br_133 wl_189 vdd gnd cell_6t
Xbit_r190_c133 bl_133 br_133 wl_190 vdd gnd cell_6t
Xbit_r191_c133 bl_133 br_133 wl_191 vdd gnd cell_6t
Xbit_r192_c133 bl_133 br_133 wl_192 vdd gnd cell_6t
Xbit_r193_c133 bl_133 br_133 wl_193 vdd gnd cell_6t
Xbit_r194_c133 bl_133 br_133 wl_194 vdd gnd cell_6t
Xbit_r195_c133 bl_133 br_133 wl_195 vdd gnd cell_6t
Xbit_r196_c133 bl_133 br_133 wl_196 vdd gnd cell_6t
Xbit_r197_c133 bl_133 br_133 wl_197 vdd gnd cell_6t
Xbit_r198_c133 bl_133 br_133 wl_198 vdd gnd cell_6t
Xbit_r199_c133 bl_133 br_133 wl_199 vdd gnd cell_6t
Xbit_r200_c133 bl_133 br_133 wl_200 vdd gnd cell_6t
Xbit_r201_c133 bl_133 br_133 wl_201 vdd gnd cell_6t
Xbit_r202_c133 bl_133 br_133 wl_202 vdd gnd cell_6t
Xbit_r203_c133 bl_133 br_133 wl_203 vdd gnd cell_6t
Xbit_r204_c133 bl_133 br_133 wl_204 vdd gnd cell_6t
Xbit_r205_c133 bl_133 br_133 wl_205 vdd gnd cell_6t
Xbit_r206_c133 bl_133 br_133 wl_206 vdd gnd cell_6t
Xbit_r207_c133 bl_133 br_133 wl_207 vdd gnd cell_6t
Xbit_r208_c133 bl_133 br_133 wl_208 vdd gnd cell_6t
Xbit_r209_c133 bl_133 br_133 wl_209 vdd gnd cell_6t
Xbit_r210_c133 bl_133 br_133 wl_210 vdd gnd cell_6t
Xbit_r211_c133 bl_133 br_133 wl_211 vdd gnd cell_6t
Xbit_r212_c133 bl_133 br_133 wl_212 vdd gnd cell_6t
Xbit_r213_c133 bl_133 br_133 wl_213 vdd gnd cell_6t
Xbit_r214_c133 bl_133 br_133 wl_214 vdd gnd cell_6t
Xbit_r215_c133 bl_133 br_133 wl_215 vdd gnd cell_6t
Xbit_r216_c133 bl_133 br_133 wl_216 vdd gnd cell_6t
Xbit_r217_c133 bl_133 br_133 wl_217 vdd gnd cell_6t
Xbit_r218_c133 bl_133 br_133 wl_218 vdd gnd cell_6t
Xbit_r219_c133 bl_133 br_133 wl_219 vdd gnd cell_6t
Xbit_r220_c133 bl_133 br_133 wl_220 vdd gnd cell_6t
Xbit_r221_c133 bl_133 br_133 wl_221 vdd gnd cell_6t
Xbit_r222_c133 bl_133 br_133 wl_222 vdd gnd cell_6t
Xbit_r223_c133 bl_133 br_133 wl_223 vdd gnd cell_6t
Xbit_r224_c133 bl_133 br_133 wl_224 vdd gnd cell_6t
Xbit_r225_c133 bl_133 br_133 wl_225 vdd gnd cell_6t
Xbit_r226_c133 bl_133 br_133 wl_226 vdd gnd cell_6t
Xbit_r227_c133 bl_133 br_133 wl_227 vdd gnd cell_6t
Xbit_r228_c133 bl_133 br_133 wl_228 vdd gnd cell_6t
Xbit_r229_c133 bl_133 br_133 wl_229 vdd gnd cell_6t
Xbit_r230_c133 bl_133 br_133 wl_230 vdd gnd cell_6t
Xbit_r231_c133 bl_133 br_133 wl_231 vdd gnd cell_6t
Xbit_r232_c133 bl_133 br_133 wl_232 vdd gnd cell_6t
Xbit_r233_c133 bl_133 br_133 wl_233 vdd gnd cell_6t
Xbit_r234_c133 bl_133 br_133 wl_234 vdd gnd cell_6t
Xbit_r235_c133 bl_133 br_133 wl_235 vdd gnd cell_6t
Xbit_r236_c133 bl_133 br_133 wl_236 vdd gnd cell_6t
Xbit_r237_c133 bl_133 br_133 wl_237 vdd gnd cell_6t
Xbit_r238_c133 bl_133 br_133 wl_238 vdd gnd cell_6t
Xbit_r239_c133 bl_133 br_133 wl_239 vdd gnd cell_6t
Xbit_r240_c133 bl_133 br_133 wl_240 vdd gnd cell_6t
Xbit_r241_c133 bl_133 br_133 wl_241 vdd gnd cell_6t
Xbit_r242_c133 bl_133 br_133 wl_242 vdd gnd cell_6t
Xbit_r243_c133 bl_133 br_133 wl_243 vdd gnd cell_6t
Xbit_r244_c133 bl_133 br_133 wl_244 vdd gnd cell_6t
Xbit_r245_c133 bl_133 br_133 wl_245 vdd gnd cell_6t
Xbit_r246_c133 bl_133 br_133 wl_246 vdd gnd cell_6t
Xbit_r247_c133 bl_133 br_133 wl_247 vdd gnd cell_6t
Xbit_r248_c133 bl_133 br_133 wl_248 vdd gnd cell_6t
Xbit_r249_c133 bl_133 br_133 wl_249 vdd gnd cell_6t
Xbit_r250_c133 bl_133 br_133 wl_250 vdd gnd cell_6t
Xbit_r251_c133 bl_133 br_133 wl_251 vdd gnd cell_6t
Xbit_r252_c133 bl_133 br_133 wl_252 vdd gnd cell_6t
Xbit_r253_c133 bl_133 br_133 wl_253 vdd gnd cell_6t
Xbit_r254_c133 bl_133 br_133 wl_254 vdd gnd cell_6t
Xbit_r255_c133 bl_133 br_133 wl_255 vdd gnd cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd cell_6t
Xbit_r1_c134 bl_134 br_134 wl_1 vdd gnd cell_6t
Xbit_r2_c134 bl_134 br_134 wl_2 vdd gnd cell_6t
Xbit_r3_c134 bl_134 br_134 wl_3 vdd gnd cell_6t
Xbit_r4_c134 bl_134 br_134 wl_4 vdd gnd cell_6t
Xbit_r5_c134 bl_134 br_134 wl_5 vdd gnd cell_6t
Xbit_r6_c134 bl_134 br_134 wl_6 vdd gnd cell_6t
Xbit_r7_c134 bl_134 br_134 wl_7 vdd gnd cell_6t
Xbit_r8_c134 bl_134 br_134 wl_8 vdd gnd cell_6t
Xbit_r9_c134 bl_134 br_134 wl_9 vdd gnd cell_6t
Xbit_r10_c134 bl_134 br_134 wl_10 vdd gnd cell_6t
Xbit_r11_c134 bl_134 br_134 wl_11 vdd gnd cell_6t
Xbit_r12_c134 bl_134 br_134 wl_12 vdd gnd cell_6t
Xbit_r13_c134 bl_134 br_134 wl_13 vdd gnd cell_6t
Xbit_r14_c134 bl_134 br_134 wl_14 vdd gnd cell_6t
Xbit_r15_c134 bl_134 br_134 wl_15 vdd gnd cell_6t
Xbit_r16_c134 bl_134 br_134 wl_16 vdd gnd cell_6t
Xbit_r17_c134 bl_134 br_134 wl_17 vdd gnd cell_6t
Xbit_r18_c134 bl_134 br_134 wl_18 vdd gnd cell_6t
Xbit_r19_c134 bl_134 br_134 wl_19 vdd gnd cell_6t
Xbit_r20_c134 bl_134 br_134 wl_20 vdd gnd cell_6t
Xbit_r21_c134 bl_134 br_134 wl_21 vdd gnd cell_6t
Xbit_r22_c134 bl_134 br_134 wl_22 vdd gnd cell_6t
Xbit_r23_c134 bl_134 br_134 wl_23 vdd gnd cell_6t
Xbit_r24_c134 bl_134 br_134 wl_24 vdd gnd cell_6t
Xbit_r25_c134 bl_134 br_134 wl_25 vdd gnd cell_6t
Xbit_r26_c134 bl_134 br_134 wl_26 vdd gnd cell_6t
Xbit_r27_c134 bl_134 br_134 wl_27 vdd gnd cell_6t
Xbit_r28_c134 bl_134 br_134 wl_28 vdd gnd cell_6t
Xbit_r29_c134 bl_134 br_134 wl_29 vdd gnd cell_6t
Xbit_r30_c134 bl_134 br_134 wl_30 vdd gnd cell_6t
Xbit_r31_c134 bl_134 br_134 wl_31 vdd gnd cell_6t
Xbit_r32_c134 bl_134 br_134 wl_32 vdd gnd cell_6t
Xbit_r33_c134 bl_134 br_134 wl_33 vdd gnd cell_6t
Xbit_r34_c134 bl_134 br_134 wl_34 vdd gnd cell_6t
Xbit_r35_c134 bl_134 br_134 wl_35 vdd gnd cell_6t
Xbit_r36_c134 bl_134 br_134 wl_36 vdd gnd cell_6t
Xbit_r37_c134 bl_134 br_134 wl_37 vdd gnd cell_6t
Xbit_r38_c134 bl_134 br_134 wl_38 vdd gnd cell_6t
Xbit_r39_c134 bl_134 br_134 wl_39 vdd gnd cell_6t
Xbit_r40_c134 bl_134 br_134 wl_40 vdd gnd cell_6t
Xbit_r41_c134 bl_134 br_134 wl_41 vdd gnd cell_6t
Xbit_r42_c134 bl_134 br_134 wl_42 vdd gnd cell_6t
Xbit_r43_c134 bl_134 br_134 wl_43 vdd gnd cell_6t
Xbit_r44_c134 bl_134 br_134 wl_44 vdd gnd cell_6t
Xbit_r45_c134 bl_134 br_134 wl_45 vdd gnd cell_6t
Xbit_r46_c134 bl_134 br_134 wl_46 vdd gnd cell_6t
Xbit_r47_c134 bl_134 br_134 wl_47 vdd gnd cell_6t
Xbit_r48_c134 bl_134 br_134 wl_48 vdd gnd cell_6t
Xbit_r49_c134 bl_134 br_134 wl_49 vdd gnd cell_6t
Xbit_r50_c134 bl_134 br_134 wl_50 vdd gnd cell_6t
Xbit_r51_c134 bl_134 br_134 wl_51 vdd gnd cell_6t
Xbit_r52_c134 bl_134 br_134 wl_52 vdd gnd cell_6t
Xbit_r53_c134 bl_134 br_134 wl_53 vdd gnd cell_6t
Xbit_r54_c134 bl_134 br_134 wl_54 vdd gnd cell_6t
Xbit_r55_c134 bl_134 br_134 wl_55 vdd gnd cell_6t
Xbit_r56_c134 bl_134 br_134 wl_56 vdd gnd cell_6t
Xbit_r57_c134 bl_134 br_134 wl_57 vdd gnd cell_6t
Xbit_r58_c134 bl_134 br_134 wl_58 vdd gnd cell_6t
Xbit_r59_c134 bl_134 br_134 wl_59 vdd gnd cell_6t
Xbit_r60_c134 bl_134 br_134 wl_60 vdd gnd cell_6t
Xbit_r61_c134 bl_134 br_134 wl_61 vdd gnd cell_6t
Xbit_r62_c134 bl_134 br_134 wl_62 vdd gnd cell_6t
Xbit_r63_c134 bl_134 br_134 wl_63 vdd gnd cell_6t
Xbit_r64_c134 bl_134 br_134 wl_64 vdd gnd cell_6t
Xbit_r65_c134 bl_134 br_134 wl_65 vdd gnd cell_6t
Xbit_r66_c134 bl_134 br_134 wl_66 vdd gnd cell_6t
Xbit_r67_c134 bl_134 br_134 wl_67 vdd gnd cell_6t
Xbit_r68_c134 bl_134 br_134 wl_68 vdd gnd cell_6t
Xbit_r69_c134 bl_134 br_134 wl_69 vdd gnd cell_6t
Xbit_r70_c134 bl_134 br_134 wl_70 vdd gnd cell_6t
Xbit_r71_c134 bl_134 br_134 wl_71 vdd gnd cell_6t
Xbit_r72_c134 bl_134 br_134 wl_72 vdd gnd cell_6t
Xbit_r73_c134 bl_134 br_134 wl_73 vdd gnd cell_6t
Xbit_r74_c134 bl_134 br_134 wl_74 vdd gnd cell_6t
Xbit_r75_c134 bl_134 br_134 wl_75 vdd gnd cell_6t
Xbit_r76_c134 bl_134 br_134 wl_76 vdd gnd cell_6t
Xbit_r77_c134 bl_134 br_134 wl_77 vdd gnd cell_6t
Xbit_r78_c134 bl_134 br_134 wl_78 vdd gnd cell_6t
Xbit_r79_c134 bl_134 br_134 wl_79 vdd gnd cell_6t
Xbit_r80_c134 bl_134 br_134 wl_80 vdd gnd cell_6t
Xbit_r81_c134 bl_134 br_134 wl_81 vdd gnd cell_6t
Xbit_r82_c134 bl_134 br_134 wl_82 vdd gnd cell_6t
Xbit_r83_c134 bl_134 br_134 wl_83 vdd gnd cell_6t
Xbit_r84_c134 bl_134 br_134 wl_84 vdd gnd cell_6t
Xbit_r85_c134 bl_134 br_134 wl_85 vdd gnd cell_6t
Xbit_r86_c134 bl_134 br_134 wl_86 vdd gnd cell_6t
Xbit_r87_c134 bl_134 br_134 wl_87 vdd gnd cell_6t
Xbit_r88_c134 bl_134 br_134 wl_88 vdd gnd cell_6t
Xbit_r89_c134 bl_134 br_134 wl_89 vdd gnd cell_6t
Xbit_r90_c134 bl_134 br_134 wl_90 vdd gnd cell_6t
Xbit_r91_c134 bl_134 br_134 wl_91 vdd gnd cell_6t
Xbit_r92_c134 bl_134 br_134 wl_92 vdd gnd cell_6t
Xbit_r93_c134 bl_134 br_134 wl_93 vdd gnd cell_6t
Xbit_r94_c134 bl_134 br_134 wl_94 vdd gnd cell_6t
Xbit_r95_c134 bl_134 br_134 wl_95 vdd gnd cell_6t
Xbit_r96_c134 bl_134 br_134 wl_96 vdd gnd cell_6t
Xbit_r97_c134 bl_134 br_134 wl_97 vdd gnd cell_6t
Xbit_r98_c134 bl_134 br_134 wl_98 vdd gnd cell_6t
Xbit_r99_c134 bl_134 br_134 wl_99 vdd gnd cell_6t
Xbit_r100_c134 bl_134 br_134 wl_100 vdd gnd cell_6t
Xbit_r101_c134 bl_134 br_134 wl_101 vdd gnd cell_6t
Xbit_r102_c134 bl_134 br_134 wl_102 vdd gnd cell_6t
Xbit_r103_c134 bl_134 br_134 wl_103 vdd gnd cell_6t
Xbit_r104_c134 bl_134 br_134 wl_104 vdd gnd cell_6t
Xbit_r105_c134 bl_134 br_134 wl_105 vdd gnd cell_6t
Xbit_r106_c134 bl_134 br_134 wl_106 vdd gnd cell_6t
Xbit_r107_c134 bl_134 br_134 wl_107 vdd gnd cell_6t
Xbit_r108_c134 bl_134 br_134 wl_108 vdd gnd cell_6t
Xbit_r109_c134 bl_134 br_134 wl_109 vdd gnd cell_6t
Xbit_r110_c134 bl_134 br_134 wl_110 vdd gnd cell_6t
Xbit_r111_c134 bl_134 br_134 wl_111 vdd gnd cell_6t
Xbit_r112_c134 bl_134 br_134 wl_112 vdd gnd cell_6t
Xbit_r113_c134 bl_134 br_134 wl_113 vdd gnd cell_6t
Xbit_r114_c134 bl_134 br_134 wl_114 vdd gnd cell_6t
Xbit_r115_c134 bl_134 br_134 wl_115 vdd gnd cell_6t
Xbit_r116_c134 bl_134 br_134 wl_116 vdd gnd cell_6t
Xbit_r117_c134 bl_134 br_134 wl_117 vdd gnd cell_6t
Xbit_r118_c134 bl_134 br_134 wl_118 vdd gnd cell_6t
Xbit_r119_c134 bl_134 br_134 wl_119 vdd gnd cell_6t
Xbit_r120_c134 bl_134 br_134 wl_120 vdd gnd cell_6t
Xbit_r121_c134 bl_134 br_134 wl_121 vdd gnd cell_6t
Xbit_r122_c134 bl_134 br_134 wl_122 vdd gnd cell_6t
Xbit_r123_c134 bl_134 br_134 wl_123 vdd gnd cell_6t
Xbit_r124_c134 bl_134 br_134 wl_124 vdd gnd cell_6t
Xbit_r125_c134 bl_134 br_134 wl_125 vdd gnd cell_6t
Xbit_r126_c134 bl_134 br_134 wl_126 vdd gnd cell_6t
Xbit_r127_c134 bl_134 br_134 wl_127 vdd gnd cell_6t
Xbit_r128_c134 bl_134 br_134 wl_128 vdd gnd cell_6t
Xbit_r129_c134 bl_134 br_134 wl_129 vdd gnd cell_6t
Xbit_r130_c134 bl_134 br_134 wl_130 vdd gnd cell_6t
Xbit_r131_c134 bl_134 br_134 wl_131 vdd gnd cell_6t
Xbit_r132_c134 bl_134 br_134 wl_132 vdd gnd cell_6t
Xbit_r133_c134 bl_134 br_134 wl_133 vdd gnd cell_6t
Xbit_r134_c134 bl_134 br_134 wl_134 vdd gnd cell_6t
Xbit_r135_c134 bl_134 br_134 wl_135 vdd gnd cell_6t
Xbit_r136_c134 bl_134 br_134 wl_136 vdd gnd cell_6t
Xbit_r137_c134 bl_134 br_134 wl_137 vdd gnd cell_6t
Xbit_r138_c134 bl_134 br_134 wl_138 vdd gnd cell_6t
Xbit_r139_c134 bl_134 br_134 wl_139 vdd gnd cell_6t
Xbit_r140_c134 bl_134 br_134 wl_140 vdd gnd cell_6t
Xbit_r141_c134 bl_134 br_134 wl_141 vdd gnd cell_6t
Xbit_r142_c134 bl_134 br_134 wl_142 vdd gnd cell_6t
Xbit_r143_c134 bl_134 br_134 wl_143 vdd gnd cell_6t
Xbit_r144_c134 bl_134 br_134 wl_144 vdd gnd cell_6t
Xbit_r145_c134 bl_134 br_134 wl_145 vdd gnd cell_6t
Xbit_r146_c134 bl_134 br_134 wl_146 vdd gnd cell_6t
Xbit_r147_c134 bl_134 br_134 wl_147 vdd gnd cell_6t
Xbit_r148_c134 bl_134 br_134 wl_148 vdd gnd cell_6t
Xbit_r149_c134 bl_134 br_134 wl_149 vdd gnd cell_6t
Xbit_r150_c134 bl_134 br_134 wl_150 vdd gnd cell_6t
Xbit_r151_c134 bl_134 br_134 wl_151 vdd gnd cell_6t
Xbit_r152_c134 bl_134 br_134 wl_152 vdd gnd cell_6t
Xbit_r153_c134 bl_134 br_134 wl_153 vdd gnd cell_6t
Xbit_r154_c134 bl_134 br_134 wl_154 vdd gnd cell_6t
Xbit_r155_c134 bl_134 br_134 wl_155 vdd gnd cell_6t
Xbit_r156_c134 bl_134 br_134 wl_156 vdd gnd cell_6t
Xbit_r157_c134 bl_134 br_134 wl_157 vdd gnd cell_6t
Xbit_r158_c134 bl_134 br_134 wl_158 vdd gnd cell_6t
Xbit_r159_c134 bl_134 br_134 wl_159 vdd gnd cell_6t
Xbit_r160_c134 bl_134 br_134 wl_160 vdd gnd cell_6t
Xbit_r161_c134 bl_134 br_134 wl_161 vdd gnd cell_6t
Xbit_r162_c134 bl_134 br_134 wl_162 vdd gnd cell_6t
Xbit_r163_c134 bl_134 br_134 wl_163 vdd gnd cell_6t
Xbit_r164_c134 bl_134 br_134 wl_164 vdd gnd cell_6t
Xbit_r165_c134 bl_134 br_134 wl_165 vdd gnd cell_6t
Xbit_r166_c134 bl_134 br_134 wl_166 vdd gnd cell_6t
Xbit_r167_c134 bl_134 br_134 wl_167 vdd gnd cell_6t
Xbit_r168_c134 bl_134 br_134 wl_168 vdd gnd cell_6t
Xbit_r169_c134 bl_134 br_134 wl_169 vdd gnd cell_6t
Xbit_r170_c134 bl_134 br_134 wl_170 vdd gnd cell_6t
Xbit_r171_c134 bl_134 br_134 wl_171 vdd gnd cell_6t
Xbit_r172_c134 bl_134 br_134 wl_172 vdd gnd cell_6t
Xbit_r173_c134 bl_134 br_134 wl_173 vdd gnd cell_6t
Xbit_r174_c134 bl_134 br_134 wl_174 vdd gnd cell_6t
Xbit_r175_c134 bl_134 br_134 wl_175 vdd gnd cell_6t
Xbit_r176_c134 bl_134 br_134 wl_176 vdd gnd cell_6t
Xbit_r177_c134 bl_134 br_134 wl_177 vdd gnd cell_6t
Xbit_r178_c134 bl_134 br_134 wl_178 vdd gnd cell_6t
Xbit_r179_c134 bl_134 br_134 wl_179 vdd gnd cell_6t
Xbit_r180_c134 bl_134 br_134 wl_180 vdd gnd cell_6t
Xbit_r181_c134 bl_134 br_134 wl_181 vdd gnd cell_6t
Xbit_r182_c134 bl_134 br_134 wl_182 vdd gnd cell_6t
Xbit_r183_c134 bl_134 br_134 wl_183 vdd gnd cell_6t
Xbit_r184_c134 bl_134 br_134 wl_184 vdd gnd cell_6t
Xbit_r185_c134 bl_134 br_134 wl_185 vdd gnd cell_6t
Xbit_r186_c134 bl_134 br_134 wl_186 vdd gnd cell_6t
Xbit_r187_c134 bl_134 br_134 wl_187 vdd gnd cell_6t
Xbit_r188_c134 bl_134 br_134 wl_188 vdd gnd cell_6t
Xbit_r189_c134 bl_134 br_134 wl_189 vdd gnd cell_6t
Xbit_r190_c134 bl_134 br_134 wl_190 vdd gnd cell_6t
Xbit_r191_c134 bl_134 br_134 wl_191 vdd gnd cell_6t
Xbit_r192_c134 bl_134 br_134 wl_192 vdd gnd cell_6t
Xbit_r193_c134 bl_134 br_134 wl_193 vdd gnd cell_6t
Xbit_r194_c134 bl_134 br_134 wl_194 vdd gnd cell_6t
Xbit_r195_c134 bl_134 br_134 wl_195 vdd gnd cell_6t
Xbit_r196_c134 bl_134 br_134 wl_196 vdd gnd cell_6t
Xbit_r197_c134 bl_134 br_134 wl_197 vdd gnd cell_6t
Xbit_r198_c134 bl_134 br_134 wl_198 vdd gnd cell_6t
Xbit_r199_c134 bl_134 br_134 wl_199 vdd gnd cell_6t
Xbit_r200_c134 bl_134 br_134 wl_200 vdd gnd cell_6t
Xbit_r201_c134 bl_134 br_134 wl_201 vdd gnd cell_6t
Xbit_r202_c134 bl_134 br_134 wl_202 vdd gnd cell_6t
Xbit_r203_c134 bl_134 br_134 wl_203 vdd gnd cell_6t
Xbit_r204_c134 bl_134 br_134 wl_204 vdd gnd cell_6t
Xbit_r205_c134 bl_134 br_134 wl_205 vdd gnd cell_6t
Xbit_r206_c134 bl_134 br_134 wl_206 vdd gnd cell_6t
Xbit_r207_c134 bl_134 br_134 wl_207 vdd gnd cell_6t
Xbit_r208_c134 bl_134 br_134 wl_208 vdd gnd cell_6t
Xbit_r209_c134 bl_134 br_134 wl_209 vdd gnd cell_6t
Xbit_r210_c134 bl_134 br_134 wl_210 vdd gnd cell_6t
Xbit_r211_c134 bl_134 br_134 wl_211 vdd gnd cell_6t
Xbit_r212_c134 bl_134 br_134 wl_212 vdd gnd cell_6t
Xbit_r213_c134 bl_134 br_134 wl_213 vdd gnd cell_6t
Xbit_r214_c134 bl_134 br_134 wl_214 vdd gnd cell_6t
Xbit_r215_c134 bl_134 br_134 wl_215 vdd gnd cell_6t
Xbit_r216_c134 bl_134 br_134 wl_216 vdd gnd cell_6t
Xbit_r217_c134 bl_134 br_134 wl_217 vdd gnd cell_6t
Xbit_r218_c134 bl_134 br_134 wl_218 vdd gnd cell_6t
Xbit_r219_c134 bl_134 br_134 wl_219 vdd gnd cell_6t
Xbit_r220_c134 bl_134 br_134 wl_220 vdd gnd cell_6t
Xbit_r221_c134 bl_134 br_134 wl_221 vdd gnd cell_6t
Xbit_r222_c134 bl_134 br_134 wl_222 vdd gnd cell_6t
Xbit_r223_c134 bl_134 br_134 wl_223 vdd gnd cell_6t
Xbit_r224_c134 bl_134 br_134 wl_224 vdd gnd cell_6t
Xbit_r225_c134 bl_134 br_134 wl_225 vdd gnd cell_6t
Xbit_r226_c134 bl_134 br_134 wl_226 vdd gnd cell_6t
Xbit_r227_c134 bl_134 br_134 wl_227 vdd gnd cell_6t
Xbit_r228_c134 bl_134 br_134 wl_228 vdd gnd cell_6t
Xbit_r229_c134 bl_134 br_134 wl_229 vdd gnd cell_6t
Xbit_r230_c134 bl_134 br_134 wl_230 vdd gnd cell_6t
Xbit_r231_c134 bl_134 br_134 wl_231 vdd gnd cell_6t
Xbit_r232_c134 bl_134 br_134 wl_232 vdd gnd cell_6t
Xbit_r233_c134 bl_134 br_134 wl_233 vdd gnd cell_6t
Xbit_r234_c134 bl_134 br_134 wl_234 vdd gnd cell_6t
Xbit_r235_c134 bl_134 br_134 wl_235 vdd gnd cell_6t
Xbit_r236_c134 bl_134 br_134 wl_236 vdd gnd cell_6t
Xbit_r237_c134 bl_134 br_134 wl_237 vdd gnd cell_6t
Xbit_r238_c134 bl_134 br_134 wl_238 vdd gnd cell_6t
Xbit_r239_c134 bl_134 br_134 wl_239 vdd gnd cell_6t
Xbit_r240_c134 bl_134 br_134 wl_240 vdd gnd cell_6t
Xbit_r241_c134 bl_134 br_134 wl_241 vdd gnd cell_6t
Xbit_r242_c134 bl_134 br_134 wl_242 vdd gnd cell_6t
Xbit_r243_c134 bl_134 br_134 wl_243 vdd gnd cell_6t
Xbit_r244_c134 bl_134 br_134 wl_244 vdd gnd cell_6t
Xbit_r245_c134 bl_134 br_134 wl_245 vdd gnd cell_6t
Xbit_r246_c134 bl_134 br_134 wl_246 vdd gnd cell_6t
Xbit_r247_c134 bl_134 br_134 wl_247 vdd gnd cell_6t
Xbit_r248_c134 bl_134 br_134 wl_248 vdd gnd cell_6t
Xbit_r249_c134 bl_134 br_134 wl_249 vdd gnd cell_6t
Xbit_r250_c134 bl_134 br_134 wl_250 vdd gnd cell_6t
Xbit_r251_c134 bl_134 br_134 wl_251 vdd gnd cell_6t
Xbit_r252_c134 bl_134 br_134 wl_252 vdd gnd cell_6t
Xbit_r253_c134 bl_134 br_134 wl_253 vdd gnd cell_6t
Xbit_r254_c134 bl_134 br_134 wl_254 vdd gnd cell_6t
Xbit_r255_c134 bl_134 br_134 wl_255 vdd gnd cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd cell_6t
Xbit_r1_c135 bl_135 br_135 wl_1 vdd gnd cell_6t
Xbit_r2_c135 bl_135 br_135 wl_2 vdd gnd cell_6t
Xbit_r3_c135 bl_135 br_135 wl_3 vdd gnd cell_6t
Xbit_r4_c135 bl_135 br_135 wl_4 vdd gnd cell_6t
Xbit_r5_c135 bl_135 br_135 wl_5 vdd gnd cell_6t
Xbit_r6_c135 bl_135 br_135 wl_6 vdd gnd cell_6t
Xbit_r7_c135 bl_135 br_135 wl_7 vdd gnd cell_6t
Xbit_r8_c135 bl_135 br_135 wl_8 vdd gnd cell_6t
Xbit_r9_c135 bl_135 br_135 wl_9 vdd gnd cell_6t
Xbit_r10_c135 bl_135 br_135 wl_10 vdd gnd cell_6t
Xbit_r11_c135 bl_135 br_135 wl_11 vdd gnd cell_6t
Xbit_r12_c135 bl_135 br_135 wl_12 vdd gnd cell_6t
Xbit_r13_c135 bl_135 br_135 wl_13 vdd gnd cell_6t
Xbit_r14_c135 bl_135 br_135 wl_14 vdd gnd cell_6t
Xbit_r15_c135 bl_135 br_135 wl_15 vdd gnd cell_6t
Xbit_r16_c135 bl_135 br_135 wl_16 vdd gnd cell_6t
Xbit_r17_c135 bl_135 br_135 wl_17 vdd gnd cell_6t
Xbit_r18_c135 bl_135 br_135 wl_18 vdd gnd cell_6t
Xbit_r19_c135 bl_135 br_135 wl_19 vdd gnd cell_6t
Xbit_r20_c135 bl_135 br_135 wl_20 vdd gnd cell_6t
Xbit_r21_c135 bl_135 br_135 wl_21 vdd gnd cell_6t
Xbit_r22_c135 bl_135 br_135 wl_22 vdd gnd cell_6t
Xbit_r23_c135 bl_135 br_135 wl_23 vdd gnd cell_6t
Xbit_r24_c135 bl_135 br_135 wl_24 vdd gnd cell_6t
Xbit_r25_c135 bl_135 br_135 wl_25 vdd gnd cell_6t
Xbit_r26_c135 bl_135 br_135 wl_26 vdd gnd cell_6t
Xbit_r27_c135 bl_135 br_135 wl_27 vdd gnd cell_6t
Xbit_r28_c135 bl_135 br_135 wl_28 vdd gnd cell_6t
Xbit_r29_c135 bl_135 br_135 wl_29 vdd gnd cell_6t
Xbit_r30_c135 bl_135 br_135 wl_30 vdd gnd cell_6t
Xbit_r31_c135 bl_135 br_135 wl_31 vdd gnd cell_6t
Xbit_r32_c135 bl_135 br_135 wl_32 vdd gnd cell_6t
Xbit_r33_c135 bl_135 br_135 wl_33 vdd gnd cell_6t
Xbit_r34_c135 bl_135 br_135 wl_34 vdd gnd cell_6t
Xbit_r35_c135 bl_135 br_135 wl_35 vdd gnd cell_6t
Xbit_r36_c135 bl_135 br_135 wl_36 vdd gnd cell_6t
Xbit_r37_c135 bl_135 br_135 wl_37 vdd gnd cell_6t
Xbit_r38_c135 bl_135 br_135 wl_38 vdd gnd cell_6t
Xbit_r39_c135 bl_135 br_135 wl_39 vdd gnd cell_6t
Xbit_r40_c135 bl_135 br_135 wl_40 vdd gnd cell_6t
Xbit_r41_c135 bl_135 br_135 wl_41 vdd gnd cell_6t
Xbit_r42_c135 bl_135 br_135 wl_42 vdd gnd cell_6t
Xbit_r43_c135 bl_135 br_135 wl_43 vdd gnd cell_6t
Xbit_r44_c135 bl_135 br_135 wl_44 vdd gnd cell_6t
Xbit_r45_c135 bl_135 br_135 wl_45 vdd gnd cell_6t
Xbit_r46_c135 bl_135 br_135 wl_46 vdd gnd cell_6t
Xbit_r47_c135 bl_135 br_135 wl_47 vdd gnd cell_6t
Xbit_r48_c135 bl_135 br_135 wl_48 vdd gnd cell_6t
Xbit_r49_c135 bl_135 br_135 wl_49 vdd gnd cell_6t
Xbit_r50_c135 bl_135 br_135 wl_50 vdd gnd cell_6t
Xbit_r51_c135 bl_135 br_135 wl_51 vdd gnd cell_6t
Xbit_r52_c135 bl_135 br_135 wl_52 vdd gnd cell_6t
Xbit_r53_c135 bl_135 br_135 wl_53 vdd gnd cell_6t
Xbit_r54_c135 bl_135 br_135 wl_54 vdd gnd cell_6t
Xbit_r55_c135 bl_135 br_135 wl_55 vdd gnd cell_6t
Xbit_r56_c135 bl_135 br_135 wl_56 vdd gnd cell_6t
Xbit_r57_c135 bl_135 br_135 wl_57 vdd gnd cell_6t
Xbit_r58_c135 bl_135 br_135 wl_58 vdd gnd cell_6t
Xbit_r59_c135 bl_135 br_135 wl_59 vdd gnd cell_6t
Xbit_r60_c135 bl_135 br_135 wl_60 vdd gnd cell_6t
Xbit_r61_c135 bl_135 br_135 wl_61 vdd gnd cell_6t
Xbit_r62_c135 bl_135 br_135 wl_62 vdd gnd cell_6t
Xbit_r63_c135 bl_135 br_135 wl_63 vdd gnd cell_6t
Xbit_r64_c135 bl_135 br_135 wl_64 vdd gnd cell_6t
Xbit_r65_c135 bl_135 br_135 wl_65 vdd gnd cell_6t
Xbit_r66_c135 bl_135 br_135 wl_66 vdd gnd cell_6t
Xbit_r67_c135 bl_135 br_135 wl_67 vdd gnd cell_6t
Xbit_r68_c135 bl_135 br_135 wl_68 vdd gnd cell_6t
Xbit_r69_c135 bl_135 br_135 wl_69 vdd gnd cell_6t
Xbit_r70_c135 bl_135 br_135 wl_70 vdd gnd cell_6t
Xbit_r71_c135 bl_135 br_135 wl_71 vdd gnd cell_6t
Xbit_r72_c135 bl_135 br_135 wl_72 vdd gnd cell_6t
Xbit_r73_c135 bl_135 br_135 wl_73 vdd gnd cell_6t
Xbit_r74_c135 bl_135 br_135 wl_74 vdd gnd cell_6t
Xbit_r75_c135 bl_135 br_135 wl_75 vdd gnd cell_6t
Xbit_r76_c135 bl_135 br_135 wl_76 vdd gnd cell_6t
Xbit_r77_c135 bl_135 br_135 wl_77 vdd gnd cell_6t
Xbit_r78_c135 bl_135 br_135 wl_78 vdd gnd cell_6t
Xbit_r79_c135 bl_135 br_135 wl_79 vdd gnd cell_6t
Xbit_r80_c135 bl_135 br_135 wl_80 vdd gnd cell_6t
Xbit_r81_c135 bl_135 br_135 wl_81 vdd gnd cell_6t
Xbit_r82_c135 bl_135 br_135 wl_82 vdd gnd cell_6t
Xbit_r83_c135 bl_135 br_135 wl_83 vdd gnd cell_6t
Xbit_r84_c135 bl_135 br_135 wl_84 vdd gnd cell_6t
Xbit_r85_c135 bl_135 br_135 wl_85 vdd gnd cell_6t
Xbit_r86_c135 bl_135 br_135 wl_86 vdd gnd cell_6t
Xbit_r87_c135 bl_135 br_135 wl_87 vdd gnd cell_6t
Xbit_r88_c135 bl_135 br_135 wl_88 vdd gnd cell_6t
Xbit_r89_c135 bl_135 br_135 wl_89 vdd gnd cell_6t
Xbit_r90_c135 bl_135 br_135 wl_90 vdd gnd cell_6t
Xbit_r91_c135 bl_135 br_135 wl_91 vdd gnd cell_6t
Xbit_r92_c135 bl_135 br_135 wl_92 vdd gnd cell_6t
Xbit_r93_c135 bl_135 br_135 wl_93 vdd gnd cell_6t
Xbit_r94_c135 bl_135 br_135 wl_94 vdd gnd cell_6t
Xbit_r95_c135 bl_135 br_135 wl_95 vdd gnd cell_6t
Xbit_r96_c135 bl_135 br_135 wl_96 vdd gnd cell_6t
Xbit_r97_c135 bl_135 br_135 wl_97 vdd gnd cell_6t
Xbit_r98_c135 bl_135 br_135 wl_98 vdd gnd cell_6t
Xbit_r99_c135 bl_135 br_135 wl_99 vdd gnd cell_6t
Xbit_r100_c135 bl_135 br_135 wl_100 vdd gnd cell_6t
Xbit_r101_c135 bl_135 br_135 wl_101 vdd gnd cell_6t
Xbit_r102_c135 bl_135 br_135 wl_102 vdd gnd cell_6t
Xbit_r103_c135 bl_135 br_135 wl_103 vdd gnd cell_6t
Xbit_r104_c135 bl_135 br_135 wl_104 vdd gnd cell_6t
Xbit_r105_c135 bl_135 br_135 wl_105 vdd gnd cell_6t
Xbit_r106_c135 bl_135 br_135 wl_106 vdd gnd cell_6t
Xbit_r107_c135 bl_135 br_135 wl_107 vdd gnd cell_6t
Xbit_r108_c135 bl_135 br_135 wl_108 vdd gnd cell_6t
Xbit_r109_c135 bl_135 br_135 wl_109 vdd gnd cell_6t
Xbit_r110_c135 bl_135 br_135 wl_110 vdd gnd cell_6t
Xbit_r111_c135 bl_135 br_135 wl_111 vdd gnd cell_6t
Xbit_r112_c135 bl_135 br_135 wl_112 vdd gnd cell_6t
Xbit_r113_c135 bl_135 br_135 wl_113 vdd gnd cell_6t
Xbit_r114_c135 bl_135 br_135 wl_114 vdd gnd cell_6t
Xbit_r115_c135 bl_135 br_135 wl_115 vdd gnd cell_6t
Xbit_r116_c135 bl_135 br_135 wl_116 vdd gnd cell_6t
Xbit_r117_c135 bl_135 br_135 wl_117 vdd gnd cell_6t
Xbit_r118_c135 bl_135 br_135 wl_118 vdd gnd cell_6t
Xbit_r119_c135 bl_135 br_135 wl_119 vdd gnd cell_6t
Xbit_r120_c135 bl_135 br_135 wl_120 vdd gnd cell_6t
Xbit_r121_c135 bl_135 br_135 wl_121 vdd gnd cell_6t
Xbit_r122_c135 bl_135 br_135 wl_122 vdd gnd cell_6t
Xbit_r123_c135 bl_135 br_135 wl_123 vdd gnd cell_6t
Xbit_r124_c135 bl_135 br_135 wl_124 vdd gnd cell_6t
Xbit_r125_c135 bl_135 br_135 wl_125 vdd gnd cell_6t
Xbit_r126_c135 bl_135 br_135 wl_126 vdd gnd cell_6t
Xbit_r127_c135 bl_135 br_135 wl_127 vdd gnd cell_6t
Xbit_r128_c135 bl_135 br_135 wl_128 vdd gnd cell_6t
Xbit_r129_c135 bl_135 br_135 wl_129 vdd gnd cell_6t
Xbit_r130_c135 bl_135 br_135 wl_130 vdd gnd cell_6t
Xbit_r131_c135 bl_135 br_135 wl_131 vdd gnd cell_6t
Xbit_r132_c135 bl_135 br_135 wl_132 vdd gnd cell_6t
Xbit_r133_c135 bl_135 br_135 wl_133 vdd gnd cell_6t
Xbit_r134_c135 bl_135 br_135 wl_134 vdd gnd cell_6t
Xbit_r135_c135 bl_135 br_135 wl_135 vdd gnd cell_6t
Xbit_r136_c135 bl_135 br_135 wl_136 vdd gnd cell_6t
Xbit_r137_c135 bl_135 br_135 wl_137 vdd gnd cell_6t
Xbit_r138_c135 bl_135 br_135 wl_138 vdd gnd cell_6t
Xbit_r139_c135 bl_135 br_135 wl_139 vdd gnd cell_6t
Xbit_r140_c135 bl_135 br_135 wl_140 vdd gnd cell_6t
Xbit_r141_c135 bl_135 br_135 wl_141 vdd gnd cell_6t
Xbit_r142_c135 bl_135 br_135 wl_142 vdd gnd cell_6t
Xbit_r143_c135 bl_135 br_135 wl_143 vdd gnd cell_6t
Xbit_r144_c135 bl_135 br_135 wl_144 vdd gnd cell_6t
Xbit_r145_c135 bl_135 br_135 wl_145 vdd gnd cell_6t
Xbit_r146_c135 bl_135 br_135 wl_146 vdd gnd cell_6t
Xbit_r147_c135 bl_135 br_135 wl_147 vdd gnd cell_6t
Xbit_r148_c135 bl_135 br_135 wl_148 vdd gnd cell_6t
Xbit_r149_c135 bl_135 br_135 wl_149 vdd gnd cell_6t
Xbit_r150_c135 bl_135 br_135 wl_150 vdd gnd cell_6t
Xbit_r151_c135 bl_135 br_135 wl_151 vdd gnd cell_6t
Xbit_r152_c135 bl_135 br_135 wl_152 vdd gnd cell_6t
Xbit_r153_c135 bl_135 br_135 wl_153 vdd gnd cell_6t
Xbit_r154_c135 bl_135 br_135 wl_154 vdd gnd cell_6t
Xbit_r155_c135 bl_135 br_135 wl_155 vdd gnd cell_6t
Xbit_r156_c135 bl_135 br_135 wl_156 vdd gnd cell_6t
Xbit_r157_c135 bl_135 br_135 wl_157 vdd gnd cell_6t
Xbit_r158_c135 bl_135 br_135 wl_158 vdd gnd cell_6t
Xbit_r159_c135 bl_135 br_135 wl_159 vdd gnd cell_6t
Xbit_r160_c135 bl_135 br_135 wl_160 vdd gnd cell_6t
Xbit_r161_c135 bl_135 br_135 wl_161 vdd gnd cell_6t
Xbit_r162_c135 bl_135 br_135 wl_162 vdd gnd cell_6t
Xbit_r163_c135 bl_135 br_135 wl_163 vdd gnd cell_6t
Xbit_r164_c135 bl_135 br_135 wl_164 vdd gnd cell_6t
Xbit_r165_c135 bl_135 br_135 wl_165 vdd gnd cell_6t
Xbit_r166_c135 bl_135 br_135 wl_166 vdd gnd cell_6t
Xbit_r167_c135 bl_135 br_135 wl_167 vdd gnd cell_6t
Xbit_r168_c135 bl_135 br_135 wl_168 vdd gnd cell_6t
Xbit_r169_c135 bl_135 br_135 wl_169 vdd gnd cell_6t
Xbit_r170_c135 bl_135 br_135 wl_170 vdd gnd cell_6t
Xbit_r171_c135 bl_135 br_135 wl_171 vdd gnd cell_6t
Xbit_r172_c135 bl_135 br_135 wl_172 vdd gnd cell_6t
Xbit_r173_c135 bl_135 br_135 wl_173 vdd gnd cell_6t
Xbit_r174_c135 bl_135 br_135 wl_174 vdd gnd cell_6t
Xbit_r175_c135 bl_135 br_135 wl_175 vdd gnd cell_6t
Xbit_r176_c135 bl_135 br_135 wl_176 vdd gnd cell_6t
Xbit_r177_c135 bl_135 br_135 wl_177 vdd gnd cell_6t
Xbit_r178_c135 bl_135 br_135 wl_178 vdd gnd cell_6t
Xbit_r179_c135 bl_135 br_135 wl_179 vdd gnd cell_6t
Xbit_r180_c135 bl_135 br_135 wl_180 vdd gnd cell_6t
Xbit_r181_c135 bl_135 br_135 wl_181 vdd gnd cell_6t
Xbit_r182_c135 bl_135 br_135 wl_182 vdd gnd cell_6t
Xbit_r183_c135 bl_135 br_135 wl_183 vdd gnd cell_6t
Xbit_r184_c135 bl_135 br_135 wl_184 vdd gnd cell_6t
Xbit_r185_c135 bl_135 br_135 wl_185 vdd gnd cell_6t
Xbit_r186_c135 bl_135 br_135 wl_186 vdd gnd cell_6t
Xbit_r187_c135 bl_135 br_135 wl_187 vdd gnd cell_6t
Xbit_r188_c135 bl_135 br_135 wl_188 vdd gnd cell_6t
Xbit_r189_c135 bl_135 br_135 wl_189 vdd gnd cell_6t
Xbit_r190_c135 bl_135 br_135 wl_190 vdd gnd cell_6t
Xbit_r191_c135 bl_135 br_135 wl_191 vdd gnd cell_6t
Xbit_r192_c135 bl_135 br_135 wl_192 vdd gnd cell_6t
Xbit_r193_c135 bl_135 br_135 wl_193 vdd gnd cell_6t
Xbit_r194_c135 bl_135 br_135 wl_194 vdd gnd cell_6t
Xbit_r195_c135 bl_135 br_135 wl_195 vdd gnd cell_6t
Xbit_r196_c135 bl_135 br_135 wl_196 vdd gnd cell_6t
Xbit_r197_c135 bl_135 br_135 wl_197 vdd gnd cell_6t
Xbit_r198_c135 bl_135 br_135 wl_198 vdd gnd cell_6t
Xbit_r199_c135 bl_135 br_135 wl_199 vdd gnd cell_6t
Xbit_r200_c135 bl_135 br_135 wl_200 vdd gnd cell_6t
Xbit_r201_c135 bl_135 br_135 wl_201 vdd gnd cell_6t
Xbit_r202_c135 bl_135 br_135 wl_202 vdd gnd cell_6t
Xbit_r203_c135 bl_135 br_135 wl_203 vdd gnd cell_6t
Xbit_r204_c135 bl_135 br_135 wl_204 vdd gnd cell_6t
Xbit_r205_c135 bl_135 br_135 wl_205 vdd gnd cell_6t
Xbit_r206_c135 bl_135 br_135 wl_206 vdd gnd cell_6t
Xbit_r207_c135 bl_135 br_135 wl_207 vdd gnd cell_6t
Xbit_r208_c135 bl_135 br_135 wl_208 vdd gnd cell_6t
Xbit_r209_c135 bl_135 br_135 wl_209 vdd gnd cell_6t
Xbit_r210_c135 bl_135 br_135 wl_210 vdd gnd cell_6t
Xbit_r211_c135 bl_135 br_135 wl_211 vdd gnd cell_6t
Xbit_r212_c135 bl_135 br_135 wl_212 vdd gnd cell_6t
Xbit_r213_c135 bl_135 br_135 wl_213 vdd gnd cell_6t
Xbit_r214_c135 bl_135 br_135 wl_214 vdd gnd cell_6t
Xbit_r215_c135 bl_135 br_135 wl_215 vdd gnd cell_6t
Xbit_r216_c135 bl_135 br_135 wl_216 vdd gnd cell_6t
Xbit_r217_c135 bl_135 br_135 wl_217 vdd gnd cell_6t
Xbit_r218_c135 bl_135 br_135 wl_218 vdd gnd cell_6t
Xbit_r219_c135 bl_135 br_135 wl_219 vdd gnd cell_6t
Xbit_r220_c135 bl_135 br_135 wl_220 vdd gnd cell_6t
Xbit_r221_c135 bl_135 br_135 wl_221 vdd gnd cell_6t
Xbit_r222_c135 bl_135 br_135 wl_222 vdd gnd cell_6t
Xbit_r223_c135 bl_135 br_135 wl_223 vdd gnd cell_6t
Xbit_r224_c135 bl_135 br_135 wl_224 vdd gnd cell_6t
Xbit_r225_c135 bl_135 br_135 wl_225 vdd gnd cell_6t
Xbit_r226_c135 bl_135 br_135 wl_226 vdd gnd cell_6t
Xbit_r227_c135 bl_135 br_135 wl_227 vdd gnd cell_6t
Xbit_r228_c135 bl_135 br_135 wl_228 vdd gnd cell_6t
Xbit_r229_c135 bl_135 br_135 wl_229 vdd gnd cell_6t
Xbit_r230_c135 bl_135 br_135 wl_230 vdd gnd cell_6t
Xbit_r231_c135 bl_135 br_135 wl_231 vdd gnd cell_6t
Xbit_r232_c135 bl_135 br_135 wl_232 vdd gnd cell_6t
Xbit_r233_c135 bl_135 br_135 wl_233 vdd gnd cell_6t
Xbit_r234_c135 bl_135 br_135 wl_234 vdd gnd cell_6t
Xbit_r235_c135 bl_135 br_135 wl_235 vdd gnd cell_6t
Xbit_r236_c135 bl_135 br_135 wl_236 vdd gnd cell_6t
Xbit_r237_c135 bl_135 br_135 wl_237 vdd gnd cell_6t
Xbit_r238_c135 bl_135 br_135 wl_238 vdd gnd cell_6t
Xbit_r239_c135 bl_135 br_135 wl_239 vdd gnd cell_6t
Xbit_r240_c135 bl_135 br_135 wl_240 vdd gnd cell_6t
Xbit_r241_c135 bl_135 br_135 wl_241 vdd gnd cell_6t
Xbit_r242_c135 bl_135 br_135 wl_242 vdd gnd cell_6t
Xbit_r243_c135 bl_135 br_135 wl_243 vdd gnd cell_6t
Xbit_r244_c135 bl_135 br_135 wl_244 vdd gnd cell_6t
Xbit_r245_c135 bl_135 br_135 wl_245 vdd gnd cell_6t
Xbit_r246_c135 bl_135 br_135 wl_246 vdd gnd cell_6t
Xbit_r247_c135 bl_135 br_135 wl_247 vdd gnd cell_6t
Xbit_r248_c135 bl_135 br_135 wl_248 vdd gnd cell_6t
Xbit_r249_c135 bl_135 br_135 wl_249 vdd gnd cell_6t
Xbit_r250_c135 bl_135 br_135 wl_250 vdd gnd cell_6t
Xbit_r251_c135 bl_135 br_135 wl_251 vdd gnd cell_6t
Xbit_r252_c135 bl_135 br_135 wl_252 vdd gnd cell_6t
Xbit_r253_c135 bl_135 br_135 wl_253 vdd gnd cell_6t
Xbit_r254_c135 bl_135 br_135 wl_254 vdd gnd cell_6t
Xbit_r255_c135 bl_135 br_135 wl_255 vdd gnd cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd cell_6t
Xbit_r1_c136 bl_136 br_136 wl_1 vdd gnd cell_6t
Xbit_r2_c136 bl_136 br_136 wl_2 vdd gnd cell_6t
Xbit_r3_c136 bl_136 br_136 wl_3 vdd gnd cell_6t
Xbit_r4_c136 bl_136 br_136 wl_4 vdd gnd cell_6t
Xbit_r5_c136 bl_136 br_136 wl_5 vdd gnd cell_6t
Xbit_r6_c136 bl_136 br_136 wl_6 vdd gnd cell_6t
Xbit_r7_c136 bl_136 br_136 wl_7 vdd gnd cell_6t
Xbit_r8_c136 bl_136 br_136 wl_8 vdd gnd cell_6t
Xbit_r9_c136 bl_136 br_136 wl_9 vdd gnd cell_6t
Xbit_r10_c136 bl_136 br_136 wl_10 vdd gnd cell_6t
Xbit_r11_c136 bl_136 br_136 wl_11 vdd gnd cell_6t
Xbit_r12_c136 bl_136 br_136 wl_12 vdd gnd cell_6t
Xbit_r13_c136 bl_136 br_136 wl_13 vdd gnd cell_6t
Xbit_r14_c136 bl_136 br_136 wl_14 vdd gnd cell_6t
Xbit_r15_c136 bl_136 br_136 wl_15 vdd gnd cell_6t
Xbit_r16_c136 bl_136 br_136 wl_16 vdd gnd cell_6t
Xbit_r17_c136 bl_136 br_136 wl_17 vdd gnd cell_6t
Xbit_r18_c136 bl_136 br_136 wl_18 vdd gnd cell_6t
Xbit_r19_c136 bl_136 br_136 wl_19 vdd gnd cell_6t
Xbit_r20_c136 bl_136 br_136 wl_20 vdd gnd cell_6t
Xbit_r21_c136 bl_136 br_136 wl_21 vdd gnd cell_6t
Xbit_r22_c136 bl_136 br_136 wl_22 vdd gnd cell_6t
Xbit_r23_c136 bl_136 br_136 wl_23 vdd gnd cell_6t
Xbit_r24_c136 bl_136 br_136 wl_24 vdd gnd cell_6t
Xbit_r25_c136 bl_136 br_136 wl_25 vdd gnd cell_6t
Xbit_r26_c136 bl_136 br_136 wl_26 vdd gnd cell_6t
Xbit_r27_c136 bl_136 br_136 wl_27 vdd gnd cell_6t
Xbit_r28_c136 bl_136 br_136 wl_28 vdd gnd cell_6t
Xbit_r29_c136 bl_136 br_136 wl_29 vdd gnd cell_6t
Xbit_r30_c136 bl_136 br_136 wl_30 vdd gnd cell_6t
Xbit_r31_c136 bl_136 br_136 wl_31 vdd gnd cell_6t
Xbit_r32_c136 bl_136 br_136 wl_32 vdd gnd cell_6t
Xbit_r33_c136 bl_136 br_136 wl_33 vdd gnd cell_6t
Xbit_r34_c136 bl_136 br_136 wl_34 vdd gnd cell_6t
Xbit_r35_c136 bl_136 br_136 wl_35 vdd gnd cell_6t
Xbit_r36_c136 bl_136 br_136 wl_36 vdd gnd cell_6t
Xbit_r37_c136 bl_136 br_136 wl_37 vdd gnd cell_6t
Xbit_r38_c136 bl_136 br_136 wl_38 vdd gnd cell_6t
Xbit_r39_c136 bl_136 br_136 wl_39 vdd gnd cell_6t
Xbit_r40_c136 bl_136 br_136 wl_40 vdd gnd cell_6t
Xbit_r41_c136 bl_136 br_136 wl_41 vdd gnd cell_6t
Xbit_r42_c136 bl_136 br_136 wl_42 vdd gnd cell_6t
Xbit_r43_c136 bl_136 br_136 wl_43 vdd gnd cell_6t
Xbit_r44_c136 bl_136 br_136 wl_44 vdd gnd cell_6t
Xbit_r45_c136 bl_136 br_136 wl_45 vdd gnd cell_6t
Xbit_r46_c136 bl_136 br_136 wl_46 vdd gnd cell_6t
Xbit_r47_c136 bl_136 br_136 wl_47 vdd gnd cell_6t
Xbit_r48_c136 bl_136 br_136 wl_48 vdd gnd cell_6t
Xbit_r49_c136 bl_136 br_136 wl_49 vdd gnd cell_6t
Xbit_r50_c136 bl_136 br_136 wl_50 vdd gnd cell_6t
Xbit_r51_c136 bl_136 br_136 wl_51 vdd gnd cell_6t
Xbit_r52_c136 bl_136 br_136 wl_52 vdd gnd cell_6t
Xbit_r53_c136 bl_136 br_136 wl_53 vdd gnd cell_6t
Xbit_r54_c136 bl_136 br_136 wl_54 vdd gnd cell_6t
Xbit_r55_c136 bl_136 br_136 wl_55 vdd gnd cell_6t
Xbit_r56_c136 bl_136 br_136 wl_56 vdd gnd cell_6t
Xbit_r57_c136 bl_136 br_136 wl_57 vdd gnd cell_6t
Xbit_r58_c136 bl_136 br_136 wl_58 vdd gnd cell_6t
Xbit_r59_c136 bl_136 br_136 wl_59 vdd gnd cell_6t
Xbit_r60_c136 bl_136 br_136 wl_60 vdd gnd cell_6t
Xbit_r61_c136 bl_136 br_136 wl_61 vdd gnd cell_6t
Xbit_r62_c136 bl_136 br_136 wl_62 vdd gnd cell_6t
Xbit_r63_c136 bl_136 br_136 wl_63 vdd gnd cell_6t
Xbit_r64_c136 bl_136 br_136 wl_64 vdd gnd cell_6t
Xbit_r65_c136 bl_136 br_136 wl_65 vdd gnd cell_6t
Xbit_r66_c136 bl_136 br_136 wl_66 vdd gnd cell_6t
Xbit_r67_c136 bl_136 br_136 wl_67 vdd gnd cell_6t
Xbit_r68_c136 bl_136 br_136 wl_68 vdd gnd cell_6t
Xbit_r69_c136 bl_136 br_136 wl_69 vdd gnd cell_6t
Xbit_r70_c136 bl_136 br_136 wl_70 vdd gnd cell_6t
Xbit_r71_c136 bl_136 br_136 wl_71 vdd gnd cell_6t
Xbit_r72_c136 bl_136 br_136 wl_72 vdd gnd cell_6t
Xbit_r73_c136 bl_136 br_136 wl_73 vdd gnd cell_6t
Xbit_r74_c136 bl_136 br_136 wl_74 vdd gnd cell_6t
Xbit_r75_c136 bl_136 br_136 wl_75 vdd gnd cell_6t
Xbit_r76_c136 bl_136 br_136 wl_76 vdd gnd cell_6t
Xbit_r77_c136 bl_136 br_136 wl_77 vdd gnd cell_6t
Xbit_r78_c136 bl_136 br_136 wl_78 vdd gnd cell_6t
Xbit_r79_c136 bl_136 br_136 wl_79 vdd gnd cell_6t
Xbit_r80_c136 bl_136 br_136 wl_80 vdd gnd cell_6t
Xbit_r81_c136 bl_136 br_136 wl_81 vdd gnd cell_6t
Xbit_r82_c136 bl_136 br_136 wl_82 vdd gnd cell_6t
Xbit_r83_c136 bl_136 br_136 wl_83 vdd gnd cell_6t
Xbit_r84_c136 bl_136 br_136 wl_84 vdd gnd cell_6t
Xbit_r85_c136 bl_136 br_136 wl_85 vdd gnd cell_6t
Xbit_r86_c136 bl_136 br_136 wl_86 vdd gnd cell_6t
Xbit_r87_c136 bl_136 br_136 wl_87 vdd gnd cell_6t
Xbit_r88_c136 bl_136 br_136 wl_88 vdd gnd cell_6t
Xbit_r89_c136 bl_136 br_136 wl_89 vdd gnd cell_6t
Xbit_r90_c136 bl_136 br_136 wl_90 vdd gnd cell_6t
Xbit_r91_c136 bl_136 br_136 wl_91 vdd gnd cell_6t
Xbit_r92_c136 bl_136 br_136 wl_92 vdd gnd cell_6t
Xbit_r93_c136 bl_136 br_136 wl_93 vdd gnd cell_6t
Xbit_r94_c136 bl_136 br_136 wl_94 vdd gnd cell_6t
Xbit_r95_c136 bl_136 br_136 wl_95 vdd gnd cell_6t
Xbit_r96_c136 bl_136 br_136 wl_96 vdd gnd cell_6t
Xbit_r97_c136 bl_136 br_136 wl_97 vdd gnd cell_6t
Xbit_r98_c136 bl_136 br_136 wl_98 vdd gnd cell_6t
Xbit_r99_c136 bl_136 br_136 wl_99 vdd gnd cell_6t
Xbit_r100_c136 bl_136 br_136 wl_100 vdd gnd cell_6t
Xbit_r101_c136 bl_136 br_136 wl_101 vdd gnd cell_6t
Xbit_r102_c136 bl_136 br_136 wl_102 vdd gnd cell_6t
Xbit_r103_c136 bl_136 br_136 wl_103 vdd gnd cell_6t
Xbit_r104_c136 bl_136 br_136 wl_104 vdd gnd cell_6t
Xbit_r105_c136 bl_136 br_136 wl_105 vdd gnd cell_6t
Xbit_r106_c136 bl_136 br_136 wl_106 vdd gnd cell_6t
Xbit_r107_c136 bl_136 br_136 wl_107 vdd gnd cell_6t
Xbit_r108_c136 bl_136 br_136 wl_108 vdd gnd cell_6t
Xbit_r109_c136 bl_136 br_136 wl_109 vdd gnd cell_6t
Xbit_r110_c136 bl_136 br_136 wl_110 vdd gnd cell_6t
Xbit_r111_c136 bl_136 br_136 wl_111 vdd gnd cell_6t
Xbit_r112_c136 bl_136 br_136 wl_112 vdd gnd cell_6t
Xbit_r113_c136 bl_136 br_136 wl_113 vdd gnd cell_6t
Xbit_r114_c136 bl_136 br_136 wl_114 vdd gnd cell_6t
Xbit_r115_c136 bl_136 br_136 wl_115 vdd gnd cell_6t
Xbit_r116_c136 bl_136 br_136 wl_116 vdd gnd cell_6t
Xbit_r117_c136 bl_136 br_136 wl_117 vdd gnd cell_6t
Xbit_r118_c136 bl_136 br_136 wl_118 vdd gnd cell_6t
Xbit_r119_c136 bl_136 br_136 wl_119 vdd gnd cell_6t
Xbit_r120_c136 bl_136 br_136 wl_120 vdd gnd cell_6t
Xbit_r121_c136 bl_136 br_136 wl_121 vdd gnd cell_6t
Xbit_r122_c136 bl_136 br_136 wl_122 vdd gnd cell_6t
Xbit_r123_c136 bl_136 br_136 wl_123 vdd gnd cell_6t
Xbit_r124_c136 bl_136 br_136 wl_124 vdd gnd cell_6t
Xbit_r125_c136 bl_136 br_136 wl_125 vdd gnd cell_6t
Xbit_r126_c136 bl_136 br_136 wl_126 vdd gnd cell_6t
Xbit_r127_c136 bl_136 br_136 wl_127 vdd gnd cell_6t
Xbit_r128_c136 bl_136 br_136 wl_128 vdd gnd cell_6t
Xbit_r129_c136 bl_136 br_136 wl_129 vdd gnd cell_6t
Xbit_r130_c136 bl_136 br_136 wl_130 vdd gnd cell_6t
Xbit_r131_c136 bl_136 br_136 wl_131 vdd gnd cell_6t
Xbit_r132_c136 bl_136 br_136 wl_132 vdd gnd cell_6t
Xbit_r133_c136 bl_136 br_136 wl_133 vdd gnd cell_6t
Xbit_r134_c136 bl_136 br_136 wl_134 vdd gnd cell_6t
Xbit_r135_c136 bl_136 br_136 wl_135 vdd gnd cell_6t
Xbit_r136_c136 bl_136 br_136 wl_136 vdd gnd cell_6t
Xbit_r137_c136 bl_136 br_136 wl_137 vdd gnd cell_6t
Xbit_r138_c136 bl_136 br_136 wl_138 vdd gnd cell_6t
Xbit_r139_c136 bl_136 br_136 wl_139 vdd gnd cell_6t
Xbit_r140_c136 bl_136 br_136 wl_140 vdd gnd cell_6t
Xbit_r141_c136 bl_136 br_136 wl_141 vdd gnd cell_6t
Xbit_r142_c136 bl_136 br_136 wl_142 vdd gnd cell_6t
Xbit_r143_c136 bl_136 br_136 wl_143 vdd gnd cell_6t
Xbit_r144_c136 bl_136 br_136 wl_144 vdd gnd cell_6t
Xbit_r145_c136 bl_136 br_136 wl_145 vdd gnd cell_6t
Xbit_r146_c136 bl_136 br_136 wl_146 vdd gnd cell_6t
Xbit_r147_c136 bl_136 br_136 wl_147 vdd gnd cell_6t
Xbit_r148_c136 bl_136 br_136 wl_148 vdd gnd cell_6t
Xbit_r149_c136 bl_136 br_136 wl_149 vdd gnd cell_6t
Xbit_r150_c136 bl_136 br_136 wl_150 vdd gnd cell_6t
Xbit_r151_c136 bl_136 br_136 wl_151 vdd gnd cell_6t
Xbit_r152_c136 bl_136 br_136 wl_152 vdd gnd cell_6t
Xbit_r153_c136 bl_136 br_136 wl_153 vdd gnd cell_6t
Xbit_r154_c136 bl_136 br_136 wl_154 vdd gnd cell_6t
Xbit_r155_c136 bl_136 br_136 wl_155 vdd gnd cell_6t
Xbit_r156_c136 bl_136 br_136 wl_156 vdd gnd cell_6t
Xbit_r157_c136 bl_136 br_136 wl_157 vdd gnd cell_6t
Xbit_r158_c136 bl_136 br_136 wl_158 vdd gnd cell_6t
Xbit_r159_c136 bl_136 br_136 wl_159 vdd gnd cell_6t
Xbit_r160_c136 bl_136 br_136 wl_160 vdd gnd cell_6t
Xbit_r161_c136 bl_136 br_136 wl_161 vdd gnd cell_6t
Xbit_r162_c136 bl_136 br_136 wl_162 vdd gnd cell_6t
Xbit_r163_c136 bl_136 br_136 wl_163 vdd gnd cell_6t
Xbit_r164_c136 bl_136 br_136 wl_164 vdd gnd cell_6t
Xbit_r165_c136 bl_136 br_136 wl_165 vdd gnd cell_6t
Xbit_r166_c136 bl_136 br_136 wl_166 vdd gnd cell_6t
Xbit_r167_c136 bl_136 br_136 wl_167 vdd gnd cell_6t
Xbit_r168_c136 bl_136 br_136 wl_168 vdd gnd cell_6t
Xbit_r169_c136 bl_136 br_136 wl_169 vdd gnd cell_6t
Xbit_r170_c136 bl_136 br_136 wl_170 vdd gnd cell_6t
Xbit_r171_c136 bl_136 br_136 wl_171 vdd gnd cell_6t
Xbit_r172_c136 bl_136 br_136 wl_172 vdd gnd cell_6t
Xbit_r173_c136 bl_136 br_136 wl_173 vdd gnd cell_6t
Xbit_r174_c136 bl_136 br_136 wl_174 vdd gnd cell_6t
Xbit_r175_c136 bl_136 br_136 wl_175 vdd gnd cell_6t
Xbit_r176_c136 bl_136 br_136 wl_176 vdd gnd cell_6t
Xbit_r177_c136 bl_136 br_136 wl_177 vdd gnd cell_6t
Xbit_r178_c136 bl_136 br_136 wl_178 vdd gnd cell_6t
Xbit_r179_c136 bl_136 br_136 wl_179 vdd gnd cell_6t
Xbit_r180_c136 bl_136 br_136 wl_180 vdd gnd cell_6t
Xbit_r181_c136 bl_136 br_136 wl_181 vdd gnd cell_6t
Xbit_r182_c136 bl_136 br_136 wl_182 vdd gnd cell_6t
Xbit_r183_c136 bl_136 br_136 wl_183 vdd gnd cell_6t
Xbit_r184_c136 bl_136 br_136 wl_184 vdd gnd cell_6t
Xbit_r185_c136 bl_136 br_136 wl_185 vdd gnd cell_6t
Xbit_r186_c136 bl_136 br_136 wl_186 vdd gnd cell_6t
Xbit_r187_c136 bl_136 br_136 wl_187 vdd gnd cell_6t
Xbit_r188_c136 bl_136 br_136 wl_188 vdd gnd cell_6t
Xbit_r189_c136 bl_136 br_136 wl_189 vdd gnd cell_6t
Xbit_r190_c136 bl_136 br_136 wl_190 vdd gnd cell_6t
Xbit_r191_c136 bl_136 br_136 wl_191 vdd gnd cell_6t
Xbit_r192_c136 bl_136 br_136 wl_192 vdd gnd cell_6t
Xbit_r193_c136 bl_136 br_136 wl_193 vdd gnd cell_6t
Xbit_r194_c136 bl_136 br_136 wl_194 vdd gnd cell_6t
Xbit_r195_c136 bl_136 br_136 wl_195 vdd gnd cell_6t
Xbit_r196_c136 bl_136 br_136 wl_196 vdd gnd cell_6t
Xbit_r197_c136 bl_136 br_136 wl_197 vdd gnd cell_6t
Xbit_r198_c136 bl_136 br_136 wl_198 vdd gnd cell_6t
Xbit_r199_c136 bl_136 br_136 wl_199 vdd gnd cell_6t
Xbit_r200_c136 bl_136 br_136 wl_200 vdd gnd cell_6t
Xbit_r201_c136 bl_136 br_136 wl_201 vdd gnd cell_6t
Xbit_r202_c136 bl_136 br_136 wl_202 vdd gnd cell_6t
Xbit_r203_c136 bl_136 br_136 wl_203 vdd gnd cell_6t
Xbit_r204_c136 bl_136 br_136 wl_204 vdd gnd cell_6t
Xbit_r205_c136 bl_136 br_136 wl_205 vdd gnd cell_6t
Xbit_r206_c136 bl_136 br_136 wl_206 vdd gnd cell_6t
Xbit_r207_c136 bl_136 br_136 wl_207 vdd gnd cell_6t
Xbit_r208_c136 bl_136 br_136 wl_208 vdd gnd cell_6t
Xbit_r209_c136 bl_136 br_136 wl_209 vdd gnd cell_6t
Xbit_r210_c136 bl_136 br_136 wl_210 vdd gnd cell_6t
Xbit_r211_c136 bl_136 br_136 wl_211 vdd gnd cell_6t
Xbit_r212_c136 bl_136 br_136 wl_212 vdd gnd cell_6t
Xbit_r213_c136 bl_136 br_136 wl_213 vdd gnd cell_6t
Xbit_r214_c136 bl_136 br_136 wl_214 vdd gnd cell_6t
Xbit_r215_c136 bl_136 br_136 wl_215 vdd gnd cell_6t
Xbit_r216_c136 bl_136 br_136 wl_216 vdd gnd cell_6t
Xbit_r217_c136 bl_136 br_136 wl_217 vdd gnd cell_6t
Xbit_r218_c136 bl_136 br_136 wl_218 vdd gnd cell_6t
Xbit_r219_c136 bl_136 br_136 wl_219 vdd gnd cell_6t
Xbit_r220_c136 bl_136 br_136 wl_220 vdd gnd cell_6t
Xbit_r221_c136 bl_136 br_136 wl_221 vdd gnd cell_6t
Xbit_r222_c136 bl_136 br_136 wl_222 vdd gnd cell_6t
Xbit_r223_c136 bl_136 br_136 wl_223 vdd gnd cell_6t
Xbit_r224_c136 bl_136 br_136 wl_224 vdd gnd cell_6t
Xbit_r225_c136 bl_136 br_136 wl_225 vdd gnd cell_6t
Xbit_r226_c136 bl_136 br_136 wl_226 vdd gnd cell_6t
Xbit_r227_c136 bl_136 br_136 wl_227 vdd gnd cell_6t
Xbit_r228_c136 bl_136 br_136 wl_228 vdd gnd cell_6t
Xbit_r229_c136 bl_136 br_136 wl_229 vdd gnd cell_6t
Xbit_r230_c136 bl_136 br_136 wl_230 vdd gnd cell_6t
Xbit_r231_c136 bl_136 br_136 wl_231 vdd gnd cell_6t
Xbit_r232_c136 bl_136 br_136 wl_232 vdd gnd cell_6t
Xbit_r233_c136 bl_136 br_136 wl_233 vdd gnd cell_6t
Xbit_r234_c136 bl_136 br_136 wl_234 vdd gnd cell_6t
Xbit_r235_c136 bl_136 br_136 wl_235 vdd gnd cell_6t
Xbit_r236_c136 bl_136 br_136 wl_236 vdd gnd cell_6t
Xbit_r237_c136 bl_136 br_136 wl_237 vdd gnd cell_6t
Xbit_r238_c136 bl_136 br_136 wl_238 vdd gnd cell_6t
Xbit_r239_c136 bl_136 br_136 wl_239 vdd gnd cell_6t
Xbit_r240_c136 bl_136 br_136 wl_240 vdd gnd cell_6t
Xbit_r241_c136 bl_136 br_136 wl_241 vdd gnd cell_6t
Xbit_r242_c136 bl_136 br_136 wl_242 vdd gnd cell_6t
Xbit_r243_c136 bl_136 br_136 wl_243 vdd gnd cell_6t
Xbit_r244_c136 bl_136 br_136 wl_244 vdd gnd cell_6t
Xbit_r245_c136 bl_136 br_136 wl_245 vdd gnd cell_6t
Xbit_r246_c136 bl_136 br_136 wl_246 vdd gnd cell_6t
Xbit_r247_c136 bl_136 br_136 wl_247 vdd gnd cell_6t
Xbit_r248_c136 bl_136 br_136 wl_248 vdd gnd cell_6t
Xbit_r249_c136 bl_136 br_136 wl_249 vdd gnd cell_6t
Xbit_r250_c136 bl_136 br_136 wl_250 vdd gnd cell_6t
Xbit_r251_c136 bl_136 br_136 wl_251 vdd gnd cell_6t
Xbit_r252_c136 bl_136 br_136 wl_252 vdd gnd cell_6t
Xbit_r253_c136 bl_136 br_136 wl_253 vdd gnd cell_6t
Xbit_r254_c136 bl_136 br_136 wl_254 vdd gnd cell_6t
Xbit_r255_c136 bl_136 br_136 wl_255 vdd gnd cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd cell_6t
Xbit_r1_c137 bl_137 br_137 wl_1 vdd gnd cell_6t
Xbit_r2_c137 bl_137 br_137 wl_2 vdd gnd cell_6t
Xbit_r3_c137 bl_137 br_137 wl_3 vdd gnd cell_6t
Xbit_r4_c137 bl_137 br_137 wl_4 vdd gnd cell_6t
Xbit_r5_c137 bl_137 br_137 wl_5 vdd gnd cell_6t
Xbit_r6_c137 bl_137 br_137 wl_6 vdd gnd cell_6t
Xbit_r7_c137 bl_137 br_137 wl_7 vdd gnd cell_6t
Xbit_r8_c137 bl_137 br_137 wl_8 vdd gnd cell_6t
Xbit_r9_c137 bl_137 br_137 wl_9 vdd gnd cell_6t
Xbit_r10_c137 bl_137 br_137 wl_10 vdd gnd cell_6t
Xbit_r11_c137 bl_137 br_137 wl_11 vdd gnd cell_6t
Xbit_r12_c137 bl_137 br_137 wl_12 vdd gnd cell_6t
Xbit_r13_c137 bl_137 br_137 wl_13 vdd gnd cell_6t
Xbit_r14_c137 bl_137 br_137 wl_14 vdd gnd cell_6t
Xbit_r15_c137 bl_137 br_137 wl_15 vdd gnd cell_6t
Xbit_r16_c137 bl_137 br_137 wl_16 vdd gnd cell_6t
Xbit_r17_c137 bl_137 br_137 wl_17 vdd gnd cell_6t
Xbit_r18_c137 bl_137 br_137 wl_18 vdd gnd cell_6t
Xbit_r19_c137 bl_137 br_137 wl_19 vdd gnd cell_6t
Xbit_r20_c137 bl_137 br_137 wl_20 vdd gnd cell_6t
Xbit_r21_c137 bl_137 br_137 wl_21 vdd gnd cell_6t
Xbit_r22_c137 bl_137 br_137 wl_22 vdd gnd cell_6t
Xbit_r23_c137 bl_137 br_137 wl_23 vdd gnd cell_6t
Xbit_r24_c137 bl_137 br_137 wl_24 vdd gnd cell_6t
Xbit_r25_c137 bl_137 br_137 wl_25 vdd gnd cell_6t
Xbit_r26_c137 bl_137 br_137 wl_26 vdd gnd cell_6t
Xbit_r27_c137 bl_137 br_137 wl_27 vdd gnd cell_6t
Xbit_r28_c137 bl_137 br_137 wl_28 vdd gnd cell_6t
Xbit_r29_c137 bl_137 br_137 wl_29 vdd gnd cell_6t
Xbit_r30_c137 bl_137 br_137 wl_30 vdd gnd cell_6t
Xbit_r31_c137 bl_137 br_137 wl_31 vdd gnd cell_6t
Xbit_r32_c137 bl_137 br_137 wl_32 vdd gnd cell_6t
Xbit_r33_c137 bl_137 br_137 wl_33 vdd gnd cell_6t
Xbit_r34_c137 bl_137 br_137 wl_34 vdd gnd cell_6t
Xbit_r35_c137 bl_137 br_137 wl_35 vdd gnd cell_6t
Xbit_r36_c137 bl_137 br_137 wl_36 vdd gnd cell_6t
Xbit_r37_c137 bl_137 br_137 wl_37 vdd gnd cell_6t
Xbit_r38_c137 bl_137 br_137 wl_38 vdd gnd cell_6t
Xbit_r39_c137 bl_137 br_137 wl_39 vdd gnd cell_6t
Xbit_r40_c137 bl_137 br_137 wl_40 vdd gnd cell_6t
Xbit_r41_c137 bl_137 br_137 wl_41 vdd gnd cell_6t
Xbit_r42_c137 bl_137 br_137 wl_42 vdd gnd cell_6t
Xbit_r43_c137 bl_137 br_137 wl_43 vdd gnd cell_6t
Xbit_r44_c137 bl_137 br_137 wl_44 vdd gnd cell_6t
Xbit_r45_c137 bl_137 br_137 wl_45 vdd gnd cell_6t
Xbit_r46_c137 bl_137 br_137 wl_46 vdd gnd cell_6t
Xbit_r47_c137 bl_137 br_137 wl_47 vdd gnd cell_6t
Xbit_r48_c137 bl_137 br_137 wl_48 vdd gnd cell_6t
Xbit_r49_c137 bl_137 br_137 wl_49 vdd gnd cell_6t
Xbit_r50_c137 bl_137 br_137 wl_50 vdd gnd cell_6t
Xbit_r51_c137 bl_137 br_137 wl_51 vdd gnd cell_6t
Xbit_r52_c137 bl_137 br_137 wl_52 vdd gnd cell_6t
Xbit_r53_c137 bl_137 br_137 wl_53 vdd gnd cell_6t
Xbit_r54_c137 bl_137 br_137 wl_54 vdd gnd cell_6t
Xbit_r55_c137 bl_137 br_137 wl_55 vdd gnd cell_6t
Xbit_r56_c137 bl_137 br_137 wl_56 vdd gnd cell_6t
Xbit_r57_c137 bl_137 br_137 wl_57 vdd gnd cell_6t
Xbit_r58_c137 bl_137 br_137 wl_58 vdd gnd cell_6t
Xbit_r59_c137 bl_137 br_137 wl_59 vdd gnd cell_6t
Xbit_r60_c137 bl_137 br_137 wl_60 vdd gnd cell_6t
Xbit_r61_c137 bl_137 br_137 wl_61 vdd gnd cell_6t
Xbit_r62_c137 bl_137 br_137 wl_62 vdd gnd cell_6t
Xbit_r63_c137 bl_137 br_137 wl_63 vdd gnd cell_6t
Xbit_r64_c137 bl_137 br_137 wl_64 vdd gnd cell_6t
Xbit_r65_c137 bl_137 br_137 wl_65 vdd gnd cell_6t
Xbit_r66_c137 bl_137 br_137 wl_66 vdd gnd cell_6t
Xbit_r67_c137 bl_137 br_137 wl_67 vdd gnd cell_6t
Xbit_r68_c137 bl_137 br_137 wl_68 vdd gnd cell_6t
Xbit_r69_c137 bl_137 br_137 wl_69 vdd gnd cell_6t
Xbit_r70_c137 bl_137 br_137 wl_70 vdd gnd cell_6t
Xbit_r71_c137 bl_137 br_137 wl_71 vdd gnd cell_6t
Xbit_r72_c137 bl_137 br_137 wl_72 vdd gnd cell_6t
Xbit_r73_c137 bl_137 br_137 wl_73 vdd gnd cell_6t
Xbit_r74_c137 bl_137 br_137 wl_74 vdd gnd cell_6t
Xbit_r75_c137 bl_137 br_137 wl_75 vdd gnd cell_6t
Xbit_r76_c137 bl_137 br_137 wl_76 vdd gnd cell_6t
Xbit_r77_c137 bl_137 br_137 wl_77 vdd gnd cell_6t
Xbit_r78_c137 bl_137 br_137 wl_78 vdd gnd cell_6t
Xbit_r79_c137 bl_137 br_137 wl_79 vdd gnd cell_6t
Xbit_r80_c137 bl_137 br_137 wl_80 vdd gnd cell_6t
Xbit_r81_c137 bl_137 br_137 wl_81 vdd gnd cell_6t
Xbit_r82_c137 bl_137 br_137 wl_82 vdd gnd cell_6t
Xbit_r83_c137 bl_137 br_137 wl_83 vdd gnd cell_6t
Xbit_r84_c137 bl_137 br_137 wl_84 vdd gnd cell_6t
Xbit_r85_c137 bl_137 br_137 wl_85 vdd gnd cell_6t
Xbit_r86_c137 bl_137 br_137 wl_86 vdd gnd cell_6t
Xbit_r87_c137 bl_137 br_137 wl_87 vdd gnd cell_6t
Xbit_r88_c137 bl_137 br_137 wl_88 vdd gnd cell_6t
Xbit_r89_c137 bl_137 br_137 wl_89 vdd gnd cell_6t
Xbit_r90_c137 bl_137 br_137 wl_90 vdd gnd cell_6t
Xbit_r91_c137 bl_137 br_137 wl_91 vdd gnd cell_6t
Xbit_r92_c137 bl_137 br_137 wl_92 vdd gnd cell_6t
Xbit_r93_c137 bl_137 br_137 wl_93 vdd gnd cell_6t
Xbit_r94_c137 bl_137 br_137 wl_94 vdd gnd cell_6t
Xbit_r95_c137 bl_137 br_137 wl_95 vdd gnd cell_6t
Xbit_r96_c137 bl_137 br_137 wl_96 vdd gnd cell_6t
Xbit_r97_c137 bl_137 br_137 wl_97 vdd gnd cell_6t
Xbit_r98_c137 bl_137 br_137 wl_98 vdd gnd cell_6t
Xbit_r99_c137 bl_137 br_137 wl_99 vdd gnd cell_6t
Xbit_r100_c137 bl_137 br_137 wl_100 vdd gnd cell_6t
Xbit_r101_c137 bl_137 br_137 wl_101 vdd gnd cell_6t
Xbit_r102_c137 bl_137 br_137 wl_102 vdd gnd cell_6t
Xbit_r103_c137 bl_137 br_137 wl_103 vdd gnd cell_6t
Xbit_r104_c137 bl_137 br_137 wl_104 vdd gnd cell_6t
Xbit_r105_c137 bl_137 br_137 wl_105 vdd gnd cell_6t
Xbit_r106_c137 bl_137 br_137 wl_106 vdd gnd cell_6t
Xbit_r107_c137 bl_137 br_137 wl_107 vdd gnd cell_6t
Xbit_r108_c137 bl_137 br_137 wl_108 vdd gnd cell_6t
Xbit_r109_c137 bl_137 br_137 wl_109 vdd gnd cell_6t
Xbit_r110_c137 bl_137 br_137 wl_110 vdd gnd cell_6t
Xbit_r111_c137 bl_137 br_137 wl_111 vdd gnd cell_6t
Xbit_r112_c137 bl_137 br_137 wl_112 vdd gnd cell_6t
Xbit_r113_c137 bl_137 br_137 wl_113 vdd gnd cell_6t
Xbit_r114_c137 bl_137 br_137 wl_114 vdd gnd cell_6t
Xbit_r115_c137 bl_137 br_137 wl_115 vdd gnd cell_6t
Xbit_r116_c137 bl_137 br_137 wl_116 vdd gnd cell_6t
Xbit_r117_c137 bl_137 br_137 wl_117 vdd gnd cell_6t
Xbit_r118_c137 bl_137 br_137 wl_118 vdd gnd cell_6t
Xbit_r119_c137 bl_137 br_137 wl_119 vdd gnd cell_6t
Xbit_r120_c137 bl_137 br_137 wl_120 vdd gnd cell_6t
Xbit_r121_c137 bl_137 br_137 wl_121 vdd gnd cell_6t
Xbit_r122_c137 bl_137 br_137 wl_122 vdd gnd cell_6t
Xbit_r123_c137 bl_137 br_137 wl_123 vdd gnd cell_6t
Xbit_r124_c137 bl_137 br_137 wl_124 vdd gnd cell_6t
Xbit_r125_c137 bl_137 br_137 wl_125 vdd gnd cell_6t
Xbit_r126_c137 bl_137 br_137 wl_126 vdd gnd cell_6t
Xbit_r127_c137 bl_137 br_137 wl_127 vdd gnd cell_6t
Xbit_r128_c137 bl_137 br_137 wl_128 vdd gnd cell_6t
Xbit_r129_c137 bl_137 br_137 wl_129 vdd gnd cell_6t
Xbit_r130_c137 bl_137 br_137 wl_130 vdd gnd cell_6t
Xbit_r131_c137 bl_137 br_137 wl_131 vdd gnd cell_6t
Xbit_r132_c137 bl_137 br_137 wl_132 vdd gnd cell_6t
Xbit_r133_c137 bl_137 br_137 wl_133 vdd gnd cell_6t
Xbit_r134_c137 bl_137 br_137 wl_134 vdd gnd cell_6t
Xbit_r135_c137 bl_137 br_137 wl_135 vdd gnd cell_6t
Xbit_r136_c137 bl_137 br_137 wl_136 vdd gnd cell_6t
Xbit_r137_c137 bl_137 br_137 wl_137 vdd gnd cell_6t
Xbit_r138_c137 bl_137 br_137 wl_138 vdd gnd cell_6t
Xbit_r139_c137 bl_137 br_137 wl_139 vdd gnd cell_6t
Xbit_r140_c137 bl_137 br_137 wl_140 vdd gnd cell_6t
Xbit_r141_c137 bl_137 br_137 wl_141 vdd gnd cell_6t
Xbit_r142_c137 bl_137 br_137 wl_142 vdd gnd cell_6t
Xbit_r143_c137 bl_137 br_137 wl_143 vdd gnd cell_6t
Xbit_r144_c137 bl_137 br_137 wl_144 vdd gnd cell_6t
Xbit_r145_c137 bl_137 br_137 wl_145 vdd gnd cell_6t
Xbit_r146_c137 bl_137 br_137 wl_146 vdd gnd cell_6t
Xbit_r147_c137 bl_137 br_137 wl_147 vdd gnd cell_6t
Xbit_r148_c137 bl_137 br_137 wl_148 vdd gnd cell_6t
Xbit_r149_c137 bl_137 br_137 wl_149 vdd gnd cell_6t
Xbit_r150_c137 bl_137 br_137 wl_150 vdd gnd cell_6t
Xbit_r151_c137 bl_137 br_137 wl_151 vdd gnd cell_6t
Xbit_r152_c137 bl_137 br_137 wl_152 vdd gnd cell_6t
Xbit_r153_c137 bl_137 br_137 wl_153 vdd gnd cell_6t
Xbit_r154_c137 bl_137 br_137 wl_154 vdd gnd cell_6t
Xbit_r155_c137 bl_137 br_137 wl_155 vdd gnd cell_6t
Xbit_r156_c137 bl_137 br_137 wl_156 vdd gnd cell_6t
Xbit_r157_c137 bl_137 br_137 wl_157 vdd gnd cell_6t
Xbit_r158_c137 bl_137 br_137 wl_158 vdd gnd cell_6t
Xbit_r159_c137 bl_137 br_137 wl_159 vdd gnd cell_6t
Xbit_r160_c137 bl_137 br_137 wl_160 vdd gnd cell_6t
Xbit_r161_c137 bl_137 br_137 wl_161 vdd gnd cell_6t
Xbit_r162_c137 bl_137 br_137 wl_162 vdd gnd cell_6t
Xbit_r163_c137 bl_137 br_137 wl_163 vdd gnd cell_6t
Xbit_r164_c137 bl_137 br_137 wl_164 vdd gnd cell_6t
Xbit_r165_c137 bl_137 br_137 wl_165 vdd gnd cell_6t
Xbit_r166_c137 bl_137 br_137 wl_166 vdd gnd cell_6t
Xbit_r167_c137 bl_137 br_137 wl_167 vdd gnd cell_6t
Xbit_r168_c137 bl_137 br_137 wl_168 vdd gnd cell_6t
Xbit_r169_c137 bl_137 br_137 wl_169 vdd gnd cell_6t
Xbit_r170_c137 bl_137 br_137 wl_170 vdd gnd cell_6t
Xbit_r171_c137 bl_137 br_137 wl_171 vdd gnd cell_6t
Xbit_r172_c137 bl_137 br_137 wl_172 vdd gnd cell_6t
Xbit_r173_c137 bl_137 br_137 wl_173 vdd gnd cell_6t
Xbit_r174_c137 bl_137 br_137 wl_174 vdd gnd cell_6t
Xbit_r175_c137 bl_137 br_137 wl_175 vdd gnd cell_6t
Xbit_r176_c137 bl_137 br_137 wl_176 vdd gnd cell_6t
Xbit_r177_c137 bl_137 br_137 wl_177 vdd gnd cell_6t
Xbit_r178_c137 bl_137 br_137 wl_178 vdd gnd cell_6t
Xbit_r179_c137 bl_137 br_137 wl_179 vdd gnd cell_6t
Xbit_r180_c137 bl_137 br_137 wl_180 vdd gnd cell_6t
Xbit_r181_c137 bl_137 br_137 wl_181 vdd gnd cell_6t
Xbit_r182_c137 bl_137 br_137 wl_182 vdd gnd cell_6t
Xbit_r183_c137 bl_137 br_137 wl_183 vdd gnd cell_6t
Xbit_r184_c137 bl_137 br_137 wl_184 vdd gnd cell_6t
Xbit_r185_c137 bl_137 br_137 wl_185 vdd gnd cell_6t
Xbit_r186_c137 bl_137 br_137 wl_186 vdd gnd cell_6t
Xbit_r187_c137 bl_137 br_137 wl_187 vdd gnd cell_6t
Xbit_r188_c137 bl_137 br_137 wl_188 vdd gnd cell_6t
Xbit_r189_c137 bl_137 br_137 wl_189 vdd gnd cell_6t
Xbit_r190_c137 bl_137 br_137 wl_190 vdd gnd cell_6t
Xbit_r191_c137 bl_137 br_137 wl_191 vdd gnd cell_6t
Xbit_r192_c137 bl_137 br_137 wl_192 vdd gnd cell_6t
Xbit_r193_c137 bl_137 br_137 wl_193 vdd gnd cell_6t
Xbit_r194_c137 bl_137 br_137 wl_194 vdd gnd cell_6t
Xbit_r195_c137 bl_137 br_137 wl_195 vdd gnd cell_6t
Xbit_r196_c137 bl_137 br_137 wl_196 vdd gnd cell_6t
Xbit_r197_c137 bl_137 br_137 wl_197 vdd gnd cell_6t
Xbit_r198_c137 bl_137 br_137 wl_198 vdd gnd cell_6t
Xbit_r199_c137 bl_137 br_137 wl_199 vdd gnd cell_6t
Xbit_r200_c137 bl_137 br_137 wl_200 vdd gnd cell_6t
Xbit_r201_c137 bl_137 br_137 wl_201 vdd gnd cell_6t
Xbit_r202_c137 bl_137 br_137 wl_202 vdd gnd cell_6t
Xbit_r203_c137 bl_137 br_137 wl_203 vdd gnd cell_6t
Xbit_r204_c137 bl_137 br_137 wl_204 vdd gnd cell_6t
Xbit_r205_c137 bl_137 br_137 wl_205 vdd gnd cell_6t
Xbit_r206_c137 bl_137 br_137 wl_206 vdd gnd cell_6t
Xbit_r207_c137 bl_137 br_137 wl_207 vdd gnd cell_6t
Xbit_r208_c137 bl_137 br_137 wl_208 vdd gnd cell_6t
Xbit_r209_c137 bl_137 br_137 wl_209 vdd gnd cell_6t
Xbit_r210_c137 bl_137 br_137 wl_210 vdd gnd cell_6t
Xbit_r211_c137 bl_137 br_137 wl_211 vdd gnd cell_6t
Xbit_r212_c137 bl_137 br_137 wl_212 vdd gnd cell_6t
Xbit_r213_c137 bl_137 br_137 wl_213 vdd gnd cell_6t
Xbit_r214_c137 bl_137 br_137 wl_214 vdd gnd cell_6t
Xbit_r215_c137 bl_137 br_137 wl_215 vdd gnd cell_6t
Xbit_r216_c137 bl_137 br_137 wl_216 vdd gnd cell_6t
Xbit_r217_c137 bl_137 br_137 wl_217 vdd gnd cell_6t
Xbit_r218_c137 bl_137 br_137 wl_218 vdd gnd cell_6t
Xbit_r219_c137 bl_137 br_137 wl_219 vdd gnd cell_6t
Xbit_r220_c137 bl_137 br_137 wl_220 vdd gnd cell_6t
Xbit_r221_c137 bl_137 br_137 wl_221 vdd gnd cell_6t
Xbit_r222_c137 bl_137 br_137 wl_222 vdd gnd cell_6t
Xbit_r223_c137 bl_137 br_137 wl_223 vdd gnd cell_6t
Xbit_r224_c137 bl_137 br_137 wl_224 vdd gnd cell_6t
Xbit_r225_c137 bl_137 br_137 wl_225 vdd gnd cell_6t
Xbit_r226_c137 bl_137 br_137 wl_226 vdd gnd cell_6t
Xbit_r227_c137 bl_137 br_137 wl_227 vdd gnd cell_6t
Xbit_r228_c137 bl_137 br_137 wl_228 vdd gnd cell_6t
Xbit_r229_c137 bl_137 br_137 wl_229 vdd gnd cell_6t
Xbit_r230_c137 bl_137 br_137 wl_230 vdd gnd cell_6t
Xbit_r231_c137 bl_137 br_137 wl_231 vdd gnd cell_6t
Xbit_r232_c137 bl_137 br_137 wl_232 vdd gnd cell_6t
Xbit_r233_c137 bl_137 br_137 wl_233 vdd gnd cell_6t
Xbit_r234_c137 bl_137 br_137 wl_234 vdd gnd cell_6t
Xbit_r235_c137 bl_137 br_137 wl_235 vdd gnd cell_6t
Xbit_r236_c137 bl_137 br_137 wl_236 vdd gnd cell_6t
Xbit_r237_c137 bl_137 br_137 wl_237 vdd gnd cell_6t
Xbit_r238_c137 bl_137 br_137 wl_238 vdd gnd cell_6t
Xbit_r239_c137 bl_137 br_137 wl_239 vdd gnd cell_6t
Xbit_r240_c137 bl_137 br_137 wl_240 vdd gnd cell_6t
Xbit_r241_c137 bl_137 br_137 wl_241 vdd gnd cell_6t
Xbit_r242_c137 bl_137 br_137 wl_242 vdd gnd cell_6t
Xbit_r243_c137 bl_137 br_137 wl_243 vdd gnd cell_6t
Xbit_r244_c137 bl_137 br_137 wl_244 vdd gnd cell_6t
Xbit_r245_c137 bl_137 br_137 wl_245 vdd gnd cell_6t
Xbit_r246_c137 bl_137 br_137 wl_246 vdd gnd cell_6t
Xbit_r247_c137 bl_137 br_137 wl_247 vdd gnd cell_6t
Xbit_r248_c137 bl_137 br_137 wl_248 vdd gnd cell_6t
Xbit_r249_c137 bl_137 br_137 wl_249 vdd gnd cell_6t
Xbit_r250_c137 bl_137 br_137 wl_250 vdd gnd cell_6t
Xbit_r251_c137 bl_137 br_137 wl_251 vdd gnd cell_6t
Xbit_r252_c137 bl_137 br_137 wl_252 vdd gnd cell_6t
Xbit_r253_c137 bl_137 br_137 wl_253 vdd gnd cell_6t
Xbit_r254_c137 bl_137 br_137 wl_254 vdd gnd cell_6t
Xbit_r255_c137 bl_137 br_137 wl_255 vdd gnd cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd cell_6t
Xbit_r1_c138 bl_138 br_138 wl_1 vdd gnd cell_6t
Xbit_r2_c138 bl_138 br_138 wl_2 vdd gnd cell_6t
Xbit_r3_c138 bl_138 br_138 wl_3 vdd gnd cell_6t
Xbit_r4_c138 bl_138 br_138 wl_4 vdd gnd cell_6t
Xbit_r5_c138 bl_138 br_138 wl_5 vdd gnd cell_6t
Xbit_r6_c138 bl_138 br_138 wl_6 vdd gnd cell_6t
Xbit_r7_c138 bl_138 br_138 wl_7 vdd gnd cell_6t
Xbit_r8_c138 bl_138 br_138 wl_8 vdd gnd cell_6t
Xbit_r9_c138 bl_138 br_138 wl_9 vdd gnd cell_6t
Xbit_r10_c138 bl_138 br_138 wl_10 vdd gnd cell_6t
Xbit_r11_c138 bl_138 br_138 wl_11 vdd gnd cell_6t
Xbit_r12_c138 bl_138 br_138 wl_12 vdd gnd cell_6t
Xbit_r13_c138 bl_138 br_138 wl_13 vdd gnd cell_6t
Xbit_r14_c138 bl_138 br_138 wl_14 vdd gnd cell_6t
Xbit_r15_c138 bl_138 br_138 wl_15 vdd gnd cell_6t
Xbit_r16_c138 bl_138 br_138 wl_16 vdd gnd cell_6t
Xbit_r17_c138 bl_138 br_138 wl_17 vdd gnd cell_6t
Xbit_r18_c138 bl_138 br_138 wl_18 vdd gnd cell_6t
Xbit_r19_c138 bl_138 br_138 wl_19 vdd gnd cell_6t
Xbit_r20_c138 bl_138 br_138 wl_20 vdd gnd cell_6t
Xbit_r21_c138 bl_138 br_138 wl_21 vdd gnd cell_6t
Xbit_r22_c138 bl_138 br_138 wl_22 vdd gnd cell_6t
Xbit_r23_c138 bl_138 br_138 wl_23 vdd gnd cell_6t
Xbit_r24_c138 bl_138 br_138 wl_24 vdd gnd cell_6t
Xbit_r25_c138 bl_138 br_138 wl_25 vdd gnd cell_6t
Xbit_r26_c138 bl_138 br_138 wl_26 vdd gnd cell_6t
Xbit_r27_c138 bl_138 br_138 wl_27 vdd gnd cell_6t
Xbit_r28_c138 bl_138 br_138 wl_28 vdd gnd cell_6t
Xbit_r29_c138 bl_138 br_138 wl_29 vdd gnd cell_6t
Xbit_r30_c138 bl_138 br_138 wl_30 vdd gnd cell_6t
Xbit_r31_c138 bl_138 br_138 wl_31 vdd gnd cell_6t
Xbit_r32_c138 bl_138 br_138 wl_32 vdd gnd cell_6t
Xbit_r33_c138 bl_138 br_138 wl_33 vdd gnd cell_6t
Xbit_r34_c138 bl_138 br_138 wl_34 vdd gnd cell_6t
Xbit_r35_c138 bl_138 br_138 wl_35 vdd gnd cell_6t
Xbit_r36_c138 bl_138 br_138 wl_36 vdd gnd cell_6t
Xbit_r37_c138 bl_138 br_138 wl_37 vdd gnd cell_6t
Xbit_r38_c138 bl_138 br_138 wl_38 vdd gnd cell_6t
Xbit_r39_c138 bl_138 br_138 wl_39 vdd gnd cell_6t
Xbit_r40_c138 bl_138 br_138 wl_40 vdd gnd cell_6t
Xbit_r41_c138 bl_138 br_138 wl_41 vdd gnd cell_6t
Xbit_r42_c138 bl_138 br_138 wl_42 vdd gnd cell_6t
Xbit_r43_c138 bl_138 br_138 wl_43 vdd gnd cell_6t
Xbit_r44_c138 bl_138 br_138 wl_44 vdd gnd cell_6t
Xbit_r45_c138 bl_138 br_138 wl_45 vdd gnd cell_6t
Xbit_r46_c138 bl_138 br_138 wl_46 vdd gnd cell_6t
Xbit_r47_c138 bl_138 br_138 wl_47 vdd gnd cell_6t
Xbit_r48_c138 bl_138 br_138 wl_48 vdd gnd cell_6t
Xbit_r49_c138 bl_138 br_138 wl_49 vdd gnd cell_6t
Xbit_r50_c138 bl_138 br_138 wl_50 vdd gnd cell_6t
Xbit_r51_c138 bl_138 br_138 wl_51 vdd gnd cell_6t
Xbit_r52_c138 bl_138 br_138 wl_52 vdd gnd cell_6t
Xbit_r53_c138 bl_138 br_138 wl_53 vdd gnd cell_6t
Xbit_r54_c138 bl_138 br_138 wl_54 vdd gnd cell_6t
Xbit_r55_c138 bl_138 br_138 wl_55 vdd gnd cell_6t
Xbit_r56_c138 bl_138 br_138 wl_56 vdd gnd cell_6t
Xbit_r57_c138 bl_138 br_138 wl_57 vdd gnd cell_6t
Xbit_r58_c138 bl_138 br_138 wl_58 vdd gnd cell_6t
Xbit_r59_c138 bl_138 br_138 wl_59 vdd gnd cell_6t
Xbit_r60_c138 bl_138 br_138 wl_60 vdd gnd cell_6t
Xbit_r61_c138 bl_138 br_138 wl_61 vdd gnd cell_6t
Xbit_r62_c138 bl_138 br_138 wl_62 vdd gnd cell_6t
Xbit_r63_c138 bl_138 br_138 wl_63 vdd gnd cell_6t
Xbit_r64_c138 bl_138 br_138 wl_64 vdd gnd cell_6t
Xbit_r65_c138 bl_138 br_138 wl_65 vdd gnd cell_6t
Xbit_r66_c138 bl_138 br_138 wl_66 vdd gnd cell_6t
Xbit_r67_c138 bl_138 br_138 wl_67 vdd gnd cell_6t
Xbit_r68_c138 bl_138 br_138 wl_68 vdd gnd cell_6t
Xbit_r69_c138 bl_138 br_138 wl_69 vdd gnd cell_6t
Xbit_r70_c138 bl_138 br_138 wl_70 vdd gnd cell_6t
Xbit_r71_c138 bl_138 br_138 wl_71 vdd gnd cell_6t
Xbit_r72_c138 bl_138 br_138 wl_72 vdd gnd cell_6t
Xbit_r73_c138 bl_138 br_138 wl_73 vdd gnd cell_6t
Xbit_r74_c138 bl_138 br_138 wl_74 vdd gnd cell_6t
Xbit_r75_c138 bl_138 br_138 wl_75 vdd gnd cell_6t
Xbit_r76_c138 bl_138 br_138 wl_76 vdd gnd cell_6t
Xbit_r77_c138 bl_138 br_138 wl_77 vdd gnd cell_6t
Xbit_r78_c138 bl_138 br_138 wl_78 vdd gnd cell_6t
Xbit_r79_c138 bl_138 br_138 wl_79 vdd gnd cell_6t
Xbit_r80_c138 bl_138 br_138 wl_80 vdd gnd cell_6t
Xbit_r81_c138 bl_138 br_138 wl_81 vdd gnd cell_6t
Xbit_r82_c138 bl_138 br_138 wl_82 vdd gnd cell_6t
Xbit_r83_c138 bl_138 br_138 wl_83 vdd gnd cell_6t
Xbit_r84_c138 bl_138 br_138 wl_84 vdd gnd cell_6t
Xbit_r85_c138 bl_138 br_138 wl_85 vdd gnd cell_6t
Xbit_r86_c138 bl_138 br_138 wl_86 vdd gnd cell_6t
Xbit_r87_c138 bl_138 br_138 wl_87 vdd gnd cell_6t
Xbit_r88_c138 bl_138 br_138 wl_88 vdd gnd cell_6t
Xbit_r89_c138 bl_138 br_138 wl_89 vdd gnd cell_6t
Xbit_r90_c138 bl_138 br_138 wl_90 vdd gnd cell_6t
Xbit_r91_c138 bl_138 br_138 wl_91 vdd gnd cell_6t
Xbit_r92_c138 bl_138 br_138 wl_92 vdd gnd cell_6t
Xbit_r93_c138 bl_138 br_138 wl_93 vdd gnd cell_6t
Xbit_r94_c138 bl_138 br_138 wl_94 vdd gnd cell_6t
Xbit_r95_c138 bl_138 br_138 wl_95 vdd gnd cell_6t
Xbit_r96_c138 bl_138 br_138 wl_96 vdd gnd cell_6t
Xbit_r97_c138 bl_138 br_138 wl_97 vdd gnd cell_6t
Xbit_r98_c138 bl_138 br_138 wl_98 vdd gnd cell_6t
Xbit_r99_c138 bl_138 br_138 wl_99 vdd gnd cell_6t
Xbit_r100_c138 bl_138 br_138 wl_100 vdd gnd cell_6t
Xbit_r101_c138 bl_138 br_138 wl_101 vdd gnd cell_6t
Xbit_r102_c138 bl_138 br_138 wl_102 vdd gnd cell_6t
Xbit_r103_c138 bl_138 br_138 wl_103 vdd gnd cell_6t
Xbit_r104_c138 bl_138 br_138 wl_104 vdd gnd cell_6t
Xbit_r105_c138 bl_138 br_138 wl_105 vdd gnd cell_6t
Xbit_r106_c138 bl_138 br_138 wl_106 vdd gnd cell_6t
Xbit_r107_c138 bl_138 br_138 wl_107 vdd gnd cell_6t
Xbit_r108_c138 bl_138 br_138 wl_108 vdd gnd cell_6t
Xbit_r109_c138 bl_138 br_138 wl_109 vdd gnd cell_6t
Xbit_r110_c138 bl_138 br_138 wl_110 vdd gnd cell_6t
Xbit_r111_c138 bl_138 br_138 wl_111 vdd gnd cell_6t
Xbit_r112_c138 bl_138 br_138 wl_112 vdd gnd cell_6t
Xbit_r113_c138 bl_138 br_138 wl_113 vdd gnd cell_6t
Xbit_r114_c138 bl_138 br_138 wl_114 vdd gnd cell_6t
Xbit_r115_c138 bl_138 br_138 wl_115 vdd gnd cell_6t
Xbit_r116_c138 bl_138 br_138 wl_116 vdd gnd cell_6t
Xbit_r117_c138 bl_138 br_138 wl_117 vdd gnd cell_6t
Xbit_r118_c138 bl_138 br_138 wl_118 vdd gnd cell_6t
Xbit_r119_c138 bl_138 br_138 wl_119 vdd gnd cell_6t
Xbit_r120_c138 bl_138 br_138 wl_120 vdd gnd cell_6t
Xbit_r121_c138 bl_138 br_138 wl_121 vdd gnd cell_6t
Xbit_r122_c138 bl_138 br_138 wl_122 vdd gnd cell_6t
Xbit_r123_c138 bl_138 br_138 wl_123 vdd gnd cell_6t
Xbit_r124_c138 bl_138 br_138 wl_124 vdd gnd cell_6t
Xbit_r125_c138 bl_138 br_138 wl_125 vdd gnd cell_6t
Xbit_r126_c138 bl_138 br_138 wl_126 vdd gnd cell_6t
Xbit_r127_c138 bl_138 br_138 wl_127 vdd gnd cell_6t
Xbit_r128_c138 bl_138 br_138 wl_128 vdd gnd cell_6t
Xbit_r129_c138 bl_138 br_138 wl_129 vdd gnd cell_6t
Xbit_r130_c138 bl_138 br_138 wl_130 vdd gnd cell_6t
Xbit_r131_c138 bl_138 br_138 wl_131 vdd gnd cell_6t
Xbit_r132_c138 bl_138 br_138 wl_132 vdd gnd cell_6t
Xbit_r133_c138 bl_138 br_138 wl_133 vdd gnd cell_6t
Xbit_r134_c138 bl_138 br_138 wl_134 vdd gnd cell_6t
Xbit_r135_c138 bl_138 br_138 wl_135 vdd gnd cell_6t
Xbit_r136_c138 bl_138 br_138 wl_136 vdd gnd cell_6t
Xbit_r137_c138 bl_138 br_138 wl_137 vdd gnd cell_6t
Xbit_r138_c138 bl_138 br_138 wl_138 vdd gnd cell_6t
Xbit_r139_c138 bl_138 br_138 wl_139 vdd gnd cell_6t
Xbit_r140_c138 bl_138 br_138 wl_140 vdd gnd cell_6t
Xbit_r141_c138 bl_138 br_138 wl_141 vdd gnd cell_6t
Xbit_r142_c138 bl_138 br_138 wl_142 vdd gnd cell_6t
Xbit_r143_c138 bl_138 br_138 wl_143 vdd gnd cell_6t
Xbit_r144_c138 bl_138 br_138 wl_144 vdd gnd cell_6t
Xbit_r145_c138 bl_138 br_138 wl_145 vdd gnd cell_6t
Xbit_r146_c138 bl_138 br_138 wl_146 vdd gnd cell_6t
Xbit_r147_c138 bl_138 br_138 wl_147 vdd gnd cell_6t
Xbit_r148_c138 bl_138 br_138 wl_148 vdd gnd cell_6t
Xbit_r149_c138 bl_138 br_138 wl_149 vdd gnd cell_6t
Xbit_r150_c138 bl_138 br_138 wl_150 vdd gnd cell_6t
Xbit_r151_c138 bl_138 br_138 wl_151 vdd gnd cell_6t
Xbit_r152_c138 bl_138 br_138 wl_152 vdd gnd cell_6t
Xbit_r153_c138 bl_138 br_138 wl_153 vdd gnd cell_6t
Xbit_r154_c138 bl_138 br_138 wl_154 vdd gnd cell_6t
Xbit_r155_c138 bl_138 br_138 wl_155 vdd gnd cell_6t
Xbit_r156_c138 bl_138 br_138 wl_156 vdd gnd cell_6t
Xbit_r157_c138 bl_138 br_138 wl_157 vdd gnd cell_6t
Xbit_r158_c138 bl_138 br_138 wl_158 vdd gnd cell_6t
Xbit_r159_c138 bl_138 br_138 wl_159 vdd gnd cell_6t
Xbit_r160_c138 bl_138 br_138 wl_160 vdd gnd cell_6t
Xbit_r161_c138 bl_138 br_138 wl_161 vdd gnd cell_6t
Xbit_r162_c138 bl_138 br_138 wl_162 vdd gnd cell_6t
Xbit_r163_c138 bl_138 br_138 wl_163 vdd gnd cell_6t
Xbit_r164_c138 bl_138 br_138 wl_164 vdd gnd cell_6t
Xbit_r165_c138 bl_138 br_138 wl_165 vdd gnd cell_6t
Xbit_r166_c138 bl_138 br_138 wl_166 vdd gnd cell_6t
Xbit_r167_c138 bl_138 br_138 wl_167 vdd gnd cell_6t
Xbit_r168_c138 bl_138 br_138 wl_168 vdd gnd cell_6t
Xbit_r169_c138 bl_138 br_138 wl_169 vdd gnd cell_6t
Xbit_r170_c138 bl_138 br_138 wl_170 vdd gnd cell_6t
Xbit_r171_c138 bl_138 br_138 wl_171 vdd gnd cell_6t
Xbit_r172_c138 bl_138 br_138 wl_172 vdd gnd cell_6t
Xbit_r173_c138 bl_138 br_138 wl_173 vdd gnd cell_6t
Xbit_r174_c138 bl_138 br_138 wl_174 vdd gnd cell_6t
Xbit_r175_c138 bl_138 br_138 wl_175 vdd gnd cell_6t
Xbit_r176_c138 bl_138 br_138 wl_176 vdd gnd cell_6t
Xbit_r177_c138 bl_138 br_138 wl_177 vdd gnd cell_6t
Xbit_r178_c138 bl_138 br_138 wl_178 vdd gnd cell_6t
Xbit_r179_c138 bl_138 br_138 wl_179 vdd gnd cell_6t
Xbit_r180_c138 bl_138 br_138 wl_180 vdd gnd cell_6t
Xbit_r181_c138 bl_138 br_138 wl_181 vdd gnd cell_6t
Xbit_r182_c138 bl_138 br_138 wl_182 vdd gnd cell_6t
Xbit_r183_c138 bl_138 br_138 wl_183 vdd gnd cell_6t
Xbit_r184_c138 bl_138 br_138 wl_184 vdd gnd cell_6t
Xbit_r185_c138 bl_138 br_138 wl_185 vdd gnd cell_6t
Xbit_r186_c138 bl_138 br_138 wl_186 vdd gnd cell_6t
Xbit_r187_c138 bl_138 br_138 wl_187 vdd gnd cell_6t
Xbit_r188_c138 bl_138 br_138 wl_188 vdd gnd cell_6t
Xbit_r189_c138 bl_138 br_138 wl_189 vdd gnd cell_6t
Xbit_r190_c138 bl_138 br_138 wl_190 vdd gnd cell_6t
Xbit_r191_c138 bl_138 br_138 wl_191 vdd gnd cell_6t
Xbit_r192_c138 bl_138 br_138 wl_192 vdd gnd cell_6t
Xbit_r193_c138 bl_138 br_138 wl_193 vdd gnd cell_6t
Xbit_r194_c138 bl_138 br_138 wl_194 vdd gnd cell_6t
Xbit_r195_c138 bl_138 br_138 wl_195 vdd gnd cell_6t
Xbit_r196_c138 bl_138 br_138 wl_196 vdd gnd cell_6t
Xbit_r197_c138 bl_138 br_138 wl_197 vdd gnd cell_6t
Xbit_r198_c138 bl_138 br_138 wl_198 vdd gnd cell_6t
Xbit_r199_c138 bl_138 br_138 wl_199 vdd gnd cell_6t
Xbit_r200_c138 bl_138 br_138 wl_200 vdd gnd cell_6t
Xbit_r201_c138 bl_138 br_138 wl_201 vdd gnd cell_6t
Xbit_r202_c138 bl_138 br_138 wl_202 vdd gnd cell_6t
Xbit_r203_c138 bl_138 br_138 wl_203 vdd gnd cell_6t
Xbit_r204_c138 bl_138 br_138 wl_204 vdd gnd cell_6t
Xbit_r205_c138 bl_138 br_138 wl_205 vdd gnd cell_6t
Xbit_r206_c138 bl_138 br_138 wl_206 vdd gnd cell_6t
Xbit_r207_c138 bl_138 br_138 wl_207 vdd gnd cell_6t
Xbit_r208_c138 bl_138 br_138 wl_208 vdd gnd cell_6t
Xbit_r209_c138 bl_138 br_138 wl_209 vdd gnd cell_6t
Xbit_r210_c138 bl_138 br_138 wl_210 vdd gnd cell_6t
Xbit_r211_c138 bl_138 br_138 wl_211 vdd gnd cell_6t
Xbit_r212_c138 bl_138 br_138 wl_212 vdd gnd cell_6t
Xbit_r213_c138 bl_138 br_138 wl_213 vdd gnd cell_6t
Xbit_r214_c138 bl_138 br_138 wl_214 vdd gnd cell_6t
Xbit_r215_c138 bl_138 br_138 wl_215 vdd gnd cell_6t
Xbit_r216_c138 bl_138 br_138 wl_216 vdd gnd cell_6t
Xbit_r217_c138 bl_138 br_138 wl_217 vdd gnd cell_6t
Xbit_r218_c138 bl_138 br_138 wl_218 vdd gnd cell_6t
Xbit_r219_c138 bl_138 br_138 wl_219 vdd gnd cell_6t
Xbit_r220_c138 bl_138 br_138 wl_220 vdd gnd cell_6t
Xbit_r221_c138 bl_138 br_138 wl_221 vdd gnd cell_6t
Xbit_r222_c138 bl_138 br_138 wl_222 vdd gnd cell_6t
Xbit_r223_c138 bl_138 br_138 wl_223 vdd gnd cell_6t
Xbit_r224_c138 bl_138 br_138 wl_224 vdd gnd cell_6t
Xbit_r225_c138 bl_138 br_138 wl_225 vdd gnd cell_6t
Xbit_r226_c138 bl_138 br_138 wl_226 vdd gnd cell_6t
Xbit_r227_c138 bl_138 br_138 wl_227 vdd gnd cell_6t
Xbit_r228_c138 bl_138 br_138 wl_228 vdd gnd cell_6t
Xbit_r229_c138 bl_138 br_138 wl_229 vdd gnd cell_6t
Xbit_r230_c138 bl_138 br_138 wl_230 vdd gnd cell_6t
Xbit_r231_c138 bl_138 br_138 wl_231 vdd gnd cell_6t
Xbit_r232_c138 bl_138 br_138 wl_232 vdd gnd cell_6t
Xbit_r233_c138 bl_138 br_138 wl_233 vdd gnd cell_6t
Xbit_r234_c138 bl_138 br_138 wl_234 vdd gnd cell_6t
Xbit_r235_c138 bl_138 br_138 wl_235 vdd gnd cell_6t
Xbit_r236_c138 bl_138 br_138 wl_236 vdd gnd cell_6t
Xbit_r237_c138 bl_138 br_138 wl_237 vdd gnd cell_6t
Xbit_r238_c138 bl_138 br_138 wl_238 vdd gnd cell_6t
Xbit_r239_c138 bl_138 br_138 wl_239 vdd gnd cell_6t
Xbit_r240_c138 bl_138 br_138 wl_240 vdd gnd cell_6t
Xbit_r241_c138 bl_138 br_138 wl_241 vdd gnd cell_6t
Xbit_r242_c138 bl_138 br_138 wl_242 vdd gnd cell_6t
Xbit_r243_c138 bl_138 br_138 wl_243 vdd gnd cell_6t
Xbit_r244_c138 bl_138 br_138 wl_244 vdd gnd cell_6t
Xbit_r245_c138 bl_138 br_138 wl_245 vdd gnd cell_6t
Xbit_r246_c138 bl_138 br_138 wl_246 vdd gnd cell_6t
Xbit_r247_c138 bl_138 br_138 wl_247 vdd gnd cell_6t
Xbit_r248_c138 bl_138 br_138 wl_248 vdd gnd cell_6t
Xbit_r249_c138 bl_138 br_138 wl_249 vdd gnd cell_6t
Xbit_r250_c138 bl_138 br_138 wl_250 vdd gnd cell_6t
Xbit_r251_c138 bl_138 br_138 wl_251 vdd gnd cell_6t
Xbit_r252_c138 bl_138 br_138 wl_252 vdd gnd cell_6t
Xbit_r253_c138 bl_138 br_138 wl_253 vdd gnd cell_6t
Xbit_r254_c138 bl_138 br_138 wl_254 vdd gnd cell_6t
Xbit_r255_c138 bl_138 br_138 wl_255 vdd gnd cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd cell_6t
Xbit_r1_c139 bl_139 br_139 wl_1 vdd gnd cell_6t
Xbit_r2_c139 bl_139 br_139 wl_2 vdd gnd cell_6t
Xbit_r3_c139 bl_139 br_139 wl_3 vdd gnd cell_6t
Xbit_r4_c139 bl_139 br_139 wl_4 vdd gnd cell_6t
Xbit_r5_c139 bl_139 br_139 wl_5 vdd gnd cell_6t
Xbit_r6_c139 bl_139 br_139 wl_6 vdd gnd cell_6t
Xbit_r7_c139 bl_139 br_139 wl_7 vdd gnd cell_6t
Xbit_r8_c139 bl_139 br_139 wl_8 vdd gnd cell_6t
Xbit_r9_c139 bl_139 br_139 wl_9 vdd gnd cell_6t
Xbit_r10_c139 bl_139 br_139 wl_10 vdd gnd cell_6t
Xbit_r11_c139 bl_139 br_139 wl_11 vdd gnd cell_6t
Xbit_r12_c139 bl_139 br_139 wl_12 vdd gnd cell_6t
Xbit_r13_c139 bl_139 br_139 wl_13 vdd gnd cell_6t
Xbit_r14_c139 bl_139 br_139 wl_14 vdd gnd cell_6t
Xbit_r15_c139 bl_139 br_139 wl_15 vdd gnd cell_6t
Xbit_r16_c139 bl_139 br_139 wl_16 vdd gnd cell_6t
Xbit_r17_c139 bl_139 br_139 wl_17 vdd gnd cell_6t
Xbit_r18_c139 bl_139 br_139 wl_18 vdd gnd cell_6t
Xbit_r19_c139 bl_139 br_139 wl_19 vdd gnd cell_6t
Xbit_r20_c139 bl_139 br_139 wl_20 vdd gnd cell_6t
Xbit_r21_c139 bl_139 br_139 wl_21 vdd gnd cell_6t
Xbit_r22_c139 bl_139 br_139 wl_22 vdd gnd cell_6t
Xbit_r23_c139 bl_139 br_139 wl_23 vdd gnd cell_6t
Xbit_r24_c139 bl_139 br_139 wl_24 vdd gnd cell_6t
Xbit_r25_c139 bl_139 br_139 wl_25 vdd gnd cell_6t
Xbit_r26_c139 bl_139 br_139 wl_26 vdd gnd cell_6t
Xbit_r27_c139 bl_139 br_139 wl_27 vdd gnd cell_6t
Xbit_r28_c139 bl_139 br_139 wl_28 vdd gnd cell_6t
Xbit_r29_c139 bl_139 br_139 wl_29 vdd gnd cell_6t
Xbit_r30_c139 bl_139 br_139 wl_30 vdd gnd cell_6t
Xbit_r31_c139 bl_139 br_139 wl_31 vdd gnd cell_6t
Xbit_r32_c139 bl_139 br_139 wl_32 vdd gnd cell_6t
Xbit_r33_c139 bl_139 br_139 wl_33 vdd gnd cell_6t
Xbit_r34_c139 bl_139 br_139 wl_34 vdd gnd cell_6t
Xbit_r35_c139 bl_139 br_139 wl_35 vdd gnd cell_6t
Xbit_r36_c139 bl_139 br_139 wl_36 vdd gnd cell_6t
Xbit_r37_c139 bl_139 br_139 wl_37 vdd gnd cell_6t
Xbit_r38_c139 bl_139 br_139 wl_38 vdd gnd cell_6t
Xbit_r39_c139 bl_139 br_139 wl_39 vdd gnd cell_6t
Xbit_r40_c139 bl_139 br_139 wl_40 vdd gnd cell_6t
Xbit_r41_c139 bl_139 br_139 wl_41 vdd gnd cell_6t
Xbit_r42_c139 bl_139 br_139 wl_42 vdd gnd cell_6t
Xbit_r43_c139 bl_139 br_139 wl_43 vdd gnd cell_6t
Xbit_r44_c139 bl_139 br_139 wl_44 vdd gnd cell_6t
Xbit_r45_c139 bl_139 br_139 wl_45 vdd gnd cell_6t
Xbit_r46_c139 bl_139 br_139 wl_46 vdd gnd cell_6t
Xbit_r47_c139 bl_139 br_139 wl_47 vdd gnd cell_6t
Xbit_r48_c139 bl_139 br_139 wl_48 vdd gnd cell_6t
Xbit_r49_c139 bl_139 br_139 wl_49 vdd gnd cell_6t
Xbit_r50_c139 bl_139 br_139 wl_50 vdd gnd cell_6t
Xbit_r51_c139 bl_139 br_139 wl_51 vdd gnd cell_6t
Xbit_r52_c139 bl_139 br_139 wl_52 vdd gnd cell_6t
Xbit_r53_c139 bl_139 br_139 wl_53 vdd gnd cell_6t
Xbit_r54_c139 bl_139 br_139 wl_54 vdd gnd cell_6t
Xbit_r55_c139 bl_139 br_139 wl_55 vdd gnd cell_6t
Xbit_r56_c139 bl_139 br_139 wl_56 vdd gnd cell_6t
Xbit_r57_c139 bl_139 br_139 wl_57 vdd gnd cell_6t
Xbit_r58_c139 bl_139 br_139 wl_58 vdd gnd cell_6t
Xbit_r59_c139 bl_139 br_139 wl_59 vdd gnd cell_6t
Xbit_r60_c139 bl_139 br_139 wl_60 vdd gnd cell_6t
Xbit_r61_c139 bl_139 br_139 wl_61 vdd gnd cell_6t
Xbit_r62_c139 bl_139 br_139 wl_62 vdd gnd cell_6t
Xbit_r63_c139 bl_139 br_139 wl_63 vdd gnd cell_6t
Xbit_r64_c139 bl_139 br_139 wl_64 vdd gnd cell_6t
Xbit_r65_c139 bl_139 br_139 wl_65 vdd gnd cell_6t
Xbit_r66_c139 bl_139 br_139 wl_66 vdd gnd cell_6t
Xbit_r67_c139 bl_139 br_139 wl_67 vdd gnd cell_6t
Xbit_r68_c139 bl_139 br_139 wl_68 vdd gnd cell_6t
Xbit_r69_c139 bl_139 br_139 wl_69 vdd gnd cell_6t
Xbit_r70_c139 bl_139 br_139 wl_70 vdd gnd cell_6t
Xbit_r71_c139 bl_139 br_139 wl_71 vdd gnd cell_6t
Xbit_r72_c139 bl_139 br_139 wl_72 vdd gnd cell_6t
Xbit_r73_c139 bl_139 br_139 wl_73 vdd gnd cell_6t
Xbit_r74_c139 bl_139 br_139 wl_74 vdd gnd cell_6t
Xbit_r75_c139 bl_139 br_139 wl_75 vdd gnd cell_6t
Xbit_r76_c139 bl_139 br_139 wl_76 vdd gnd cell_6t
Xbit_r77_c139 bl_139 br_139 wl_77 vdd gnd cell_6t
Xbit_r78_c139 bl_139 br_139 wl_78 vdd gnd cell_6t
Xbit_r79_c139 bl_139 br_139 wl_79 vdd gnd cell_6t
Xbit_r80_c139 bl_139 br_139 wl_80 vdd gnd cell_6t
Xbit_r81_c139 bl_139 br_139 wl_81 vdd gnd cell_6t
Xbit_r82_c139 bl_139 br_139 wl_82 vdd gnd cell_6t
Xbit_r83_c139 bl_139 br_139 wl_83 vdd gnd cell_6t
Xbit_r84_c139 bl_139 br_139 wl_84 vdd gnd cell_6t
Xbit_r85_c139 bl_139 br_139 wl_85 vdd gnd cell_6t
Xbit_r86_c139 bl_139 br_139 wl_86 vdd gnd cell_6t
Xbit_r87_c139 bl_139 br_139 wl_87 vdd gnd cell_6t
Xbit_r88_c139 bl_139 br_139 wl_88 vdd gnd cell_6t
Xbit_r89_c139 bl_139 br_139 wl_89 vdd gnd cell_6t
Xbit_r90_c139 bl_139 br_139 wl_90 vdd gnd cell_6t
Xbit_r91_c139 bl_139 br_139 wl_91 vdd gnd cell_6t
Xbit_r92_c139 bl_139 br_139 wl_92 vdd gnd cell_6t
Xbit_r93_c139 bl_139 br_139 wl_93 vdd gnd cell_6t
Xbit_r94_c139 bl_139 br_139 wl_94 vdd gnd cell_6t
Xbit_r95_c139 bl_139 br_139 wl_95 vdd gnd cell_6t
Xbit_r96_c139 bl_139 br_139 wl_96 vdd gnd cell_6t
Xbit_r97_c139 bl_139 br_139 wl_97 vdd gnd cell_6t
Xbit_r98_c139 bl_139 br_139 wl_98 vdd gnd cell_6t
Xbit_r99_c139 bl_139 br_139 wl_99 vdd gnd cell_6t
Xbit_r100_c139 bl_139 br_139 wl_100 vdd gnd cell_6t
Xbit_r101_c139 bl_139 br_139 wl_101 vdd gnd cell_6t
Xbit_r102_c139 bl_139 br_139 wl_102 vdd gnd cell_6t
Xbit_r103_c139 bl_139 br_139 wl_103 vdd gnd cell_6t
Xbit_r104_c139 bl_139 br_139 wl_104 vdd gnd cell_6t
Xbit_r105_c139 bl_139 br_139 wl_105 vdd gnd cell_6t
Xbit_r106_c139 bl_139 br_139 wl_106 vdd gnd cell_6t
Xbit_r107_c139 bl_139 br_139 wl_107 vdd gnd cell_6t
Xbit_r108_c139 bl_139 br_139 wl_108 vdd gnd cell_6t
Xbit_r109_c139 bl_139 br_139 wl_109 vdd gnd cell_6t
Xbit_r110_c139 bl_139 br_139 wl_110 vdd gnd cell_6t
Xbit_r111_c139 bl_139 br_139 wl_111 vdd gnd cell_6t
Xbit_r112_c139 bl_139 br_139 wl_112 vdd gnd cell_6t
Xbit_r113_c139 bl_139 br_139 wl_113 vdd gnd cell_6t
Xbit_r114_c139 bl_139 br_139 wl_114 vdd gnd cell_6t
Xbit_r115_c139 bl_139 br_139 wl_115 vdd gnd cell_6t
Xbit_r116_c139 bl_139 br_139 wl_116 vdd gnd cell_6t
Xbit_r117_c139 bl_139 br_139 wl_117 vdd gnd cell_6t
Xbit_r118_c139 bl_139 br_139 wl_118 vdd gnd cell_6t
Xbit_r119_c139 bl_139 br_139 wl_119 vdd gnd cell_6t
Xbit_r120_c139 bl_139 br_139 wl_120 vdd gnd cell_6t
Xbit_r121_c139 bl_139 br_139 wl_121 vdd gnd cell_6t
Xbit_r122_c139 bl_139 br_139 wl_122 vdd gnd cell_6t
Xbit_r123_c139 bl_139 br_139 wl_123 vdd gnd cell_6t
Xbit_r124_c139 bl_139 br_139 wl_124 vdd gnd cell_6t
Xbit_r125_c139 bl_139 br_139 wl_125 vdd gnd cell_6t
Xbit_r126_c139 bl_139 br_139 wl_126 vdd gnd cell_6t
Xbit_r127_c139 bl_139 br_139 wl_127 vdd gnd cell_6t
Xbit_r128_c139 bl_139 br_139 wl_128 vdd gnd cell_6t
Xbit_r129_c139 bl_139 br_139 wl_129 vdd gnd cell_6t
Xbit_r130_c139 bl_139 br_139 wl_130 vdd gnd cell_6t
Xbit_r131_c139 bl_139 br_139 wl_131 vdd gnd cell_6t
Xbit_r132_c139 bl_139 br_139 wl_132 vdd gnd cell_6t
Xbit_r133_c139 bl_139 br_139 wl_133 vdd gnd cell_6t
Xbit_r134_c139 bl_139 br_139 wl_134 vdd gnd cell_6t
Xbit_r135_c139 bl_139 br_139 wl_135 vdd gnd cell_6t
Xbit_r136_c139 bl_139 br_139 wl_136 vdd gnd cell_6t
Xbit_r137_c139 bl_139 br_139 wl_137 vdd gnd cell_6t
Xbit_r138_c139 bl_139 br_139 wl_138 vdd gnd cell_6t
Xbit_r139_c139 bl_139 br_139 wl_139 vdd gnd cell_6t
Xbit_r140_c139 bl_139 br_139 wl_140 vdd gnd cell_6t
Xbit_r141_c139 bl_139 br_139 wl_141 vdd gnd cell_6t
Xbit_r142_c139 bl_139 br_139 wl_142 vdd gnd cell_6t
Xbit_r143_c139 bl_139 br_139 wl_143 vdd gnd cell_6t
Xbit_r144_c139 bl_139 br_139 wl_144 vdd gnd cell_6t
Xbit_r145_c139 bl_139 br_139 wl_145 vdd gnd cell_6t
Xbit_r146_c139 bl_139 br_139 wl_146 vdd gnd cell_6t
Xbit_r147_c139 bl_139 br_139 wl_147 vdd gnd cell_6t
Xbit_r148_c139 bl_139 br_139 wl_148 vdd gnd cell_6t
Xbit_r149_c139 bl_139 br_139 wl_149 vdd gnd cell_6t
Xbit_r150_c139 bl_139 br_139 wl_150 vdd gnd cell_6t
Xbit_r151_c139 bl_139 br_139 wl_151 vdd gnd cell_6t
Xbit_r152_c139 bl_139 br_139 wl_152 vdd gnd cell_6t
Xbit_r153_c139 bl_139 br_139 wl_153 vdd gnd cell_6t
Xbit_r154_c139 bl_139 br_139 wl_154 vdd gnd cell_6t
Xbit_r155_c139 bl_139 br_139 wl_155 vdd gnd cell_6t
Xbit_r156_c139 bl_139 br_139 wl_156 vdd gnd cell_6t
Xbit_r157_c139 bl_139 br_139 wl_157 vdd gnd cell_6t
Xbit_r158_c139 bl_139 br_139 wl_158 vdd gnd cell_6t
Xbit_r159_c139 bl_139 br_139 wl_159 vdd gnd cell_6t
Xbit_r160_c139 bl_139 br_139 wl_160 vdd gnd cell_6t
Xbit_r161_c139 bl_139 br_139 wl_161 vdd gnd cell_6t
Xbit_r162_c139 bl_139 br_139 wl_162 vdd gnd cell_6t
Xbit_r163_c139 bl_139 br_139 wl_163 vdd gnd cell_6t
Xbit_r164_c139 bl_139 br_139 wl_164 vdd gnd cell_6t
Xbit_r165_c139 bl_139 br_139 wl_165 vdd gnd cell_6t
Xbit_r166_c139 bl_139 br_139 wl_166 vdd gnd cell_6t
Xbit_r167_c139 bl_139 br_139 wl_167 vdd gnd cell_6t
Xbit_r168_c139 bl_139 br_139 wl_168 vdd gnd cell_6t
Xbit_r169_c139 bl_139 br_139 wl_169 vdd gnd cell_6t
Xbit_r170_c139 bl_139 br_139 wl_170 vdd gnd cell_6t
Xbit_r171_c139 bl_139 br_139 wl_171 vdd gnd cell_6t
Xbit_r172_c139 bl_139 br_139 wl_172 vdd gnd cell_6t
Xbit_r173_c139 bl_139 br_139 wl_173 vdd gnd cell_6t
Xbit_r174_c139 bl_139 br_139 wl_174 vdd gnd cell_6t
Xbit_r175_c139 bl_139 br_139 wl_175 vdd gnd cell_6t
Xbit_r176_c139 bl_139 br_139 wl_176 vdd gnd cell_6t
Xbit_r177_c139 bl_139 br_139 wl_177 vdd gnd cell_6t
Xbit_r178_c139 bl_139 br_139 wl_178 vdd gnd cell_6t
Xbit_r179_c139 bl_139 br_139 wl_179 vdd gnd cell_6t
Xbit_r180_c139 bl_139 br_139 wl_180 vdd gnd cell_6t
Xbit_r181_c139 bl_139 br_139 wl_181 vdd gnd cell_6t
Xbit_r182_c139 bl_139 br_139 wl_182 vdd gnd cell_6t
Xbit_r183_c139 bl_139 br_139 wl_183 vdd gnd cell_6t
Xbit_r184_c139 bl_139 br_139 wl_184 vdd gnd cell_6t
Xbit_r185_c139 bl_139 br_139 wl_185 vdd gnd cell_6t
Xbit_r186_c139 bl_139 br_139 wl_186 vdd gnd cell_6t
Xbit_r187_c139 bl_139 br_139 wl_187 vdd gnd cell_6t
Xbit_r188_c139 bl_139 br_139 wl_188 vdd gnd cell_6t
Xbit_r189_c139 bl_139 br_139 wl_189 vdd gnd cell_6t
Xbit_r190_c139 bl_139 br_139 wl_190 vdd gnd cell_6t
Xbit_r191_c139 bl_139 br_139 wl_191 vdd gnd cell_6t
Xbit_r192_c139 bl_139 br_139 wl_192 vdd gnd cell_6t
Xbit_r193_c139 bl_139 br_139 wl_193 vdd gnd cell_6t
Xbit_r194_c139 bl_139 br_139 wl_194 vdd gnd cell_6t
Xbit_r195_c139 bl_139 br_139 wl_195 vdd gnd cell_6t
Xbit_r196_c139 bl_139 br_139 wl_196 vdd gnd cell_6t
Xbit_r197_c139 bl_139 br_139 wl_197 vdd gnd cell_6t
Xbit_r198_c139 bl_139 br_139 wl_198 vdd gnd cell_6t
Xbit_r199_c139 bl_139 br_139 wl_199 vdd gnd cell_6t
Xbit_r200_c139 bl_139 br_139 wl_200 vdd gnd cell_6t
Xbit_r201_c139 bl_139 br_139 wl_201 vdd gnd cell_6t
Xbit_r202_c139 bl_139 br_139 wl_202 vdd gnd cell_6t
Xbit_r203_c139 bl_139 br_139 wl_203 vdd gnd cell_6t
Xbit_r204_c139 bl_139 br_139 wl_204 vdd gnd cell_6t
Xbit_r205_c139 bl_139 br_139 wl_205 vdd gnd cell_6t
Xbit_r206_c139 bl_139 br_139 wl_206 vdd gnd cell_6t
Xbit_r207_c139 bl_139 br_139 wl_207 vdd gnd cell_6t
Xbit_r208_c139 bl_139 br_139 wl_208 vdd gnd cell_6t
Xbit_r209_c139 bl_139 br_139 wl_209 vdd gnd cell_6t
Xbit_r210_c139 bl_139 br_139 wl_210 vdd gnd cell_6t
Xbit_r211_c139 bl_139 br_139 wl_211 vdd gnd cell_6t
Xbit_r212_c139 bl_139 br_139 wl_212 vdd gnd cell_6t
Xbit_r213_c139 bl_139 br_139 wl_213 vdd gnd cell_6t
Xbit_r214_c139 bl_139 br_139 wl_214 vdd gnd cell_6t
Xbit_r215_c139 bl_139 br_139 wl_215 vdd gnd cell_6t
Xbit_r216_c139 bl_139 br_139 wl_216 vdd gnd cell_6t
Xbit_r217_c139 bl_139 br_139 wl_217 vdd gnd cell_6t
Xbit_r218_c139 bl_139 br_139 wl_218 vdd gnd cell_6t
Xbit_r219_c139 bl_139 br_139 wl_219 vdd gnd cell_6t
Xbit_r220_c139 bl_139 br_139 wl_220 vdd gnd cell_6t
Xbit_r221_c139 bl_139 br_139 wl_221 vdd gnd cell_6t
Xbit_r222_c139 bl_139 br_139 wl_222 vdd gnd cell_6t
Xbit_r223_c139 bl_139 br_139 wl_223 vdd gnd cell_6t
Xbit_r224_c139 bl_139 br_139 wl_224 vdd gnd cell_6t
Xbit_r225_c139 bl_139 br_139 wl_225 vdd gnd cell_6t
Xbit_r226_c139 bl_139 br_139 wl_226 vdd gnd cell_6t
Xbit_r227_c139 bl_139 br_139 wl_227 vdd gnd cell_6t
Xbit_r228_c139 bl_139 br_139 wl_228 vdd gnd cell_6t
Xbit_r229_c139 bl_139 br_139 wl_229 vdd gnd cell_6t
Xbit_r230_c139 bl_139 br_139 wl_230 vdd gnd cell_6t
Xbit_r231_c139 bl_139 br_139 wl_231 vdd gnd cell_6t
Xbit_r232_c139 bl_139 br_139 wl_232 vdd gnd cell_6t
Xbit_r233_c139 bl_139 br_139 wl_233 vdd gnd cell_6t
Xbit_r234_c139 bl_139 br_139 wl_234 vdd gnd cell_6t
Xbit_r235_c139 bl_139 br_139 wl_235 vdd gnd cell_6t
Xbit_r236_c139 bl_139 br_139 wl_236 vdd gnd cell_6t
Xbit_r237_c139 bl_139 br_139 wl_237 vdd gnd cell_6t
Xbit_r238_c139 bl_139 br_139 wl_238 vdd gnd cell_6t
Xbit_r239_c139 bl_139 br_139 wl_239 vdd gnd cell_6t
Xbit_r240_c139 bl_139 br_139 wl_240 vdd gnd cell_6t
Xbit_r241_c139 bl_139 br_139 wl_241 vdd gnd cell_6t
Xbit_r242_c139 bl_139 br_139 wl_242 vdd gnd cell_6t
Xbit_r243_c139 bl_139 br_139 wl_243 vdd gnd cell_6t
Xbit_r244_c139 bl_139 br_139 wl_244 vdd gnd cell_6t
Xbit_r245_c139 bl_139 br_139 wl_245 vdd gnd cell_6t
Xbit_r246_c139 bl_139 br_139 wl_246 vdd gnd cell_6t
Xbit_r247_c139 bl_139 br_139 wl_247 vdd gnd cell_6t
Xbit_r248_c139 bl_139 br_139 wl_248 vdd gnd cell_6t
Xbit_r249_c139 bl_139 br_139 wl_249 vdd gnd cell_6t
Xbit_r250_c139 bl_139 br_139 wl_250 vdd gnd cell_6t
Xbit_r251_c139 bl_139 br_139 wl_251 vdd gnd cell_6t
Xbit_r252_c139 bl_139 br_139 wl_252 vdd gnd cell_6t
Xbit_r253_c139 bl_139 br_139 wl_253 vdd gnd cell_6t
Xbit_r254_c139 bl_139 br_139 wl_254 vdd gnd cell_6t
Xbit_r255_c139 bl_139 br_139 wl_255 vdd gnd cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd cell_6t
Xbit_r1_c140 bl_140 br_140 wl_1 vdd gnd cell_6t
Xbit_r2_c140 bl_140 br_140 wl_2 vdd gnd cell_6t
Xbit_r3_c140 bl_140 br_140 wl_3 vdd gnd cell_6t
Xbit_r4_c140 bl_140 br_140 wl_4 vdd gnd cell_6t
Xbit_r5_c140 bl_140 br_140 wl_5 vdd gnd cell_6t
Xbit_r6_c140 bl_140 br_140 wl_6 vdd gnd cell_6t
Xbit_r7_c140 bl_140 br_140 wl_7 vdd gnd cell_6t
Xbit_r8_c140 bl_140 br_140 wl_8 vdd gnd cell_6t
Xbit_r9_c140 bl_140 br_140 wl_9 vdd gnd cell_6t
Xbit_r10_c140 bl_140 br_140 wl_10 vdd gnd cell_6t
Xbit_r11_c140 bl_140 br_140 wl_11 vdd gnd cell_6t
Xbit_r12_c140 bl_140 br_140 wl_12 vdd gnd cell_6t
Xbit_r13_c140 bl_140 br_140 wl_13 vdd gnd cell_6t
Xbit_r14_c140 bl_140 br_140 wl_14 vdd gnd cell_6t
Xbit_r15_c140 bl_140 br_140 wl_15 vdd gnd cell_6t
Xbit_r16_c140 bl_140 br_140 wl_16 vdd gnd cell_6t
Xbit_r17_c140 bl_140 br_140 wl_17 vdd gnd cell_6t
Xbit_r18_c140 bl_140 br_140 wl_18 vdd gnd cell_6t
Xbit_r19_c140 bl_140 br_140 wl_19 vdd gnd cell_6t
Xbit_r20_c140 bl_140 br_140 wl_20 vdd gnd cell_6t
Xbit_r21_c140 bl_140 br_140 wl_21 vdd gnd cell_6t
Xbit_r22_c140 bl_140 br_140 wl_22 vdd gnd cell_6t
Xbit_r23_c140 bl_140 br_140 wl_23 vdd gnd cell_6t
Xbit_r24_c140 bl_140 br_140 wl_24 vdd gnd cell_6t
Xbit_r25_c140 bl_140 br_140 wl_25 vdd gnd cell_6t
Xbit_r26_c140 bl_140 br_140 wl_26 vdd gnd cell_6t
Xbit_r27_c140 bl_140 br_140 wl_27 vdd gnd cell_6t
Xbit_r28_c140 bl_140 br_140 wl_28 vdd gnd cell_6t
Xbit_r29_c140 bl_140 br_140 wl_29 vdd gnd cell_6t
Xbit_r30_c140 bl_140 br_140 wl_30 vdd gnd cell_6t
Xbit_r31_c140 bl_140 br_140 wl_31 vdd gnd cell_6t
Xbit_r32_c140 bl_140 br_140 wl_32 vdd gnd cell_6t
Xbit_r33_c140 bl_140 br_140 wl_33 vdd gnd cell_6t
Xbit_r34_c140 bl_140 br_140 wl_34 vdd gnd cell_6t
Xbit_r35_c140 bl_140 br_140 wl_35 vdd gnd cell_6t
Xbit_r36_c140 bl_140 br_140 wl_36 vdd gnd cell_6t
Xbit_r37_c140 bl_140 br_140 wl_37 vdd gnd cell_6t
Xbit_r38_c140 bl_140 br_140 wl_38 vdd gnd cell_6t
Xbit_r39_c140 bl_140 br_140 wl_39 vdd gnd cell_6t
Xbit_r40_c140 bl_140 br_140 wl_40 vdd gnd cell_6t
Xbit_r41_c140 bl_140 br_140 wl_41 vdd gnd cell_6t
Xbit_r42_c140 bl_140 br_140 wl_42 vdd gnd cell_6t
Xbit_r43_c140 bl_140 br_140 wl_43 vdd gnd cell_6t
Xbit_r44_c140 bl_140 br_140 wl_44 vdd gnd cell_6t
Xbit_r45_c140 bl_140 br_140 wl_45 vdd gnd cell_6t
Xbit_r46_c140 bl_140 br_140 wl_46 vdd gnd cell_6t
Xbit_r47_c140 bl_140 br_140 wl_47 vdd gnd cell_6t
Xbit_r48_c140 bl_140 br_140 wl_48 vdd gnd cell_6t
Xbit_r49_c140 bl_140 br_140 wl_49 vdd gnd cell_6t
Xbit_r50_c140 bl_140 br_140 wl_50 vdd gnd cell_6t
Xbit_r51_c140 bl_140 br_140 wl_51 vdd gnd cell_6t
Xbit_r52_c140 bl_140 br_140 wl_52 vdd gnd cell_6t
Xbit_r53_c140 bl_140 br_140 wl_53 vdd gnd cell_6t
Xbit_r54_c140 bl_140 br_140 wl_54 vdd gnd cell_6t
Xbit_r55_c140 bl_140 br_140 wl_55 vdd gnd cell_6t
Xbit_r56_c140 bl_140 br_140 wl_56 vdd gnd cell_6t
Xbit_r57_c140 bl_140 br_140 wl_57 vdd gnd cell_6t
Xbit_r58_c140 bl_140 br_140 wl_58 vdd gnd cell_6t
Xbit_r59_c140 bl_140 br_140 wl_59 vdd gnd cell_6t
Xbit_r60_c140 bl_140 br_140 wl_60 vdd gnd cell_6t
Xbit_r61_c140 bl_140 br_140 wl_61 vdd gnd cell_6t
Xbit_r62_c140 bl_140 br_140 wl_62 vdd gnd cell_6t
Xbit_r63_c140 bl_140 br_140 wl_63 vdd gnd cell_6t
Xbit_r64_c140 bl_140 br_140 wl_64 vdd gnd cell_6t
Xbit_r65_c140 bl_140 br_140 wl_65 vdd gnd cell_6t
Xbit_r66_c140 bl_140 br_140 wl_66 vdd gnd cell_6t
Xbit_r67_c140 bl_140 br_140 wl_67 vdd gnd cell_6t
Xbit_r68_c140 bl_140 br_140 wl_68 vdd gnd cell_6t
Xbit_r69_c140 bl_140 br_140 wl_69 vdd gnd cell_6t
Xbit_r70_c140 bl_140 br_140 wl_70 vdd gnd cell_6t
Xbit_r71_c140 bl_140 br_140 wl_71 vdd gnd cell_6t
Xbit_r72_c140 bl_140 br_140 wl_72 vdd gnd cell_6t
Xbit_r73_c140 bl_140 br_140 wl_73 vdd gnd cell_6t
Xbit_r74_c140 bl_140 br_140 wl_74 vdd gnd cell_6t
Xbit_r75_c140 bl_140 br_140 wl_75 vdd gnd cell_6t
Xbit_r76_c140 bl_140 br_140 wl_76 vdd gnd cell_6t
Xbit_r77_c140 bl_140 br_140 wl_77 vdd gnd cell_6t
Xbit_r78_c140 bl_140 br_140 wl_78 vdd gnd cell_6t
Xbit_r79_c140 bl_140 br_140 wl_79 vdd gnd cell_6t
Xbit_r80_c140 bl_140 br_140 wl_80 vdd gnd cell_6t
Xbit_r81_c140 bl_140 br_140 wl_81 vdd gnd cell_6t
Xbit_r82_c140 bl_140 br_140 wl_82 vdd gnd cell_6t
Xbit_r83_c140 bl_140 br_140 wl_83 vdd gnd cell_6t
Xbit_r84_c140 bl_140 br_140 wl_84 vdd gnd cell_6t
Xbit_r85_c140 bl_140 br_140 wl_85 vdd gnd cell_6t
Xbit_r86_c140 bl_140 br_140 wl_86 vdd gnd cell_6t
Xbit_r87_c140 bl_140 br_140 wl_87 vdd gnd cell_6t
Xbit_r88_c140 bl_140 br_140 wl_88 vdd gnd cell_6t
Xbit_r89_c140 bl_140 br_140 wl_89 vdd gnd cell_6t
Xbit_r90_c140 bl_140 br_140 wl_90 vdd gnd cell_6t
Xbit_r91_c140 bl_140 br_140 wl_91 vdd gnd cell_6t
Xbit_r92_c140 bl_140 br_140 wl_92 vdd gnd cell_6t
Xbit_r93_c140 bl_140 br_140 wl_93 vdd gnd cell_6t
Xbit_r94_c140 bl_140 br_140 wl_94 vdd gnd cell_6t
Xbit_r95_c140 bl_140 br_140 wl_95 vdd gnd cell_6t
Xbit_r96_c140 bl_140 br_140 wl_96 vdd gnd cell_6t
Xbit_r97_c140 bl_140 br_140 wl_97 vdd gnd cell_6t
Xbit_r98_c140 bl_140 br_140 wl_98 vdd gnd cell_6t
Xbit_r99_c140 bl_140 br_140 wl_99 vdd gnd cell_6t
Xbit_r100_c140 bl_140 br_140 wl_100 vdd gnd cell_6t
Xbit_r101_c140 bl_140 br_140 wl_101 vdd gnd cell_6t
Xbit_r102_c140 bl_140 br_140 wl_102 vdd gnd cell_6t
Xbit_r103_c140 bl_140 br_140 wl_103 vdd gnd cell_6t
Xbit_r104_c140 bl_140 br_140 wl_104 vdd gnd cell_6t
Xbit_r105_c140 bl_140 br_140 wl_105 vdd gnd cell_6t
Xbit_r106_c140 bl_140 br_140 wl_106 vdd gnd cell_6t
Xbit_r107_c140 bl_140 br_140 wl_107 vdd gnd cell_6t
Xbit_r108_c140 bl_140 br_140 wl_108 vdd gnd cell_6t
Xbit_r109_c140 bl_140 br_140 wl_109 vdd gnd cell_6t
Xbit_r110_c140 bl_140 br_140 wl_110 vdd gnd cell_6t
Xbit_r111_c140 bl_140 br_140 wl_111 vdd gnd cell_6t
Xbit_r112_c140 bl_140 br_140 wl_112 vdd gnd cell_6t
Xbit_r113_c140 bl_140 br_140 wl_113 vdd gnd cell_6t
Xbit_r114_c140 bl_140 br_140 wl_114 vdd gnd cell_6t
Xbit_r115_c140 bl_140 br_140 wl_115 vdd gnd cell_6t
Xbit_r116_c140 bl_140 br_140 wl_116 vdd gnd cell_6t
Xbit_r117_c140 bl_140 br_140 wl_117 vdd gnd cell_6t
Xbit_r118_c140 bl_140 br_140 wl_118 vdd gnd cell_6t
Xbit_r119_c140 bl_140 br_140 wl_119 vdd gnd cell_6t
Xbit_r120_c140 bl_140 br_140 wl_120 vdd gnd cell_6t
Xbit_r121_c140 bl_140 br_140 wl_121 vdd gnd cell_6t
Xbit_r122_c140 bl_140 br_140 wl_122 vdd gnd cell_6t
Xbit_r123_c140 bl_140 br_140 wl_123 vdd gnd cell_6t
Xbit_r124_c140 bl_140 br_140 wl_124 vdd gnd cell_6t
Xbit_r125_c140 bl_140 br_140 wl_125 vdd gnd cell_6t
Xbit_r126_c140 bl_140 br_140 wl_126 vdd gnd cell_6t
Xbit_r127_c140 bl_140 br_140 wl_127 vdd gnd cell_6t
Xbit_r128_c140 bl_140 br_140 wl_128 vdd gnd cell_6t
Xbit_r129_c140 bl_140 br_140 wl_129 vdd gnd cell_6t
Xbit_r130_c140 bl_140 br_140 wl_130 vdd gnd cell_6t
Xbit_r131_c140 bl_140 br_140 wl_131 vdd gnd cell_6t
Xbit_r132_c140 bl_140 br_140 wl_132 vdd gnd cell_6t
Xbit_r133_c140 bl_140 br_140 wl_133 vdd gnd cell_6t
Xbit_r134_c140 bl_140 br_140 wl_134 vdd gnd cell_6t
Xbit_r135_c140 bl_140 br_140 wl_135 vdd gnd cell_6t
Xbit_r136_c140 bl_140 br_140 wl_136 vdd gnd cell_6t
Xbit_r137_c140 bl_140 br_140 wl_137 vdd gnd cell_6t
Xbit_r138_c140 bl_140 br_140 wl_138 vdd gnd cell_6t
Xbit_r139_c140 bl_140 br_140 wl_139 vdd gnd cell_6t
Xbit_r140_c140 bl_140 br_140 wl_140 vdd gnd cell_6t
Xbit_r141_c140 bl_140 br_140 wl_141 vdd gnd cell_6t
Xbit_r142_c140 bl_140 br_140 wl_142 vdd gnd cell_6t
Xbit_r143_c140 bl_140 br_140 wl_143 vdd gnd cell_6t
Xbit_r144_c140 bl_140 br_140 wl_144 vdd gnd cell_6t
Xbit_r145_c140 bl_140 br_140 wl_145 vdd gnd cell_6t
Xbit_r146_c140 bl_140 br_140 wl_146 vdd gnd cell_6t
Xbit_r147_c140 bl_140 br_140 wl_147 vdd gnd cell_6t
Xbit_r148_c140 bl_140 br_140 wl_148 vdd gnd cell_6t
Xbit_r149_c140 bl_140 br_140 wl_149 vdd gnd cell_6t
Xbit_r150_c140 bl_140 br_140 wl_150 vdd gnd cell_6t
Xbit_r151_c140 bl_140 br_140 wl_151 vdd gnd cell_6t
Xbit_r152_c140 bl_140 br_140 wl_152 vdd gnd cell_6t
Xbit_r153_c140 bl_140 br_140 wl_153 vdd gnd cell_6t
Xbit_r154_c140 bl_140 br_140 wl_154 vdd gnd cell_6t
Xbit_r155_c140 bl_140 br_140 wl_155 vdd gnd cell_6t
Xbit_r156_c140 bl_140 br_140 wl_156 vdd gnd cell_6t
Xbit_r157_c140 bl_140 br_140 wl_157 vdd gnd cell_6t
Xbit_r158_c140 bl_140 br_140 wl_158 vdd gnd cell_6t
Xbit_r159_c140 bl_140 br_140 wl_159 vdd gnd cell_6t
Xbit_r160_c140 bl_140 br_140 wl_160 vdd gnd cell_6t
Xbit_r161_c140 bl_140 br_140 wl_161 vdd gnd cell_6t
Xbit_r162_c140 bl_140 br_140 wl_162 vdd gnd cell_6t
Xbit_r163_c140 bl_140 br_140 wl_163 vdd gnd cell_6t
Xbit_r164_c140 bl_140 br_140 wl_164 vdd gnd cell_6t
Xbit_r165_c140 bl_140 br_140 wl_165 vdd gnd cell_6t
Xbit_r166_c140 bl_140 br_140 wl_166 vdd gnd cell_6t
Xbit_r167_c140 bl_140 br_140 wl_167 vdd gnd cell_6t
Xbit_r168_c140 bl_140 br_140 wl_168 vdd gnd cell_6t
Xbit_r169_c140 bl_140 br_140 wl_169 vdd gnd cell_6t
Xbit_r170_c140 bl_140 br_140 wl_170 vdd gnd cell_6t
Xbit_r171_c140 bl_140 br_140 wl_171 vdd gnd cell_6t
Xbit_r172_c140 bl_140 br_140 wl_172 vdd gnd cell_6t
Xbit_r173_c140 bl_140 br_140 wl_173 vdd gnd cell_6t
Xbit_r174_c140 bl_140 br_140 wl_174 vdd gnd cell_6t
Xbit_r175_c140 bl_140 br_140 wl_175 vdd gnd cell_6t
Xbit_r176_c140 bl_140 br_140 wl_176 vdd gnd cell_6t
Xbit_r177_c140 bl_140 br_140 wl_177 vdd gnd cell_6t
Xbit_r178_c140 bl_140 br_140 wl_178 vdd gnd cell_6t
Xbit_r179_c140 bl_140 br_140 wl_179 vdd gnd cell_6t
Xbit_r180_c140 bl_140 br_140 wl_180 vdd gnd cell_6t
Xbit_r181_c140 bl_140 br_140 wl_181 vdd gnd cell_6t
Xbit_r182_c140 bl_140 br_140 wl_182 vdd gnd cell_6t
Xbit_r183_c140 bl_140 br_140 wl_183 vdd gnd cell_6t
Xbit_r184_c140 bl_140 br_140 wl_184 vdd gnd cell_6t
Xbit_r185_c140 bl_140 br_140 wl_185 vdd gnd cell_6t
Xbit_r186_c140 bl_140 br_140 wl_186 vdd gnd cell_6t
Xbit_r187_c140 bl_140 br_140 wl_187 vdd gnd cell_6t
Xbit_r188_c140 bl_140 br_140 wl_188 vdd gnd cell_6t
Xbit_r189_c140 bl_140 br_140 wl_189 vdd gnd cell_6t
Xbit_r190_c140 bl_140 br_140 wl_190 vdd gnd cell_6t
Xbit_r191_c140 bl_140 br_140 wl_191 vdd gnd cell_6t
Xbit_r192_c140 bl_140 br_140 wl_192 vdd gnd cell_6t
Xbit_r193_c140 bl_140 br_140 wl_193 vdd gnd cell_6t
Xbit_r194_c140 bl_140 br_140 wl_194 vdd gnd cell_6t
Xbit_r195_c140 bl_140 br_140 wl_195 vdd gnd cell_6t
Xbit_r196_c140 bl_140 br_140 wl_196 vdd gnd cell_6t
Xbit_r197_c140 bl_140 br_140 wl_197 vdd gnd cell_6t
Xbit_r198_c140 bl_140 br_140 wl_198 vdd gnd cell_6t
Xbit_r199_c140 bl_140 br_140 wl_199 vdd gnd cell_6t
Xbit_r200_c140 bl_140 br_140 wl_200 vdd gnd cell_6t
Xbit_r201_c140 bl_140 br_140 wl_201 vdd gnd cell_6t
Xbit_r202_c140 bl_140 br_140 wl_202 vdd gnd cell_6t
Xbit_r203_c140 bl_140 br_140 wl_203 vdd gnd cell_6t
Xbit_r204_c140 bl_140 br_140 wl_204 vdd gnd cell_6t
Xbit_r205_c140 bl_140 br_140 wl_205 vdd gnd cell_6t
Xbit_r206_c140 bl_140 br_140 wl_206 vdd gnd cell_6t
Xbit_r207_c140 bl_140 br_140 wl_207 vdd gnd cell_6t
Xbit_r208_c140 bl_140 br_140 wl_208 vdd gnd cell_6t
Xbit_r209_c140 bl_140 br_140 wl_209 vdd gnd cell_6t
Xbit_r210_c140 bl_140 br_140 wl_210 vdd gnd cell_6t
Xbit_r211_c140 bl_140 br_140 wl_211 vdd gnd cell_6t
Xbit_r212_c140 bl_140 br_140 wl_212 vdd gnd cell_6t
Xbit_r213_c140 bl_140 br_140 wl_213 vdd gnd cell_6t
Xbit_r214_c140 bl_140 br_140 wl_214 vdd gnd cell_6t
Xbit_r215_c140 bl_140 br_140 wl_215 vdd gnd cell_6t
Xbit_r216_c140 bl_140 br_140 wl_216 vdd gnd cell_6t
Xbit_r217_c140 bl_140 br_140 wl_217 vdd gnd cell_6t
Xbit_r218_c140 bl_140 br_140 wl_218 vdd gnd cell_6t
Xbit_r219_c140 bl_140 br_140 wl_219 vdd gnd cell_6t
Xbit_r220_c140 bl_140 br_140 wl_220 vdd gnd cell_6t
Xbit_r221_c140 bl_140 br_140 wl_221 vdd gnd cell_6t
Xbit_r222_c140 bl_140 br_140 wl_222 vdd gnd cell_6t
Xbit_r223_c140 bl_140 br_140 wl_223 vdd gnd cell_6t
Xbit_r224_c140 bl_140 br_140 wl_224 vdd gnd cell_6t
Xbit_r225_c140 bl_140 br_140 wl_225 vdd gnd cell_6t
Xbit_r226_c140 bl_140 br_140 wl_226 vdd gnd cell_6t
Xbit_r227_c140 bl_140 br_140 wl_227 vdd gnd cell_6t
Xbit_r228_c140 bl_140 br_140 wl_228 vdd gnd cell_6t
Xbit_r229_c140 bl_140 br_140 wl_229 vdd gnd cell_6t
Xbit_r230_c140 bl_140 br_140 wl_230 vdd gnd cell_6t
Xbit_r231_c140 bl_140 br_140 wl_231 vdd gnd cell_6t
Xbit_r232_c140 bl_140 br_140 wl_232 vdd gnd cell_6t
Xbit_r233_c140 bl_140 br_140 wl_233 vdd gnd cell_6t
Xbit_r234_c140 bl_140 br_140 wl_234 vdd gnd cell_6t
Xbit_r235_c140 bl_140 br_140 wl_235 vdd gnd cell_6t
Xbit_r236_c140 bl_140 br_140 wl_236 vdd gnd cell_6t
Xbit_r237_c140 bl_140 br_140 wl_237 vdd gnd cell_6t
Xbit_r238_c140 bl_140 br_140 wl_238 vdd gnd cell_6t
Xbit_r239_c140 bl_140 br_140 wl_239 vdd gnd cell_6t
Xbit_r240_c140 bl_140 br_140 wl_240 vdd gnd cell_6t
Xbit_r241_c140 bl_140 br_140 wl_241 vdd gnd cell_6t
Xbit_r242_c140 bl_140 br_140 wl_242 vdd gnd cell_6t
Xbit_r243_c140 bl_140 br_140 wl_243 vdd gnd cell_6t
Xbit_r244_c140 bl_140 br_140 wl_244 vdd gnd cell_6t
Xbit_r245_c140 bl_140 br_140 wl_245 vdd gnd cell_6t
Xbit_r246_c140 bl_140 br_140 wl_246 vdd gnd cell_6t
Xbit_r247_c140 bl_140 br_140 wl_247 vdd gnd cell_6t
Xbit_r248_c140 bl_140 br_140 wl_248 vdd gnd cell_6t
Xbit_r249_c140 bl_140 br_140 wl_249 vdd gnd cell_6t
Xbit_r250_c140 bl_140 br_140 wl_250 vdd gnd cell_6t
Xbit_r251_c140 bl_140 br_140 wl_251 vdd gnd cell_6t
Xbit_r252_c140 bl_140 br_140 wl_252 vdd gnd cell_6t
Xbit_r253_c140 bl_140 br_140 wl_253 vdd gnd cell_6t
Xbit_r254_c140 bl_140 br_140 wl_254 vdd gnd cell_6t
Xbit_r255_c140 bl_140 br_140 wl_255 vdd gnd cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd cell_6t
Xbit_r1_c141 bl_141 br_141 wl_1 vdd gnd cell_6t
Xbit_r2_c141 bl_141 br_141 wl_2 vdd gnd cell_6t
Xbit_r3_c141 bl_141 br_141 wl_3 vdd gnd cell_6t
Xbit_r4_c141 bl_141 br_141 wl_4 vdd gnd cell_6t
Xbit_r5_c141 bl_141 br_141 wl_5 vdd gnd cell_6t
Xbit_r6_c141 bl_141 br_141 wl_6 vdd gnd cell_6t
Xbit_r7_c141 bl_141 br_141 wl_7 vdd gnd cell_6t
Xbit_r8_c141 bl_141 br_141 wl_8 vdd gnd cell_6t
Xbit_r9_c141 bl_141 br_141 wl_9 vdd gnd cell_6t
Xbit_r10_c141 bl_141 br_141 wl_10 vdd gnd cell_6t
Xbit_r11_c141 bl_141 br_141 wl_11 vdd gnd cell_6t
Xbit_r12_c141 bl_141 br_141 wl_12 vdd gnd cell_6t
Xbit_r13_c141 bl_141 br_141 wl_13 vdd gnd cell_6t
Xbit_r14_c141 bl_141 br_141 wl_14 vdd gnd cell_6t
Xbit_r15_c141 bl_141 br_141 wl_15 vdd gnd cell_6t
Xbit_r16_c141 bl_141 br_141 wl_16 vdd gnd cell_6t
Xbit_r17_c141 bl_141 br_141 wl_17 vdd gnd cell_6t
Xbit_r18_c141 bl_141 br_141 wl_18 vdd gnd cell_6t
Xbit_r19_c141 bl_141 br_141 wl_19 vdd gnd cell_6t
Xbit_r20_c141 bl_141 br_141 wl_20 vdd gnd cell_6t
Xbit_r21_c141 bl_141 br_141 wl_21 vdd gnd cell_6t
Xbit_r22_c141 bl_141 br_141 wl_22 vdd gnd cell_6t
Xbit_r23_c141 bl_141 br_141 wl_23 vdd gnd cell_6t
Xbit_r24_c141 bl_141 br_141 wl_24 vdd gnd cell_6t
Xbit_r25_c141 bl_141 br_141 wl_25 vdd gnd cell_6t
Xbit_r26_c141 bl_141 br_141 wl_26 vdd gnd cell_6t
Xbit_r27_c141 bl_141 br_141 wl_27 vdd gnd cell_6t
Xbit_r28_c141 bl_141 br_141 wl_28 vdd gnd cell_6t
Xbit_r29_c141 bl_141 br_141 wl_29 vdd gnd cell_6t
Xbit_r30_c141 bl_141 br_141 wl_30 vdd gnd cell_6t
Xbit_r31_c141 bl_141 br_141 wl_31 vdd gnd cell_6t
Xbit_r32_c141 bl_141 br_141 wl_32 vdd gnd cell_6t
Xbit_r33_c141 bl_141 br_141 wl_33 vdd gnd cell_6t
Xbit_r34_c141 bl_141 br_141 wl_34 vdd gnd cell_6t
Xbit_r35_c141 bl_141 br_141 wl_35 vdd gnd cell_6t
Xbit_r36_c141 bl_141 br_141 wl_36 vdd gnd cell_6t
Xbit_r37_c141 bl_141 br_141 wl_37 vdd gnd cell_6t
Xbit_r38_c141 bl_141 br_141 wl_38 vdd gnd cell_6t
Xbit_r39_c141 bl_141 br_141 wl_39 vdd gnd cell_6t
Xbit_r40_c141 bl_141 br_141 wl_40 vdd gnd cell_6t
Xbit_r41_c141 bl_141 br_141 wl_41 vdd gnd cell_6t
Xbit_r42_c141 bl_141 br_141 wl_42 vdd gnd cell_6t
Xbit_r43_c141 bl_141 br_141 wl_43 vdd gnd cell_6t
Xbit_r44_c141 bl_141 br_141 wl_44 vdd gnd cell_6t
Xbit_r45_c141 bl_141 br_141 wl_45 vdd gnd cell_6t
Xbit_r46_c141 bl_141 br_141 wl_46 vdd gnd cell_6t
Xbit_r47_c141 bl_141 br_141 wl_47 vdd gnd cell_6t
Xbit_r48_c141 bl_141 br_141 wl_48 vdd gnd cell_6t
Xbit_r49_c141 bl_141 br_141 wl_49 vdd gnd cell_6t
Xbit_r50_c141 bl_141 br_141 wl_50 vdd gnd cell_6t
Xbit_r51_c141 bl_141 br_141 wl_51 vdd gnd cell_6t
Xbit_r52_c141 bl_141 br_141 wl_52 vdd gnd cell_6t
Xbit_r53_c141 bl_141 br_141 wl_53 vdd gnd cell_6t
Xbit_r54_c141 bl_141 br_141 wl_54 vdd gnd cell_6t
Xbit_r55_c141 bl_141 br_141 wl_55 vdd gnd cell_6t
Xbit_r56_c141 bl_141 br_141 wl_56 vdd gnd cell_6t
Xbit_r57_c141 bl_141 br_141 wl_57 vdd gnd cell_6t
Xbit_r58_c141 bl_141 br_141 wl_58 vdd gnd cell_6t
Xbit_r59_c141 bl_141 br_141 wl_59 vdd gnd cell_6t
Xbit_r60_c141 bl_141 br_141 wl_60 vdd gnd cell_6t
Xbit_r61_c141 bl_141 br_141 wl_61 vdd gnd cell_6t
Xbit_r62_c141 bl_141 br_141 wl_62 vdd gnd cell_6t
Xbit_r63_c141 bl_141 br_141 wl_63 vdd gnd cell_6t
Xbit_r64_c141 bl_141 br_141 wl_64 vdd gnd cell_6t
Xbit_r65_c141 bl_141 br_141 wl_65 vdd gnd cell_6t
Xbit_r66_c141 bl_141 br_141 wl_66 vdd gnd cell_6t
Xbit_r67_c141 bl_141 br_141 wl_67 vdd gnd cell_6t
Xbit_r68_c141 bl_141 br_141 wl_68 vdd gnd cell_6t
Xbit_r69_c141 bl_141 br_141 wl_69 vdd gnd cell_6t
Xbit_r70_c141 bl_141 br_141 wl_70 vdd gnd cell_6t
Xbit_r71_c141 bl_141 br_141 wl_71 vdd gnd cell_6t
Xbit_r72_c141 bl_141 br_141 wl_72 vdd gnd cell_6t
Xbit_r73_c141 bl_141 br_141 wl_73 vdd gnd cell_6t
Xbit_r74_c141 bl_141 br_141 wl_74 vdd gnd cell_6t
Xbit_r75_c141 bl_141 br_141 wl_75 vdd gnd cell_6t
Xbit_r76_c141 bl_141 br_141 wl_76 vdd gnd cell_6t
Xbit_r77_c141 bl_141 br_141 wl_77 vdd gnd cell_6t
Xbit_r78_c141 bl_141 br_141 wl_78 vdd gnd cell_6t
Xbit_r79_c141 bl_141 br_141 wl_79 vdd gnd cell_6t
Xbit_r80_c141 bl_141 br_141 wl_80 vdd gnd cell_6t
Xbit_r81_c141 bl_141 br_141 wl_81 vdd gnd cell_6t
Xbit_r82_c141 bl_141 br_141 wl_82 vdd gnd cell_6t
Xbit_r83_c141 bl_141 br_141 wl_83 vdd gnd cell_6t
Xbit_r84_c141 bl_141 br_141 wl_84 vdd gnd cell_6t
Xbit_r85_c141 bl_141 br_141 wl_85 vdd gnd cell_6t
Xbit_r86_c141 bl_141 br_141 wl_86 vdd gnd cell_6t
Xbit_r87_c141 bl_141 br_141 wl_87 vdd gnd cell_6t
Xbit_r88_c141 bl_141 br_141 wl_88 vdd gnd cell_6t
Xbit_r89_c141 bl_141 br_141 wl_89 vdd gnd cell_6t
Xbit_r90_c141 bl_141 br_141 wl_90 vdd gnd cell_6t
Xbit_r91_c141 bl_141 br_141 wl_91 vdd gnd cell_6t
Xbit_r92_c141 bl_141 br_141 wl_92 vdd gnd cell_6t
Xbit_r93_c141 bl_141 br_141 wl_93 vdd gnd cell_6t
Xbit_r94_c141 bl_141 br_141 wl_94 vdd gnd cell_6t
Xbit_r95_c141 bl_141 br_141 wl_95 vdd gnd cell_6t
Xbit_r96_c141 bl_141 br_141 wl_96 vdd gnd cell_6t
Xbit_r97_c141 bl_141 br_141 wl_97 vdd gnd cell_6t
Xbit_r98_c141 bl_141 br_141 wl_98 vdd gnd cell_6t
Xbit_r99_c141 bl_141 br_141 wl_99 vdd gnd cell_6t
Xbit_r100_c141 bl_141 br_141 wl_100 vdd gnd cell_6t
Xbit_r101_c141 bl_141 br_141 wl_101 vdd gnd cell_6t
Xbit_r102_c141 bl_141 br_141 wl_102 vdd gnd cell_6t
Xbit_r103_c141 bl_141 br_141 wl_103 vdd gnd cell_6t
Xbit_r104_c141 bl_141 br_141 wl_104 vdd gnd cell_6t
Xbit_r105_c141 bl_141 br_141 wl_105 vdd gnd cell_6t
Xbit_r106_c141 bl_141 br_141 wl_106 vdd gnd cell_6t
Xbit_r107_c141 bl_141 br_141 wl_107 vdd gnd cell_6t
Xbit_r108_c141 bl_141 br_141 wl_108 vdd gnd cell_6t
Xbit_r109_c141 bl_141 br_141 wl_109 vdd gnd cell_6t
Xbit_r110_c141 bl_141 br_141 wl_110 vdd gnd cell_6t
Xbit_r111_c141 bl_141 br_141 wl_111 vdd gnd cell_6t
Xbit_r112_c141 bl_141 br_141 wl_112 vdd gnd cell_6t
Xbit_r113_c141 bl_141 br_141 wl_113 vdd gnd cell_6t
Xbit_r114_c141 bl_141 br_141 wl_114 vdd gnd cell_6t
Xbit_r115_c141 bl_141 br_141 wl_115 vdd gnd cell_6t
Xbit_r116_c141 bl_141 br_141 wl_116 vdd gnd cell_6t
Xbit_r117_c141 bl_141 br_141 wl_117 vdd gnd cell_6t
Xbit_r118_c141 bl_141 br_141 wl_118 vdd gnd cell_6t
Xbit_r119_c141 bl_141 br_141 wl_119 vdd gnd cell_6t
Xbit_r120_c141 bl_141 br_141 wl_120 vdd gnd cell_6t
Xbit_r121_c141 bl_141 br_141 wl_121 vdd gnd cell_6t
Xbit_r122_c141 bl_141 br_141 wl_122 vdd gnd cell_6t
Xbit_r123_c141 bl_141 br_141 wl_123 vdd gnd cell_6t
Xbit_r124_c141 bl_141 br_141 wl_124 vdd gnd cell_6t
Xbit_r125_c141 bl_141 br_141 wl_125 vdd gnd cell_6t
Xbit_r126_c141 bl_141 br_141 wl_126 vdd gnd cell_6t
Xbit_r127_c141 bl_141 br_141 wl_127 vdd gnd cell_6t
Xbit_r128_c141 bl_141 br_141 wl_128 vdd gnd cell_6t
Xbit_r129_c141 bl_141 br_141 wl_129 vdd gnd cell_6t
Xbit_r130_c141 bl_141 br_141 wl_130 vdd gnd cell_6t
Xbit_r131_c141 bl_141 br_141 wl_131 vdd gnd cell_6t
Xbit_r132_c141 bl_141 br_141 wl_132 vdd gnd cell_6t
Xbit_r133_c141 bl_141 br_141 wl_133 vdd gnd cell_6t
Xbit_r134_c141 bl_141 br_141 wl_134 vdd gnd cell_6t
Xbit_r135_c141 bl_141 br_141 wl_135 vdd gnd cell_6t
Xbit_r136_c141 bl_141 br_141 wl_136 vdd gnd cell_6t
Xbit_r137_c141 bl_141 br_141 wl_137 vdd gnd cell_6t
Xbit_r138_c141 bl_141 br_141 wl_138 vdd gnd cell_6t
Xbit_r139_c141 bl_141 br_141 wl_139 vdd gnd cell_6t
Xbit_r140_c141 bl_141 br_141 wl_140 vdd gnd cell_6t
Xbit_r141_c141 bl_141 br_141 wl_141 vdd gnd cell_6t
Xbit_r142_c141 bl_141 br_141 wl_142 vdd gnd cell_6t
Xbit_r143_c141 bl_141 br_141 wl_143 vdd gnd cell_6t
Xbit_r144_c141 bl_141 br_141 wl_144 vdd gnd cell_6t
Xbit_r145_c141 bl_141 br_141 wl_145 vdd gnd cell_6t
Xbit_r146_c141 bl_141 br_141 wl_146 vdd gnd cell_6t
Xbit_r147_c141 bl_141 br_141 wl_147 vdd gnd cell_6t
Xbit_r148_c141 bl_141 br_141 wl_148 vdd gnd cell_6t
Xbit_r149_c141 bl_141 br_141 wl_149 vdd gnd cell_6t
Xbit_r150_c141 bl_141 br_141 wl_150 vdd gnd cell_6t
Xbit_r151_c141 bl_141 br_141 wl_151 vdd gnd cell_6t
Xbit_r152_c141 bl_141 br_141 wl_152 vdd gnd cell_6t
Xbit_r153_c141 bl_141 br_141 wl_153 vdd gnd cell_6t
Xbit_r154_c141 bl_141 br_141 wl_154 vdd gnd cell_6t
Xbit_r155_c141 bl_141 br_141 wl_155 vdd gnd cell_6t
Xbit_r156_c141 bl_141 br_141 wl_156 vdd gnd cell_6t
Xbit_r157_c141 bl_141 br_141 wl_157 vdd gnd cell_6t
Xbit_r158_c141 bl_141 br_141 wl_158 vdd gnd cell_6t
Xbit_r159_c141 bl_141 br_141 wl_159 vdd gnd cell_6t
Xbit_r160_c141 bl_141 br_141 wl_160 vdd gnd cell_6t
Xbit_r161_c141 bl_141 br_141 wl_161 vdd gnd cell_6t
Xbit_r162_c141 bl_141 br_141 wl_162 vdd gnd cell_6t
Xbit_r163_c141 bl_141 br_141 wl_163 vdd gnd cell_6t
Xbit_r164_c141 bl_141 br_141 wl_164 vdd gnd cell_6t
Xbit_r165_c141 bl_141 br_141 wl_165 vdd gnd cell_6t
Xbit_r166_c141 bl_141 br_141 wl_166 vdd gnd cell_6t
Xbit_r167_c141 bl_141 br_141 wl_167 vdd gnd cell_6t
Xbit_r168_c141 bl_141 br_141 wl_168 vdd gnd cell_6t
Xbit_r169_c141 bl_141 br_141 wl_169 vdd gnd cell_6t
Xbit_r170_c141 bl_141 br_141 wl_170 vdd gnd cell_6t
Xbit_r171_c141 bl_141 br_141 wl_171 vdd gnd cell_6t
Xbit_r172_c141 bl_141 br_141 wl_172 vdd gnd cell_6t
Xbit_r173_c141 bl_141 br_141 wl_173 vdd gnd cell_6t
Xbit_r174_c141 bl_141 br_141 wl_174 vdd gnd cell_6t
Xbit_r175_c141 bl_141 br_141 wl_175 vdd gnd cell_6t
Xbit_r176_c141 bl_141 br_141 wl_176 vdd gnd cell_6t
Xbit_r177_c141 bl_141 br_141 wl_177 vdd gnd cell_6t
Xbit_r178_c141 bl_141 br_141 wl_178 vdd gnd cell_6t
Xbit_r179_c141 bl_141 br_141 wl_179 vdd gnd cell_6t
Xbit_r180_c141 bl_141 br_141 wl_180 vdd gnd cell_6t
Xbit_r181_c141 bl_141 br_141 wl_181 vdd gnd cell_6t
Xbit_r182_c141 bl_141 br_141 wl_182 vdd gnd cell_6t
Xbit_r183_c141 bl_141 br_141 wl_183 vdd gnd cell_6t
Xbit_r184_c141 bl_141 br_141 wl_184 vdd gnd cell_6t
Xbit_r185_c141 bl_141 br_141 wl_185 vdd gnd cell_6t
Xbit_r186_c141 bl_141 br_141 wl_186 vdd gnd cell_6t
Xbit_r187_c141 bl_141 br_141 wl_187 vdd gnd cell_6t
Xbit_r188_c141 bl_141 br_141 wl_188 vdd gnd cell_6t
Xbit_r189_c141 bl_141 br_141 wl_189 vdd gnd cell_6t
Xbit_r190_c141 bl_141 br_141 wl_190 vdd gnd cell_6t
Xbit_r191_c141 bl_141 br_141 wl_191 vdd gnd cell_6t
Xbit_r192_c141 bl_141 br_141 wl_192 vdd gnd cell_6t
Xbit_r193_c141 bl_141 br_141 wl_193 vdd gnd cell_6t
Xbit_r194_c141 bl_141 br_141 wl_194 vdd gnd cell_6t
Xbit_r195_c141 bl_141 br_141 wl_195 vdd gnd cell_6t
Xbit_r196_c141 bl_141 br_141 wl_196 vdd gnd cell_6t
Xbit_r197_c141 bl_141 br_141 wl_197 vdd gnd cell_6t
Xbit_r198_c141 bl_141 br_141 wl_198 vdd gnd cell_6t
Xbit_r199_c141 bl_141 br_141 wl_199 vdd gnd cell_6t
Xbit_r200_c141 bl_141 br_141 wl_200 vdd gnd cell_6t
Xbit_r201_c141 bl_141 br_141 wl_201 vdd gnd cell_6t
Xbit_r202_c141 bl_141 br_141 wl_202 vdd gnd cell_6t
Xbit_r203_c141 bl_141 br_141 wl_203 vdd gnd cell_6t
Xbit_r204_c141 bl_141 br_141 wl_204 vdd gnd cell_6t
Xbit_r205_c141 bl_141 br_141 wl_205 vdd gnd cell_6t
Xbit_r206_c141 bl_141 br_141 wl_206 vdd gnd cell_6t
Xbit_r207_c141 bl_141 br_141 wl_207 vdd gnd cell_6t
Xbit_r208_c141 bl_141 br_141 wl_208 vdd gnd cell_6t
Xbit_r209_c141 bl_141 br_141 wl_209 vdd gnd cell_6t
Xbit_r210_c141 bl_141 br_141 wl_210 vdd gnd cell_6t
Xbit_r211_c141 bl_141 br_141 wl_211 vdd gnd cell_6t
Xbit_r212_c141 bl_141 br_141 wl_212 vdd gnd cell_6t
Xbit_r213_c141 bl_141 br_141 wl_213 vdd gnd cell_6t
Xbit_r214_c141 bl_141 br_141 wl_214 vdd gnd cell_6t
Xbit_r215_c141 bl_141 br_141 wl_215 vdd gnd cell_6t
Xbit_r216_c141 bl_141 br_141 wl_216 vdd gnd cell_6t
Xbit_r217_c141 bl_141 br_141 wl_217 vdd gnd cell_6t
Xbit_r218_c141 bl_141 br_141 wl_218 vdd gnd cell_6t
Xbit_r219_c141 bl_141 br_141 wl_219 vdd gnd cell_6t
Xbit_r220_c141 bl_141 br_141 wl_220 vdd gnd cell_6t
Xbit_r221_c141 bl_141 br_141 wl_221 vdd gnd cell_6t
Xbit_r222_c141 bl_141 br_141 wl_222 vdd gnd cell_6t
Xbit_r223_c141 bl_141 br_141 wl_223 vdd gnd cell_6t
Xbit_r224_c141 bl_141 br_141 wl_224 vdd gnd cell_6t
Xbit_r225_c141 bl_141 br_141 wl_225 vdd gnd cell_6t
Xbit_r226_c141 bl_141 br_141 wl_226 vdd gnd cell_6t
Xbit_r227_c141 bl_141 br_141 wl_227 vdd gnd cell_6t
Xbit_r228_c141 bl_141 br_141 wl_228 vdd gnd cell_6t
Xbit_r229_c141 bl_141 br_141 wl_229 vdd gnd cell_6t
Xbit_r230_c141 bl_141 br_141 wl_230 vdd gnd cell_6t
Xbit_r231_c141 bl_141 br_141 wl_231 vdd gnd cell_6t
Xbit_r232_c141 bl_141 br_141 wl_232 vdd gnd cell_6t
Xbit_r233_c141 bl_141 br_141 wl_233 vdd gnd cell_6t
Xbit_r234_c141 bl_141 br_141 wl_234 vdd gnd cell_6t
Xbit_r235_c141 bl_141 br_141 wl_235 vdd gnd cell_6t
Xbit_r236_c141 bl_141 br_141 wl_236 vdd gnd cell_6t
Xbit_r237_c141 bl_141 br_141 wl_237 vdd gnd cell_6t
Xbit_r238_c141 bl_141 br_141 wl_238 vdd gnd cell_6t
Xbit_r239_c141 bl_141 br_141 wl_239 vdd gnd cell_6t
Xbit_r240_c141 bl_141 br_141 wl_240 vdd gnd cell_6t
Xbit_r241_c141 bl_141 br_141 wl_241 vdd gnd cell_6t
Xbit_r242_c141 bl_141 br_141 wl_242 vdd gnd cell_6t
Xbit_r243_c141 bl_141 br_141 wl_243 vdd gnd cell_6t
Xbit_r244_c141 bl_141 br_141 wl_244 vdd gnd cell_6t
Xbit_r245_c141 bl_141 br_141 wl_245 vdd gnd cell_6t
Xbit_r246_c141 bl_141 br_141 wl_246 vdd gnd cell_6t
Xbit_r247_c141 bl_141 br_141 wl_247 vdd gnd cell_6t
Xbit_r248_c141 bl_141 br_141 wl_248 vdd gnd cell_6t
Xbit_r249_c141 bl_141 br_141 wl_249 vdd gnd cell_6t
Xbit_r250_c141 bl_141 br_141 wl_250 vdd gnd cell_6t
Xbit_r251_c141 bl_141 br_141 wl_251 vdd gnd cell_6t
Xbit_r252_c141 bl_141 br_141 wl_252 vdd gnd cell_6t
Xbit_r253_c141 bl_141 br_141 wl_253 vdd gnd cell_6t
Xbit_r254_c141 bl_141 br_141 wl_254 vdd gnd cell_6t
Xbit_r255_c141 bl_141 br_141 wl_255 vdd gnd cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd cell_6t
Xbit_r1_c142 bl_142 br_142 wl_1 vdd gnd cell_6t
Xbit_r2_c142 bl_142 br_142 wl_2 vdd gnd cell_6t
Xbit_r3_c142 bl_142 br_142 wl_3 vdd gnd cell_6t
Xbit_r4_c142 bl_142 br_142 wl_4 vdd gnd cell_6t
Xbit_r5_c142 bl_142 br_142 wl_5 vdd gnd cell_6t
Xbit_r6_c142 bl_142 br_142 wl_6 vdd gnd cell_6t
Xbit_r7_c142 bl_142 br_142 wl_7 vdd gnd cell_6t
Xbit_r8_c142 bl_142 br_142 wl_8 vdd gnd cell_6t
Xbit_r9_c142 bl_142 br_142 wl_9 vdd gnd cell_6t
Xbit_r10_c142 bl_142 br_142 wl_10 vdd gnd cell_6t
Xbit_r11_c142 bl_142 br_142 wl_11 vdd gnd cell_6t
Xbit_r12_c142 bl_142 br_142 wl_12 vdd gnd cell_6t
Xbit_r13_c142 bl_142 br_142 wl_13 vdd gnd cell_6t
Xbit_r14_c142 bl_142 br_142 wl_14 vdd gnd cell_6t
Xbit_r15_c142 bl_142 br_142 wl_15 vdd gnd cell_6t
Xbit_r16_c142 bl_142 br_142 wl_16 vdd gnd cell_6t
Xbit_r17_c142 bl_142 br_142 wl_17 vdd gnd cell_6t
Xbit_r18_c142 bl_142 br_142 wl_18 vdd gnd cell_6t
Xbit_r19_c142 bl_142 br_142 wl_19 vdd gnd cell_6t
Xbit_r20_c142 bl_142 br_142 wl_20 vdd gnd cell_6t
Xbit_r21_c142 bl_142 br_142 wl_21 vdd gnd cell_6t
Xbit_r22_c142 bl_142 br_142 wl_22 vdd gnd cell_6t
Xbit_r23_c142 bl_142 br_142 wl_23 vdd gnd cell_6t
Xbit_r24_c142 bl_142 br_142 wl_24 vdd gnd cell_6t
Xbit_r25_c142 bl_142 br_142 wl_25 vdd gnd cell_6t
Xbit_r26_c142 bl_142 br_142 wl_26 vdd gnd cell_6t
Xbit_r27_c142 bl_142 br_142 wl_27 vdd gnd cell_6t
Xbit_r28_c142 bl_142 br_142 wl_28 vdd gnd cell_6t
Xbit_r29_c142 bl_142 br_142 wl_29 vdd gnd cell_6t
Xbit_r30_c142 bl_142 br_142 wl_30 vdd gnd cell_6t
Xbit_r31_c142 bl_142 br_142 wl_31 vdd gnd cell_6t
Xbit_r32_c142 bl_142 br_142 wl_32 vdd gnd cell_6t
Xbit_r33_c142 bl_142 br_142 wl_33 vdd gnd cell_6t
Xbit_r34_c142 bl_142 br_142 wl_34 vdd gnd cell_6t
Xbit_r35_c142 bl_142 br_142 wl_35 vdd gnd cell_6t
Xbit_r36_c142 bl_142 br_142 wl_36 vdd gnd cell_6t
Xbit_r37_c142 bl_142 br_142 wl_37 vdd gnd cell_6t
Xbit_r38_c142 bl_142 br_142 wl_38 vdd gnd cell_6t
Xbit_r39_c142 bl_142 br_142 wl_39 vdd gnd cell_6t
Xbit_r40_c142 bl_142 br_142 wl_40 vdd gnd cell_6t
Xbit_r41_c142 bl_142 br_142 wl_41 vdd gnd cell_6t
Xbit_r42_c142 bl_142 br_142 wl_42 vdd gnd cell_6t
Xbit_r43_c142 bl_142 br_142 wl_43 vdd gnd cell_6t
Xbit_r44_c142 bl_142 br_142 wl_44 vdd gnd cell_6t
Xbit_r45_c142 bl_142 br_142 wl_45 vdd gnd cell_6t
Xbit_r46_c142 bl_142 br_142 wl_46 vdd gnd cell_6t
Xbit_r47_c142 bl_142 br_142 wl_47 vdd gnd cell_6t
Xbit_r48_c142 bl_142 br_142 wl_48 vdd gnd cell_6t
Xbit_r49_c142 bl_142 br_142 wl_49 vdd gnd cell_6t
Xbit_r50_c142 bl_142 br_142 wl_50 vdd gnd cell_6t
Xbit_r51_c142 bl_142 br_142 wl_51 vdd gnd cell_6t
Xbit_r52_c142 bl_142 br_142 wl_52 vdd gnd cell_6t
Xbit_r53_c142 bl_142 br_142 wl_53 vdd gnd cell_6t
Xbit_r54_c142 bl_142 br_142 wl_54 vdd gnd cell_6t
Xbit_r55_c142 bl_142 br_142 wl_55 vdd gnd cell_6t
Xbit_r56_c142 bl_142 br_142 wl_56 vdd gnd cell_6t
Xbit_r57_c142 bl_142 br_142 wl_57 vdd gnd cell_6t
Xbit_r58_c142 bl_142 br_142 wl_58 vdd gnd cell_6t
Xbit_r59_c142 bl_142 br_142 wl_59 vdd gnd cell_6t
Xbit_r60_c142 bl_142 br_142 wl_60 vdd gnd cell_6t
Xbit_r61_c142 bl_142 br_142 wl_61 vdd gnd cell_6t
Xbit_r62_c142 bl_142 br_142 wl_62 vdd gnd cell_6t
Xbit_r63_c142 bl_142 br_142 wl_63 vdd gnd cell_6t
Xbit_r64_c142 bl_142 br_142 wl_64 vdd gnd cell_6t
Xbit_r65_c142 bl_142 br_142 wl_65 vdd gnd cell_6t
Xbit_r66_c142 bl_142 br_142 wl_66 vdd gnd cell_6t
Xbit_r67_c142 bl_142 br_142 wl_67 vdd gnd cell_6t
Xbit_r68_c142 bl_142 br_142 wl_68 vdd gnd cell_6t
Xbit_r69_c142 bl_142 br_142 wl_69 vdd gnd cell_6t
Xbit_r70_c142 bl_142 br_142 wl_70 vdd gnd cell_6t
Xbit_r71_c142 bl_142 br_142 wl_71 vdd gnd cell_6t
Xbit_r72_c142 bl_142 br_142 wl_72 vdd gnd cell_6t
Xbit_r73_c142 bl_142 br_142 wl_73 vdd gnd cell_6t
Xbit_r74_c142 bl_142 br_142 wl_74 vdd gnd cell_6t
Xbit_r75_c142 bl_142 br_142 wl_75 vdd gnd cell_6t
Xbit_r76_c142 bl_142 br_142 wl_76 vdd gnd cell_6t
Xbit_r77_c142 bl_142 br_142 wl_77 vdd gnd cell_6t
Xbit_r78_c142 bl_142 br_142 wl_78 vdd gnd cell_6t
Xbit_r79_c142 bl_142 br_142 wl_79 vdd gnd cell_6t
Xbit_r80_c142 bl_142 br_142 wl_80 vdd gnd cell_6t
Xbit_r81_c142 bl_142 br_142 wl_81 vdd gnd cell_6t
Xbit_r82_c142 bl_142 br_142 wl_82 vdd gnd cell_6t
Xbit_r83_c142 bl_142 br_142 wl_83 vdd gnd cell_6t
Xbit_r84_c142 bl_142 br_142 wl_84 vdd gnd cell_6t
Xbit_r85_c142 bl_142 br_142 wl_85 vdd gnd cell_6t
Xbit_r86_c142 bl_142 br_142 wl_86 vdd gnd cell_6t
Xbit_r87_c142 bl_142 br_142 wl_87 vdd gnd cell_6t
Xbit_r88_c142 bl_142 br_142 wl_88 vdd gnd cell_6t
Xbit_r89_c142 bl_142 br_142 wl_89 vdd gnd cell_6t
Xbit_r90_c142 bl_142 br_142 wl_90 vdd gnd cell_6t
Xbit_r91_c142 bl_142 br_142 wl_91 vdd gnd cell_6t
Xbit_r92_c142 bl_142 br_142 wl_92 vdd gnd cell_6t
Xbit_r93_c142 bl_142 br_142 wl_93 vdd gnd cell_6t
Xbit_r94_c142 bl_142 br_142 wl_94 vdd gnd cell_6t
Xbit_r95_c142 bl_142 br_142 wl_95 vdd gnd cell_6t
Xbit_r96_c142 bl_142 br_142 wl_96 vdd gnd cell_6t
Xbit_r97_c142 bl_142 br_142 wl_97 vdd gnd cell_6t
Xbit_r98_c142 bl_142 br_142 wl_98 vdd gnd cell_6t
Xbit_r99_c142 bl_142 br_142 wl_99 vdd gnd cell_6t
Xbit_r100_c142 bl_142 br_142 wl_100 vdd gnd cell_6t
Xbit_r101_c142 bl_142 br_142 wl_101 vdd gnd cell_6t
Xbit_r102_c142 bl_142 br_142 wl_102 vdd gnd cell_6t
Xbit_r103_c142 bl_142 br_142 wl_103 vdd gnd cell_6t
Xbit_r104_c142 bl_142 br_142 wl_104 vdd gnd cell_6t
Xbit_r105_c142 bl_142 br_142 wl_105 vdd gnd cell_6t
Xbit_r106_c142 bl_142 br_142 wl_106 vdd gnd cell_6t
Xbit_r107_c142 bl_142 br_142 wl_107 vdd gnd cell_6t
Xbit_r108_c142 bl_142 br_142 wl_108 vdd gnd cell_6t
Xbit_r109_c142 bl_142 br_142 wl_109 vdd gnd cell_6t
Xbit_r110_c142 bl_142 br_142 wl_110 vdd gnd cell_6t
Xbit_r111_c142 bl_142 br_142 wl_111 vdd gnd cell_6t
Xbit_r112_c142 bl_142 br_142 wl_112 vdd gnd cell_6t
Xbit_r113_c142 bl_142 br_142 wl_113 vdd gnd cell_6t
Xbit_r114_c142 bl_142 br_142 wl_114 vdd gnd cell_6t
Xbit_r115_c142 bl_142 br_142 wl_115 vdd gnd cell_6t
Xbit_r116_c142 bl_142 br_142 wl_116 vdd gnd cell_6t
Xbit_r117_c142 bl_142 br_142 wl_117 vdd gnd cell_6t
Xbit_r118_c142 bl_142 br_142 wl_118 vdd gnd cell_6t
Xbit_r119_c142 bl_142 br_142 wl_119 vdd gnd cell_6t
Xbit_r120_c142 bl_142 br_142 wl_120 vdd gnd cell_6t
Xbit_r121_c142 bl_142 br_142 wl_121 vdd gnd cell_6t
Xbit_r122_c142 bl_142 br_142 wl_122 vdd gnd cell_6t
Xbit_r123_c142 bl_142 br_142 wl_123 vdd gnd cell_6t
Xbit_r124_c142 bl_142 br_142 wl_124 vdd gnd cell_6t
Xbit_r125_c142 bl_142 br_142 wl_125 vdd gnd cell_6t
Xbit_r126_c142 bl_142 br_142 wl_126 vdd gnd cell_6t
Xbit_r127_c142 bl_142 br_142 wl_127 vdd gnd cell_6t
Xbit_r128_c142 bl_142 br_142 wl_128 vdd gnd cell_6t
Xbit_r129_c142 bl_142 br_142 wl_129 vdd gnd cell_6t
Xbit_r130_c142 bl_142 br_142 wl_130 vdd gnd cell_6t
Xbit_r131_c142 bl_142 br_142 wl_131 vdd gnd cell_6t
Xbit_r132_c142 bl_142 br_142 wl_132 vdd gnd cell_6t
Xbit_r133_c142 bl_142 br_142 wl_133 vdd gnd cell_6t
Xbit_r134_c142 bl_142 br_142 wl_134 vdd gnd cell_6t
Xbit_r135_c142 bl_142 br_142 wl_135 vdd gnd cell_6t
Xbit_r136_c142 bl_142 br_142 wl_136 vdd gnd cell_6t
Xbit_r137_c142 bl_142 br_142 wl_137 vdd gnd cell_6t
Xbit_r138_c142 bl_142 br_142 wl_138 vdd gnd cell_6t
Xbit_r139_c142 bl_142 br_142 wl_139 vdd gnd cell_6t
Xbit_r140_c142 bl_142 br_142 wl_140 vdd gnd cell_6t
Xbit_r141_c142 bl_142 br_142 wl_141 vdd gnd cell_6t
Xbit_r142_c142 bl_142 br_142 wl_142 vdd gnd cell_6t
Xbit_r143_c142 bl_142 br_142 wl_143 vdd gnd cell_6t
Xbit_r144_c142 bl_142 br_142 wl_144 vdd gnd cell_6t
Xbit_r145_c142 bl_142 br_142 wl_145 vdd gnd cell_6t
Xbit_r146_c142 bl_142 br_142 wl_146 vdd gnd cell_6t
Xbit_r147_c142 bl_142 br_142 wl_147 vdd gnd cell_6t
Xbit_r148_c142 bl_142 br_142 wl_148 vdd gnd cell_6t
Xbit_r149_c142 bl_142 br_142 wl_149 vdd gnd cell_6t
Xbit_r150_c142 bl_142 br_142 wl_150 vdd gnd cell_6t
Xbit_r151_c142 bl_142 br_142 wl_151 vdd gnd cell_6t
Xbit_r152_c142 bl_142 br_142 wl_152 vdd gnd cell_6t
Xbit_r153_c142 bl_142 br_142 wl_153 vdd gnd cell_6t
Xbit_r154_c142 bl_142 br_142 wl_154 vdd gnd cell_6t
Xbit_r155_c142 bl_142 br_142 wl_155 vdd gnd cell_6t
Xbit_r156_c142 bl_142 br_142 wl_156 vdd gnd cell_6t
Xbit_r157_c142 bl_142 br_142 wl_157 vdd gnd cell_6t
Xbit_r158_c142 bl_142 br_142 wl_158 vdd gnd cell_6t
Xbit_r159_c142 bl_142 br_142 wl_159 vdd gnd cell_6t
Xbit_r160_c142 bl_142 br_142 wl_160 vdd gnd cell_6t
Xbit_r161_c142 bl_142 br_142 wl_161 vdd gnd cell_6t
Xbit_r162_c142 bl_142 br_142 wl_162 vdd gnd cell_6t
Xbit_r163_c142 bl_142 br_142 wl_163 vdd gnd cell_6t
Xbit_r164_c142 bl_142 br_142 wl_164 vdd gnd cell_6t
Xbit_r165_c142 bl_142 br_142 wl_165 vdd gnd cell_6t
Xbit_r166_c142 bl_142 br_142 wl_166 vdd gnd cell_6t
Xbit_r167_c142 bl_142 br_142 wl_167 vdd gnd cell_6t
Xbit_r168_c142 bl_142 br_142 wl_168 vdd gnd cell_6t
Xbit_r169_c142 bl_142 br_142 wl_169 vdd gnd cell_6t
Xbit_r170_c142 bl_142 br_142 wl_170 vdd gnd cell_6t
Xbit_r171_c142 bl_142 br_142 wl_171 vdd gnd cell_6t
Xbit_r172_c142 bl_142 br_142 wl_172 vdd gnd cell_6t
Xbit_r173_c142 bl_142 br_142 wl_173 vdd gnd cell_6t
Xbit_r174_c142 bl_142 br_142 wl_174 vdd gnd cell_6t
Xbit_r175_c142 bl_142 br_142 wl_175 vdd gnd cell_6t
Xbit_r176_c142 bl_142 br_142 wl_176 vdd gnd cell_6t
Xbit_r177_c142 bl_142 br_142 wl_177 vdd gnd cell_6t
Xbit_r178_c142 bl_142 br_142 wl_178 vdd gnd cell_6t
Xbit_r179_c142 bl_142 br_142 wl_179 vdd gnd cell_6t
Xbit_r180_c142 bl_142 br_142 wl_180 vdd gnd cell_6t
Xbit_r181_c142 bl_142 br_142 wl_181 vdd gnd cell_6t
Xbit_r182_c142 bl_142 br_142 wl_182 vdd gnd cell_6t
Xbit_r183_c142 bl_142 br_142 wl_183 vdd gnd cell_6t
Xbit_r184_c142 bl_142 br_142 wl_184 vdd gnd cell_6t
Xbit_r185_c142 bl_142 br_142 wl_185 vdd gnd cell_6t
Xbit_r186_c142 bl_142 br_142 wl_186 vdd gnd cell_6t
Xbit_r187_c142 bl_142 br_142 wl_187 vdd gnd cell_6t
Xbit_r188_c142 bl_142 br_142 wl_188 vdd gnd cell_6t
Xbit_r189_c142 bl_142 br_142 wl_189 vdd gnd cell_6t
Xbit_r190_c142 bl_142 br_142 wl_190 vdd gnd cell_6t
Xbit_r191_c142 bl_142 br_142 wl_191 vdd gnd cell_6t
Xbit_r192_c142 bl_142 br_142 wl_192 vdd gnd cell_6t
Xbit_r193_c142 bl_142 br_142 wl_193 vdd gnd cell_6t
Xbit_r194_c142 bl_142 br_142 wl_194 vdd gnd cell_6t
Xbit_r195_c142 bl_142 br_142 wl_195 vdd gnd cell_6t
Xbit_r196_c142 bl_142 br_142 wl_196 vdd gnd cell_6t
Xbit_r197_c142 bl_142 br_142 wl_197 vdd gnd cell_6t
Xbit_r198_c142 bl_142 br_142 wl_198 vdd gnd cell_6t
Xbit_r199_c142 bl_142 br_142 wl_199 vdd gnd cell_6t
Xbit_r200_c142 bl_142 br_142 wl_200 vdd gnd cell_6t
Xbit_r201_c142 bl_142 br_142 wl_201 vdd gnd cell_6t
Xbit_r202_c142 bl_142 br_142 wl_202 vdd gnd cell_6t
Xbit_r203_c142 bl_142 br_142 wl_203 vdd gnd cell_6t
Xbit_r204_c142 bl_142 br_142 wl_204 vdd gnd cell_6t
Xbit_r205_c142 bl_142 br_142 wl_205 vdd gnd cell_6t
Xbit_r206_c142 bl_142 br_142 wl_206 vdd gnd cell_6t
Xbit_r207_c142 bl_142 br_142 wl_207 vdd gnd cell_6t
Xbit_r208_c142 bl_142 br_142 wl_208 vdd gnd cell_6t
Xbit_r209_c142 bl_142 br_142 wl_209 vdd gnd cell_6t
Xbit_r210_c142 bl_142 br_142 wl_210 vdd gnd cell_6t
Xbit_r211_c142 bl_142 br_142 wl_211 vdd gnd cell_6t
Xbit_r212_c142 bl_142 br_142 wl_212 vdd gnd cell_6t
Xbit_r213_c142 bl_142 br_142 wl_213 vdd gnd cell_6t
Xbit_r214_c142 bl_142 br_142 wl_214 vdd gnd cell_6t
Xbit_r215_c142 bl_142 br_142 wl_215 vdd gnd cell_6t
Xbit_r216_c142 bl_142 br_142 wl_216 vdd gnd cell_6t
Xbit_r217_c142 bl_142 br_142 wl_217 vdd gnd cell_6t
Xbit_r218_c142 bl_142 br_142 wl_218 vdd gnd cell_6t
Xbit_r219_c142 bl_142 br_142 wl_219 vdd gnd cell_6t
Xbit_r220_c142 bl_142 br_142 wl_220 vdd gnd cell_6t
Xbit_r221_c142 bl_142 br_142 wl_221 vdd gnd cell_6t
Xbit_r222_c142 bl_142 br_142 wl_222 vdd gnd cell_6t
Xbit_r223_c142 bl_142 br_142 wl_223 vdd gnd cell_6t
Xbit_r224_c142 bl_142 br_142 wl_224 vdd gnd cell_6t
Xbit_r225_c142 bl_142 br_142 wl_225 vdd gnd cell_6t
Xbit_r226_c142 bl_142 br_142 wl_226 vdd gnd cell_6t
Xbit_r227_c142 bl_142 br_142 wl_227 vdd gnd cell_6t
Xbit_r228_c142 bl_142 br_142 wl_228 vdd gnd cell_6t
Xbit_r229_c142 bl_142 br_142 wl_229 vdd gnd cell_6t
Xbit_r230_c142 bl_142 br_142 wl_230 vdd gnd cell_6t
Xbit_r231_c142 bl_142 br_142 wl_231 vdd gnd cell_6t
Xbit_r232_c142 bl_142 br_142 wl_232 vdd gnd cell_6t
Xbit_r233_c142 bl_142 br_142 wl_233 vdd gnd cell_6t
Xbit_r234_c142 bl_142 br_142 wl_234 vdd gnd cell_6t
Xbit_r235_c142 bl_142 br_142 wl_235 vdd gnd cell_6t
Xbit_r236_c142 bl_142 br_142 wl_236 vdd gnd cell_6t
Xbit_r237_c142 bl_142 br_142 wl_237 vdd gnd cell_6t
Xbit_r238_c142 bl_142 br_142 wl_238 vdd gnd cell_6t
Xbit_r239_c142 bl_142 br_142 wl_239 vdd gnd cell_6t
Xbit_r240_c142 bl_142 br_142 wl_240 vdd gnd cell_6t
Xbit_r241_c142 bl_142 br_142 wl_241 vdd gnd cell_6t
Xbit_r242_c142 bl_142 br_142 wl_242 vdd gnd cell_6t
Xbit_r243_c142 bl_142 br_142 wl_243 vdd gnd cell_6t
Xbit_r244_c142 bl_142 br_142 wl_244 vdd gnd cell_6t
Xbit_r245_c142 bl_142 br_142 wl_245 vdd gnd cell_6t
Xbit_r246_c142 bl_142 br_142 wl_246 vdd gnd cell_6t
Xbit_r247_c142 bl_142 br_142 wl_247 vdd gnd cell_6t
Xbit_r248_c142 bl_142 br_142 wl_248 vdd gnd cell_6t
Xbit_r249_c142 bl_142 br_142 wl_249 vdd gnd cell_6t
Xbit_r250_c142 bl_142 br_142 wl_250 vdd gnd cell_6t
Xbit_r251_c142 bl_142 br_142 wl_251 vdd gnd cell_6t
Xbit_r252_c142 bl_142 br_142 wl_252 vdd gnd cell_6t
Xbit_r253_c142 bl_142 br_142 wl_253 vdd gnd cell_6t
Xbit_r254_c142 bl_142 br_142 wl_254 vdd gnd cell_6t
Xbit_r255_c142 bl_142 br_142 wl_255 vdd gnd cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd cell_6t
Xbit_r1_c143 bl_143 br_143 wl_1 vdd gnd cell_6t
Xbit_r2_c143 bl_143 br_143 wl_2 vdd gnd cell_6t
Xbit_r3_c143 bl_143 br_143 wl_3 vdd gnd cell_6t
Xbit_r4_c143 bl_143 br_143 wl_4 vdd gnd cell_6t
Xbit_r5_c143 bl_143 br_143 wl_5 vdd gnd cell_6t
Xbit_r6_c143 bl_143 br_143 wl_6 vdd gnd cell_6t
Xbit_r7_c143 bl_143 br_143 wl_7 vdd gnd cell_6t
Xbit_r8_c143 bl_143 br_143 wl_8 vdd gnd cell_6t
Xbit_r9_c143 bl_143 br_143 wl_9 vdd gnd cell_6t
Xbit_r10_c143 bl_143 br_143 wl_10 vdd gnd cell_6t
Xbit_r11_c143 bl_143 br_143 wl_11 vdd gnd cell_6t
Xbit_r12_c143 bl_143 br_143 wl_12 vdd gnd cell_6t
Xbit_r13_c143 bl_143 br_143 wl_13 vdd gnd cell_6t
Xbit_r14_c143 bl_143 br_143 wl_14 vdd gnd cell_6t
Xbit_r15_c143 bl_143 br_143 wl_15 vdd gnd cell_6t
Xbit_r16_c143 bl_143 br_143 wl_16 vdd gnd cell_6t
Xbit_r17_c143 bl_143 br_143 wl_17 vdd gnd cell_6t
Xbit_r18_c143 bl_143 br_143 wl_18 vdd gnd cell_6t
Xbit_r19_c143 bl_143 br_143 wl_19 vdd gnd cell_6t
Xbit_r20_c143 bl_143 br_143 wl_20 vdd gnd cell_6t
Xbit_r21_c143 bl_143 br_143 wl_21 vdd gnd cell_6t
Xbit_r22_c143 bl_143 br_143 wl_22 vdd gnd cell_6t
Xbit_r23_c143 bl_143 br_143 wl_23 vdd gnd cell_6t
Xbit_r24_c143 bl_143 br_143 wl_24 vdd gnd cell_6t
Xbit_r25_c143 bl_143 br_143 wl_25 vdd gnd cell_6t
Xbit_r26_c143 bl_143 br_143 wl_26 vdd gnd cell_6t
Xbit_r27_c143 bl_143 br_143 wl_27 vdd gnd cell_6t
Xbit_r28_c143 bl_143 br_143 wl_28 vdd gnd cell_6t
Xbit_r29_c143 bl_143 br_143 wl_29 vdd gnd cell_6t
Xbit_r30_c143 bl_143 br_143 wl_30 vdd gnd cell_6t
Xbit_r31_c143 bl_143 br_143 wl_31 vdd gnd cell_6t
Xbit_r32_c143 bl_143 br_143 wl_32 vdd gnd cell_6t
Xbit_r33_c143 bl_143 br_143 wl_33 vdd gnd cell_6t
Xbit_r34_c143 bl_143 br_143 wl_34 vdd gnd cell_6t
Xbit_r35_c143 bl_143 br_143 wl_35 vdd gnd cell_6t
Xbit_r36_c143 bl_143 br_143 wl_36 vdd gnd cell_6t
Xbit_r37_c143 bl_143 br_143 wl_37 vdd gnd cell_6t
Xbit_r38_c143 bl_143 br_143 wl_38 vdd gnd cell_6t
Xbit_r39_c143 bl_143 br_143 wl_39 vdd gnd cell_6t
Xbit_r40_c143 bl_143 br_143 wl_40 vdd gnd cell_6t
Xbit_r41_c143 bl_143 br_143 wl_41 vdd gnd cell_6t
Xbit_r42_c143 bl_143 br_143 wl_42 vdd gnd cell_6t
Xbit_r43_c143 bl_143 br_143 wl_43 vdd gnd cell_6t
Xbit_r44_c143 bl_143 br_143 wl_44 vdd gnd cell_6t
Xbit_r45_c143 bl_143 br_143 wl_45 vdd gnd cell_6t
Xbit_r46_c143 bl_143 br_143 wl_46 vdd gnd cell_6t
Xbit_r47_c143 bl_143 br_143 wl_47 vdd gnd cell_6t
Xbit_r48_c143 bl_143 br_143 wl_48 vdd gnd cell_6t
Xbit_r49_c143 bl_143 br_143 wl_49 vdd gnd cell_6t
Xbit_r50_c143 bl_143 br_143 wl_50 vdd gnd cell_6t
Xbit_r51_c143 bl_143 br_143 wl_51 vdd gnd cell_6t
Xbit_r52_c143 bl_143 br_143 wl_52 vdd gnd cell_6t
Xbit_r53_c143 bl_143 br_143 wl_53 vdd gnd cell_6t
Xbit_r54_c143 bl_143 br_143 wl_54 vdd gnd cell_6t
Xbit_r55_c143 bl_143 br_143 wl_55 vdd gnd cell_6t
Xbit_r56_c143 bl_143 br_143 wl_56 vdd gnd cell_6t
Xbit_r57_c143 bl_143 br_143 wl_57 vdd gnd cell_6t
Xbit_r58_c143 bl_143 br_143 wl_58 vdd gnd cell_6t
Xbit_r59_c143 bl_143 br_143 wl_59 vdd gnd cell_6t
Xbit_r60_c143 bl_143 br_143 wl_60 vdd gnd cell_6t
Xbit_r61_c143 bl_143 br_143 wl_61 vdd gnd cell_6t
Xbit_r62_c143 bl_143 br_143 wl_62 vdd gnd cell_6t
Xbit_r63_c143 bl_143 br_143 wl_63 vdd gnd cell_6t
Xbit_r64_c143 bl_143 br_143 wl_64 vdd gnd cell_6t
Xbit_r65_c143 bl_143 br_143 wl_65 vdd gnd cell_6t
Xbit_r66_c143 bl_143 br_143 wl_66 vdd gnd cell_6t
Xbit_r67_c143 bl_143 br_143 wl_67 vdd gnd cell_6t
Xbit_r68_c143 bl_143 br_143 wl_68 vdd gnd cell_6t
Xbit_r69_c143 bl_143 br_143 wl_69 vdd gnd cell_6t
Xbit_r70_c143 bl_143 br_143 wl_70 vdd gnd cell_6t
Xbit_r71_c143 bl_143 br_143 wl_71 vdd gnd cell_6t
Xbit_r72_c143 bl_143 br_143 wl_72 vdd gnd cell_6t
Xbit_r73_c143 bl_143 br_143 wl_73 vdd gnd cell_6t
Xbit_r74_c143 bl_143 br_143 wl_74 vdd gnd cell_6t
Xbit_r75_c143 bl_143 br_143 wl_75 vdd gnd cell_6t
Xbit_r76_c143 bl_143 br_143 wl_76 vdd gnd cell_6t
Xbit_r77_c143 bl_143 br_143 wl_77 vdd gnd cell_6t
Xbit_r78_c143 bl_143 br_143 wl_78 vdd gnd cell_6t
Xbit_r79_c143 bl_143 br_143 wl_79 vdd gnd cell_6t
Xbit_r80_c143 bl_143 br_143 wl_80 vdd gnd cell_6t
Xbit_r81_c143 bl_143 br_143 wl_81 vdd gnd cell_6t
Xbit_r82_c143 bl_143 br_143 wl_82 vdd gnd cell_6t
Xbit_r83_c143 bl_143 br_143 wl_83 vdd gnd cell_6t
Xbit_r84_c143 bl_143 br_143 wl_84 vdd gnd cell_6t
Xbit_r85_c143 bl_143 br_143 wl_85 vdd gnd cell_6t
Xbit_r86_c143 bl_143 br_143 wl_86 vdd gnd cell_6t
Xbit_r87_c143 bl_143 br_143 wl_87 vdd gnd cell_6t
Xbit_r88_c143 bl_143 br_143 wl_88 vdd gnd cell_6t
Xbit_r89_c143 bl_143 br_143 wl_89 vdd gnd cell_6t
Xbit_r90_c143 bl_143 br_143 wl_90 vdd gnd cell_6t
Xbit_r91_c143 bl_143 br_143 wl_91 vdd gnd cell_6t
Xbit_r92_c143 bl_143 br_143 wl_92 vdd gnd cell_6t
Xbit_r93_c143 bl_143 br_143 wl_93 vdd gnd cell_6t
Xbit_r94_c143 bl_143 br_143 wl_94 vdd gnd cell_6t
Xbit_r95_c143 bl_143 br_143 wl_95 vdd gnd cell_6t
Xbit_r96_c143 bl_143 br_143 wl_96 vdd gnd cell_6t
Xbit_r97_c143 bl_143 br_143 wl_97 vdd gnd cell_6t
Xbit_r98_c143 bl_143 br_143 wl_98 vdd gnd cell_6t
Xbit_r99_c143 bl_143 br_143 wl_99 vdd gnd cell_6t
Xbit_r100_c143 bl_143 br_143 wl_100 vdd gnd cell_6t
Xbit_r101_c143 bl_143 br_143 wl_101 vdd gnd cell_6t
Xbit_r102_c143 bl_143 br_143 wl_102 vdd gnd cell_6t
Xbit_r103_c143 bl_143 br_143 wl_103 vdd gnd cell_6t
Xbit_r104_c143 bl_143 br_143 wl_104 vdd gnd cell_6t
Xbit_r105_c143 bl_143 br_143 wl_105 vdd gnd cell_6t
Xbit_r106_c143 bl_143 br_143 wl_106 vdd gnd cell_6t
Xbit_r107_c143 bl_143 br_143 wl_107 vdd gnd cell_6t
Xbit_r108_c143 bl_143 br_143 wl_108 vdd gnd cell_6t
Xbit_r109_c143 bl_143 br_143 wl_109 vdd gnd cell_6t
Xbit_r110_c143 bl_143 br_143 wl_110 vdd gnd cell_6t
Xbit_r111_c143 bl_143 br_143 wl_111 vdd gnd cell_6t
Xbit_r112_c143 bl_143 br_143 wl_112 vdd gnd cell_6t
Xbit_r113_c143 bl_143 br_143 wl_113 vdd gnd cell_6t
Xbit_r114_c143 bl_143 br_143 wl_114 vdd gnd cell_6t
Xbit_r115_c143 bl_143 br_143 wl_115 vdd gnd cell_6t
Xbit_r116_c143 bl_143 br_143 wl_116 vdd gnd cell_6t
Xbit_r117_c143 bl_143 br_143 wl_117 vdd gnd cell_6t
Xbit_r118_c143 bl_143 br_143 wl_118 vdd gnd cell_6t
Xbit_r119_c143 bl_143 br_143 wl_119 vdd gnd cell_6t
Xbit_r120_c143 bl_143 br_143 wl_120 vdd gnd cell_6t
Xbit_r121_c143 bl_143 br_143 wl_121 vdd gnd cell_6t
Xbit_r122_c143 bl_143 br_143 wl_122 vdd gnd cell_6t
Xbit_r123_c143 bl_143 br_143 wl_123 vdd gnd cell_6t
Xbit_r124_c143 bl_143 br_143 wl_124 vdd gnd cell_6t
Xbit_r125_c143 bl_143 br_143 wl_125 vdd gnd cell_6t
Xbit_r126_c143 bl_143 br_143 wl_126 vdd gnd cell_6t
Xbit_r127_c143 bl_143 br_143 wl_127 vdd gnd cell_6t
Xbit_r128_c143 bl_143 br_143 wl_128 vdd gnd cell_6t
Xbit_r129_c143 bl_143 br_143 wl_129 vdd gnd cell_6t
Xbit_r130_c143 bl_143 br_143 wl_130 vdd gnd cell_6t
Xbit_r131_c143 bl_143 br_143 wl_131 vdd gnd cell_6t
Xbit_r132_c143 bl_143 br_143 wl_132 vdd gnd cell_6t
Xbit_r133_c143 bl_143 br_143 wl_133 vdd gnd cell_6t
Xbit_r134_c143 bl_143 br_143 wl_134 vdd gnd cell_6t
Xbit_r135_c143 bl_143 br_143 wl_135 vdd gnd cell_6t
Xbit_r136_c143 bl_143 br_143 wl_136 vdd gnd cell_6t
Xbit_r137_c143 bl_143 br_143 wl_137 vdd gnd cell_6t
Xbit_r138_c143 bl_143 br_143 wl_138 vdd gnd cell_6t
Xbit_r139_c143 bl_143 br_143 wl_139 vdd gnd cell_6t
Xbit_r140_c143 bl_143 br_143 wl_140 vdd gnd cell_6t
Xbit_r141_c143 bl_143 br_143 wl_141 vdd gnd cell_6t
Xbit_r142_c143 bl_143 br_143 wl_142 vdd gnd cell_6t
Xbit_r143_c143 bl_143 br_143 wl_143 vdd gnd cell_6t
Xbit_r144_c143 bl_143 br_143 wl_144 vdd gnd cell_6t
Xbit_r145_c143 bl_143 br_143 wl_145 vdd gnd cell_6t
Xbit_r146_c143 bl_143 br_143 wl_146 vdd gnd cell_6t
Xbit_r147_c143 bl_143 br_143 wl_147 vdd gnd cell_6t
Xbit_r148_c143 bl_143 br_143 wl_148 vdd gnd cell_6t
Xbit_r149_c143 bl_143 br_143 wl_149 vdd gnd cell_6t
Xbit_r150_c143 bl_143 br_143 wl_150 vdd gnd cell_6t
Xbit_r151_c143 bl_143 br_143 wl_151 vdd gnd cell_6t
Xbit_r152_c143 bl_143 br_143 wl_152 vdd gnd cell_6t
Xbit_r153_c143 bl_143 br_143 wl_153 vdd gnd cell_6t
Xbit_r154_c143 bl_143 br_143 wl_154 vdd gnd cell_6t
Xbit_r155_c143 bl_143 br_143 wl_155 vdd gnd cell_6t
Xbit_r156_c143 bl_143 br_143 wl_156 vdd gnd cell_6t
Xbit_r157_c143 bl_143 br_143 wl_157 vdd gnd cell_6t
Xbit_r158_c143 bl_143 br_143 wl_158 vdd gnd cell_6t
Xbit_r159_c143 bl_143 br_143 wl_159 vdd gnd cell_6t
Xbit_r160_c143 bl_143 br_143 wl_160 vdd gnd cell_6t
Xbit_r161_c143 bl_143 br_143 wl_161 vdd gnd cell_6t
Xbit_r162_c143 bl_143 br_143 wl_162 vdd gnd cell_6t
Xbit_r163_c143 bl_143 br_143 wl_163 vdd gnd cell_6t
Xbit_r164_c143 bl_143 br_143 wl_164 vdd gnd cell_6t
Xbit_r165_c143 bl_143 br_143 wl_165 vdd gnd cell_6t
Xbit_r166_c143 bl_143 br_143 wl_166 vdd gnd cell_6t
Xbit_r167_c143 bl_143 br_143 wl_167 vdd gnd cell_6t
Xbit_r168_c143 bl_143 br_143 wl_168 vdd gnd cell_6t
Xbit_r169_c143 bl_143 br_143 wl_169 vdd gnd cell_6t
Xbit_r170_c143 bl_143 br_143 wl_170 vdd gnd cell_6t
Xbit_r171_c143 bl_143 br_143 wl_171 vdd gnd cell_6t
Xbit_r172_c143 bl_143 br_143 wl_172 vdd gnd cell_6t
Xbit_r173_c143 bl_143 br_143 wl_173 vdd gnd cell_6t
Xbit_r174_c143 bl_143 br_143 wl_174 vdd gnd cell_6t
Xbit_r175_c143 bl_143 br_143 wl_175 vdd gnd cell_6t
Xbit_r176_c143 bl_143 br_143 wl_176 vdd gnd cell_6t
Xbit_r177_c143 bl_143 br_143 wl_177 vdd gnd cell_6t
Xbit_r178_c143 bl_143 br_143 wl_178 vdd gnd cell_6t
Xbit_r179_c143 bl_143 br_143 wl_179 vdd gnd cell_6t
Xbit_r180_c143 bl_143 br_143 wl_180 vdd gnd cell_6t
Xbit_r181_c143 bl_143 br_143 wl_181 vdd gnd cell_6t
Xbit_r182_c143 bl_143 br_143 wl_182 vdd gnd cell_6t
Xbit_r183_c143 bl_143 br_143 wl_183 vdd gnd cell_6t
Xbit_r184_c143 bl_143 br_143 wl_184 vdd gnd cell_6t
Xbit_r185_c143 bl_143 br_143 wl_185 vdd gnd cell_6t
Xbit_r186_c143 bl_143 br_143 wl_186 vdd gnd cell_6t
Xbit_r187_c143 bl_143 br_143 wl_187 vdd gnd cell_6t
Xbit_r188_c143 bl_143 br_143 wl_188 vdd gnd cell_6t
Xbit_r189_c143 bl_143 br_143 wl_189 vdd gnd cell_6t
Xbit_r190_c143 bl_143 br_143 wl_190 vdd gnd cell_6t
Xbit_r191_c143 bl_143 br_143 wl_191 vdd gnd cell_6t
Xbit_r192_c143 bl_143 br_143 wl_192 vdd gnd cell_6t
Xbit_r193_c143 bl_143 br_143 wl_193 vdd gnd cell_6t
Xbit_r194_c143 bl_143 br_143 wl_194 vdd gnd cell_6t
Xbit_r195_c143 bl_143 br_143 wl_195 vdd gnd cell_6t
Xbit_r196_c143 bl_143 br_143 wl_196 vdd gnd cell_6t
Xbit_r197_c143 bl_143 br_143 wl_197 vdd gnd cell_6t
Xbit_r198_c143 bl_143 br_143 wl_198 vdd gnd cell_6t
Xbit_r199_c143 bl_143 br_143 wl_199 vdd gnd cell_6t
Xbit_r200_c143 bl_143 br_143 wl_200 vdd gnd cell_6t
Xbit_r201_c143 bl_143 br_143 wl_201 vdd gnd cell_6t
Xbit_r202_c143 bl_143 br_143 wl_202 vdd gnd cell_6t
Xbit_r203_c143 bl_143 br_143 wl_203 vdd gnd cell_6t
Xbit_r204_c143 bl_143 br_143 wl_204 vdd gnd cell_6t
Xbit_r205_c143 bl_143 br_143 wl_205 vdd gnd cell_6t
Xbit_r206_c143 bl_143 br_143 wl_206 vdd gnd cell_6t
Xbit_r207_c143 bl_143 br_143 wl_207 vdd gnd cell_6t
Xbit_r208_c143 bl_143 br_143 wl_208 vdd gnd cell_6t
Xbit_r209_c143 bl_143 br_143 wl_209 vdd gnd cell_6t
Xbit_r210_c143 bl_143 br_143 wl_210 vdd gnd cell_6t
Xbit_r211_c143 bl_143 br_143 wl_211 vdd gnd cell_6t
Xbit_r212_c143 bl_143 br_143 wl_212 vdd gnd cell_6t
Xbit_r213_c143 bl_143 br_143 wl_213 vdd gnd cell_6t
Xbit_r214_c143 bl_143 br_143 wl_214 vdd gnd cell_6t
Xbit_r215_c143 bl_143 br_143 wl_215 vdd gnd cell_6t
Xbit_r216_c143 bl_143 br_143 wl_216 vdd gnd cell_6t
Xbit_r217_c143 bl_143 br_143 wl_217 vdd gnd cell_6t
Xbit_r218_c143 bl_143 br_143 wl_218 vdd gnd cell_6t
Xbit_r219_c143 bl_143 br_143 wl_219 vdd gnd cell_6t
Xbit_r220_c143 bl_143 br_143 wl_220 vdd gnd cell_6t
Xbit_r221_c143 bl_143 br_143 wl_221 vdd gnd cell_6t
Xbit_r222_c143 bl_143 br_143 wl_222 vdd gnd cell_6t
Xbit_r223_c143 bl_143 br_143 wl_223 vdd gnd cell_6t
Xbit_r224_c143 bl_143 br_143 wl_224 vdd gnd cell_6t
Xbit_r225_c143 bl_143 br_143 wl_225 vdd gnd cell_6t
Xbit_r226_c143 bl_143 br_143 wl_226 vdd gnd cell_6t
Xbit_r227_c143 bl_143 br_143 wl_227 vdd gnd cell_6t
Xbit_r228_c143 bl_143 br_143 wl_228 vdd gnd cell_6t
Xbit_r229_c143 bl_143 br_143 wl_229 vdd gnd cell_6t
Xbit_r230_c143 bl_143 br_143 wl_230 vdd gnd cell_6t
Xbit_r231_c143 bl_143 br_143 wl_231 vdd gnd cell_6t
Xbit_r232_c143 bl_143 br_143 wl_232 vdd gnd cell_6t
Xbit_r233_c143 bl_143 br_143 wl_233 vdd gnd cell_6t
Xbit_r234_c143 bl_143 br_143 wl_234 vdd gnd cell_6t
Xbit_r235_c143 bl_143 br_143 wl_235 vdd gnd cell_6t
Xbit_r236_c143 bl_143 br_143 wl_236 vdd gnd cell_6t
Xbit_r237_c143 bl_143 br_143 wl_237 vdd gnd cell_6t
Xbit_r238_c143 bl_143 br_143 wl_238 vdd gnd cell_6t
Xbit_r239_c143 bl_143 br_143 wl_239 vdd gnd cell_6t
Xbit_r240_c143 bl_143 br_143 wl_240 vdd gnd cell_6t
Xbit_r241_c143 bl_143 br_143 wl_241 vdd gnd cell_6t
Xbit_r242_c143 bl_143 br_143 wl_242 vdd gnd cell_6t
Xbit_r243_c143 bl_143 br_143 wl_243 vdd gnd cell_6t
Xbit_r244_c143 bl_143 br_143 wl_244 vdd gnd cell_6t
Xbit_r245_c143 bl_143 br_143 wl_245 vdd gnd cell_6t
Xbit_r246_c143 bl_143 br_143 wl_246 vdd gnd cell_6t
Xbit_r247_c143 bl_143 br_143 wl_247 vdd gnd cell_6t
Xbit_r248_c143 bl_143 br_143 wl_248 vdd gnd cell_6t
Xbit_r249_c143 bl_143 br_143 wl_249 vdd gnd cell_6t
Xbit_r250_c143 bl_143 br_143 wl_250 vdd gnd cell_6t
Xbit_r251_c143 bl_143 br_143 wl_251 vdd gnd cell_6t
Xbit_r252_c143 bl_143 br_143 wl_252 vdd gnd cell_6t
Xbit_r253_c143 bl_143 br_143 wl_253 vdd gnd cell_6t
Xbit_r254_c143 bl_143 br_143 wl_254 vdd gnd cell_6t
Xbit_r255_c143 bl_143 br_143 wl_255 vdd gnd cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd cell_6t
Xbit_r1_c144 bl_144 br_144 wl_1 vdd gnd cell_6t
Xbit_r2_c144 bl_144 br_144 wl_2 vdd gnd cell_6t
Xbit_r3_c144 bl_144 br_144 wl_3 vdd gnd cell_6t
Xbit_r4_c144 bl_144 br_144 wl_4 vdd gnd cell_6t
Xbit_r5_c144 bl_144 br_144 wl_5 vdd gnd cell_6t
Xbit_r6_c144 bl_144 br_144 wl_6 vdd gnd cell_6t
Xbit_r7_c144 bl_144 br_144 wl_7 vdd gnd cell_6t
Xbit_r8_c144 bl_144 br_144 wl_8 vdd gnd cell_6t
Xbit_r9_c144 bl_144 br_144 wl_9 vdd gnd cell_6t
Xbit_r10_c144 bl_144 br_144 wl_10 vdd gnd cell_6t
Xbit_r11_c144 bl_144 br_144 wl_11 vdd gnd cell_6t
Xbit_r12_c144 bl_144 br_144 wl_12 vdd gnd cell_6t
Xbit_r13_c144 bl_144 br_144 wl_13 vdd gnd cell_6t
Xbit_r14_c144 bl_144 br_144 wl_14 vdd gnd cell_6t
Xbit_r15_c144 bl_144 br_144 wl_15 vdd gnd cell_6t
Xbit_r16_c144 bl_144 br_144 wl_16 vdd gnd cell_6t
Xbit_r17_c144 bl_144 br_144 wl_17 vdd gnd cell_6t
Xbit_r18_c144 bl_144 br_144 wl_18 vdd gnd cell_6t
Xbit_r19_c144 bl_144 br_144 wl_19 vdd gnd cell_6t
Xbit_r20_c144 bl_144 br_144 wl_20 vdd gnd cell_6t
Xbit_r21_c144 bl_144 br_144 wl_21 vdd gnd cell_6t
Xbit_r22_c144 bl_144 br_144 wl_22 vdd gnd cell_6t
Xbit_r23_c144 bl_144 br_144 wl_23 vdd gnd cell_6t
Xbit_r24_c144 bl_144 br_144 wl_24 vdd gnd cell_6t
Xbit_r25_c144 bl_144 br_144 wl_25 vdd gnd cell_6t
Xbit_r26_c144 bl_144 br_144 wl_26 vdd gnd cell_6t
Xbit_r27_c144 bl_144 br_144 wl_27 vdd gnd cell_6t
Xbit_r28_c144 bl_144 br_144 wl_28 vdd gnd cell_6t
Xbit_r29_c144 bl_144 br_144 wl_29 vdd gnd cell_6t
Xbit_r30_c144 bl_144 br_144 wl_30 vdd gnd cell_6t
Xbit_r31_c144 bl_144 br_144 wl_31 vdd gnd cell_6t
Xbit_r32_c144 bl_144 br_144 wl_32 vdd gnd cell_6t
Xbit_r33_c144 bl_144 br_144 wl_33 vdd gnd cell_6t
Xbit_r34_c144 bl_144 br_144 wl_34 vdd gnd cell_6t
Xbit_r35_c144 bl_144 br_144 wl_35 vdd gnd cell_6t
Xbit_r36_c144 bl_144 br_144 wl_36 vdd gnd cell_6t
Xbit_r37_c144 bl_144 br_144 wl_37 vdd gnd cell_6t
Xbit_r38_c144 bl_144 br_144 wl_38 vdd gnd cell_6t
Xbit_r39_c144 bl_144 br_144 wl_39 vdd gnd cell_6t
Xbit_r40_c144 bl_144 br_144 wl_40 vdd gnd cell_6t
Xbit_r41_c144 bl_144 br_144 wl_41 vdd gnd cell_6t
Xbit_r42_c144 bl_144 br_144 wl_42 vdd gnd cell_6t
Xbit_r43_c144 bl_144 br_144 wl_43 vdd gnd cell_6t
Xbit_r44_c144 bl_144 br_144 wl_44 vdd gnd cell_6t
Xbit_r45_c144 bl_144 br_144 wl_45 vdd gnd cell_6t
Xbit_r46_c144 bl_144 br_144 wl_46 vdd gnd cell_6t
Xbit_r47_c144 bl_144 br_144 wl_47 vdd gnd cell_6t
Xbit_r48_c144 bl_144 br_144 wl_48 vdd gnd cell_6t
Xbit_r49_c144 bl_144 br_144 wl_49 vdd gnd cell_6t
Xbit_r50_c144 bl_144 br_144 wl_50 vdd gnd cell_6t
Xbit_r51_c144 bl_144 br_144 wl_51 vdd gnd cell_6t
Xbit_r52_c144 bl_144 br_144 wl_52 vdd gnd cell_6t
Xbit_r53_c144 bl_144 br_144 wl_53 vdd gnd cell_6t
Xbit_r54_c144 bl_144 br_144 wl_54 vdd gnd cell_6t
Xbit_r55_c144 bl_144 br_144 wl_55 vdd gnd cell_6t
Xbit_r56_c144 bl_144 br_144 wl_56 vdd gnd cell_6t
Xbit_r57_c144 bl_144 br_144 wl_57 vdd gnd cell_6t
Xbit_r58_c144 bl_144 br_144 wl_58 vdd gnd cell_6t
Xbit_r59_c144 bl_144 br_144 wl_59 vdd gnd cell_6t
Xbit_r60_c144 bl_144 br_144 wl_60 vdd gnd cell_6t
Xbit_r61_c144 bl_144 br_144 wl_61 vdd gnd cell_6t
Xbit_r62_c144 bl_144 br_144 wl_62 vdd gnd cell_6t
Xbit_r63_c144 bl_144 br_144 wl_63 vdd gnd cell_6t
Xbit_r64_c144 bl_144 br_144 wl_64 vdd gnd cell_6t
Xbit_r65_c144 bl_144 br_144 wl_65 vdd gnd cell_6t
Xbit_r66_c144 bl_144 br_144 wl_66 vdd gnd cell_6t
Xbit_r67_c144 bl_144 br_144 wl_67 vdd gnd cell_6t
Xbit_r68_c144 bl_144 br_144 wl_68 vdd gnd cell_6t
Xbit_r69_c144 bl_144 br_144 wl_69 vdd gnd cell_6t
Xbit_r70_c144 bl_144 br_144 wl_70 vdd gnd cell_6t
Xbit_r71_c144 bl_144 br_144 wl_71 vdd gnd cell_6t
Xbit_r72_c144 bl_144 br_144 wl_72 vdd gnd cell_6t
Xbit_r73_c144 bl_144 br_144 wl_73 vdd gnd cell_6t
Xbit_r74_c144 bl_144 br_144 wl_74 vdd gnd cell_6t
Xbit_r75_c144 bl_144 br_144 wl_75 vdd gnd cell_6t
Xbit_r76_c144 bl_144 br_144 wl_76 vdd gnd cell_6t
Xbit_r77_c144 bl_144 br_144 wl_77 vdd gnd cell_6t
Xbit_r78_c144 bl_144 br_144 wl_78 vdd gnd cell_6t
Xbit_r79_c144 bl_144 br_144 wl_79 vdd gnd cell_6t
Xbit_r80_c144 bl_144 br_144 wl_80 vdd gnd cell_6t
Xbit_r81_c144 bl_144 br_144 wl_81 vdd gnd cell_6t
Xbit_r82_c144 bl_144 br_144 wl_82 vdd gnd cell_6t
Xbit_r83_c144 bl_144 br_144 wl_83 vdd gnd cell_6t
Xbit_r84_c144 bl_144 br_144 wl_84 vdd gnd cell_6t
Xbit_r85_c144 bl_144 br_144 wl_85 vdd gnd cell_6t
Xbit_r86_c144 bl_144 br_144 wl_86 vdd gnd cell_6t
Xbit_r87_c144 bl_144 br_144 wl_87 vdd gnd cell_6t
Xbit_r88_c144 bl_144 br_144 wl_88 vdd gnd cell_6t
Xbit_r89_c144 bl_144 br_144 wl_89 vdd gnd cell_6t
Xbit_r90_c144 bl_144 br_144 wl_90 vdd gnd cell_6t
Xbit_r91_c144 bl_144 br_144 wl_91 vdd gnd cell_6t
Xbit_r92_c144 bl_144 br_144 wl_92 vdd gnd cell_6t
Xbit_r93_c144 bl_144 br_144 wl_93 vdd gnd cell_6t
Xbit_r94_c144 bl_144 br_144 wl_94 vdd gnd cell_6t
Xbit_r95_c144 bl_144 br_144 wl_95 vdd gnd cell_6t
Xbit_r96_c144 bl_144 br_144 wl_96 vdd gnd cell_6t
Xbit_r97_c144 bl_144 br_144 wl_97 vdd gnd cell_6t
Xbit_r98_c144 bl_144 br_144 wl_98 vdd gnd cell_6t
Xbit_r99_c144 bl_144 br_144 wl_99 vdd gnd cell_6t
Xbit_r100_c144 bl_144 br_144 wl_100 vdd gnd cell_6t
Xbit_r101_c144 bl_144 br_144 wl_101 vdd gnd cell_6t
Xbit_r102_c144 bl_144 br_144 wl_102 vdd gnd cell_6t
Xbit_r103_c144 bl_144 br_144 wl_103 vdd gnd cell_6t
Xbit_r104_c144 bl_144 br_144 wl_104 vdd gnd cell_6t
Xbit_r105_c144 bl_144 br_144 wl_105 vdd gnd cell_6t
Xbit_r106_c144 bl_144 br_144 wl_106 vdd gnd cell_6t
Xbit_r107_c144 bl_144 br_144 wl_107 vdd gnd cell_6t
Xbit_r108_c144 bl_144 br_144 wl_108 vdd gnd cell_6t
Xbit_r109_c144 bl_144 br_144 wl_109 vdd gnd cell_6t
Xbit_r110_c144 bl_144 br_144 wl_110 vdd gnd cell_6t
Xbit_r111_c144 bl_144 br_144 wl_111 vdd gnd cell_6t
Xbit_r112_c144 bl_144 br_144 wl_112 vdd gnd cell_6t
Xbit_r113_c144 bl_144 br_144 wl_113 vdd gnd cell_6t
Xbit_r114_c144 bl_144 br_144 wl_114 vdd gnd cell_6t
Xbit_r115_c144 bl_144 br_144 wl_115 vdd gnd cell_6t
Xbit_r116_c144 bl_144 br_144 wl_116 vdd gnd cell_6t
Xbit_r117_c144 bl_144 br_144 wl_117 vdd gnd cell_6t
Xbit_r118_c144 bl_144 br_144 wl_118 vdd gnd cell_6t
Xbit_r119_c144 bl_144 br_144 wl_119 vdd gnd cell_6t
Xbit_r120_c144 bl_144 br_144 wl_120 vdd gnd cell_6t
Xbit_r121_c144 bl_144 br_144 wl_121 vdd gnd cell_6t
Xbit_r122_c144 bl_144 br_144 wl_122 vdd gnd cell_6t
Xbit_r123_c144 bl_144 br_144 wl_123 vdd gnd cell_6t
Xbit_r124_c144 bl_144 br_144 wl_124 vdd gnd cell_6t
Xbit_r125_c144 bl_144 br_144 wl_125 vdd gnd cell_6t
Xbit_r126_c144 bl_144 br_144 wl_126 vdd gnd cell_6t
Xbit_r127_c144 bl_144 br_144 wl_127 vdd gnd cell_6t
Xbit_r128_c144 bl_144 br_144 wl_128 vdd gnd cell_6t
Xbit_r129_c144 bl_144 br_144 wl_129 vdd gnd cell_6t
Xbit_r130_c144 bl_144 br_144 wl_130 vdd gnd cell_6t
Xbit_r131_c144 bl_144 br_144 wl_131 vdd gnd cell_6t
Xbit_r132_c144 bl_144 br_144 wl_132 vdd gnd cell_6t
Xbit_r133_c144 bl_144 br_144 wl_133 vdd gnd cell_6t
Xbit_r134_c144 bl_144 br_144 wl_134 vdd gnd cell_6t
Xbit_r135_c144 bl_144 br_144 wl_135 vdd gnd cell_6t
Xbit_r136_c144 bl_144 br_144 wl_136 vdd gnd cell_6t
Xbit_r137_c144 bl_144 br_144 wl_137 vdd gnd cell_6t
Xbit_r138_c144 bl_144 br_144 wl_138 vdd gnd cell_6t
Xbit_r139_c144 bl_144 br_144 wl_139 vdd gnd cell_6t
Xbit_r140_c144 bl_144 br_144 wl_140 vdd gnd cell_6t
Xbit_r141_c144 bl_144 br_144 wl_141 vdd gnd cell_6t
Xbit_r142_c144 bl_144 br_144 wl_142 vdd gnd cell_6t
Xbit_r143_c144 bl_144 br_144 wl_143 vdd gnd cell_6t
Xbit_r144_c144 bl_144 br_144 wl_144 vdd gnd cell_6t
Xbit_r145_c144 bl_144 br_144 wl_145 vdd gnd cell_6t
Xbit_r146_c144 bl_144 br_144 wl_146 vdd gnd cell_6t
Xbit_r147_c144 bl_144 br_144 wl_147 vdd gnd cell_6t
Xbit_r148_c144 bl_144 br_144 wl_148 vdd gnd cell_6t
Xbit_r149_c144 bl_144 br_144 wl_149 vdd gnd cell_6t
Xbit_r150_c144 bl_144 br_144 wl_150 vdd gnd cell_6t
Xbit_r151_c144 bl_144 br_144 wl_151 vdd gnd cell_6t
Xbit_r152_c144 bl_144 br_144 wl_152 vdd gnd cell_6t
Xbit_r153_c144 bl_144 br_144 wl_153 vdd gnd cell_6t
Xbit_r154_c144 bl_144 br_144 wl_154 vdd gnd cell_6t
Xbit_r155_c144 bl_144 br_144 wl_155 vdd gnd cell_6t
Xbit_r156_c144 bl_144 br_144 wl_156 vdd gnd cell_6t
Xbit_r157_c144 bl_144 br_144 wl_157 vdd gnd cell_6t
Xbit_r158_c144 bl_144 br_144 wl_158 vdd gnd cell_6t
Xbit_r159_c144 bl_144 br_144 wl_159 vdd gnd cell_6t
Xbit_r160_c144 bl_144 br_144 wl_160 vdd gnd cell_6t
Xbit_r161_c144 bl_144 br_144 wl_161 vdd gnd cell_6t
Xbit_r162_c144 bl_144 br_144 wl_162 vdd gnd cell_6t
Xbit_r163_c144 bl_144 br_144 wl_163 vdd gnd cell_6t
Xbit_r164_c144 bl_144 br_144 wl_164 vdd gnd cell_6t
Xbit_r165_c144 bl_144 br_144 wl_165 vdd gnd cell_6t
Xbit_r166_c144 bl_144 br_144 wl_166 vdd gnd cell_6t
Xbit_r167_c144 bl_144 br_144 wl_167 vdd gnd cell_6t
Xbit_r168_c144 bl_144 br_144 wl_168 vdd gnd cell_6t
Xbit_r169_c144 bl_144 br_144 wl_169 vdd gnd cell_6t
Xbit_r170_c144 bl_144 br_144 wl_170 vdd gnd cell_6t
Xbit_r171_c144 bl_144 br_144 wl_171 vdd gnd cell_6t
Xbit_r172_c144 bl_144 br_144 wl_172 vdd gnd cell_6t
Xbit_r173_c144 bl_144 br_144 wl_173 vdd gnd cell_6t
Xbit_r174_c144 bl_144 br_144 wl_174 vdd gnd cell_6t
Xbit_r175_c144 bl_144 br_144 wl_175 vdd gnd cell_6t
Xbit_r176_c144 bl_144 br_144 wl_176 vdd gnd cell_6t
Xbit_r177_c144 bl_144 br_144 wl_177 vdd gnd cell_6t
Xbit_r178_c144 bl_144 br_144 wl_178 vdd gnd cell_6t
Xbit_r179_c144 bl_144 br_144 wl_179 vdd gnd cell_6t
Xbit_r180_c144 bl_144 br_144 wl_180 vdd gnd cell_6t
Xbit_r181_c144 bl_144 br_144 wl_181 vdd gnd cell_6t
Xbit_r182_c144 bl_144 br_144 wl_182 vdd gnd cell_6t
Xbit_r183_c144 bl_144 br_144 wl_183 vdd gnd cell_6t
Xbit_r184_c144 bl_144 br_144 wl_184 vdd gnd cell_6t
Xbit_r185_c144 bl_144 br_144 wl_185 vdd gnd cell_6t
Xbit_r186_c144 bl_144 br_144 wl_186 vdd gnd cell_6t
Xbit_r187_c144 bl_144 br_144 wl_187 vdd gnd cell_6t
Xbit_r188_c144 bl_144 br_144 wl_188 vdd gnd cell_6t
Xbit_r189_c144 bl_144 br_144 wl_189 vdd gnd cell_6t
Xbit_r190_c144 bl_144 br_144 wl_190 vdd gnd cell_6t
Xbit_r191_c144 bl_144 br_144 wl_191 vdd gnd cell_6t
Xbit_r192_c144 bl_144 br_144 wl_192 vdd gnd cell_6t
Xbit_r193_c144 bl_144 br_144 wl_193 vdd gnd cell_6t
Xbit_r194_c144 bl_144 br_144 wl_194 vdd gnd cell_6t
Xbit_r195_c144 bl_144 br_144 wl_195 vdd gnd cell_6t
Xbit_r196_c144 bl_144 br_144 wl_196 vdd gnd cell_6t
Xbit_r197_c144 bl_144 br_144 wl_197 vdd gnd cell_6t
Xbit_r198_c144 bl_144 br_144 wl_198 vdd gnd cell_6t
Xbit_r199_c144 bl_144 br_144 wl_199 vdd gnd cell_6t
Xbit_r200_c144 bl_144 br_144 wl_200 vdd gnd cell_6t
Xbit_r201_c144 bl_144 br_144 wl_201 vdd gnd cell_6t
Xbit_r202_c144 bl_144 br_144 wl_202 vdd gnd cell_6t
Xbit_r203_c144 bl_144 br_144 wl_203 vdd gnd cell_6t
Xbit_r204_c144 bl_144 br_144 wl_204 vdd gnd cell_6t
Xbit_r205_c144 bl_144 br_144 wl_205 vdd gnd cell_6t
Xbit_r206_c144 bl_144 br_144 wl_206 vdd gnd cell_6t
Xbit_r207_c144 bl_144 br_144 wl_207 vdd gnd cell_6t
Xbit_r208_c144 bl_144 br_144 wl_208 vdd gnd cell_6t
Xbit_r209_c144 bl_144 br_144 wl_209 vdd gnd cell_6t
Xbit_r210_c144 bl_144 br_144 wl_210 vdd gnd cell_6t
Xbit_r211_c144 bl_144 br_144 wl_211 vdd gnd cell_6t
Xbit_r212_c144 bl_144 br_144 wl_212 vdd gnd cell_6t
Xbit_r213_c144 bl_144 br_144 wl_213 vdd gnd cell_6t
Xbit_r214_c144 bl_144 br_144 wl_214 vdd gnd cell_6t
Xbit_r215_c144 bl_144 br_144 wl_215 vdd gnd cell_6t
Xbit_r216_c144 bl_144 br_144 wl_216 vdd gnd cell_6t
Xbit_r217_c144 bl_144 br_144 wl_217 vdd gnd cell_6t
Xbit_r218_c144 bl_144 br_144 wl_218 vdd gnd cell_6t
Xbit_r219_c144 bl_144 br_144 wl_219 vdd gnd cell_6t
Xbit_r220_c144 bl_144 br_144 wl_220 vdd gnd cell_6t
Xbit_r221_c144 bl_144 br_144 wl_221 vdd gnd cell_6t
Xbit_r222_c144 bl_144 br_144 wl_222 vdd gnd cell_6t
Xbit_r223_c144 bl_144 br_144 wl_223 vdd gnd cell_6t
Xbit_r224_c144 bl_144 br_144 wl_224 vdd gnd cell_6t
Xbit_r225_c144 bl_144 br_144 wl_225 vdd gnd cell_6t
Xbit_r226_c144 bl_144 br_144 wl_226 vdd gnd cell_6t
Xbit_r227_c144 bl_144 br_144 wl_227 vdd gnd cell_6t
Xbit_r228_c144 bl_144 br_144 wl_228 vdd gnd cell_6t
Xbit_r229_c144 bl_144 br_144 wl_229 vdd gnd cell_6t
Xbit_r230_c144 bl_144 br_144 wl_230 vdd gnd cell_6t
Xbit_r231_c144 bl_144 br_144 wl_231 vdd gnd cell_6t
Xbit_r232_c144 bl_144 br_144 wl_232 vdd gnd cell_6t
Xbit_r233_c144 bl_144 br_144 wl_233 vdd gnd cell_6t
Xbit_r234_c144 bl_144 br_144 wl_234 vdd gnd cell_6t
Xbit_r235_c144 bl_144 br_144 wl_235 vdd gnd cell_6t
Xbit_r236_c144 bl_144 br_144 wl_236 vdd gnd cell_6t
Xbit_r237_c144 bl_144 br_144 wl_237 vdd gnd cell_6t
Xbit_r238_c144 bl_144 br_144 wl_238 vdd gnd cell_6t
Xbit_r239_c144 bl_144 br_144 wl_239 vdd gnd cell_6t
Xbit_r240_c144 bl_144 br_144 wl_240 vdd gnd cell_6t
Xbit_r241_c144 bl_144 br_144 wl_241 vdd gnd cell_6t
Xbit_r242_c144 bl_144 br_144 wl_242 vdd gnd cell_6t
Xbit_r243_c144 bl_144 br_144 wl_243 vdd gnd cell_6t
Xbit_r244_c144 bl_144 br_144 wl_244 vdd gnd cell_6t
Xbit_r245_c144 bl_144 br_144 wl_245 vdd gnd cell_6t
Xbit_r246_c144 bl_144 br_144 wl_246 vdd gnd cell_6t
Xbit_r247_c144 bl_144 br_144 wl_247 vdd gnd cell_6t
Xbit_r248_c144 bl_144 br_144 wl_248 vdd gnd cell_6t
Xbit_r249_c144 bl_144 br_144 wl_249 vdd gnd cell_6t
Xbit_r250_c144 bl_144 br_144 wl_250 vdd gnd cell_6t
Xbit_r251_c144 bl_144 br_144 wl_251 vdd gnd cell_6t
Xbit_r252_c144 bl_144 br_144 wl_252 vdd gnd cell_6t
Xbit_r253_c144 bl_144 br_144 wl_253 vdd gnd cell_6t
Xbit_r254_c144 bl_144 br_144 wl_254 vdd gnd cell_6t
Xbit_r255_c144 bl_144 br_144 wl_255 vdd gnd cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd cell_6t
Xbit_r1_c145 bl_145 br_145 wl_1 vdd gnd cell_6t
Xbit_r2_c145 bl_145 br_145 wl_2 vdd gnd cell_6t
Xbit_r3_c145 bl_145 br_145 wl_3 vdd gnd cell_6t
Xbit_r4_c145 bl_145 br_145 wl_4 vdd gnd cell_6t
Xbit_r5_c145 bl_145 br_145 wl_5 vdd gnd cell_6t
Xbit_r6_c145 bl_145 br_145 wl_6 vdd gnd cell_6t
Xbit_r7_c145 bl_145 br_145 wl_7 vdd gnd cell_6t
Xbit_r8_c145 bl_145 br_145 wl_8 vdd gnd cell_6t
Xbit_r9_c145 bl_145 br_145 wl_9 vdd gnd cell_6t
Xbit_r10_c145 bl_145 br_145 wl_10 vdd gnd cell_6t
Xbit_r11_c145 bl_145 br_145 wl_11 vdd gnd cell_6t
Xbit_r12_c145 bl_145 br_145 wl_12 vdd gnd cell_6t
Xbit_r13_c145 bl_145 br_145 wl_13 vdd gnd cell_6t
Xbit_r14_c145 bl_145 br_145 wl_14 vdd gnd cell_6t
Xbit_r15_c145 bl_145 br_145 wl_15 vdd gnd cell_6t
Xbit_r16_c145 bl_145 br_145 wl_16 vdd gnd cell_6t
Xbit_r17_c145 bl_145 br_145 wl_17 vdd gnd cell_6t
Xbit_r18_c145 bl_145 br_145 wl_18 vdd gnd cell_6t
Xbit_r19_c145 bl_145 br_145 wl_19 vdd gnd cell_6t
Xbit_r20_c145 bl_145 br_145 wl_20 vdd gnd cell_6t
Xbit_r21_c145 bl_145 br_145 wl_21 vdd gnd cell_6t
Xbit_r22_c145 bl_145 br_145 wl_22 vdd gnd cell_6t
Xbit_r23_c145 bl_145 br_145 wl_23 vdd gnd cell_6t
Xbit_r24_c145 bl_145 br_145 wl_24 vdd gnd cell_6t
Xbit_r25_c145 bl_145 br_145 wl_25 vdd gnd cell_6t
Xbit_r26_c145 bl_145 br_145 wl_26 vdd gnd cell_6t
Xbit_r27_c145 bl_145 br_145 wl_27 vdd gnd cell_6t
Xbit_r28_c145 bl_145 br_145 wl_28 vdd gnd cell_6t
Xbit_r29_c145 bl_145 br_145 wl_29 vdd gnd cell_6t
Xbit_r30_c145 bl_145 br_145 wl_30 vdd gnd cell_6t
Xbit_r31_c145 bl_145 br_145 wl_31 vdd gnd cell_6t
Xbit_r32_c145 bl_145 br_145 wl_32 vdd gnd cell_6t
Xbit_r33_c145 bl_145 br_145 wl_33 vdd gnd cell_6t
Xbit_r34_c145 bl_145 br_145 wl_34 vdd gnd cell_6t
Xbit_r35_c145 bl_145 br_145 wl_35 vdd gnd cell_6t
Xbit_r36_c145 bl_145 br_145 wl_36 vdd gnd cell_6t
Xbit_r37_c145 bl_145 br_145 wl_37 vdd gnd cell_6t
Xbit_r38_c145 bl_145 br_145 wl_38 vdd gnd cell_6t
Xbit_r39_c145 bl_145 br_145 wl_39 vdd gnd cell_6t
Xbit_r40_c145 bl_145 br_145 wl_40 vdd gnd cell_6t
Xbit_r41_c145 bl_145 br_145 wl_41 vdd gnd cell_6t
Xbit_r42_c145 bl_145 br_145 wl_42 vdd gnd cell_6t
Xbit_r43_c145 bl_145 br_145 wl_43 vdd gnd cell_6t
Xbit_r44_c145 bl_145 br_145 wl_44 vdd gnd cell_6t
Xbit_r45_c145 bl_145 br_145 wl_45 vdd gnd cell_6t
Xbit_r46_c145 bl_145 br_145 wl_46 vdd gnd cell_6t
Xbit_r47_c145 bl_145 br_145 wl_47 vdd gnd cell_6t
Xbit_r48_c145 bl_145 br_145 wl_48 vdd gnd cell_6t
Xbit_r49_c145 bl_145 br_145 wl_49 vdd gnd cell_6t
Xbit_r50_c145 bl_145 br_145 wl_50 vdd gnd cell_6t
Xbit_r51_c145 bl_145 br_145 wl_51 vdd gnd cell_6t
Xbit_r52_c145 bl_145 br_145 wl_52 vdd gnd cell_6t
Xbit_r53_c145 bl_145 br_145 wl_53 vdd gnd cell_6t
Xbit_r54_c145 bl_145 br_145 wl_54 vdd gnd cell_6t
Xbit_r55_c145 bl_145 br_145 wl_55 vdd gnd cell_6t
Xbit_r56_c145 bl_145 br_145 wl_56 vdd gnd cell_6t
Xbit_r57_c145 bl_145 br_145 wl_57 vdd gnd cell_6t
Xbit_r58_c145 bl_145 br_145 wl_58 vdd gnd cell_6t
Xbit_r59_c145 bl_145 br_145 wl_59 vdd gnd cell_6t
Xbit_r60_c145 bl_145 br_145 wl_60 vdd gnd cell_6t
Xbit_r61_c145 bl_145 br_145 wl_61 vdd gnd cell_6t
Xbit_r62_c145 bl_145 br_145 wl_62 vdd gnd cell_6t
Xbit_r63_c145 bl_145 br_145 wl_63 vdd gnd cell_6t
Xbit_r64_c145 bl_145 br_145 wl_64 vdd gnd cell_6t
Xbit_r65_c145 bl_145 br_145 wl_65 vdd gnd cell_6t
Xbit_r66_c145 bl_145 br_145 wl_66 vdd gnd cell_6t
Xbit_r67_c145 bl_145 br_145 wl_67 vdd gnd cell_6t
Xbit_r68_c145 bl_145 br_145 wl_68 vdd gnd cell_6t
Xbit_r69_c145 bl_145 br_145 wl_69 vdd gnd cell_6t
Xbit_r70_c145 bl_145 br_145 wl_70 vdd gnd cell_6t
Xbit_r71_c145 bl_145 br_145 wl_71 vdd gnd cell_6t
Xbit_r72_c145 bl_145 br_145 wl_72 vdd gnd cell_6t
Xbit_r73_c145 bl_145 br_145 wl_73 vdd gnd cell_6t
Xbit_r74_c145 bl_145 br_145 wl_74 vdd gnd cell_6t
Xbit_r75_c145 bl_145 br_145 wl_75 vdd gnd cell_6t
Xbit_r76_c145 bl_145 br_145 wl_76 vdd gnd cell_6t
Xbit_r77_c145 bl_145 br_145 wl_77 vdd gnd cell_6t
Xbit_r78_c145 bl_145 br_145 wl_78 vdd gnd cell_6t
Xbit_r79_c145 bl_145 br_145 wl_79 vdd gnd cell_6t
Xbit_r80_c145 bl_145 br_145 wl_80 vdd gnd cell_6t
Xbit_r81_c145 bl_145 br_145 wl_81 vdd gnd cell_6t
Xbit_r82_c145 bl_145 br_145 wl_82 vdd gnd cell_6t
Xbit_r83_c145 bl_145 br_145 wl_83 vdd gnd cell_6t
Xbit_r84_c145 bl_145 br_145 wl_84 vdd gnd cell_6t
Xbit_r85_c145 bl_145 br_145 wl_85 vdd gnd cell_6t
Xbit_r86_c145 bl_145 br_145 wl_86 vdd gnd cell_6t
Xbit_r87_c145 bl_145 br_145 wl_87 vdd gnd cell_6t
Xbit_r88_c145 bl_145 br_145 wl_88 vdd gnd cell_6t
Xbit_r89_c145 bl_145 br_145 wl_89 vdd gnd cell_6t
Xbit_r90_c145 bl_145 br_145 wl_90 vdd gnd cell_6t
Xbit_r91_c145 bl_145 br_145 wl_91 vdd gnd cell_6t
Xbit_r92_c145 bl_145 br_145 wl_92 vdd gnd cell_6t
Xbit_r93_c145 bl_145 br_145 wl_93 vdd gnd cell_6t
Xbit_r94_c145 bl_145 br_145 wl_94 vdd gnd cell_6t
Xbit_r95_c145 bl_145 br_145 wl_95 vdd gnd cell_6t
Xbit_r96_c145 bl_145 br_145 wl_96 vdd gnd cell_6t
Xbit_r97_c145 bl_145 br_145 wl_97 vdd gnd cell_6t
Xbit_r98_c145 bl_145 br_145 wl_98 vdd gnd cell_6t
Xbit_r99_c145 bl_145 br_145 wl_99 vdd gnd cell_6t
Xbit_r100_c145 bl_145 br_145 wl_100 vdd gnd cell_6t
Xbit_r101_c145 bl_145 br_145 wl_101 vdd gnd cell_6t
Xbit_r102_c145 bl_145 br_145 wl_102 vdd gnd cell_6t
Xbit_r103_c145 bl_145 br_145 wl_103 vdd gnd cell_6t
Xbit_r104_c145 bl_145 br_145 wl_104 vdd gnd cell_6t
Xbit_r105_c145 bl_145 br_145 wl_105 vdd gnd cell_6t
Xbit_r106_c145 bl_145 br_145 wl_106 vdd gnd cell_6t
Xbit_r107_c145 bl_145 br_145 wl_107 vdd gnd cell_6t
Xbit_r108_c145 bl_145 br_145 wl_108 vdd gnd cell_6t
Xbit_r109_c145 bl_145 br_145 wl_109 vdd gnd cell_6t
Xbit_r110_c145 bl_145 br_145 wl_110 vdd gnd cell_6t
Xbit_r111_c145 bl_145 br_145 wl_111 vdd gnd cell_6t
Xbit_r112_c145 bl_145 br_145 wl_112 vdd gnd cell_6t
Xbit_r113_c145 bl_145 br_145 wl_113 vdd gnd cell_6t
Xbit_r114_c145 bl_145 br_145 wl_114 vdd gnd cell_6t
Xbit_r115_c145 bl_145 br_145 wl_115 vdd gnd cell_6t
Xbit_r116_c145 bl_145 br_145 wl_116 vdd gnd cell_6t
Xbit_r117_c145 bl_145 br_145 wl_117 vdd gnd cell_6t
Xbit_r118_c145 bl_145 br_145 wl_118 vdd gnd cell_6t
Xbit_r119_c145 bl_145 br_145 wl_119 vdd gnd cell_6t
Xbit_r120_c145 bl_145 br_145 wl_120 vdd gnd cell_6t
Xbit_r121_c145 bl_145 br_145 wl_121 vdd gnd cell_6t
Xbit_r122_c145 bl_145 br_145 wl_122 vdd gnd cell_6t
Xbit_r123_c145 bl_145 br_145 wl_123 vdd gnd cell_6t
Xbit_r124_c145 bl_145 br_145 wl_124 vdd gnd cell_6t
Xbit_r125_c145 bl_145 br_145 wl_125 vdd gnd cell_6t
Xbit_r126_c145 bl_145 br_145 wl_126 vdd gnd cell_6t
Xbit_r127_c145 bl_145 br_145 wl_127 vdd gnd cell_6t
Xbit_r128_c145 bl_145 br_145 wl_128 vdd gnd cell_6t
Xbit_r129_c145 bl_145 br_145 wl_129 vdd gnd cell_6t
Xbit_r130_c145 bl_145 br_145 wl_130 vdd gnd cell_6t
Xbit_r131_c145 bl_145 br_145 wl_131 vdd gnd cell_6t
Xbit_r132_c145 bl_145 br_145 wl_132 vdd gnd cell_6t
Xbit_r133_c145 bl_145 br_145 wl_133 vdd gnd cell_6t
Xbit_r134_c145 bl_145 br_145 wl_134 vdd gnd cell_6t
Xbit_r135_c145 bl_145 br_145 wl_135 vdd gnd cell_6t
Xbit_r136_c145 bl_145 br_145 wl_136 vdd gnd cell_6t
Xbit_r137_c145 bl_145 br_145 wl_137 vdd gnd cell_6t
Xbit_r138_c145 bl_145 br_145 wl_138 vdd gnd cell_6t
Xbit_r139_c145 bl_145 br_145 wl_139 vdd gnd cell_6t
Xbit_r140_c145 bl_145 br_145 wl_140 vdd gnd cell_6t
Xbit_r141_c145 bl_145 br_145 wl_141 vdd gnd cell_6t
Xbit_r142_c145 bl_145 br_145 wl_142 vdd gnd cell_6t
Xbit_r143_c145 bl_145 br_145 wl_143 vdd gnd cell_6t
Xbit_r144_c145 bl_145 br_145 wl_144 vdd gnd cell_6t
Xbit_r145_c145 bl_145 br_145 wl_145 vdd gnd cell_6t
Xbit_r146_c145 bl_145 br_145 wl_146 vdd gnd cell_6t
Xbit_r147_c145 bl_145 br_145 wl_147 vdd gnd cell_6t
Xbit_r148_c145 bl_145 br_145 wl_148 vdd gnd cell_6t
Xbit_r149_c145 bl_145 br_145 wl_149 vdd gnd cell_6t
Xbit_r150_c145 bl_145 br_145 wl_150 vdd gnd cell_6t
Xbit_r151_c145 bl_145 br_145 wl_151 vdd gnd cell_6t
Xbit_r152_c145 bl_145 br_145 wl_152 vdd gnd cell_6t
Xbit_r153_c145 bl_145 br_145 wl_153 vdd gnd cell_6t
Xbit_r154_c145 bl_145 br_145 wl_154 vdd gnd cell_6t
Xbit_r155_c145 bl_145 br_145 wl_155 vdd gnd cell_6t
Xbit_r156_c145 bl_145 br_145 wl_156 vdd gnd cell_6t
Xbit_r157_c145 bl_145 br_145 wl_157 vdd gnd cell_6t
Xbit_r158_c145 bl_145 br_145 wl_158 vdd gnd cell_6t
Xbit_r159_c145 bl_145 br_145 wl_159 vdd gnd cell_6t
Xbit_r160_c145 bl_145 br_145 wl_160 vdd gnd cell_6t
Xbit_r161_c145 bl_145 br_145 wl_161 vdd gnd cell_6t
Xbit_r162_c145 bl_145 br_145 wl_162 vdd gnd cell_6t
Xbit_r163_c145 bl_145 br_145 wl_163 vdd gnd cell_6t
Xbit_r164_c145 bl_145 br_145 wl_164 vdd gnd cell_6t
Xbit_r165_c145 bl_145 br_145 wl_165 vdd gnd cell_6t
Xbit_r166_c145 bl_145 br_145 wl_166 vdd gnd cell_6t
Xbit_r167_c145 bl_145 br_145 wl_167 vdd gnd cell_6t
Xbit_r168_c145 bl_145 br_145 wl_168 vdd gnd cell_6t
Xbit_r169_c145 bl_145 br_145 wl_169 vdd gnd cell_6t
Xbit_r170_c145 bl_145 br_145 wl_170 vdd gnd cell_6t
Xbit_r171_c145 bl_145 br_145 wl_171 vdd gnd cell_6t
Xbit_r172_c145 bl_145 br_145 wl_172 vdd gnd cell_6t
Xbit_r173_c145 bl_145 br_145 wl_173 vdd gnd cell_6t
Xbit_r174_c145 bl_145 br_145 wl_174 vdd gnd cell_6t
Xbit_r175_c145 bl_145 br_145 wl_175 vdd gnd cell_6t
Xbit_r176_c145 bl_145 br_145 wl_176 vdd gnd cell_6t
Xbit_r177_c145 bl_145 br_145 wl_177 vdd gnd cell_6t
Xbit_r178_c145 bl_145 br_145 wl_178 vdd gnd cell_6t
Xbit_r179_c145 bl_145 br_145 wl_179 vdd gnd cell_6t
Xbit_r180_c145 bl_145 br_145 wl_180 vdd gnd cell_6t
Xbit_r181_c145 bl_145 br_145 wl_181 vdd gnd cell_6t
Xbit_r182_c145 bl_145 br_145 wl_182 vdd gnd cell_6t
Xbit_r183_c145 bl_145 br_145 wl_183 vdd gnd cell_6t
Xbit_r184_c145 bl_145 br_145 wl_184 vdd gnd cell_6t
Xbit_r185_c145 bl_145 br_145 wl_185 vdd gnd cell_6t
Xbit_r186_c145 bl_145 br_145 wl_186 vdd gnd cell_6t
Xbit_r187_c145 bl_145 br_145 wl_187 vdd gnd cell_6t
Xbit_r188_c145 bl_145 br_145 wl_188 vdd gnd cell_6t
Xbit_r189_c145 bl_145 br_145 wl_189 vdd gnd cell_6t
Xbit_r190_c145 bl_145 br_145 wl_190 vdd gnd cell_6t
Xbit_r191_c145 bl_145 br_145 wl_191 vdd gnd cell_6t
Xbit_r192_c145 bl_145 br_145 wl_192 vdd gnd cell_6t
Xbit_r193_c145 bl_145 br_145 wl_193 vdd gnd cell_6t
Xbit_r194_c145 bl_145 br_145 wl_194 vdd gnd cell_6t
Xbit_r195_c145 bl_145 br_145 wl_195 vdd gnd cell_6t
Xbit_r196_c145 bl_145 br_145 wl_196 vdd gnd cell_6t
Xbit_r197_c145 bl_145 br_145 wl_197 vdd gnd cell_6t
Xbit_r198_c145 bl_145 br_145 wl_198 vdd gnd cell_6t
Xbit_r199_c145 bl_145 br_145 wl_199 vdd gnd cell_6t
Xbit_r200_c145 bl_145 br_145 wl_200 vdd gnd cell_6t
Xbit_r201_c145 bl_145 br_145 wl_201 vdd gnd cell_6t
Xbit_r202_c145 bl_145 br_145 wl_202 vdd gnd cell_6t
Xbit_r203_c145 bl_145 br_145 wl_203 vdd gnd cell_6t
Xbit_r204_c145 bl_145 br_145 wl_204 vdd gnd cell_6t
Xbit_r205_c145 bl_145 br_145 wl_205 vdd gnd cell_6t
Xbit_r206_c145 bl_145 br_145 wl_206 vdd gnd cell_6t
Xbit_r207_c145 bl_145 br_145 wl_207 vdd gnd cell_6t
Xbit_r208_c145 bl_145 br_145 wl_208 vdd gnd cell_6t
Xbit_r209_c145 bl_145 br_145 wl_209 vdd gnd cell_6t
Xbit_r210_c145 bl_145 br_145 wl_210 vdd gnd cell_6t
Xbit_r211_c145 bl_145 br_145 wl_211 vdd gnd cell_6t
Xbit_r212_c145 bl_145 br_145 wl_212 vdd gnd cell_6t
Xbit_r213_c145 bl_145 br_145 wl_213 vdd gnd cell_6t
Xbit_r214_c145 bl_145 br_145 wl_214 vdd gnd cell_6t
Xbit_r215_c145 bl_145 br_145 wl_215 vdd gnd cell_6t
Xbit_r216_c145 bl_145 br_145 wl_216 vdd gnd cell_6t
Xbit_r217_c145 bl_145 br_145 wl_217 vdd gnd cell_6t
Xbit_r218_c145 bl_145 br_145 wl_218 vdd gnd cell_6t
Xbit_r219_c145 bl_145 br_145 wl_219 vdd gnd cell_6t
Xbit_r220_c145 bl_145 br_145 wl_220 vdd gnd cell_6t
Xbit_r221_c145 bl_145 br_145 wl_221 vdd gnd cell_6t
Xbit_r222_c145 bl_145 br_145 wl_222 vdd gnd cell_6t
Xbit_r223_c145 bl_145 br_145 wl_223 vdd gnd cell_6t
Xbit_r224_c145 bl_145 br_145 wl_224 vdd gnd cell_6t
Xbit_r225_c145 bl_145 br_145 wl_225 vdd gnd cell_6t
Xbit_r226_c145 bl_145 br_145 wl_226 vdd gnd cell_6t
Xbit_r227_c145 bl_145 br_145 wl_227 vdd gnd cell_6t
Xbit_r228_c145 bl_145 br_145 wl_228 vdd gnd cell_6t
Xbit_r229_c145 bl_145 br_145 wl_229 vdd gnd cell_6t
Xbit_r230_c145 bl_145 br_145 wl_230 vdd gnd cell_6t
Xbit_r231_c145 bl_145 br_145 wl_231 vdd gnd cell_6t
Xbit_r232_c145 bl_145 br_145 wl_232 vdd gnd cell_6t
Xbit_r233_c145 bl_145 br_145 wl_233 vdd gnd cell_6t
Xbit_r234_c145 bl_145 br_145 wl_234 vdd gnd cell_6t
Xbit_r235_c145 bl_145 br_145 wl_235 vdd gnd cell_6t
Xbit_r236_c145 bl_145 br_145 wl_236 vdd gnd cell_6t
Xbit_r237_c145 bl_145 br_145 wl_237 vdd gnd cell_6t
Xbit_r238_c145 bl_145 br_145 wl_238 vdd gnd cell_6t
Xbit_r239_c145 bl_145 br_145 wl_239 vdd gnd cell_6t
Xbit_r240_c145 bl_145 br_145 wl_240 vdd gnd cell_6t
Xbit_r241_c145 bl_145 br_145 wl_241 vdd gnd cell_6t
Xbit_r242_c145 bl_145 br_145 wl_242 vdd gnd cell_6t
Xbit_r243_c145 bl_145 br_145 wl_243 vdd gnd cell_6t
Xbit_r244_c145 bl_145 br_145 wl_244 vdd gnd cell_6t
Xbit_r245_c145 bl_145 br_145 wl_245 vdd gnd cell_6t
Xbit_r246_c145 bl_145 br_145 wl_246 vdd gnd cell_6t
Xbit_r247_c145 bl_145 br_145 wl_247 vdd gnd cell_6t
Xbit_r248_c145 bl_145 br_145 wl_248 vdd gnd cell_6t
Xbit_r249_c145 bl_145 br_145 wl_249 vdd gnd cell_6t
Xbit_r250_c145 bl_145 br_145 wl_250 vdd gnd cell_6t
Xbit_r251_c145 bl_145 br_145 wl_251 vdd gnd cell_6t
Xbit_r252_c145 bl_145 br_145 wl_252 vdd gnd cell_6t
Xbit_r253_c145 bl_145 br_145 wl_253 vdd gnd cell_6t
Xbit_r254_c145 bl_145 br_145 wl_254 vdd gnd cell_6t
Xbit_r255_c145 bl_145 br_145 wl_255 vdd gnd cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd cell_6t
Xbit_r1_c146 bl_146 br_146 wl_1 vdd gnd cell_6t
Xbit_r2_c146 bl_146 br_146 wl_2 vdd gnd cell_6t
Xbit_r3_c146 bl_146 br_146 wl_3 vdd gnd cell_6t
Xbit_r4_c146 bl_146 br_146 wl_4 vdd gnd cell_6t
Xbit_r5_c146 bl_146 br_146 wl_5 vdd gnd cell_6t
Xbit_r6_c146 bl_146 br_146 wl_6 vdd gnd cell_6t
Xbit_r7_c146 bl_146 br_146 wl_7 vdd gnd cell_6t
Xbit_r8_c146 bl_146 br_146 wl_8 vdd gnd cell_6t
Xbit_r9_c146 bl_146 br_146 wl_9 vdd gnd cell_6t
Xbit_r10_c146 bl_146 br_146 wl_10 vdd gnd cell_6t
Xbit_r11_c146 bl_146 br_146 wl_11 vdd gnd cell_6t
Xbit_r12_c146 bl_146 br_146 wl_12 vdd gnd cell_6t
Xbit_r13_c146 bl_146 br_146 wl_13 vdd gnd cell_6t
Xbit_r14_c146 bl_146 br_146 wl_14 vdd gnd cell_6t
Xbit_r15_c146 bl_146 br_146 wl_15 vdd gnd cell_6t
Xbit_r16_c146 bl_146 br_146 wl_16 vdd gnd cell_6t
Xbit_r17_c146 bl_146 br_146 wl_17 vdd gnd cell_6t
Xbit_r18_c146 bl_146 br_146 wl_18 vdd gnd cell_6t
Xbit_r19_c146 bl_146 br_146 wl_19 vdd gnd cell_6t
Xbit_r20_c146 bl_146 br_146 wl_20 vdd gnd cell_6t
Xbit_r21_c146 bl_146 br_146 wl_21 vdd gnd cell_6t
Xbit_r22_c146 bl_146 br_146 wl_22 vdd gnd cell_6t
Xbit_r23_c146 bl_146 br_146 wl_23 vdd gnd cell_6t
Xbit_r24_c146 bl_146 br_146 wl_24 vdd gnd cell_6t
Xbit_r25_c146 bl_146 br_146 wl_25 vdd gnd cell_6t
Xbit_r26_c146 bl_146 br_146 wl_26 vdd gnd cell_6t
Xbit_r27_c146 bl_146 br_146 wl_27 vdd gnd cell_6t
Xbit_r28_c146 bl_146 br_146 wl_28 vdd gnd cell_6t
Xbit_r29_c146 bl_146 br_146 wl_29 vdd gnd cell_6t
Xbit_r30_c146 bl_146 br_146 wl_30 vdd gnd cell_6t
Xbit_r31_c146 bl_146 br_146 wl_31 vdd gnd cell_6t
Xbit_r32_c146 bl_146 br_146 wl_32 vdd gnd cell_6t
Xbit_r33_c146 bl_146 br_146 wl_33 vdd gnd cell_6t
Xbit_r34_c146 bl_146 br_146 wl_34 vdd gnd cell_6t
Xbit_r35_c146 bl_146 br_146 wl_35 vdd gnd cell_6t
Xbit_r36_c146 bl_146 br_146 wl_36 vdd gnd cell_6t
Xbit_r37_c146 bl_146 br_146 wl_37 vdd gnd cell_6t
Xbit_r38_c146 bl_146 br_146 wl_38 vdd gnd cell_6t
Xbit_r39_c146 bl_146 br_146 wl_39 vdd gnd cell_6t
Xbit_r40_c146 bl_146 br_146 wl_40 vdd gnd cell_6t
Xbit_r41_c146 bl_146 br_146 wl_41 vdd gnd cell_6t
Xbit_r42_c146 bl_146 br_146 wl_42 vdd gnd cell_6t
Xbit_r43_c146 bl_146 br_146 wl_43 vdd gnd cell_6t
Xbit_r44_c146 bl_146 br_146 wl_44 vdd gnd cell_6t
Xbit_r45_c146 bl_146 br_146 wl_45 vdd gnd cell_6t
Xbit_r46_c146 bl_146 br_146 wl_46 vdd gnd cell_6t
Xbit_r47_c146 bl_146 br_146 wl_47 vdd gnd cell_6t
Xbit_r48_c146 bl_146 br_146 wl_48 vdd gnd cell_6t
Xbit_r49_c146 bl_146 br_146 wl_49 vdd gnd cell_6t
Xbit_r50_c146 bl_146 br_146 wl_50 vdd gnd cell_6t
Xbit_r51_c146 bl_146 br_146 wl_51 vdd gnd cell_6t
Xbit_r52_c146 bl_146 br_146 wl_52 vdd gnd cell_6t
Xbit_r53_c146 bl_146 br_146 wl_53 vdd gnd cell_6t
Xbit_r54_c146 bl_146 br_146 wl_54 vdd gnd cell_6t
Xbit_r55_c146 bl_146 br_146 wl_55 vdd gnd cell_6t
Xbit_r56_c146 bl_146 br_146 wl_56 vdd gnd cell_6t
Xbit_r57_c146 bl_146 br_146 wl_57 vdd gnd cell_6t
Xbit_r58_c146 bl_146 br_146 wl_58 vdd gnd cell_6t
Xbit_r59_c146 bl_146 br_146 wl_59 vdd gnd cell_6t
Xbit_r60_c146 bl_146 br_146 wl_60 vdd gnd cell_6t
Xbit_r61_c146 bl_146 br_146 wl_61 vdd gnd cell_6t
Xbit_r62_c146 bl_146 br_146 wl_62 vdd gnd cell_6t
Xbit_r63_c146 bl_146 br_146 wl_63 vdd gnd cell_6t
Xbit_r64_c146 bl_146 br_146 wl_64 vdd gnd cell_6t
Xbit_r65_c146 bl_146 br_146 wl_65 vdd gnd cell_6t
Xbit_r66_c146 bl_146 br_146 wl_66 vdd gnd cell_6t
Xbit_r67_c146 bl_146 br_146 wl_67 vdd gnd cell_6t
Xbit_r68_c146 bl_146 br_146 wl_68 vdd gnd cell_6t
Xbit_r69_c146 bl_146 br_146 wl_69 vdd gnd cell_6t
Xbit_r70_c146 bl_146 br_146 wl_70 vdd gnd cell_6t
Xbit_r71_c146 bl_146 br_146 wl_71 vdd gnd cell_6t
Xbit_r72_c146 bl_146 br_146 wl_72 vdd gnd cell_6t
Xbit_r73_c146 bl_146 br_146 wl_73 vdd gnd cell_6t
Xbit_r74_c146 bl_146 br_146 wl_74 vdd gnd cell_6t
Xbit_r75_c146 bl_146 br_146 wl_75 vdd gnd cell_6t
Xbit_r76_c146 bl_146 br_146 wl_76 vdd gnd cell_6t
Xbit_r77_c146 bl_146 br_146 wl_77 vdd gnd cell_6t
Xbit_r78_c146 bl_146 br_146 wl_78 vdd gnd cell_6t
Xbit_r79_c146 bl_146 br_146 wl_79 vdd gnd cell_6t
Xbit_r80_c146 bl_146 br_146 wl_80 vdd gnd cell_6t
Xbit_r81_c146 bl_146 br_146 wl_81 vdd gnd cell_6t
Xbit_r82_c146 bl_146 br_146 wl_82 vdd gnd cell_6t
Xbit_r83_c146 bl_146 br_146 wl_83 vdd gnd cell_6t
Xbit_r84_c146 bl_146 br_146 wl_84 vdd gnd cell_6t
Xbit_r85_c146 bl_146 br_146 wl_85 vdd gnd cell_6t
Xbit_r86_c146 bl_146 br_146 wl_86 vdd gnd cell_6t
Xbit_r87_c146 bl_146 br_146 wl_87 vdd gnd cell_6t
Xbit_r88_c146 bl_146 br_146 wl_88 vdd gnd cell_6t
Xbit_r89_c146 bl_146 br_146 wl_89 vdd gnd cell_6t
Xbit_r90_c146 bl_146 br_146 wl_90 vdd gnd cell_6t
Xbit_r91_c146 bl_146 br_146 wl_91 vdd gnd cell_6t
Xbit_r92_c146 bl_146 br_146 wl_92 vdd gnd cell_6t
Xbit_r93_c146 bl_146 br_146 wl_93 vdd gnd cell_6t
Xbit_r94_c146 bl_146 br_146 wl_94 vdd gnd cell_6t
Xbit_r95_c146 bl_146 br_146 wl_95 vdd gnd cell_6t
Xbit_r96_c146 bl_146 br_146 wl_96 vdd gnd cell_6t
Xbit_r97_c146 bl_146 br_146 wl_97 vdd gnd cell_6t
Xbit_r98_c146 bl_146 br_146 wl_98 vdd gnd cell_6t
Xbit_r99_c146 bl_146 br_146 wl_99 vdd gnd cell_6t
Xbit_r100_c146 bl_146 br_146 wl_100 vdd gnd cell_6t
Xbit_r101_c146 bl_146 br_146 wl_101 vdd gnd cell_6t
Xbit_r102_c146 bl_146 br_146 wl_102 vdd gnd cell_6t
Xbit_r103_c146 bl_146 br_146 wl_103 vdd gnd cell_6t
Xbit_r104_c146 bl_146 br_146 wl_104 vdd gnd cell_6t
Xbit_r105_c146 bl_146 br_146 wl_105 vdd gnd cell_6t
Xbit_r106_c146 bl_146 br_146 wl_106 vdd gnd cell_6t
Xbit_r107_c146 bl_146 br_146 wl_107 vdd gnd cell_6t
Xbit_r108_c146 bl_146 br_146 wl_108 vdd gnd cell_6t
Xbit_r109_c146 bl_146 br_146 wl_109 vdd gnd cell_6t
Xbit_r110_c146 bl_146 br_146 wl_110 vdd gnd cell_6t
Xbit_r111_c146 bl_146 br_146 wl_111 vdd gnd cell_6t
Xbit_r112_c146 bl_146 br_146 wl_112 vdd gnd cell_6t
Xbit_r113_c146 bl_146 br_146 wl_113 vdd gnd cell_6t
Xbit_r114_c146 bl_146 br_146 wl_114 vdd gnd cell_6t
Xbit_r115_c146 bl_146 br_146 wl_115 vdd gnd cell_6t
Xbit_r116_c146 bl_146 br_146 wl_116 vdd gnd cell_6t
Xbit_r117_c146 bl_146 br_146 wl_117 vdd gnd cell_6t
Xbit_r118_c146 bl_146 br_146 wl_118 vdd gnd cell_6t
Xbit_r119_c146 bl_146 br_146 wl_119 vdd gnd cell_6t
Xbit_r120_c146 bl_146 br_146 wl_120 vdd gnd cell_6t
Xbit_r121_c146 bl_146 br_146 wl_121 vdd gnd cell_6t
Xbit_r122_c146 bl_146 br_146 wl_122 vdd gnd cell_6t
Xbit_r123_c146 bl_146 br_146 wl_123 vdd gnd cell_6t
Xbit_r124_c146 bl_146 br_146 wl_124 vdd gnd cell_6t
Xbit_r125_c146 bl_146 br_146 wl_125 vdd gnd cell_6t
Xbit_r126_c146 bl_146 br_146 wl_126 vdd gnd cell_6t
Xbit_r127_c146 bl_146 br_146 wl_127 vdd gnd cell_6t
Xbit_r128_c146 bl_146 br_146 wl_128 vdd gnd cell_6t
Xbit_r129_c146 bl_146 br_146 wl_129 vdd gnd cell_6t
Xbit_r130_c146 bl_146 br_146 wl_130 vdd gnd cell_6t
Xbit_r131_c146 bl_146 br_146 wl_131 vdd gnd cell_6t
Xbit_r132_c146 bl_146 br_146 wl_132 vdd gnd cell_6t
Xbit_r133_c146 bl_146 br_146 wl_133 vdd gnd cell_6t
Xbit_r134_c146 bl_146 br_146 wl_134 vdd gnd cell_6t
Xbit_r135_c146 bl_146 br_146 wl_135 vdd gnd cell_6t
Xbit_r136_c146 bl_146 br_146 wl_136 vdd gnd cell_6t
Xbit_r137_c146 bl_146 br_146 wl_137 vdd gnd cell_6t
Xbit_r138_c146 bl_146 br_146 wl_138 vdd gnd cell_6t
Xbit_r139_c146 bl_146 br_146 wl_139 vdd gnd cell_6t
Xbit_r140_c146 bl_146 br_146 wl_140 vdd gnd cell_6t
Xbit_r141_c146 bl_146 br_146 wl_141 vdd gnd cell_6t
Xbit_r142_c146 bl_146 br_146 wl_142 vdd gnd cell_6t
Xbit_r143_c146 bl_146 br_146 wl_143 vdd gnd cell_6t
Xbit_r144_c146 bl_146 br_146 wl_144 vdd gnd cell_6t
Xbit_r145_c146 bl_146 br_146 wl_145 vdd gnd cell_6t
Xbit_r146_c146 bl_146 br_146 wl_146 vdd gnd cell_6t
Xbit_r147_c146 bl_146 br_146 wl_147 vdd gnd cell_6t
Xbit_r148_c146 bl_146 br_146 wl_148 vdd gnd cell_6t
Xbit_r149_c146 bl_146 br_146 wl_149 vdd gnd cell_6t
Xbit_r150_c146 bl_146 br_146 wl_150 vdd gnd cell_6t
Xbit_r151_c146 bl_146 br_146 wl_151 vdd gnd cell_6t
Xbit_r152_c146 bl_146 br_146 wl_152 vdd gnd cell_6t
Xbit_r153_c146 bl_146 br_146 wl_153 vdd gnd cell_6t
Xbit_r154_c146 bl_146 br_146 wl_154 vdd gnd cell_6t
Xbit_r155_c146 bl_146 br_146 wl_155 vdd gnd cell_6t
Xbit_r156_c146 bl_146 br_146 wl_156 vdd gnd cell_6t
Xbit_r157_c146 bl_146 br_146 wl_157 vdd gnd cell_6t
Xbit_r158_c146 bl_146 br_146 wl_158 vdd gnd cell_6t
Xbit_r159_c146 bl_146 br_146 wl_159 vdd gnd cell_6t
Xbit_r160_c146 bl_146 br_146 wl_160 vdd gnd cell_6t
Xbit_r161_c146 bl_146 br_146 wl_161 vdd gnd cell_6t
Xbit_r162_c146 bl_146 br_146 wl_162 vdd gnd cell_6t
Xbit_r163_c146 bl_146 br_146 wl_163 vdd gnd cell_6t
Xbit_r164_c146 bl_146 br_146 wl_164 vdd gnd cell_6t
Xbit_r165_c146 bl_146 br_146 wl_165 vdd gnd cell_6t
Xbit_r166_c146 bl_146 br_146 wl_166 vdd gnd cell_6t
Xbit_r167_c146 bl_146 br_146 wl_167 vdd gnd cell_6t
Xbit_r168_c146 bl_146 br_146 wl_168 vdd gnd cell_6t
Xbit_r169_c146 bl_146 br_146 wl_169 vdd gnd cell_6t
Xbit_r170_c146 bl_146 br_146 wl_170 vdd gnd cell_6t
Xbit_r171_c146 bl_146 br_146 wl_171 vdd gnd cell_6t
Xbit_r172_c146 bl_146 br_146 wl_172 vdd gnd cell_6t
Xbit_r173_c146 bl_146 br_146 wl_173 vdd gnd cell_6t
Xbit_r174_c146 bl_146 br_146 wl_174 vdd gnd cell_6t
Xbit_r175_c146 bl_146 br_146 wl_175 vdd gnd cell_6t
Xbit_r176_c146 bl_146 br_146 wl_176 vdd gnd cell_6t
Xbit_r177_c146 bl_146 br_146 wl_177 vdd gnd cell_6t
Xbit_r178_c146 bl_146 br_146 wl_178 vdd gnd cell_6t
Xbit_r179_c146 bl_146 br_146 wl_179 vdd gnd cell_6t
Xbit_r180_c146 bl_146 br_146 wl_180 vdd gnd cell_6t
Xbit_r181_c146 bl_146 br_146 wl_181 vdd gnd cell_6t
Xbit_r182_c146 bl_146 br_146 wl_182 vdd gnd cell_6t
Xbit_r183_c146 bl_146 br_146 wl_183 vdd gnd cell_6t
Xbit_r184_c146 bl_146 br_146 wl_184 vdd gnd cell_6t
Xbit_r185_c146 bl_146 br_146 wl_185 vdd gnd cell_6t
Xbit_r186_c146 bl_146 br_146 wl_186 vdd gnd cell_6t
Xbit_r187_c146 bl_146 br_146 wl_187 vdd gnd cell_6t
Xbit_r188_c146 bl_146 br_146 wl_188 vdd gnd cell_6t
Xbit_r189_c146 bl_146 br_146 wl_189 vdd gnd cell_6t
Xbit_r190_c146 bl_146 br_146 wl_190 vdd gnd cell_6t
Xbit_r191_c146 bl_146 br_146 wl_191 vdd gnd cell_6t
Xbit_r192_c146 bl_146 br_146 wl_192 vdd gnd cell_6t
Xbit_r193_c146 bl_146 br_146 wl_193 vdd gnd cell_6t
Xbit_r194_c146 bl_146 br_146 wl_194 vdd gnd cell_6t
Xbit_r195_c146 bl_146 br_146 wl_195 vdd gnd cell_6t
Xbit_r196_c146 bl_146 br_146 wl_196 vdd gnd cell_6t
Xbit_r197_c146 bl_146 br_146 wl_197 vdd gnd cell_6t
Xbit_r198_c146 bl_146 br_146 wl_198 vdd gnd cell_6t
Xbit_r199_c146 bl_146 br_146 wl_199 vdd gnd cell_6t
Xbit_r200_c146 bl_146 br_146 wl_200 vdd gnd cell_6t
Xbit_r201_c146 bl_146 br_146 wl_201 vdd gnd cell_6t
Xbit_r202_c146 bl_146 br_146 wl_202 vdd gnd cell_6t
Xbit_r203_c146 bl_146 br_146 wl_203 vdd gnd cell_6t
Xbit_r204_c146 bl_146 br_146 wl_204 vdd gnd cell_6t
Xbit_r205_c146 bl_146 br_146 wl_205 vdd gnd cell_6t
Xbit_r206_c146 bl_146 br_146 wl_206 vdd gnd cell_6t
Xbit_r207_c146 bl_146 br_146 wl_207 vdd gnd cell_6t
Xbit_r208_c146 bl_146 br_146 wl_208 vdd gnd cell_6t
Xbit_r209_c146 bl_146 br_146 wl_209 vdd gnd cell_6t
Xbit_r210_c146 bl_146 br_146 wl_210 vdd gnd cell_6t
Xbit_r211_c146 bl_146 br_146 wl_211 vdd gnd cell_6t
Xbit_r212_c146 bl_146 br_146 wl_212 vdd gnd cell_6t
Xbit_r213_c146 bl_146 br_146 wl_213 vdd gnd cell_6t
Xbit_r214_c146 bl_146 br_146 wl_214 vdd gnd cell_6t
Xbit_r215_c146 bl_146 br_146 wl_215 vdd gnd cell_6t
Xbit_r216_c146 bl_146 br_146 wl_216 vdd gnd cell_6t
Xbit_r217_c146 bl_146 br_146 wl_217 vdd gnd cell_6t
Xbit_r218_c146 bl_146 br_146 wl_218 vdd gnd cell_6t
Xbit_r219_c146 bl_146 br_146 wl_219 vdd gnd cell_6t
Xbit_r220_c146 bl_146 br_146 wl_220 vdd gnd cell_6t
Xbit_r221_c146 bl_146 br_146 wl_221 vdd gnd cell_6t
Xbit_r222_c146 bl_146 br_146 wl_222 vdd gnd cell_6t
Xbit_r223_c146 bl_146 br_146 wl_223 vdd gnd cell_6t
Xbit_r224_c146 bl_146 br_146 wl_224 vdd gnd cell_6t
Xbit_r225_c146 bl_146 br_146 wl_225 vdd gnd cell_6t
Xbit_r226_c146 bl_146 br_146 wl_226 vdd gnd cell_6t
Xbit_r227_c146 bl_146 br_146 wl_227 vdd gnd cell_6t
Xbit_r228_c146 bl_146 br_146 wl_228 vdd gnd cell_6t
Xbit_r229_c146 bl_146 br_146 wl_229 vdd gnd cell_6t
Xbit_r230_c146 bl_146 br_146 wl_230 vdd gnd cell_6t
Xbit_r231_c146 bl_146 br_146 wl_231 vdd gnd cell_6t
Xbit_r232_c146 bl_146 br_146 wl_232 vdd gnd cell_6t
Xbit_r233_c146 bl_146 br_146 wl_233 vdd gnd cell_6t
Xbit_r234_c146 bl_146 br_146 wl_234 vdd gnd cell_6t
Xbit_r235_c146 bl_146 br_146 wl_235 vdd gnd cell_6t
Xbit_r236_c146 bl_146 br_146 wl_236 vdd gnd cell_6t
Xbit_r237_c146 bl_146 br_146 wl_237 vdd gnd cell_6t
Xbit_r238_c146 bl_146 br_146 wl_238 vdd gnd cell_6t
Xbit_r239_c146 bl_146 br_146 wl_239 vdd gnd cell_6t
Xbit_r240_c146 bl_146 br_146 wl_240 vdd gnd cell_6t
Xbit_r241_c146 bl_146 br_146 wl_241 vdd gnd cell_6t
Xbit_r242_c146 bl_146 br_146 wl_242 vdd gnd cell_6t
Xbit_r243_c146 bl_146 br_146 wl_243 vdd gnd cell_6t
Xbit_r244_c146 bl_146 br_146 wl_244 vdd gnd cell_6t
Xbit_r245_c146 bl_146 br_146 wl_245 vdd gnd cell_6t
Xbit_r246_c146 bl_146 br_146 wl_246 vdd gnd cell_6t
Xbit_r247_c146 bl_146 br_146 wl_247 vdd gnd cell_6t
Xbit_r248_c146 bl_146 br_146 wl_248 vdd gnd cell_6t
Xbit_r249_c146 bl_146 br_146 wl_249 vdd gnd cell_6t
Xbit_r250_c146 bl_146 br_146 wl_250 vdd gnd cell_6t
Xbit_r251_c146 bl_146 br_146 wl_251 vdd gnd cell_6t
Xbit_r252_c146 bl_146 br_146 wl_252 vdd gnd cell_6t
Xbit_r253_c146 bl_146 br_146 wl_253 vdd gnd cell_6t
Xbit_r254_c146 bl_146 br_146 wl_254 vdd gnd cell_6t
Xbit_r255_c146 bl_146 br_146 wl_255 vdd gnd cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd cell_6t
Xbit_r1_c147 bl_147 br_147 wl_1 vdd gnd cell_6t
Xbit_r2_c147 bl_147 br_147 wl_2 vdd gnd cell_6t
Xbit_r3_c147 bl_147 br_147 wl_3 vdd gnd cell_6t
Xbit_r4_c147 bl_147 br_147 wl_4 vdd gnd cell_6t
Xbit_r5_c147 bl_147 br_147 wl_5 vdd gnd cell_6t
Xbit_r6_c147 bl_147 br_147 wl_6 vdd gnd cell_6t
Xbit_r7_c147 bl_147 br_147 wl_7 vdd gnd cell_6t
Xbit_r8_c147 bl_147 br_147 wl_8 vdd gnd cell_6t
Xbit_r9_c147 bl_147 br_147 wl_9 vdd gnd cell_6t
Xbit_r10_c147 bl_147 br_147 wl_10 vdd gnd cell_6t
Xbit_r11_c147 bl_147 br_147 wl_11 vdd gnd cell_6t
Xbit_r12_c147 bl_147 br_147 wl_12 vdd gnd cell_6t
Xbit_r13_c147 bl_147 br_147 wl_13 vdd gnd cell_6t
Xbit_r14_c147 bl_147 br_147 wl_14 vdd gnd cell_6t
Xbit_r15_c147 bl_147 br_147 wl_15 vdd gnd cell_6t
Xbit_r16_c147 bl_147 br_147 wl_16 vdd gnd cell_6t
Xbit_r17_c147 bl_147 br_147 wl_17 vdd gnd cell_6t
Xbit_r18_c147 bl_147 br_147 wl_18 vdd gnd cell_6t
Xbit_r19_c147 bl_147 br_147 wl_19 vdd gnd cell_6t
Xbit_r20_c147 bl_147 br_147 wl_20 vdd gnd cell_6t
Xbit_r21_c147 bl_147 br_147 wl_21 vdd gnd cell_6t
Xbit_r22_c147 bl_147 br_147 wl_22 vdd gnd cell_6t
Xbit_r23_c147 bl_147 br_147 wl_23 vdd gnd cell_6t
Xbit_r24_c147 bl_147 br_147 wl_24 vdd gnd cell_6t
Xbit_r25_c147 bl_147 br_147 wl_25 vdd gnd cell_6t
Xbit_r26_c147 bl_147 br_147 wl_26 vdd gnd cell_6t
Xbit_r27_c147 bl_147 br_147 wl_27 vdd gnd cell_6t
Xbit_r28_c147 bl_147 br_147 wl_28 vdd gnd cell_6t
Xbit_r29_c147 bl_147 br_147 wl_29 vdd gnd cell_6t
Xbit_r30_c147 bl_147 br_147 wl_30 vdd gnd cell_6t
Xbit_r31_c147 bl_147 br_147 wl_31 vdd gnd cell_6t
Xbit_r32_c147 bl_147 br_147 wl_32 vdd gnd cell_6t
Xbit_r33_c147 bl_147 br_147 wl_33 vdd gnd cell_6t
Xbit_r34_c147 bl_147 br_147 wl_34 vdd gnd cell_6t
Xbit_r35_c147 bl_147 br_147 wl_35 vdd gnd cell_6t
Xbit_r36_c147 bl_147 br_147 wl_36 vdd gnd cell_6t
Xbit_r37_c147 bl_147 br_147 wl_37 vdd gnd cell_6t
Xbit_r38_c147 bl_147 br_147 wl_38 vdd gnd cell_6t
Xbit_r39_c147 bl_147 br_147 wl_39 vdd gnd cell_6t
Xbit_r40_c147 bl_147 br_147 wl_40 vdd gnd cell_6t
Xbit_r41_c147 bl_147 br_147 wl_41 vdd gnd cell_6t
Xbit_r42_c147 bl_147 br_147 wl_42 vdd gnd cell_6t
Xbit_r43_c147 bl_147 br_147 wl_43 vdd gnd cell_6t
Xbit_r44_c147 bl_147 br_147 wl_44 vdd gnd cell_6t
Xbit_r45_c147 bl_147 br_147 wl_45 vdd gnd cell_6t
Xbit_r46_c147 bl_147 br_147 wl_46 vdd gnd cell_6t
Xbit_r47_c147 bl_147 br_147 wl_47 vdd gnd cell_6t
Xbit_r48_c147 bl_147 br_147 wl_48 vdd gnd cell_6t
Xbit_r49_c147 bl_147 br_147 wl_49 vdd gnd cell_6t
Xbit_r50_c147 bl_147 br_147 wl_50 vdd gnd cell_6t
Xbit_r51_c147 bl_147 br_147 wl_51 vdd gnd cell_6t
Xbit_r52_c147 bl_147 br_147 wl_52 vdd gnd cell_6t
Xbit_r53_c147 bl_147 br_147 wl_53 vdd gnd cell_6t
Xbit_r54_c147 bl_147 br_147 wl_54 vdd gnd cell_6t
Xbit_r55_c147 bl_147 br_147 wl_55 vdd gnd cell_6t
Xbit_r56_c147 bl_147 br_147 wl_56 vdd gnd cell_6t
Xbit_r57_c147 bl_147 br_147 wl_57 vdd gnd cell_6t
Xbit_r58_c147 bl_147 br_147 wl_58 vdd gnd cell_6t
Xbit_r59_c147 bl_147 br_147 wl_59 vdd gnd cell_6t
Xbit_r60_c147 bl_147 br_147 wl_60 vdd gnd cell_6t
Xbit_r61_c147 bl_147 br_147 wl_61 vdd gnd cell_6t
Xbit_r62_c147 bl_147 br_147 wl_62 vdd gnd cell_6t
Xbit_r63_c147 bl_147 br_147 wl_63 vdd gnd cell_6t
Xbit_r64_c147 bl_147 br_147 wl_64 vdd gnd cell_6t
Xbit_r65_c147 bl_147 br_147 wl_65 vdd gnd cell_6t
Xbit_r66_c147 bl_147 br_147 wl_66 vdd gnd cell_6t
Xbit_r67_c147 bl_147 br_147 wl_67 vdd gnd cell_6t
Xbit_r68_c147 bl_147 br_147 wl_68 vdd gnd cell_6t
Xbit_r69_c147 bl_147 br_147 wl_69 vdd gnd cell_6t
Xbit_r70_c147 bl_147 br_147 wl_70 vdd gnd cell_6t
Xbit_r71_c147 bl_147 br_147 wl_71 vdd gnd cell_6t
Xbit_r72_c147 bl_147 br_147 wl_72 vdd gnd cell_6t
Xbit_r73_c147 bl_147 br_147 wl_73 vdd gnd cell_6t
Xbit_r74_c147 bl_147 br_147 wl_74 vdd gnd cell_6t
Xbit_r75_c147 bl_147 br_147 wl_75 vdd gnd cell_6t
Xbit_r76_c147 bl_147 br_147 wl_76 vdd gnd cell_6t
Xbit_r77_c147 bl_147 br_147 wl_77 vdd gnd cell_6t
Xbit_r78_c147 bl_147 br_147 wl_78 vdd gnd cell_6t
Xbit_r79_c147 bl_147 br_147 wl_79 vdd gnd cell_6t
Xbit_r80_c147 bl_147 br_147 wl_80 vdd gnd cell_6t
Xbit_r81_c147 bl_147 br_147 wl_81 vdd gnd cell_6t
Xbit_r82_c147 bl_147 br_147 wl_82 vdd gnd cell_6t
Xbit_r83_c147 bl_147 br_147 wl_83 vdd gnd cell_6t
Xbit_r84_c147 bl_147 br_147 wl_84 vdd gnd cell_6t
Xbit_r85_c147 bl_147 br_147 wl_85 vdd gnd cell_6t
Xbit_r86_c147 bl_147 br_147 wl_86 vdd gnd cell_6t
Xbit_r87_c147 bl_147 br_147 wl_87 vdd gnd cell_6t
Xbit_r88_c147 bl_147 br_147 wl_88 vdd gnd cell_6t
Xbit_r89_c147 bl_147 br_147 wl_89 vdd gnd cell_6t
Xbit_r90_c147 bl_147 br_147 wl_90 vdd gnd cell_6t
Xbit_r91_c147 bl_147 br_147 wl_91 vdd gnd cell_6t
Xbit_r92_c147 bl_147 br_147 wl_92 vdd gnd cell_6t
Xbit_r93_c147 bl_147 br_147 wl_93 vdd gnd cell_6t
Xbit_r94_c147 bl_147 br_147 wl_94 vdd gnd cell_6t
Xbit_r95_c147 bl_147 br_147 wl_95 vdd gnd cell_6t
Xbit_r96_c147 bl_147 br_147 wl_96 vdd gnd cell_6t
Xbit_r97_c147 bl_147 br_147 wl_97 vdd gnd cell_6t
Xbit_r98_c147 bl_147 br_147 wl_98 vdd gnd cell_6t
Xbit_r99_c147 bl_147 br_147 wl_99 vdd gnd cell_6t
Xbit_r100_c147 bl_147 br_147 wl_100 vdd gnd cell_6t
Xbit_r101_c147 bl_147 br_147 wl_101 vdd gnd cell_6t
Xbit_r102_c147 bl_147 br_147 wl_102 vdd gnd cell_6t
Xbit_r103_c147 bl_147 br_147 wl_103 vdd gnd cell_6t
Xbit_r104_c147 bl_147 br_147 wl_104 vdd gnd cell_6t
Xbit_r105_c147 bl_147 br_147 wl_105 vdd gnd cell_6t
Xbit_r106_c147 bl_147 br_147 wl_106 vdd gnd cell_6t
Xbit_r107_c147 bl_147 br_147 wl_107 vdd gnd cell_6t
Xbit_r108_c147 bl_147 br_147 wl_108 vdd gnd cell_6t
Xbit_r109_c147 bl_147 br_147 wl_109 vdd gnd cell_6t
Xbit_r110_c147 bl_147 br_147 wl_110 vdd gnd cell_6t
Xbit_r111_c147 bl_147 br_147 wl_111 vdd gnd cell_6t
Xbit_r112_c147 bl_147 br_147 wl_112 vdd gnd cell_6t
Xbit_r113_c147 bl_147 br_147 wl_113 vdd gnd cell_6t
Xbit_r114_c147 bl_147 br_147 wl_114 vdd gnd cell_6t
Xbit_r115_c147 bl_147 br_147 wl_115 vdd gnd cell_6t
Xbit_r116_c147 bl_147 br_147 wl_116 vdd gnd cell_6t
Xbit_r117_c147 bl_147 br_147 wl_117 vdd gnd cell_6t
Xbit_r118_c147 bl_147 br_147 wl_118 vdd gnd cell_6t
Xbit_r119_c147 bl_147 br_147 wl_119 vdd gnd cell_6t
Xbit_r120_c147 bl_147 br_147 wl_120 vdd gnd cell_6t
Xbit_r121_c147 bl_147 br_147 wl_121 vdd gnd cell_6t
Xbit_r122_c147 bl_147 br_147 wl_122 vdd gnd cell_6t
Xbit_r123_c147 bl_147 br_147 wl_123 vdd gnd cell_6t
Xbit_r124_c147 bl_147 br_147 wl_124 vdd gnd cell_6t
Xbit_r125_c147 bl_147 br_147 wl_125 vdd gnd cell_6t
Xbit_r126_c147 bl_147 br_147 wl_126 vdd gnd cell_6t
Xbit_r127_c147 bl_147 br_147 wl_127 vdd gnd cell_6t
Xbit_r128_c147 bl_147 br_147 wl_128 vdd gnd cell_6t
Xbit_r129_c147 bl_147 br_147 wl_129 vdd gnd cell_6t
Xbit_r130_c147 bl_147 br_147 wl_130 vdd gnd cell_6t
Xbit_r131_c147 bl_147 br_147 wl_131 vdd gnd cell_6t
Xbit_r132_c147 bl_147 br_147 wl_132 vdd gnd cell_6t
Xbit_r133_c147 bl_147 br_147 wl_133 vdd gnd cell_6t
Xbit_r134_c147 bl_147 br_147 wl_134 vdd gnd cell_6t
Xbit_r135_c147 bl_147 br_147 wl_135 vdd gnd cell_6t
Xbit_r136_c147 bl_147 br_147 wl_136 vdd gnd cell_6t
Xbit_r137_c147 bl_147 br_147 wl_137 vdd gnd cell_6t
Xbit_r138_c147 bl_147 br_147 wl_138 vdd gnd cell_6t
Xbit_r139_c147 bl_147 br_147 wl_139 vdd gnd cell_6t
Xbit_r140_c147 bl_147 br_147 wl_140 vdd gnd cell_6t
Xbit_r141_c147 bl_147 br_147 wl_141 vdd gnd cell_6t
Xbit_r142_c147 bl_147 br_147 wl_142 vdd gnd cell_6t
Xbit_r143_c147 bl_147 br_147 wl_143 vdd gnd cell_6t
Xbit_r144_c147 bl_147 br_147 wl_144 vdd gnd cell_6t
Xbit_r145_c147 bl_147 br_147 wl_145 vdd gnd cell_6t
Xbit_r146_c147 bl_147 br_147 wl_146 vdd gnd cell_6t
Xbit_r147_c147 bl_147 br_147 wl_147 vdd gnd cell_6t
Xbit_r148_c147 bl_147 br_147 wl_148 vdd gnd cell_6t
Xbit_r149_c147 bl_147 br_147 wl_149 vdd gnd cell_6t
Xbit_r150_c147 bl_147 br_147 wl_150 vdd gnd cell_6t
Xbit_r151_c147 bl_147 br_147 wl_151 vdd gnd cell_6t
Xbit_r152_c147 bl_147 br_147 wl_152 vdd gnd cell_6t
Xbit_r153_c147 bl_147 br_147 wl_153 vdd gnd cell_6t
Xbit_r154_c147 bl_147 br_147 wl_154 vdd gnd cell_6t
Xbit_r155_c147 bl_147 br_147 wl_155 vdd gnd cell_6t
Xbit_r156_c147 bl_147 br_147 wl_156 vdd gnd cell_6t
Xbit_r157_c147 bl_147 br_147 wl_157 vdd gnd cell_6t
Xbit_r158_c147 bl_147 br_147 wl_158 vdd gnd cell_6t
Xbit_r159_c147 bl_147 br_147 wl_159 vdd gnd cell_6t
Xbit_r160_c147 bl_147 br_147 wl_160 vdd gnd cell_6t
Xbit_r161_c147 bl_147 br_147 wl_161 vdd gnd cell_6t
Xbit_r162_c147 bl_147 br_147 wl_162 vdd gnd cell_6t
Xbit_r163_c147 bl_147 br_147 wl_163 vdd gnd cell_6t
Xbit_r164_c147 bl_147 br_147 wl_164 vdd gnd cell_6t
Xbit_r165_c147 bl_147 br_147 wl_165 vdd gnd cell_6t
Xbit_r166_c147 bl_147 br_147 wl_166 vdd gnd cell_6t
Xbit_r167_c147 bl_147 br_147 wl_167 vdd gnd cell_6t
Xbit_r168_c147 bl_147 br_147 wl_168 vdd gnd cell_6t
Xbit_r169_c147 bl_147 br_147 wl_169 vdd gnd cell_6t
Xbit_r170_c147 bl_147 br_147 wl_170 vdd gnd cell_6t
Xbit_r171_c147 bl_147 br_147 wl_171 vdd gnd cell_6t
Xbit_r172_c147 bl_147 br_147 wl_172 vdd gnd cell_6t
Xbit_r173_c147 bl_147 br_147 wl_173 vdd gnd cell_6t
Xbit_r174_c147 bl_147 br_147 wl_174 vdd gnd cell_6t
Xbit_r175_c147 bl_147 br_147 wl_175 vdd gnd cell_6t
Xbit_r176_c147 bl_147 br_147 wl_176 vdd gnd cell_6t
Xbit_r177_c147 bl_147 br_147 wl_177 vdd gnd cell_6t
Xbit_r178_c147 bl_147 br_147 wl_178 vdd gnd cell_6t
Xbit_r179_c147 bl_147 br_147 wl_179 vdd gnd cell_6t
Xbit_r180_c147 bl_147 br_147 wl_180 vdd gnd cell_6t
Xbit_r181_c147 bl_147 br_147 wl_181 vdd gnd cell_6t
Xbit_r182_c147 bl_147 br_147 wl_182 vdd gnd cell_6t
Xbit_r183_c147 bl_147 br_147 wl_183 vdd gnd cell_6t
Xbit_r184_c147 bl_147 br_147 wl_184 vdd gnd cell_6t
Xbit_r185_c147 bl_147 br_147 wl_185 vdd gnd cell_6t
Xbit_r186_c147 bl_147 br_147 wl_186 vdd gnd cell_6t
Xbit_r187_c147 bl_147 br_147 wl_187 vdd gnd cell_6t
Xbit_r188_c147 bl_147 br_147 wl_188 vdd gnd cell_6t
Xbit_r189_c147 bl_147 br_147 wl_189 vdd gnd cell_6t
Xbit_r190_c147 bl_147 br_147 wl_190 vdd gnd cell_6t
Xbit_r191_c147 bl_147 br_147 wl_191 vdd gnd cell_6t
Xbit_r192_c147 bl_147 br_147 wl_192 vdd gnd cell_6t
Xbit_r193_c147 bl_147 br_147 wl_193 vdd gnd cell_6t
Xbit_r194_c147 bl_147 br_147 wl_194 vdd gnd cell_6t
Xbit_r195_c147 bl_147 br_147 wl_195 vdd gnd cell_6t
Xbit_r196_c147 bl_147 br_147 wl_196 vdd gnd cell_6t
Xbit_r197_c147 bl_147 br_147 wl_197 vdd gnd cell_6t
Xbit_r198_c147 bl_147 br_147 wl_198 vdd gnd cell_6t
Xbit_r199_c147 bl_147 br_147 wl_199 vdd gnd cell_6t
Xbit_r200_c147 bl_147 br_147 wl_200 vdd gnd cell_6t
Xbit_r201_c147 bl_147 br_147 wl_201 vdd gnd cell_6t
Xbit_r202_c147 bl_147 br_147 wl_202 vdd gnd cell_6t
Xbit_r203_c147 bl_147 br_147 wl_203 vdd gnd cell_6t
Xbit_r204_c147 bl_147 br_147 wl_204 vdd gnd cell_6t
Xbit_r205_c147 bl_147 br_147 wl_205 vdd gnd cell_6t
Xbit_r206_c147 bl_147 br_147 wl_206 vdd gnd cell_6t
Xbit_r207_c147 bl_147 br_147 wl_207 vdd gnd cell_6t
Xbit_r208_c147 bl_147 br_147 wl_208 vdd gnd cell_6t
Xbit_r209_c147 bl_147 br_147 wl_209 vdd gnd cell_6t
Xbit_r210_c147 bl_147 br_147 wl_210 vdd gnd cell_6t
Xbit_r211_c147 bl_147 br_147 wl_211 vdd gnd cell_6t
Xbit_r212_c147 bl_147 br_147 wl_212 vdd gnd cell_6t
Xbit_r213_c147 bl_147 br_147 wl_213 vdd gnd cell_6t
Xbit_r214_c147 bl_147 br_147 wl_214 vdd gnd cell_6t
Xbit_r215_c147 bl_147 br_147 wl_215 vdd gnd cell_6t
Xbit_r216_c147 bl_147 br_147 wl_216 vdd gnd cell_6t
Xbit_r217_c147 bl_147 br_147 wl_217 vdd gnd cell_6t
Xbit_r218_c147 bl_147 br_147 wl_218 vdd gnd cell_6t
Xbit_r219_c147 bl_147 br_147 wl_219 vdd gnd cell_6t
Xbit_r220_c147 bl_147 br_147 wl_220 vdd gnd cell_6t
Xbit_r221_c147 bl_147 br_147 wl_221 vdd gnd cell_6t
Xbit_r222_c147 bl_147 br_147 wl_222 vdd gnd cell_6t
Xbit_r223_c147 bl_147 br_147 wl_223 vdd gnd cell_6t
Xbit_r224_c147 bl_147 br_147 wl_224 vdd gnd cell_6t
Xbit_r225_c147 bl_147 br_147 wl_225 vdd gnd cell_6t
Xbit_r226_c147 bl_147 br_147 wl_226 vdd gnd cell_6t
Xbit_r227_c147 bl_147 br_147 wl_227 vdd gnd cell_6t
Xbit_r228_c147 bl_147 br_147 wl_228 vdd gnd cell_6t
Xbit_r229_c147 bl_147 br_147 wl_229 vdd gnd cell_6t
Xbit_r230_c147 bl_147 br_147 wl_230 vdd gnd cell_6t
Xbit_r231_c147 bl_147 br_147 wl_231 vdd gnd cell_6t
Xbit_r232_c147 bl_147 br_147 wl_232 vdd gnd cell_6t
Xbit_r233_c147 bl_147 br_147 wl_233 vdd gnd cell_6t
Xbit_r234_c147 bl_147 br_147 wl_234 vdd gnd cell_6t
Xbit_r235_c147 bl_147 br_147 wl_235 vdd gnd cell_6t
Xbit_r236_c147 bl_147 br_147 wl_236 vdd gnd cell_6t
Xbit_r237_c147 bl_147 br_147 wl_237 vdd gnd cell_6t
Xbit_r238_c147 bl_147 br_147 wl_238 vdd gnd cell_6t
Xbit_r239_c147 bl_147 br_147 wl_239 vdd gnd cell_6t
Xbit_r240_c147 bl_147 br_147 wl_240 vdd gnd cell_6t
Xbit_r241_c147 bl_147 br_147 wl_241 vdd gnd cell_6t
Xbit_r242_c147 bl_147 br_147 wl_242 vdd gnd cell_6t
Xbit_r243_c147 bl_147 br_147 wl_243 vdd gnd cell_6t
Xbit_r244_c147 bl_147 br_147 wl_244 vdd gnd cell_6t
Xbit_r245_c147 bl_147 br_147 wl_245 vdd gnd cell_6t
Xbit_r246_c147 bl_147 br_147 wl_246 vdd gnd cell_6t
Xbit_r247_c147 bl_147 br_147 wl_247 vdd gnd cell_6t
Xbit_r248_c147 bl_147 br_147 wl_248 vdd gnd cell_6t
Xbit_r249_c147 bl_147 br_147 wl_249 vdd gnd cell_6t
Xbit_r250_c147 bl_147 br_147 wl_250 vdd gnd cell_6t
Xbit_r251_c147 bl_147 br_147 wl_251 vdd gnd cell_6t
Xbit_r252_c147 bl_147 br_147 wl_252 vdd gnd cell_6t
Xbit_r253_c147 bl_147 br_147 wl_253 vdd gnd cell_6t
Xbit_r254_c147 bl_147 br_147 wl_254 vdd gnd cell_6t
Xbit_r255_c147 bl_147 br_147 wl_255 vdd gnd cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd cell_6t
Xbit_r1_c148 bl_148 br_148 wl_1 vdd gnd cell_6t
Xbit_r2_c148 bl_148 br_148 wl_2 vdd gnd cell_6t
Xbit_r3_c148 bl_148 br_148 wl_3 vdd gnd cell_6t
Xbit_r4_c148 bl_148 br_148 wl_4 vdd gnd cell_6t
Xbit_r5_c148 bl_148 br_148 wl_5 vdd gnd cell_6t
Xbit_r6_c148 bl_148 br_148 wl_6 vdd gnd cell_6t
Xbit_r7_c148 bl_148 br_148 wl_7 vdd gnd cell_6t
Xbit_r8_c148 bl_148 br_148 wl_8 vdd gnd cell_6t
Xbit_r9_c148 bl_148 br_148 wl_9 vdd gnd cell_6t
Xbit_r10_c148 bl_148 br_148 wl_10 vdd gnd cell_6t
Xbit_r11_c148 bl_148 br_148 wl_11 vdd gnd cell_6t
Xbit_r12_c148 bl_148 br_148 wl_12 vdd gnd cell_6t
Xbit_r13_c148 bl_148 br_148 wl_13 vdd gnd cell_6t
Xbit_r14_c148 bl_148 br_148 wl_14 vdd gnd cell_6t
Xbit_r15_c148 bl_148 br_148 wl_15 vdd gnd cell_6t
Xbit_r16_c148 bl_148 br_148 wl_16 vdd gnd cell_6t
Xbit_r17_c148 bl_148 br_148 wl_17 vdd gnd cell_6t
Xbit_r18_c148 bl_148 br_148 wl_18 vdd gnd cell_6t
Xbit_r19_c148 bl_148 br_148 wl_19 vdd gnd cell_6t
Xbit_r20_c148 bl_148 br_148 wl_20 vdd gnd cell_6t
Xbit_r21_c148 bl_148 br_148 wl_21 vdd gnd cell_6t
Xbit_r22_c148 bl_148 br_148 wl_22 vdd gnd cell_6t
Xbit_r23_c148 bl_148 br_148 wl_23 vdd gnd cell_6t
Xbit_r24_c148 bl_148 br_148 wl_24 vdd gnd cell_6t
Xbit_r25_c148 bl_148 br_148 wl_25 vdd gnd cell_6t
Xbit_r26_c148 bl_148 br_148 wl_26 vdd gnd cell_6t
Xbit_r27_c148 bl_148 br_148 wl_27 vdd gnd cell_6t
Xbit_r28_c148 bl_148 br_148 wl_28 vdd gnd cell_6t
Xbit_r29_c148 bl_148 br_148 wl_29 vdd gnd cell_6t
Xbit_r30_c148 bl_148 br_148 wl_30 vdd gnd cell_6t
Xbit_r31_c148 bl_148 br_148 wl_31 vdd gnd cell_6t
Xbit_r32_c148 bl_148 br_148 wl_32 vdd gnd cell_6t
Xbit_r33_c148 bl_148 br_148 wl_33 vdd gnd cell_6t
Xbit_r34_c148 bl_148 br_148 wl_34 vdd gnd cell_6t
Xbit_r35_c148 bl_148 br_148 wl_35 vdd gnd cell_6t
Xbit_r36_c148 bl_148 br_148 wl_36 vdd gnd cell_6t
Xbit_r37_c148 bl_148 br_148 wl_37 vdd gnd cell_6t
Xbit_r38_c148 bl_148 br_148 wl_38 vdd gnd cell_6t
Xbit_r39_c148 bl_148 br_148 wl_39 vdd gnd cell_6t
Xbit_r40_c148 bl_148 br_148 wl_40 vdd gnd cell_6t
Xbit_r41_c148 bl_148 br_148 wl_41 vdd gnd cell_6t
Xbit_r42_c148 bl_148 br_148 wl_42 vdd gnd cell_6t
Xbit_r43_c148 bl_148 br_148 wl_43 vdd gnd cell_6t
Xbit_r44_c148 bl_148 br_148 wl_44 vdd gnd cell_6t
Xbit_r45_c148 bl_148 br_148 wl_45 vdd gnd cell_6t
Xbit_r46_c148 bl_148 br_148 wl_46 vdd gnd cell_6t
Xbit_r47_c148 bl_148 br_148 wl_47 vdd gnd cell_6t
Xbit_r48_c148 bl_148 br_148 wl_48 vdd gnd cell_6t
Xbit_r49_c148 bl_148 br_148 wl_49 vdd gnd cell_6t
Xbit_r50_c148 bl_148 br_148 wl_50 vdd gnd cell_6t
Xbit_r51_c148 bl_148 br_148 wl_51 vdd gnd cell_6t
Xbit_r52_c148 bl_148 br_148 wl_52 vdd gnd cell_6t
Xbit_r53_c148 bl_148 br_148 wl_53 vdd gnd cell_6t
Xbit_r54_c148 bl_148 br_148 wl_54 vdd gnd cell_6t
Xbit_r55_c148 bl_148 br_148 wl_55 vdd gnd cell_6t
Xbit_r56_c148 bl_148 br_148 wl_56 vdd gnd cell_6t
Xbit_r57_c148 bl_148 br_148 wl_57 vdd gnd cell_6t
Xbit_r58_c148 bl_148 br_148 wl_58 vdd gnd cell_6t
Xbit_r59_c148 bl_148 br_148 wl_59 vdd gnd cell_6t
Xbit_r60_c148 bl_148 br_148 wl_60 vdd gnd cell_6t
Xbit_r61_c148 bl_148 br_148 wl_61 vdd gnd cell_6t
Xbit_r62_c148 bl_148 br_148 wl_62 vdd gnd cell_6t
Xbit_r63_c148 bl_148 br_148 wl_63 vdd gnd cell_6t
Xbit_r64_c148 bl_148 br_148 wl_64 vdd gnd cell_6t
Xbit_r65_c148 bl_148 br_148 wl_65 vdd gnd cell_6t
Xbit_r66_c148 bl_148 br_148 wl_66 vdd gnd cell_6t
Xbit_r67_c148 bl_148 br_148 wl_67 vdd gnd cell_6t
Xbit_r68_c148 bl_148 br_148 wl_68 vdd gnd cell_6t
Xbit_r69_c148 bl_148 br_148 wl_69 vdd gnd cell_6t
Xbit_r70_c148 bl_148 br_148 wl_70 vdd gnd cell_6t
Xbit_r71_c148 bl_148 br_148 wl_71 vdd gnd cell_6t
Xbit_r72_c148 bl_148 br_148 wl_72 vdd gnd cell_6t
Xbit_r73_c148 bl_148 br_148 wl_73 vdd gnd cell_6t
Xbit_r74_c148 bl_148 br_148 wl_74 vdd gnd cell_6t
Xbit_r75_c148 bl_148 br_148 wl_75 vdd gnd cell_6t
Xbit_r76_c148 bl_148 br_148 wl_76 vdd gnd cell_6t
Xbit_r77_c148 bl_148 br_148 wl_77 vdd gnd cell_6t
Xbit_r78_c148 bl_148 br_148 wl_78 vdd gnd cell_6t
Xbit_r79_c148 bl_148 br_148 wl_79 vdd gnd cell_6t
Xbit_r80_c148 bl_148 br_148 wl_80 vdd gnd cell_6t
Xbit_r81_c148 bl_148 br_148 wl_81 vdd gnd cell_6t
Xbit_r82_c148 bl_148 br_148 wl_82 vdd gnd cell_6t
Xbit_r83_c148 bl_148 br_148 wl_83 vdd gnd cell_6t
Xbit_r84_c148 bl_148 br_148 wl_84 vdd gnd cell_6t
Xbit_r85_c148 bl_148 br_148 wl_85 vdd gnd cell_6t
Xbit_r86_c148 bl_148 br_148 wl_86 vdd gnd cell_6t
Xbit_r87_c148 bl_148 br_148 wl_87 vdd gnd cell_6t
Xbit_r88_c148 bl_148 br_148 wl_88 vdd gnd cell_6t
Xbit_r89_c148 bl_148 br_148 wl_89 vdd gnd cell_6t
Xbit_r90_c148 bl_148 br_148 wl_90 vdd gnd cell_6t
Xbit_r91_c148 bl_148 br_148 wl_91 vdd gnd cell_6t
Xbit_r92_c148 bl_148 br_148 wl_92 vdd gnd cell_6t
Xbit_r93_c148 bl_148 br_148 wl_93 vdd gnd cell_6t
Xbit_r94_c148 bl_148 br_148 wl_94 vdd gnd cell_6t
Xbit_r95_c148 bl_148 br_148 wl_95 vdd gnd cell_6t
Xbit_r96_c148 bl_148 br_148 wl_96 vdd gnd cell_6t
Xbit_r97_c148 bl_148 br_148 wl_97 vdd gnd cell_6t
Xbit_r98_c148 bl_148 br_148 wl_98 vdd gnd cell_6t
Xbit_r99_c148 bl_148 br_148 wl_99 vdd gnd cell_6t
Xbit_r100_c148 bl_148 br_148 wl_100 vdd gnd cell_6t
Xbit_r101_c148 bl_148 br_148 wl_101 vdd gnd cell_6t
Xbit_r102_c148 bl_148 br_148 wl_102 vdd gnd cell_6t
Xbit_r103_c148 bl_148 br_148 wl_103 vdd gnd cell_6t
Xbit_r104_c148 bl_148 br_148 wl_104 vdd gnd cell_6t
Xbit_r105_c148 bl_148 br_148 wl_105 vdd gnd cell_6t
Xbit_r106_c148 bl_148 br_148 wl_106 vdd gnd cell_6t
Xbit_r107_c148 bl_148 br_148 wl_107 vdd gnd cell_6t
Xbit_r108_c148 bl_148 br_148 wl_108 vdd gnd cell_6t
Xbit_r109_c148 bl_148 br_148 wl_109 vdd gnd cell_6t
Xbit_r110_c148 bl_148 br_148 wl_110 vdd gnd cell_6t
Xbit_r111_c148 bl_148 br_148 wl_111 vdd gnd cell_6t
Xbit_r112_c148 bl_148 br_148 wl_112 vdd gnd cell_6t
Xbit_r113_c148 bl_148 br_148 wl_113 vdd gnd cell_6t
Xbit_r114_c148 bl_148 br_148 wl_114 vdd gnd cell_6t
Xbit_r115_c148 bl_148 br_148 wl_115 vdd gnd cell_6t
Xbit_r116_c148 bl_148 br_148 wl_116 vdd gnd cell_6t
Xbit_r117_c148 bl_148 br_148 wl_117 vdd gnd cell_6t
Xbit_r118_c148 bl_148 br_148 wl_118 vdd gnd cell_6t
Xbit_r119_c148 bl_148 br_148 wl_119 vdd gnd cell_6t
Xbit_r120_c148 bl_148 br_148 wl_120 vdd gnd cell_6t
Xbit_r121_c148 bl_148 br_148 wl_121 vdd gnd cell_6t
Xbit_r122_c148 bl_148 br_148 wl_122 vdd gnd cell_6t
Xbit_r123_c148 bl_148 br_148 wl_123 vdd gnd cell_6t
Xbit_r124_c148 bl_148 br_148 wl_124 vdd gnd cell_6t
Xbit_r125_c148 bl_148 br_148 wl_125 vdd gnd cell_6t
Xbit_r126_c148 bl_148 br_148 wl_126 vdd gnd cell_6t
Xbit_r127_c148 bl_148 br_148 wl_127 vdd gnd cell_6t
Xbit_r128_c148 bl_148 br_148 wl_128 vdd gnd cell_6t
Xbit_r129_c148 bl_148 br_148 wl_129 vdd gnd cell_6t
Xbit_r130_c148 bl_148 br_148 wl_130 vdd gnd cell_6t
Xbit_r131_c148 bl_148 br_148 wl_131 vdd gnd cell_6t
Xbit_r132_c148 bl_148 br_148 wl_132 vdd gnd cell_6t
Xbit_r133_c148 bl_148 br_148 wl_133 vdd gnd cell_6t
Xbit_r134_c148 bl_148 br_148 wl_134 vdd gnd cell_6t
Xbit_r135_c148 bl_148 br_148 wl_135 vdd gnd cell_6t
Xbit_r136_c148 bl_148 br_148 wl_136 vdd gnd cell_6t
Xbit_r137_c148 bl_148 br_148 wl_137 vdd gnd cell_6t
Xbit_r138_c148 bl_148 br_148 wl_138 vdd gnd cell_6t
Xbit_r139_c148 bl_148 br_148 wl_139 vdd gnd cell_6t
Xbit_r140_c148 bl_148 br_148 wl_140 vdd gnd cell_6t
Xbit_r141_c148 bl_148 br_148 wl_141 vdd gnd cell_6t
Xbit_r142_c148 bl_148 br_148 wl_142 vdd gnd cell_6t
Xbit_r143_c148 bl_148 br_148 wl_143 vdd gnd cell_6t
Xbit_r144_c148 bl_148 br_148 wl_144 vdd gnd cell_6t
Xbit_r145_c148 bl_148 br_148 wl_145 vdd gnd cell_6t
Xbit_r146_c148 bl_148 br_148 wl_146 vdd gnd cell_6t
Xbit_r147_c148 bl_148 br_148 wl_147 vdd gnd cell_6t
Xbit_r148_c148 bl_148 br_148 wl_148 vdd gnd cell_6t
Xbit_r149_c148 bl_148 br_148 wl_149 vdd gnd cell_6t
Xbit_r150_c148 bl_148 br_148 wl_150 vdd gnd cell_6t
Xbit_r151_c148 bl_148 br_148 wl_151 vdd gnd cell_6t
Xbit_r152_c148 bl_148 br_148 wl_152 vdd gnd cell_6t
Xbit_r153_c148 bl_148 br_148 wl_153 vdd gnd cell_6t
Xbit_r154_c148 bl_148 br_148 wl_154 vdd gnd cell_6t
Xbit_r155_c148 bl_148 br_148 wl_155 vdd gnd cell_6t
Xbit_r156_c148 bl_148 br_148 wl_156 vdd gnd cell_6t
Xbit_r157_c148 bl_148 br_148 wl_157 vdd gnd cell_6t
Xbit_r158_c148 bl_148 br_148 wl_158 vdd gnd cell_6t
Xbit_r159_c148 bl_148 br_148 wl_159 vdd gnd cell_6t
Xbit_r160_c148 bl_148 br_148 wl_160 vdd gnd cell_6t
Xbit_r161_c148 bl_148 br_148 wl_161 vdd gnd cell_6t
Xbit_r162_c148 bl_148 br_148 wl_162 vdd gnd cell_6t
Xbit_r163_c148 bl_148 br_148 wl_163 vdd gnd cell_6t
Xbit_r164_c148 bl_148 br_148 wl_164 vdd gnd cell_6t
Xbit_r165_c148 bl_148 br_148 wl_165 vdd gnd cell_6t
Xbit_r166_c148 bl_148 br_148 wl_166 vdd gnd cell_6t
Xbit_r167_c148 bl_148 br_148 wl_167 vdd gnd cell_6t
Xbit_r168_c148 bl_148 br_148 wl_168 vdd gnd cell_6t
Xbit_r169_c148 bl_148 br_148 wl_169 vdd gnd cell_6t
Xbit_r170_c148 bl_148 br_148 wl_170 vdd gnd cell_6t
Xbit_r171_c148 bl_148 br_148 wl_171 vdd gnd cell_6t
Xbit_r172_c148 bl_148 br_148 wl_172 vdd gnd cell_6t
Xbit_r173_c148 bl_148 br_148 wl_173 vdd gnd cell_6t
Xbit_r174_c148 bl_148 br_148 wl_174 vdd gnd cell_6t
Xbit_r175_c148 bl_148 br_148 wl_175 vdd gnd cell_6t
Xbit_r176_c148 bl_148 br_148 wl_176 vdd gnd cell_6t
Xbit_r177_c148 bl_148 br_148 wl_177 vdd gnd cell_6t
Xbit_r178_c148 bl_148 br_148 wl_178 vdd gnd cell_6t
Xbit_r179_c148 bl_148 br_148 wl_179 vdd gnd cell_6t
Xbit_r180_c148 bl_148 br_148 wl_180 vdd gnd cell_6t
Xbit_r181_c148 bl_148 br_148 wl_181 vdd gnd cell_6t
Xbit_r182_c148 bl_148 br_148 wl_182 vdd gnd cell_6t
Xbit_r183_c148 bl_148 br_148 wl_183 vdd gnd cell_6t
Xbit_r184_c148 bl_148 br_148 wl_184 vdd gnd cell_6t
Xbit_r185_c148 bl_148 br_148 wl_185 vdd gnd cell_6t
Xbit_r186_c148 bl_148 br_148 wl_186 vdd gnd cell_6t
Xbit_r187_c148 bl_148 br_148 wl_187 vdd gnd cell_6t
Xbit_r188_c148 bl_148 br_148 wl_188 vdd gnd cell_6t
Xbit_r189_c148 bl_148 br_148 wl_189 vdd gnd cell_6t
Xbit_r190_c148 bl_148 br_148 wl_190 vdd gnd cell_6t
Xbit_r191_c148 bl_148 br_148 wl_191 vdd gnd cell_6t
Xbit_r192_c148 bl_148 br_148 wl_192 vdd gnd cell_6t
Xbit_r193_c148 bl_148 br_148 wl_193 vdd gnd cell_6t
Xbit_r194_c148 bl_148 br_148 wl_194 vdd gnd cell_6t
Xbit_r195_c148 bl_148 br_148 wl_195 vdd gnd cell_6t
Xbit_r196_c148 bl_148 br_148 wl_196 vdd gnd cell_6t
Xbit_r197_c148 bl_148 br_148 wl_197 vdd gnd cell_6t
Xbit_r198_c148 bl_148 br_148 wl_198 vdd gnd cell_6t
Xbit_r199_c148 bl_148 br_148 wl_199 vdd gnd cell_6t
Xbit_r200_c148 bl_148 br_148 wl_200 vdd gnd cell_6t
Xbit_r201_c148 bl_148 br_148 wl_201 vdd gnd cell_6t
Xbit_r202_c148 bl_148 br_148 wl_202 vdd gnd cell_6t
Xbit_r203_c148 bl_148 br_148 wl_203 vdd gnd cell_6t
Xbit_r204_c148 bl_148 br_148 wl_204 vdd gnd cell_6t
Xbit_r205_c148 bl_148 br_148 wl_205 vdd gnd cell_6t
Xbit_r206_c148 bl_148 br_148 wl_206 vdd gnd cell_6t
Xbit_r207_c148 bl_148 br_148 wl_207 vdd gnd cell_6t
Xbit_r208_c148 bl_148 br_148 wl_208 vdd gnd cell_6t
Xbit_r209_c148 bl_148 br_148 wl_209 vdd gnd cell_6t
Xbit_r210_c148 bl_148 br_148 wl_210 vdd gnd cell_6t
Xbit_r211_c148 bl_148 br_148 wl_211 vdd gnd cell_6t
Xbit_r212_c148 bl_148 br_148 wl_212 vdd gnd cell_6t
Xbit_r213_c148 bl_148 br_148 wl_213 vdd gnd cell_6t
Xbit_r214_c148 bl_148 br_148 wl_214 vdd gnd cell_6t
Xbit_r215_c148 bl_148 br_148 wl_215 vdd gnd cell_6t
Xbit_r216_c148 bl_148 br_148 wl_216 vdd gnd cell_6t
Xbit_r217_c148 bl_148 br_148 wl_217 vdd gnd cell_6t
Xbit_r218_c148 bl_148 br_148 wl_218 vdd gnd cell_6t
Xbit_r219_c148 bl_148 br_148 wl_219 vdd gnd cell_6t
Xbit_r220_c148 bl_148 br_148 wl_220 vdd gnd cell_6t
Xbit_r221_c148 bl_148 br_148 wl_221 vdd gnd cell_6t
Xbit_r222_c148 bl_148 br_148 wl_222 vdd gnd cell_6t
Xbit_r223_c148 bl_148 br_148 wl_223 vdd gnd cell_6t
Xbit_r224_c148 bl_148 br_148 wl_224 vdd gnd cell_6t
Xbit_r225_c148 bl_148 br_148 wl_225 vdd gnd cell_6t
Xbit_r226_c148 bl_148 br_148 wl_226 vdd gnd cell_6t
Xbit_r227_c148 bl_148 br_148 wl_227 vdd gnd cell_6t
Xbit_r228_c148 bl_148 br_148 wl_228 vdd gnd cell_6t
Xbit_r229_c148 bl_148 br_148 wl_229 vdd gnd cell_6t
Xbit_r230_c148 bl_148 br_148 wl_230 vdd gnd cell_6t
Xbit_r231_c148 bl_148 br_148 wl_231 vdd gnd cell_6t
Xbit_r232_c148 bl_148 br_148 wl_232 vdd gnd cell_6t
Xbit_r233_c148 bl_148 br_148 wl_233 vdd gnd cell_6t
Xbit_r234_c148 bl_148 br_148 wl_234 vdd gnd cell_6t
Xbit_r235_c148 bl_148 br_148 wl_235 vdd gnd cell_6t
Xbit_r236_c148 bl_148 br_148 wl_236 vdd gnd cell_6t
Xbit_r237_c148 bl_148 br_148 wl_237 vdd gnd cell_6t
Xbit_r238_c148 bl_148 br_148 wl_238 vdd gnd cell_6t
Xbit_r239_c148 bl_148 br_148 wl_239 vdd gnd cell_6t
Xbit_r240_c148 bl_148 br_148 wl_240 vdd gnd cell_6t
Xbit_r241_c148 bl_148 br_148 wl_241 vdd gnd cell_6t
Xbit_r242_c148 bl_148 br_148 wl_242 vdd gnd cell_6t
Xbit_r243_c148 bl_148 br_148 wl_243 vdd gnd cell_6t
Xbit_r244_c148 bl_148 br_148 wl_244 vdd gnd cell_6t
Xbit_r245_c148 bl_148 br_148 wl_245 vdd gnd cell_6t
Xbit_r246_c148 bl_148 br_148 wl_246 vdd gnd cell_6t
Xbit_r247_c148 bl_148 br_148 wl_247 vdd gnd cell_6t
Xbit_r248_c148 bl_148 br_148 wl_248 vdd gnd cell_6t
Xbit_r249_c148 bl_148 br_148 wl_249 vdd gnd cell_6t
Xbit_r250_c148 bl_148 br_148 wl_250 vdd gnd cell_6t
Xbit_r251_c148 bl_148 br_148 wl_251 vdd gnd cell_6t
Xbit_r252_c148 bl_148 br_148 wl_252 vdd gnd cell_6t
Xbit_r253_c148 bl_148 br_148 wl_253 vdd gnd cell_6t
Xbit_r254_c148 bl_148 br_148 wl_254 vdd gnd cell_6t
Xbit_r255_c148 bl_148 br_148 wl_255 vdd gnd cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd cell_6t
Xbit_r1_c149 bl_149 br_149 wl_1 vdd gnd cell_6t
Xbit_r2_c149 bl_149 br_149 wl_2 vdd gnd cell_6t
Xbit_r3_c149 bl_149 br_149 wl_3 vdd gnd cell_6t
Xbit_r4_c149 bl_149 br_149 wl_4 vdd gnd cell_6t
Xbit_r5_c149 bl_149 br_149 wl_5 vdd gnd cell_6t
Xbit_r6_c149 bl_149 br_149 wl_6 vdd gnd cell_6t
Xbit_r7_c149 bl_149 br_149 wl_7 vdd gnd cell_6t
Xbit_r8_c149 bl_149 br_149 wl_8 vdd gnd cell_6t
Xbit_r9_c149 bl_149 br_149 wl_9 vdd gnd cell_6t
Xbit_r10_c149 bl_149 br_149 wl_10 vdd gnd cell_6t
Xbit_r11_c149 bl_149 br_149 wl_11 vdd gnd cell_6t
Xbit_r12_c149 bl_149 br_149 wl_12 vdd gnd cell_6t
Xbit_r13_c149 bl_149 br_149 wl_13 vdd gnd cell_6t
Xbit_r14_c149 bl_149 br_149 wl_14 vdd gnd cell_6t
Xbit_r15_c149 bl_149 br_149 wl_15 vdd gnd cell_6t
Xbit_r16_c149 bl_149 br_149 wl_16 vdd gnd cell_6t
Xbit_r17_c149 bl_149 br_149 wl_17 vdd gnd cell_6t
Xbit_r18_c149 bl_149 br_149 wl_18 vdd gnd cell_6t
Xbit_r19_c149 bl_149 br_149 wl_19 vdd gnd cell_6t
Xbit_r20_c149 bl_149 br_149 wl_20 vdd gnd cell_6t
Xbit_r21_c149 bl_149 br_149 wl_21 vdd gnd cell_6t
Xbit_r22_c149 bl_149 br_149 wl_22 vdd gnd cell_6t
Xbit_r23_c149 bl_149 br_149 wl_23 vdd gnd cell_6t
Xbit_r24_c149 bl_149 br_149 wl_24 vdd gnd cell_6t
Xbit_r25_c149 bl_149 br_149 wl_25 vdd gnd cell_6t
Xbit_r26_c149 bl_149 br_149 wl_26 vdd gnd cell_6t
Xbit_r27_c149 bl_149 br_149 wl_27 vdd gnd cell_6t
Xbit_r28_c149 bl_149 br_149 wl_28 vdd gnd cell_6t
Xbit_r29_c149 bl_149 br_149 wl_29 vdd gnd cell_6t
Xbit_r30_c149 bl_149 br_149 wl_30 vdd gnd cell_6t
Xbit_r31_c149 bl_149 br_149 wl_31 vdd gnd cell_6t
Xbit_r32_c149 bl_149 br_149 wl_32 vdd gnd cell_6t
Xbit_r33_c149 bl_149 br_149 wl_33 vdd gnd cell_6t
Xbit_r34_c149 bl_149 br_149 wl_34 vdd gnd cell_6t
Xbit_r35_c149 bl_149 br_149 wl_35 vdd gnd cell_6t
Xbit_r36_c149 bl_149 br_149 wl_36 vdd gnd cell_6t
Xbit_r37_c149 bl_149 br_149 wl_37 vdd gnd cell_6t
Xbit_r38_c149 bl_149 br_149 wl_38 vdd gnd cell_6t
Xbit_r39_c149 bl_149 br_149 wl_39 vdd gnd cell_6t
Xbit_r40_c149 bl_149 br_149 wl_40 vdd gnd cell_6t
Xbit_r41_c149 bl_149 br_149 wl_41 vdd gnd cell_6t
Xbit_r42_c149 bl_149 br_149 wl_42 vdd gnd cell_6t
Xbit_r43_c149 bl_149 br_149 wl_43 vdd gnd cell_6t
Xbit_r44_c149 bl_149 br_149 wl_44 vdd gnd cell_6t
Xbit_r45_c149 bl_149 br_149 wl_45 vdd gnd cell_6t
Xbit_r46_c149 bl_149 br_149 wl_46 vdd gnd cell_6t
Xbit_r47_c149 bl_149 br_149 wl_47 vdd gnd cell_6t
Xbit_r48_c149 bl_149 br_149 wl_48 vdd gnd cell_6t
Xbit_r49_c149 bl_149 br_149 wl_49 vdd gnd cell_6t
Xbit_r50_c149 bl_149 br_149 wl_50 vdd gnd cell_6t
Xbit_r51_c149 bl_149 br_149 wl_51 vdd gnd cell_6t
Xbit_r52_c149 bl_149 br_149 wl_52 vdd gnd cell_6t
Xbit_r53_c149 bl_149 br_149 wl_53 vdd gnd cell_6t
Xbit_r54_c149 bl_149 br_149 wl_54 vdd gnd cell_6t
Xbit_r55_c149 bl_149 br_149 wl_55 vdd gnd cell_6t
Xbit_r56_c149 bl_149 br_149 wl_56 vdd gnd cell_6t
Xbit_r57_c149 bl_149 br_149 wl_57 vdd gnd cell_6t
Xbit_r58_c149 bl_149 br_149 wl_58 vdd gnd cell_6t
Xbit_r59_c149 bl_149 br_149 wl_59 vdd gnd cell_6t
Xbit_r60_c149 bl_149 br_149 wl_60 vdd gnd cell_6t
Xbit_r61_c149 bl_149 br_149 wl_61 vdd gnd cell_6t
Xbit_r62_c149 bl_149 br_149 wl_62 vdd gnd cell_6t
Xbit_r63_c149 bl_149 br_149 wl_63 vdd gnd cell_6t
Xbit_r64_c149 bl_149 br_149 wl_64 vdd gnd cell_6t
Xbit_r65_c149 bl_149 br_149 wl_65 vdd gnd cell_6t
Xbit_r66_c149 bl_149 br_149 wl_66 vdd gnd cell_6t
Xbit_r67_c149 bl_149 br_149 wl_67 vdd gnd cell_6t
Xbit_r68_c149 bl_149 br_149 wl_68 vdd gnd cell_6t
Xbit_r69_c149 bl_149 br_149 wl_69 vdd gnd cell_6t
Xbit_r70_c149 bl_149 br_149 wl_70 vdd gnd cell_6t
Xbit_r71_c149 bl_149 br_149 wl_71 vdd gnd cell_6t
Xbit_r72_c149 bl_149 br_149 wl_72 vdd gnd cell_6t
Xbit_r73_c149 bl_149 br_149 wl_73 vdd gnd cell_6t
Xbit_r74_c149 bl_149 br_149 wl_74 vdd gnd cell_6t
Xbit_r75_c149 bl_149 br_149 wl_75 vdd gnd cell_6t
Xbit_r76_c149 bl_149 br_149 wl_76 vdd gnd cell_6t
Xbit_r77_c149 bl_149 br_149 wl_77 vdd gnd cell_6t
Xbit_r78_c149 bl_149 br_149 wl_78 vdd gnd cell_6t
Xbit_r79_c149 bl_149 br_149 wl_79 vdd gnd cell_6t
Xbit_r80_c149 bl_149 br_149 wl_80 vdd gnd cell_6t
Xbit_r81_c149 bl_149 br_149 wl_81 vdd gnd cell_6t
Xbit_r82_c149 bl_149 br_149 wl_82 vdd gnd cell_6t
Xbit_r83_c149 bl_149 br_149 wl_83 vdd gnd cell_6t
Xbit_r84_c149 bl_149 br_149 wl_84 vdd gnd cell_6t
Xbit_r85_c149 bl_149 br_149 wl_85 vdd gnd cell_6t
Xbit_r86_c149 bl_149 br_149 wl_86 vdd gnd cell_6t
Xbit_r87_c149 bl_149 br_149 wl_87 vdd gnd cell_6t
Xbit_r88_c149 bl_149 br_149 wl_88 vdd gnd cell_6t
Xbit_r89_c149 bl_149 br_149 wl_89 vdd gnd cell_6t
Xbit_r90_c149 bl_149 br_149 wl_90 vdd gnd cell_6t
Xbit_r91_c149 bl_149 br_149 wl_91 vdd gnd cell_6t
Xbit_r92_c149 bl_149 br_149 wl_92 vdd gnd cell_6t
Xbit_r93_c149 bl_149 br_149 wl_93 vdd gnd cell_6t
Xbit_r94_c149 bl_149 br_149 wl_94 vdd gnd cell_6t
Xbit_r95_c149 bl_149 br_149 wl_95 vdd gnd cell_6t
Xbit_r96_c149 bl_149 br_149 wl_96 vdd gnd cell_6t
Xbit_r97_c149 bl_149 br_149 wl_97 vdd gnd cell_6t
Xbit_r98_c149 bl_149 br_149 wl_98 vdd gnd cell_6t
Xbit_r99_c149 bl_149 br_149 wl_99 vdd gnd cell_6t
Xbit_r100_c149 bl_149 br_149 wl_100 vdd gnd cell_6t
Xbit_r101_c149 bl_149 br_149 wl_101 vdd gnd cell_6t
Xbit_r102_c149 bl_149 br_149 wl_102 vdd gnd cell_6t
Xbit_r103_c149 bl_149 br_149 wl_103 vdd gnd cell_6t
Xbit_r104_c149 bl_149 br_149 wl_104 vdd gnd cell_6t
Xbit_r105_c149 bl_149 br_149 wl_105 vdd gnd cell_6t
Xbit_r106_c149 bl_149 br_149 wl_106 vdd gnd cell_6t
Xbit_r107_c149 bl_149 br_149 wl_107 vdd gnd cell_6t
Xbit_r108_c149 bl_149 br_149 wl_108 vdd gnd cell_6t
Xbit_r109_c149 bl_149 br_149 wl_109 vdd gnd cell_6t
Xbit_r110_c149 bl_149 br_149 wl_110 vdd gnd cell_6t
Xbit_r111_c149 bl_149 br_149 wl_111 vdd gnd cell_6t
Xbit_r112_c149 bl_149 br_149 wl_112 vdd gnd cell_6t
Xbit_r113_c149 bl_149 br_149 wl_113 vdd gnd cell_6t
Xbit_r114_c149 bl_149 br_149 wl_114 vdd gnd cell_6t
Xbit_r115_c149 bl_149 br_149 wl_115 vdd gnd cell_6t
Xbit_r116_c149 bl_149 br_149 wl_116 vdd gnd cell_6t
Xbit_r117_c149 bl_149 br_149 wl_117 vdd gnd cell_6t
Xbit_r118_c149 bl_149 br_149 wl_118 vdd gnd cell_6t
Xbit_r119_c149 bl_149 br_149 wl_119 vdd gnd cell_6t
Xbit_r120_c149 bl_149 br_149 wl_120 vdd gnd cell_6t
Xbit_r121_c149 bl_149 br_149 wl_121 vdd gnd cell_6t
Xbit_r122_c149 bl_149 br_149 wl_122 vdd gnd cell_6t
Xbit_r123_c149 bl_149 br_149 wl_123 vdd gnd cell_6t
Xbit_r124_c149 bl_149 br_149 wl_124 vdd gnd cell_6t
Xbit_r125_c149 bl_149 br_149 wl_125 vdd gnd cell_6t
Xbit_r126_c149 bl_149 br_149 wl_126 vdd gnd cell_6t
Xbit_r127_c149 bl_149 br_149 wl_127 vdd gnd cell_6t
Xbit_r128_c149 bl_149 br_149 wl_128 vdd gnd cell_6t
Xbit_r129_c149 bl_149 br_149 wl_129 vdd gnd cell_6t
Xbit_r130_c149 bl_149 br_149 wl_130 vdd gnd cell_6t
Xbit_r131_c149 bl_149 br_149 wl_131 vdd gnd cell_6t
Xbit_r132_c149 bl_149 br_149 wl_132 vdd gnd cell_6t
Xbit_r133_c149 bl_149 br_149 wl_133 vdd gnd cell_6t
Xbit_r134_c149 bl_149 br_149 wl_134 vdd gnd cell_6t
Xbit_r135_c149 bl_149 br_149 wl_135 vdd gnd cell_6t
Xbit_r136_c149 bl_149 br_149 wl_136 vdd gnd cell_6t
Xbit_r137_c149 bl_149 br_149 wl_137 vdd gnd cell_6t
Xbit_r138_c149 bl_149 br_149 wl_138 vdd gnd cell_6t
Xbit_r139_c149 bl_149 br_149 wl_139 vdd gnd cell_6t
Xbit_r140_c149 bl_149 br_149 wl_140 vdd gnd cell_6t
Xbit_r141_c149 bl_149 br_149 wl_141 vdd gnd cell_6t
Xbit_r142_c149 bl_149 br_149 wl_142 vdd gnd cell_6t
Xbit_r143_c149 bl_149 br_149 wl_143 vdd gnd cell_6t
Xbit_r144_c149 bl_149 br_149 wl_144 vdd gnd cell_6t
Xbit_r145_c149 bl_149 br_149 wl_145 vdd gnd cell_6t
Xbit_r146_c149 bl_149 br_149 wl_146 vdd gnd cell_6t
Xbit_r147_c149 bl_149 br_149 wl_147 vdd gnd cell_6t
Xbit_r148_c149 bl_149 br_149 wl_148 vdd gnd cell_6t
Xbit_r149_c149 bl_149 br_149 wl_149 vdd gnd cell_6t
Xbit_r150_c149 bl_149 br_149 wl_150 vdd gnd cell_6t
Xbit_r151_c149 bl_149 br_149 wl_151 vdd gnd cell_6t
Xbit_r152_c149 bl_149 br_149 wl_152 vdd gnd cell_6t
Xbit_r153_c149 bl_149 br_149 wl_153 vdd gnd cell_6t
Xbit_r154_c149 bl_149 br_149 wl_154 vdd gnd cell_6t
Xbit_r155_c149 bl_149 br_149 wl_155 vdd gnd cell_6t
Xbit_r156_c149 bl_149 br_149 wl_156 vdd gnd cell_6t
Xbit_r157_c149 bl_149 br_149 wl_157 vdd gnd cell_6t
Xbit_r158_c149 bl_149 br_149 wl_158 vdd gnd cell_6t
Xbit_r159_c149 bl_149 br_149 wl_159 vdd gnd cell_6t
Xbit_r160_c149 bl_149 br_149 wl_160 vdd gnd cell_6t
Xbit_r161_c149 bl_149 br_149 wl_161 vdd gnd cell_6t
Xbit_r162_c149 bl_149 br_149 wl_162 vdd gnd cell_6t
Xbit_r163_c149 bl_149 br_149 wl_163 vdd gnd cell_6t
Xbit_r164_c149 bl_149 br_149 wl_164 vdd gnd cell_6t
Xbit_r165_c149 bl_149 br_149 wl_165 vdd gnd cell_6t
Xbit_r166_c149 bl_149 br_149 wl_166 vdd gnd cell_6t
Xbit_r167_c149 bl_149 br_149 wl_167 vdd gnd cell_6t
Xbit_r168_c149 bl_149 br_149 wl_168 vdd gnd cell_6t
Xbit_r169_c149 bl_149 br_149 wl_169 vdd gnd cell_6t
Xbit_r170_c149 bl_149 br_149 wl_170 vdd gnd cell_6t
Xbit_r171_c149 bl_149 br_149 wl_171 vdd gnd cell_6t
Xbit_r172_c149 bl_149 br_149 wl_172 vdd gnd cell_6t
Xbit_r173_c149 bl_149 br_149 wl_173 vdd gnd cell_6t
Xbit_r174_c149 bl_149 br_149 wl_174 vdd gnd cell_6t
Xbit_r175_c149 bl_149 br_149 wl_175 vdd gnd cell_6t
Xbit_r176_c149 bl_149 br_149 wl_176 vdd gnd cell_6t
Xbit_r177_c149 bl_149 br_149 wl_177 vdd gnd cell_6t
Xbit_r178_c149 bl_149 br_149 wl_178 vdd gnd cell_6t
Xbit_r179_c149 bl_149 br_149 wl_179 vdd gnd cell_6t
Xbit_r180_c149 bl_149 br_149 wl_180 vdd gnd cell_6t
Xbit_r181_c149 bl_149 br_149 wl_181 vdd gnd cell_6t
Xbit_r182_c149 bl_149 br_149 wl_182 vdd gnd cell_6t
Xbit_r183_c149 bl_149 br_149 wl_183 vdd gnd cell_6t
Xbit_r184_c149 bl_149 br_149 wl_184 vdd gnd cell_6t
Xbit_r185_c149 bl_149 br_149 wl_185 vdd gnd cell_6t
Xbit_r186_c149 bl_149 br_149 wl_186 vdd gnd cell_6t
Xbit_r187_c149 bl_149 br_149 wl_187 vdd gnd cell_6t
Xbit_r188_c149 bl_149 br_149 wl_188 vdd gnd cell_6t
Xbit_r189_c149 bl_149 br_149 wl_189 vdd gnd cell_6t
Xbit_r190_c149 bl_149 br_149 wl_190 vdd gnd cell_6t
Xbit_r191_c149 bl_149 br_149 wl_191 vdd gnd cell_6t
Xbit_r192_c149 bl_149 br_149 wl_192 vdd gnd cell_6t
Xbit_r193_c149 bl_149 br_149 wl_193 vdd gnd cell_6t
Xbit_r194_c149 bl_149 br_149 wl_194 vdd gnd cell_6t
Xbit_r195_c149 bl_149 br_149 wl_195 vdd gnd cell_6t
Xbit_r196_c149 bl_149 br_149 wl_196 vdd gnd cell_6t
Xbit_r197_c149 bl_149 br_149 wl_197 vdd gnd cell_6t
Xbit_r198_c149 bl_149 br_149 wl_198 vdd gnd cell_6t
Xbit_r199_c149 bl_149 br_149 wl_199 vdd gnd cell_6t
Xbit_r200_c149 bl_149 br_149 wl_200 vdd gnd cell_6t
Xbit_r201_c149 bl_149 br_149 wl_201 vdd gnd cell_6t
Xbit_r202_c149 bl_149 br_149 wl_202 vdd gnd cell_6t
Xbit_r203_c149 bl_149 br_149 wl_203 vdd gnd cell_6t
Xbit_r204_c149 bl_149 br_149 wl_204 vdd gnd cell_6t
Xbit_r205_c149 bl_149 br_149 wl_205 vdd gnd cell_6t
Xbit_r206_c149 bl_149 br_149 wl_206 vdd gnd cell_6t
Xbit_r207_c149 bl_149 br_149 wl_207 vdd gnd cell_6t
Xbit_r208_c149 bl_149 br_149 wl_208 vdd gnd cell_6t
Xbit_r209_c149 bl_149 br_149 wl_209 vdd gnd cell_6t
Xbit_r210_c149 bl_149 br_149 wl_210 vdd gnd cell_6t
Xbit_r211_c149 bl_149 br_149 wl_211 vdd gnd cell_6t
Xbit_r212_c149 bl_149 br_149 wl_212 vdd gnd cell_6t
Xbit_r213_c149 bl_149 br_149 wl_213 vdd gnd cell_6t
Xbit_r214_c149 bl_149 br_149 wl_214 vdd gnd cell_6t
Xbit_r215_c149 bl_149 br_149 wl_215 vdd gnd cell_6t
Xbit_r216_c149 bl_149 br_149 wl_216 vdd gnd cell_6t
Xbit_r217_c149 bl_149 br_149 wl_217 vdd gnd cell_6t
Xbit_r218_c149 bl_149 br_149 wl_218 vdd gnd cell_6t
Xbit_r219_c149 bl_149 br_149 wl_219 vdd gnd cell_6t
Xbit_r220_c149 bl_149 br_149 wl_220 vdd gnd cell_6t
Xbit_r221_c149 bl_149 br_149 wl_221 vdd gnd cell_6t
Xbit_r222_c149 bl_149 br_149 wl_222 vdd gnd cell_6t
Xbit_r223_c149 bl_149 br_149 wl_223 vdd gnd cell_6t
Xbit_r224_c149 bl_149 br_149 wl_224 vdd gnd cell_6t
Xbit_r225_c149 bl_149 br_149 wl_225 vdd gnd cell_6t
Xbit_r226_c149 bl_149 br_149 wl_226 vdd gnd cell_6t
Xbit_r227_c149 bl_149 br_149 wl_227 vdd gnd cell_6t
Xbit_r228_c149 bl_149 br_149 wl_228 vdd gnd cell_6t
Xbit_r229_c149 bl_149 br_149 wl_229 vdd gnd cell_6t
Xbit_r230_c149 bl_149 br_149 wl_230 vdd gnd cell_6t
Xbit_r231_c149 bl_149 br_149 wl_231 vdd gnd cell_6t
Xbit_r232_c149 bl_149 br_149 wl_232 vdd gnd cell_6t
Xbit_r233_c149 bl_149 br_149 wl_233 vdd gnd cell_6t
Xbit_r234_c149 bl_149 br_149 wl_234 vdd gnd cell_6t
Xbit_r235_c149 bl_149 br_149 wl_235 vdd gnd cell_6t
Xbit_r236_c149 bl_149 br_149 wl_236 vdd gnd cell_6t
Xbit_r237_c149 bl_149 br_149 wl_237 vdd gnd cell_6t
Xbit_r238_c149 bl_149 br_149 wl_238 vdd gnd cell_6t
Xbit_r239_c149 bl_149 br_149 wl_239 vdd gnd cell_6t
Xbit_r240_c149 bl_149 br_149 wl_240 vdd gnd cell_6t
Xbit_r241_c149 bl_149 br_149 wl_241 vdd gnd cell_6t
Xbit_r242_c149 bl_149 br_149 wl_242 vdd gnd cell_6t
Xbit_r243_c149 bl_149 br_149 wl_243 vdd gnd cell_6t
Xbit_r244_c149 bl_149 br_149 wl_244 vdd gnd cell_6t
Xbit_r245_c149 bl_149 br_149 wl_245 vdd gnd cell_6t
Xbit_r246_c149 bl_149 br_149 wl_246 vdd gnd cell_6t
Xbit_r247_c149 bl_149 br_149 wl_247 vdd gnd cell_6t
Xbit_r248_c149 bl_149 br_149 wl_248 vdd gnd cell_6t
Xbit_r249_c149 bl_149 br_149 wl_249 vdd gnd cell_6t
Xbit_r250_c149 bl_149 br_149 wl_250 vdd gnd cell_6t
Xbit_r251_c149 bl_149 br_149 wl_251 vdd gnd cell_6t
Xbit_r252_c149 bl_149 br_149 wl_252 vdd gnd cell_6t
Xbit_r253_c149 bl_149 br_149 wl_253 vdd gnd cell_6t
Xbit_r254_c149 bl_149 br_149 wl_254 vdd gnd cell_6t
Xbit_r255_c149 bl_149 br_149 wl_255 vdd gnd cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd cell_6t
Xbit_r1_c150 bl_150 br_150 wl_1 vdd gnd cell_6t
Xbit_r2_c150 bl_150 br_150 wl_2 vdd gnd cell_6t
Xbit_r3_c150 bl_150 br_150 wl_3 vdd gnd cell_6t
Xbit_r4_c150 bl_150 br_150 wl_4 vdd gnd cell_6t
Xbit_r5_c150 bl_150 br_150 wl_5 vdd gnd cell_6t
Xbit_r6_c150 bl_150 br_150 wl_6 vdd gnd cell_6t
Xbit_r7_c150 bl_150 br_150 wl_7 vdd gnd cell_6t
Xbit_r8_c150 bl_150 br_150 wl_8 vdd gnd cell_6t
Xbit_r9_c150 bl_150 br_150 wl_9 vdd gnd cell_6t
Xbit_r10_c150 bl_150 br_150 wl_10 vdd gnd cell_6t
Xbit_r11_c150 bl_150 br_150 wl_11 vdd gnd cell_6t
Xbit_r12_c150 bl_150 br_150 wl_12 vdd gnd cell_6t
Xbit_r13_c150 bl_150 br_150 wl_13 vdd gnd cell_6t
Xbit_r14_c150 bl_150 br_150 wl_14 vdd gnd cell_6t
Xbit_r15_c150 bl_150 br_150 wl_15 vdd gnd cell_6t
Xbit_r16_c150 bl_150 br_150 wl_16 vdd gnd cell_6t
Xbit_r17_c150 bl_150 br_150 wl_17 vdd gnd cell_6t
Xbit_r18_c150 bl_150 br_150 wl_18 vdd gnd cell_6t
Xbit_r19_c150 bl_150 br_150 wl_19 vdd gnd cell_6t
Xbit_r20_c150 bl_150 br_150 wl_20 vdd gnd cell_6t
Xbit_r21_c150 bl_150 br_150 wl_21 vdd gnd cell_6t
Xbit_r22_c150 bl_150 br_150 wl_22 vdd gnd cell_6t
Xbit_r23_c150 bl_150 br_150 wl_23 vdd gnd cell_6t
Xbit_r24_c150 bl_150 br_150 wl_24 vdd gnd cell_6t
Xbit_r25_c150 bl_150 br_150 wl_25 vdd gnd cell_6t
Xbit_r26_c150 bl_150 br_150 wl_26 vdd gnd cell_6t
Xbit_r27_c150 bl_150 br_150 wl_27 vdd gnd cell_6t
Xbit_r28_c150 bl_150 br_150 wl_28 vdd gnd cell_6t
Xbit_r29_c150 bl_150 br_150 wl_29 vdd gnd cell_6t
Xbit_r30_c150 bl_150 br_150 wl_30 vdd gnd cell_6t
Xbit_r31_c150 bl_150 br_150 wl_31 vdd gnd cell_6t
Xbit_r32_c150 bl_150 br_150 wl_32 vdd gnd cell_6t
Xbit_r33_c150 bl_150 br_150 wl_33 vdd gnd cell_6t
Xbit_r34_c150 bl_150 br_150 wl_34 vdd gnd cell_6t
Xbit_r35_c150 bl_150 br_150 wl_35 vdd gnd cell_6t
Xbit_r36_c150 bl_150 br_150 wl_36 vdd gnd cell_6t
Xbit_r37_c150 bl_150 br_150 wl_37 vdd gnd cell_6t
Xbit_r38_c150 bl_150 br_150 wl_38 vdd gnd cell_6t
Xbit_r39_c150 bl_150 br_150 wl_39 vdd gnd cell_6t
Xbit_r40_c150 bl_150 br_150 wl_40 vdd gnd cell_6t
Xbit_r41_c150 bl_150 br_150 wl_41 vdd gnd cell_6t
Xbit_r42_c150 bl_150 br_150 wl_42 vdd gnd cell_6t
Xbit_r43_c150 bl_150 br_150 wl_43 vdd gnd cell_6t
Xbit_r44_c150 bl_150 br_150 wl_44 vdd gnd cell_6t
Xbit_r45_c150 bl_150 br_150 wl_45 vdd gnd cell_6t
Xbit_r46_c150 bl_150 br_150 wl_46 vdd gnd cell_6t
Xbit_r47_c150 bl_150 br_150 wl_47 vdd gnd cell_6t
Xbit_r48_c150 bl_150 br_150 wl_48 vdd gnd cell_6t
Xbit_r49_c150 bl_150 br_150 wl_49 vdd gnd cell_6t
Xbit_r50_c150 bl_150 br_150 wl_50 vdd gnd cell_6t
Xbit_r51_c150 bl_150 br_150 wl_51 vdd gnd cell_6t
Xbit_r52_c150 bl_150 br_150 wl_52 vdd gnd cell_6t
Xbit_r53_c150 bl_150 br_150 wl_53 vdd gnd cell_6t
Xbit_r54_c150 bl_150 br_150 wl_54 vdd gnd cell_6t
Xbit_r55_c150 bl_150 br_150 wl_55 vdd gnd cell_6t
Xbit_r56_c150 bl_150 br_150 wl_56 vdd gnd cell_6t
Xbit_r57_c150 bl_150 br_150 wl_57 vdd gnd cell_6t
Xbit_r58_c150 bl_150 br_150 wl_58 vdd gnd cell_6t
Xbit_r59_c150 bl_150 br_150 wl_59 vdd gnd cell_6t
Xbit_r60_c150 bl_150 br_150 wl_60 vdd gnd cell_6t
Xbit_r61_c150 bl_150 br_150 wl_61 vdd gnd cell_6t
Xbit_r62_c150 bl_150 br_150 wl_62 vdd gnd cell_6t
Xbit_r63_c150 bl_150 br_150 wl_63 vdd gnd cell_6t
Xbit_r64_c150 bl_150 br_150 wl_64 vdd gnd cell_6t
Xbit_r65_c150 bl_150 br_150 wl_65 vdd gnd cell_6t
Xbit_r66_c150 bl_150 br_150 wl_66 vdd gnd cell_6t
Xbit_r67_c150 bl_150 br_150 wl_67 vdd gnd cell_6t
Xbit_r68_c150 bl_150 br_150 wl_68 vdd gnd cell_6t
Xbit_r69_c150 bl_150 br_150 wl_69 vdd gnd cell_6t
Xbit_r70_c150 bl_150 br_150 wl_70 vdd gnd cell_6t
Xbit_r71_c150 bl_150 br_150 wl_71 vdd gnd cell_6t
Xbit_r72_c150 bl_150 br_150 wl_72 vdd gnd cell_6t
Xbit_r73_c150 bl_150 br_150 wl_73 vdd gnd cell_6t
Xbit_r74_c150 bl_150 br_150 wl_74 vdd gnd cell_6t
Xbit_r75_c150 bl_150 br_150 wl_75 vdd gnd cell_6t
Xbit_r76_c150 bl_150 br_150 wl_76 vdd gnd cell_6t
Xbit_r77_c150 bl_150 br_150 wl_77 vdd gnd cell_6t
Xbit_r78_c150 bl_150 br_150 wl_78 vdd gnd cell_6t
Xbit_r79_c150 bl_150 br_150 wl_79 vdd gnd cell_6t
Xbit_r80_c150 bl_150 br_150 wl_80 vdd gnd cell_6t
Xbit_r81_c150 bl_150 br_150 wl_81 vdd gnd cell_6t
Xbit_r82_c150 bl_150 br_150 wl_82 vdd gnd cell_6t
Xbit_r83_c150 bl_150 br_150 wl_83 vdd gnd cell_6t
Xbit_r84_c150 bl_150 br_150 wl_84 vdd gnd cell_6t
Xbit_r85_c150 bl_150 br_150 wl_85 vdd gnd cell_6t
Xbit_r86_c150 bl_150 br_150 wl_86 vdd gnd cell_6t
Xbit_r87_c150 bl_150 br_150 wl_87 vdd gnd cell_6t
Xbit_r88_c150 bl_150 br_150 wl_88 vdd gnd cell_6t
Xbit_r89_c150 bl_150 br_150 wl_89 vdd gnd cell_6t
Xbit_r90_c150 bl_150 br_150 wl_90 vdd gnd cell_6t
Xbit_r91_c150 bl_150 br_150 wl_91 vdd gnd cell_6t
Xbit_r92_c150 bl_150 br_150 wl_92 vdd gnd cell_6t
Xbit_r93_c150 bl_150 br_150 wl_93 vdd gnd cell_6t
Xbit_r94_c150 bl_150 br_150 wl_94 vdd gnd cell_6t
Xbit_r95_c150 bl_150 br_150 wl_95 vdd gnd cell_6t
Xbit_r96_c150 bl_150 br_150 wl_96 vdd gnd cell_6t
Xbit_r97_c150 bl_150 br_150 wl_97 vdd gnd cell_6t
Xbit_r98_c150 bl_150 br_150 wl_98 vdd gnd cell_6t
Xbit_r99_c150 bl_150 br_150 wl_99 vdd gnd cell_6t
Xbit_r100_c150 bl_150 br_150 wl_100 vdd gnd cell_6t
Xbit_r101_c150 bl_150 br_150 wl_101 vdd gnd cell_6t
Xbit_r102_c150 bl_150 br_150 wl_102 vdd gnd cell_6t
Xbit_r103_c150 bl_150 br_150 wl_103 vdd gnd cell_6t
Xbit_r104_c150 bl_150 br_150 wl_104 vdd gnd cell_6t
Xbit_r105_c150 bl_150 br_150 wl_105 vdd gnd cell_6t
Xbit_r106_c150 bl_150 br_150 wl_106 vdd gnd cell_6t
Xbit_r107_c150 bl_150 br_150 wl_107 vdd gnd cell_6t
Xbit_r108_c150 bl_150 br_150 wl_108 vdd gnd cell_6t
Xbit_r109_c150 bl_150 br_150 wl_109 vdd gnd cell_6t
Xbit_r110_c150 bl_150 br_150 wl_110 vdd gnd cell_6t
Xbit_r111_c150 bl_150 br_150 wl_111 vdd gnd cell_6t
Xbit_r112_c150 bl_150 br_150 wl_112 vdd gnd cell_6t
Xbit_r113_c150 bl_150 br_150 wl_113 vdd gnd cell_6t
Xbit_r114_c150 bl_150 br_150 wl_114 vdd gnd cell_6t
Xbit_r115_c150 bl_150 br_150 wl_115 vdd gnd cell_6t
Xbit_r116_c150 bl_150 br_150 wl_116 vdd gnd cell_6t
Xbit_r117_c150 bl_150 br_150 wl_117 vdd gnd cell_6t
Xbit_r118_c150 bl_150 br_150 wl_118 vdd gnd cell_6t
Xbit_r119_c150 bl_150 br_150 wl_119 vdd gnd cell_6t
Xbit_r120_c150 bl_150 br_150 wl_120 vdd gnd cell_6t
Xbit_r121_c150 bl_150 br_150 wl_121 vdd gnd cell_6t
Xbit_r122_c150 bl_150 br_150 wl_122 vdd gnd cell_6t
Xbit_r123_c150 bl_150 br_150 wl_123 vdd gnd cell_6t
Xbit_r124_c150 bl_150 br_150 wl_124 vdd gnd cell_6t
Xbit_r125_c150 bl_150 br_150 wl_125 vdd gnd cell_6t
Xbit_r126_c150 bl_150 br_150 wl_126 vdd gnd cell_6t
Xbit_r127_c150 bl_150 br_150 wl_127 vdd gnd cell_6t
Xbit_r128_c150 bl_150 br_150 wl_128 vdd gnd cell_6t
Xbit_r129_c150 bl_150 br_150 wl_129 vdd gnd cell_6t
Xbit_r130_c150 bl_150 br_150 wl_130 vdd gnd cell_6t
Xbit_r131_c150 bl_150 br_150 wl_131 vdd gnd cell_6t
Xbit_r132_c150 bl_150 br_150 wl_132 vdd gnd cell_6t
Xbit_r133_c150 bl_150 br_150 wl_133 vdd gnd cell_6t
Xbit_r134_c150 bl_150 br_150 wl_134 vdd gnd cell_6t
Xbit_r135_c150 bl_150 br_150 wl_135 vdd gnd cell_6t
Xbit_r136_c150 bl_150 br_150 wl_136 vdd gnd cell_6t
Xbit_r137_c150 bl_150 br_150 wl_137 vdd gnd cell_6t
Xbit_r138_c150 bl_150 br_150 wl_138 vdd gnd cell_6t
Xbit_r139_c150 bl_150 br_150 wl_139 vdd gnd cell_6t
Xbit_r140_c150 bl_150 br_150 wl_140 vdd gnd cell_6t
Xbit_r141_c150 bl_150 br_150 wl_141 vdd gnd cell_6t
Xbit_r142_c150 bl_150 br_150 wl_142 vdd gnd cell_6t
Xbit_r143_c150 bl_150 br_150 wl_143 vdd gnd cell_6t
Xbit_r144_c150 bl_150 br_150 wl_144 vdd gnd cell_6t
Xbit_r145_c150 bl_150 br_150 wl_145 vdd gnd cell_6t
Xbit_r146_c150 bl_150 br_150 wl_146 vdd gnd cell_6t
Xbit_r147_c150 bl_150 br_150 wl_147 vdd gnd cell_6t
Xbit_r148_c150 bl_150 br_150 wl_148 vdd gnd cell_6t
Xbit_r149_c150 bl_150 br_150 wl_149 vdd gnd cell_6t
Xbit_r150_c150 bl_150 br_150 wl_150 vdd gnd cell_6t
Xbit_r151_c150 bl_150 br_150 wl_151 vdd gnd cell_6t
Xbit_r152_c150 bl_150 br_150 wl_152 vdd gnd cell_6t
Xbit_r153_c150 bl_150 br_150 wl_153 vdd gnd cell_6t
Xbit_r154_c150 bl_150 br_150 wl_154 vdd gnd cell_6t
Xbit_r155_c150 bl_150 br_150 wl_155 vdd gnd cell_6t
Xbit_r156_c150 bl_150 br_150 wl_156 vdd gnd cell_6t
Xbit_r157_c150 bl_150 br_150 wl_157 vdd gnd cell_6t
Xbit_r158_c150 bl_150 br_150 wl_158 vdd gnd cell_6t
Xbit_r159_c150 bl_150 br_150 wl_159 vdd gnd cell_6t
Xbit_r160_c150 bl_150 br_150 wl_160 vdd gnd cell_6t
Xbit_r161_c150 bl_150 br_150 wl_161 vdd gnd cell_6t
Xbit_r162_c150 bl_150 br_150 wl_162 vdd gnd cell_6t
Xbit_r163_c150 bl_150 br_150 wl_163 vdd gnd cell_6t
Xbit_r164_c150 bl_150 br_150 wl_164 vdd gnd cell_6t
Xbit_r165_c150 bl_150 br_150 wl_165 vdd gnd cell_6t
Xbit_r166_c150 bl_150 br_150 wl_166 vdd gnd cell_6t
Xbit_r167_c150 bl_150 br_150 wl_167 vdd gnd cell_6t
Xbit_r168_c150 bl_150 br_150 wl_168 vdd gnd cell_6t
Xbit_r169_c150 bl_150 br_150 wl_169 vdd gnd cell_6t
Xbit_r170_c150 bl_150 br_150 wl_170 vdd gnd cell_6t
Xbit_r171_c150 bl_150 br_150 wl_171 vdd gnd cell_6t
Xbit_r172_c150 bl_150 br_150 wl_172 vdd gnd cell_6t
Xbit_r173_c150 bl_150 br_150 wl_173 vdd gnd cell_6t
Xbit_r174_c150 bl_150 br_150 wl_174 vdd gnd cell_6t
Xbit_r175_c150 bl_150 br_150 wl_175 vdd gnd cell_6t
Xbit_r176_c150 bl_150 br_150 wl_176 vdd gnd cell_6t
Xbit_r177_c150 bl_150 br_150 wl_177 vdd gnd cell_6t
Xbit_r178_c150 bl_150 br_150 wl_178 vdd gnd cell_6t
Xbit_r179_c150 bl_150 br_150 wl_179 vdd gnd cell_6t
Xbit_r180_c150 bl_150 br_150 wl_180 vdd gnd cell_6t
Xbit_r181_c150 bl_150 br_150 wl_181 vdd gnd cell_6t
Xbit_r182_c150 bl_150 br_150 wl_182 vdd gnd cell_6t
Xbit_r183_c150 bl_150 br_150 wl_183 vdd gnd cell_6t
Xbit_r184_c150 bl_150 br_150 wl_184 vdd gnd cell_6t
Xbit_r185_c150 bl_150 br_150 wl_185 vdd gnd cell_6t
Xbit_r186_c150 bl_150 br_150 wl_186 vdd gnd cell_6t
Xbit_r187_c150 bl_150 br_150 wl_187 vdd gnd cell_6t
Xbit_r188_c150 bl_150 br_150 wl_188 vdd gnd cell_6t
Xbit_r189_c150 bl_150 br_150 wl_189 vdd gnd cell_6t
Xbit_r190_c150 bl_150 br_150 wl_190 vdd gnd cell_6t
Xbit_r191_c150 bl_150 br_150 wl_191 vdd gnd cell_6t
Xbit_r192_c150 bl_150 br_150 wl_192 vdd gnd cell_6t
Xbit_r193_c150 bl_150 br_150 wl_193 vdd gnd cell_6t
Xbit_r194_c150 bl_150 br_150 wl_194 vdd gnd cell_6t
Xbit_r195_c150 bl_150 br_150 wl_195 vdd gnd cell_6t
Xbit_r196_c150 bl_150 br_150 wl_196 vdd gnd cell_6t
Xbit_r197_c150 bl_150 br_150 wl_197 vdd gnd cell_6t
Xbit_r198_c150 bl_150 br_150 wl_198 vdd gnd cell_6t
Xbit_r199_c150 bl_150 br_150 wl_199 vdd gnd cell_6t
Xbit_r200_c150 bl_150 br_150 wl_200 vdd gnd cell_6t
Xbit_r201_c150 bl_150 br_150 wl_201 vdd gnd cell_6t
Xbit_r202_c150 bl_150 br_150 wl_202 vdd gnd cell_6t
Xbit_r203_c150 bl_150 br_150 wl_203 vdd gnd cell_6t
Xbit_r204_c150 bl_150 br_150 wl_204 vdd gnd cell_6t
Xbit_r205_c150 bl_150 br_150 wl_205 vdd gnd cell_6t
Xbit_r206_c150 bl_150 br_150 wl_206 vdd gnd cell_6t
Xbit_r207_c150 bl_150 br_150 wl_207 vdd gnd cell_6t
Xbit_r208_c150 bl_150 br_150 wl_208 vdd gnd cell_6t
Xbit_r209_c150 bl_150 br_150 wl_209 vdd gnd cell_6t
Xbit_r210_c150 bl_150 br_150 wl_210 vdd gnd cell_6t
Xbit_r211_c150 bl_150 br_150 wl_211 vdd gnd cell_6t
Xbit_r212_c150 bl_150 br_150 wl_212 vdd gnd cell_6t
Xbit_r213_c150 bl_150 br_150 wl_213 vdd gnd cell_6t
Xbit_r214_c150 bl_150 br_150 wl_214 vdd gnd cell_6t
Xbit_r215_c150 bl_150 br_150 wl_215 vdd gnd cell_6t
Xbit_r216_c150 bl_150 br_150 wl_216 vdd gnd cell_6t
Xbit_r217_c150 bl_150 br_150 wl_217 vdd gnd cell_6t
Xbit_r218_c150 bl_150 br_150 wl_218 vdd gnd cell_6t
Xbit_r219_c150 bl_150 br_150 wl_219 vdd gnd cell_6t
Xbit_r220_c150 bl_150 br_150 wl_220 vdd gnd cell_6t
Xbit_r221_c150 bl_150 br_150 wl_221 vdd gnd cell_6t
Xbit_r222_c150 bl_150 br_150 wl_222 vdd gnd cell_6t
Xbit_r223_c150 bl_150 br_150 wl_223 vdd gnd cell_6t
Xbit_r224_c150 bl_150 br_150 wl_224 vdd gnd cell_6t
Xbit_r225_c150 bl_150 br_150 wl_225 vdd gnd cell_6t
Xbit_r226_c150 bl_150 br_150 wl_226 vdd gnd cell_6t
Xbit_r227_c150 bl_150 br_150 wl_227 vdd gnd cell_6t
Xbit_r228_c150 bl_150 br_150 wl_228 vdd gnd cell_6t
Xbit_r229_c150 bl_150 br_150 wl_229 vdd gnd cell_6t
Xbit_r230_c150 bl_150 br_150 wl_230 vdd gnd cell_6t
Xbit_r231_c150 bl_150 br_150 wl_231 vdd gnd cell_6t
Xbit_r232_c150 bl_150 br_150 wl_232 vdd gnd cell_6t
Xbit_r233_c150 bl_150 br_150 wl_233 vdd gnd cell_6t
Xbit_r234_c150 bl_150 br_150 wl_234 vdd gnd cell_6t
Xbit_r235_c150 bl_150 br_150 wl_235 vdd gnd cell_6t
Xbit_r236_c150 bl_150 br_150 wl_236 vdd gnd cell_6t
Xbit_r237_c150 bl_150 br_150 wl_237 vdd gnd cell_6t
Xbit_r238_c150 bl_150 br_150 wl_238 vdd gnd cell_6t
Xbit_r239_c150 bl_150 br_150 wl_239 vdd gnd cell_6t
Xbit_r240_c150 bl_150 br_150 wl_240 vdd gnd cell_6t
Xbit_r241_c150 bl_150 br_150 wl_241 vdd gnd cell_6t
Xbit_r242_c150 bl_150 br_150 wl_242 vdd gnd cell_6t
Xbit_r243_c150 bl_150 br_150 wl_243 vdd gnd cell_6t
Xbit_r244_c150 bl_150 br_150 wl_244 vdd gnd cell_6t
Xbit_r245_c150 bl_150 br_150 wl_245 vdd gnd cell_6t
Xbit_r246_c150 bl_150 br_150 wl_246 vdd gnd cell_6t
Xbit_r247_c150 bl_150 br_150 wl_247 vdd gnd cell_6t
Xbit_r248_c150 bl_150 br_150 wl_248 vdd gnd cell_6t
Xbit_r249_c150 bl_150 br_150 wl_249 vdd gnd cell_6t
Xbit_r250_c150 bl_150 br_150 wl_250 vdd gnd cell_6t
Xbit_r251_c150 bl_150 br_150 wl_251 vdd gnd cell_6t
Xbit_r252_c150 bl_150 br_150 wl_252 vdd gnd cell_6t
Xbit_r253_c150 bl_150 br_150 wl_253 vdd gnd cell_6t
Xbit_r254_c150 bl_150 br_150 wl_254 vdd gnd cell_6t
Xbit_r255_c150 bl_150 br_150 wl_255 vdd gnd cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd cell_6t
Xbit_r1_c151 bl_151 br_151 wl_1 vdd gnd cell_6t
Xbit_r2_c151 bl_151 br_151 wl_2 vdd gnd cell_6t
Xbit_r3_c151 bl_151 br_151 wl_3 vdd gnd cell_6t
Xbit_r4_c151 bl_151 br_151 wl_4 vdd gnd cell_6t
Xbit_r5_c151 bl_151 br_151 wl_5 vdd gnd cell_6t
Xbit_r6_c151 bl_151 br_151 wl_6 vdd gnd cell_6t
Xbit_r7_c151 bl_151 br_151 wl_7 vdd gnd cell_6t
Xbit_r8_c151 bl_151 br_151 wl_8 vdd gnd cell_6t
Xbit_r9_c151 bl_151 br_151 wl_9 vdd gnd cell_6t
Xbit_r10_c151 bl_151 br_151 wl_10 vdd gnd cell_6t
Xbit_r11_c151 bl_151 br_151 wl_11 vdd gnd cell_6t
Xbit_r12_c151 bl_151 br_151 wl_12 vdd gnd cell_6t
Xbit_r13_c151 bl_151 br_151 wl_13 vdd gnd cell_6t
Xbit_r14_c151 bl_151 br_151 wl_14 vdd gnd cell_6t
Xbit_r15_c151 bl_151 br_151 wl_15 vdd gnd cell_6t
Xbit_r16_c151 bl_151 br_151 wl_16 vdd gnd cell_6t
Xbit_r17_c151 bl_151 br_151 wl_17 vdd gnd cell_6t
Xbit_r18_c151 bl_151 br_151 wl_18 vdd gnd cell_6t
Xbit_r19_c151 bl_151 br_151 wl_19 vdd gnd cell_6t
Xbit_r20_c151 bl_151 br_151 wl_20 vdd gnd cell_6t
Xbit_r21_c151 bl_151 br_151 wl_21 vdd gnd cell_6t
Xbit_r22_c151 bl_151 br_151 wl_22 vdd gnd cell_6t
Xbit_r23_c151 bl_151 br_151 wl_23 vdd gnd cell_6t
Xbit_r24_c151 bl_151 br_151 wl_24 vdd gnd cell_6t
Xbit_r25_c151 bl_151 br_151 wl_25 vdd gnd cell_6t
Xbit_r26_c151 bl_151 br_151 wl_26 vdd gnd cell_6t
Xbit_r27_c151 bl_151 br_151 wl_27 vdd gnd cell_6t
Xbit_r28_c151 bl_151 br_151 wl_28 vdd gnd cell_6t
Xbit_r29_c151 bl_151 br_151 wl_29 vdd gnd cell_6t
Xbit_r30_c151 bl_151 br_151 wl_30 vdd gnd cell_6t
Xbit_r31_c151 bl_151 br_151 wl_31 vdd gnd cell_6t
Xbit_r32_c151 bl_151 br_151 wl_32 vdd gnd cell_6t
Xbit_r33_c151 bl_151 br_151 wl_33 vdd gnd cell_6t
Xbit_r34_c151 bl_151 br_151 wl_34 vdd gnd cell_6t
Xbit_r35_c151 bl_151 br_151 wl_35 vdd gnd cell_6t
Xbit_r36_c151 bl_151 br_151 wl_36 vdd gnd cell_6t
Xbit_r37_c151 bl_151 br_151 wl_37 vdd gnd cell_6t
Xbit_r38_c151 bl_151 br_151 wl_38 vdd gnd cell_6t
Xbit_r39_c151 bl_151 br_151 wl_39 vdd gnd cell_6t
Xbit_r40_c151 bl_151 br_151 wl_40 vdd gnd cell_6t
Xbit_r41_c151 bl_151 br_151 wl_41 vdd gnd cell_6t
Xbit_r42_c151 bl_151 br_151 wl_42 vdd gnd cell_6t
Xbit_r43_c151 bl_151 br_151 wl_43 vdd gnd cell_6t
Xbit_r44_c151 bl_151 br_151 wl_44 vdd gnd cell_6t
Xbit_r45_c151 bl_151 br_151 wl_45 vdd gnd cell_6t
Xbit_r46_c151 bl_151 br_151 wl_46 vdd gnd cell_6t
Xbit_r47_c151 bl_151 br_151 wl_47 vdd gnd cell_6t
Xbit_r48_c151 bl_151 br_151 wl_48 vdd gnd cell_6t
Xbit_r49_c151 bl_151 br_151 wl_49 vdd gnd cell_6t
Xbit_r50_c151 bl_151 br_151 wl_50 vdd gnd cell_6t
Xbit_r51_c151 bl_151 br_151 wl_51 vdd gnd cell_6t
Xbit_r52_c151 bl_151 br_151 wl_52 vdd gnd cell_6t
Xbit_r53_c151 bl_151 br_151 wl_53 vdd gnd cell_6t
Xbit_r54_c151 bl_151 br_151 wl_54 vdd gnd cell_6t
Xbit_r55_c151 bl_151 br_151 wl_55 vdd gnd cell_6t
Xbit_r56_c151 bl_151 br_151 wl_56 vdd gnd cell_6t
Xbit_r57_c151 bl_151 br_151 wl_57 vdd gnd cell_6t
Xbit_r58_c151 bl_151 br_151 wl_58 vdd gnd cell_6t
Xbit_r59_c151 bl_151 br_151 wl_59 vdd gnd cell_6t
Xbit_r60_c151 bl_151 br_151 wl_60 vdd gnd cell_6t
Xbit_r61_c151 bl_151 br_151 wl_61 vdd gnd cell_6t
Xbit_r62_c151 bl_151 br_151 wl_62 vdd gnd cell_6t
Xbit_r63_c151 bl_151 br_151 wl_63 vdd gnd cell_6t
Xbit_r64_c151 bl_151 br_151 wl_64 vdd gnd cell_6t
Xbit_r65_c151 bl_151 br_151 wl_65 vdd gnd cell_6t
Xbit_r66_c151 bl_151 br_151 wl_66 vdd gnd cell_6t
Xbit_r67_c151 bl_151 br_151 wl_67 vdd gnd cell_6t
Xbit_r68_c151 bl_151 br_151 wl_68 vdd gnd cell_6t
Xbit_r69_c151 bl_151 br_151 wl_69 vdd gnd cell_6t
Xbit_r70_c151 bl_151 br_151 wl_70 vdd gnd cell_6t
Xbit_r71_c151 bl_151 br_151 wl_71 vdd gnd cell_6t
Xbit_r72_c151 bl_151 br_151 wl_72 vdd gnd cell_6t
Xbit_r73_c151 bl_151 br_151 wl_73 vdd gnd cell_6t
Xbit_r74_c151 bl_151 br_151 wl_74 vdd gnd cell_6t
Xbit_r75_c151 bl_151 br_151 wl_75 vdd gnd cell_6t
Xbit_r76_c151 bl_151 br_151 wl_76 vdd gnd cell_6t
Xbit_r77_c151 bl_151 br_151 wl_77 vdd gnd cell_6t
Xbit_r78_c151 bl_151 br_151 wl_78 vdd gnd cell_6t
Xbit_r79_c151 bl_151 br_151 wl_79 vdd gnd cell_6t
Xbit_r80_c151 bl_151 br_151 wl_80 vdd gnd cell_6t
Xbit_r81_c151 bl_151 br_151 wl_81 vdd gnd cell_6t
Xbit_r82_c151 bl_151 br_151 wl_82 vdd gnd cell_6t
Xbit_r83_c151 bl_151 br_151 wl_83 vdd gnd cell_6t
Xbit_r84_c151 bl_151 br_151 wl_84 vdd gnd cell_6t
Xbit_r85_c151 bl_151 br_151 wl_85 vdd gnd cell_6t
Xbit_r86_c151 bl_151 br_151 wl_86 vdd gnd cell_6t
Xbit_r87_c151 bl_151 br_151 wl_87 vdd gnd cell_6t
Xbit_r88_c151 bl_151 br_151 wl_88 vdd gnd cell_6t
Xbit_r89_c151 bl_151 br_151 wl_89 vdd gnd cell_6t
Xbit_r90_c151 bl_151 br_151 wl_90 vdd gnd cell_6t
Xbit_r91_c151 bl_151 br_151 wl_91 vdd gnd cell_6t
Xbit_r92_c151 bl_151 br_151 wl_92 vdd gnd cell_6t
Xbit_r93_c151 bl_151 br_151 wl_93 vdd gnd cell_6t
Xbit_r94_c151 bl_151 br_151 wl_94 vdd gnd cell_6t
Xbit_r95_c151 bl_151 br_151 wl_95 vdd gnd cell_6t
Xbit_r96_c151 bl_151 br_151 wl_96 vdd gnd cell_6t
Xbit_r97_c151 bl_151 br_151 wl_97 vdd gnd cell_6t
Xbit_r98_c151 bl_151 br_151 wl_98 vdd gnd cell_6t
Xbit_r99_c151 bl_151 br_151 wl_99 vdd gnd cell_6t
Xbit_r100_c151 bl_151 br_151 wl_100 vdd gnd cell_6t
Xbit_r101_c151 bl_151 br_151 wl_101 vdd gnd cell_6t
Xbit_r102_c151 bl_151 br_151 wl_102 vdd gnd cell_6t
Xbit_r103_c151 bl_151 br_151 wl_103 vdd gnd cell_6t
Xbit_r104_c151 bl_151 br_151 wl_104 vdd gnd cell_6t
Xbit_r105_c151 bl_151 br_151 wl_105 vdd gnd cell_6t
Xbit_r106_c151 bl_151 br_151 wl_106 vdd gnd cell_6t
Xbit_r107_c151 bl_151 br_151 wl_107 vdd gnd cell_6t
Xbit_r108_c151 bl_151 br_151 wl_108 vdd gnd cell_6t
Xbit_r109_c151 bl_151 br_151 wl_109 vdd gnd cell_6t
Xbit_r110_c151 bl_151 br_151 wl_110 vdd gnd cell_6t
Xbit_r111_c151 bl_151 br_151 wl_111 vdd gnd cell_6t
Xbit_r112_c151 bl_151 br_151 wl_112 vdd gnd cell_6t
Xbit_r113_c151 bl_151 br_151 wl_113 vdd gnd cell_6t
Xbit_r114_c151 bl_151 br_151 wl_114 vdd gnd cell_6t
Xbit_r115_c151 bl_151 br_151 wl_115 vdd gnd cell_6t
Xbit_r116_c151 bl_151 br_151 wl_116 vdd gnd cell_6t
Xbit_r117_c151 bl_151 br_151 wl_117 vdd gnd cell_6t
Xbit_r118_c151 bl_151 br_151 wl_118 vdd gnd cell_6t
Xbit_r119_c151 bl_151 br_151 wl_119 vdd gnd cell_6t
Xbit_r120_c151 bl_151 br_151 wl_120 vdd gnd cell_6t
Xbit_r121_c151 bl_151 br_151 wl_121 vdd gnd cell_6t
Xbit_r122_c151 bl_151 br_151 wl_122 vdd gnd cell_6t
Xbit_r123_c151 bl_151 br_151 wl_123 vdd gnd cell_6t
Xbit_r124_c151 bl_151 br_151 wl_124 vdd gnd cell_6t
Xbit_r125_c151 bl_151 br_151 wl_125 vdd gnd cell_6t
Xbit_r126_c151 bl_151 br_151 wl_126 vdd gnd cell_6t
Xbit_r127_c151 bl_151 br_151 wl_127 vdd gnd cell_6t
Xbit_r128_c151 bl_151 br_151 wl_128 vdd gnd cell_6t
Xbit_r129_c151 bl_151 br_151 wl_129 vdd gnd cell_6t
Xbit_r130_c151 bl_151 br_151 wl_130 vdd gnd cell_6t
Xbit_r131_c151 bl_151 br_151 wl_131 vdd gnd cell_6t
Xbit_r132_c151 bl_151 br_151 wl_132 vdd gnd cell_6t
Xbit_r133_c151 bl_151 br_151 wl_133 vdd gnd cell_6t
Xbit_r134_c151 bl_151 br_151 wl_134 vdd gnd cell_6t
Xbit_r135_c151 bl_151 br_151 wl_135 vdd gnd cell_6t
Xbit_r136_c151 bl_151 br_151 wl_136 vdd gnd cell_6t
Xbit_r137_c151 bl_151 br_151 wl_137 vdd gnd cell_6t
Xbit_r138_c151 bl_151 br_151 wl_138 vdd gnd cell_6t
Xbit_r139_c151 bl_151 br_151 wl_139 vdd gnd cell_6t
Xbit_r140_c151 bl_151 br_151 wl_140 vdd gnd cell_6t
Xbit_r141_c151 bl_151 br_151 wl_141 vdd gnd cell_6t
Xbit_r142_c151 bl_151 br_151 wl_142 vdd gnd cell_6t
Xbit_r143_c151 bl_151 br_151 wl_143 vdd gnd cell_6t
Xbit_r144_c151 bl_151 br_151 wl_144 vdd gnd cell_6t
Xbit_r145_c151 bl_151 br_151 wl_145 vdd gnd cell_6t
Xbit_r146_c151 bl_151 br_151 wl_146 vdd gnd cell_6t
Xbit_r147_c151 bl_151 br_151 wl_147 vdd gnd cell_6t
Xbit_r148_c151 bl_151 br_151 wl_148 vdd gnd cell_6t
Xbit_r149_c151 bl_151 br_151 wl_149 vdd gnd cell_6t
Xbit_r150_c151 bl_151 br_151 wl_150 vdd gnd cell_6t
Xbit_r151_c151 bl_151 br_151 wl_151 vdd gnd cell_6t
Xbit_r152_c151 bl_151 br_151 wl_152 vdd gnd cell_6t
Xbit_r153_c151 bl_151 br_151 wl_153 vdd gnd cell_6t
Xbit_r154_c151 bl_151 br_151 wl_154 vdd gnd cell_6t
Xbit_r155_c151 bl_151 br_151 wl_155 vdd gnd cell_6t
Xbit_r156_c151 bl_151 br_151 wl_156 vdd gnd cell_6t
Xbit_r157_c151 bl_151 br_151 wl_157 vdd gnd cell_6t
Xbit_r158_c151 bl_151 br_151 wl_158 vdd gnd cell_6t
Xbit_r159_c151 bl_151 br_151 wl_159 vdd gnd cell_6t
Xbit_r160_c151 bl_151 br_151 wl_160 vdd gnd cell_6t
Xbit_r161_c151 bl_151 br_151 wl_161 vdd gnd cell_6t
Xbit_r162_c151 bl_151 br_151 wl_162 vdd gnd cell_6t
Xbit_r163_c151 bl_151 br_151 wl_163 vdd gnd cell_6t
Xbit_r164_c151 bl_151 br_151 wl_164 vdd gnd cell_6t
Xbit_r165_c151 bl_151 br_151 wl_165 vdd gnd cell_6t
Xbit_r166_c151 bl_151 br_151 wl_166 vdd gnd cell_6t
Xbit_r167_c151 bl_151 br_151 wl_167 vdd gnd cell_6t
Xbit_r168_c151 bl_151 br_151 wl_168 vdd gnd cell_6t
Xbit_r169_c151 bl_151 br_151 wl_169 vdd gnd cell_6t
Xbit_r170_c151 bl_151 br_151 wl_170 vdd gnd cell_6t
Xbit_r171_c151 bl_151 br_151 wl_171 vdd gnd cell_6t
Xbit_r172_c151 bl_151 br_151 wl_172 vdd gnd cell_6t
Xbit_r173_c151 bl_151 br_151 wl_173 vdd gnd cell_6t
Xbit_r174_c151 bl_151 br_151 wl_174 vdd gnd cell_6t
Xbit_r175_c151 bl_151 br_151 wl_175 vdd gnd cell_6t
Xbit_r176_c151 bl_151 br_151 wl_176 vdd gnd cell_6t
Xbit_r177_c151 bl_151 br_151 wl_177 vdd gnd cell_6t
Xbit_r178_c151 bl_151 br_151 wl_178 vdd gnd cell_6t
Xbit_r179_c151 bl_151 br_151 wl_179 vdd gnd cell_6t
Xbit_r180_c151 bl_151 br_151 wl_180 vdd gnd cell_6t
Xbit_r181_c151 bl_151 br_151 wl_181 vdd gnd cell_6t
Xbit_r182_c151 bl_151 br_151 wl_182 vdd gnd cell_6t
Xbit_r183_c151 bl_151 br_151 wl_183 vdd gnd cell_6t
Xbit_r184_c151 bl_151 br_151 wl_184 vdd gnd cell_6t
Xbit_r185_c151 bl_151 br_151 wl_185 vdd gnd cell_6t
Xbit_r186_c151 bl_151 br_151 wl_186 vdd gnd cell_6t
Xbit_r187_c151 bl_151 br_151 wl_187 vdd gnd cell_6t
Xbit_r188_c151 bl_151 br_151 wl_188 vdd gnd cell_6t
Xbit_r189_c151 bl_151 br_151 wl_189 vdd gnd cell_6t
Xbit_r190_c151 bl_151 br_151 wl_190 vdd gnd cell_6t
Xbit_r191_c151 bl_151 br_151 wl_191 vdd gnd cell_6t
Xbit_r192_c151 bl_151 br_151 wl_192 vdd gnd cell_6t
Xbit_r193_c151 bl_151 br_151 wl_193 vdd gnd cell_6t
Xbit_r194_c151 bl_151 br_151 wl_194 vdd gnd cell_6t
Xbit_r195_c151 bl_151 br_151 wl_195 vdd gnd cell_6t
Xbit_r196_c151 bl_151 br_151 wl_196 vdd gnd cell_6t
Xbit_r197_c151 bl_151 br_151 wl_197 vdd gnd cell_6t
Xbit_r198_c151 bl_151 br_151 wl_198 vdd gnd cell_6t
Xbit_r199_c151 bl_151 br_151 wl_199 vdd gnd cell_6t
Xbit_r200_c151 bl_151 br_151 wl_200 vdd gnd cell_6t
Xbit_r201_c151 bl_151 br_151 wl_201 vdd gnd cell_6t
Xbit_r202_c151 bl_151 br_151 wl_202 vdd gnd cell_6t
Xbit_r203_c151 bl_151 br_151 wl_203 vdd gnd cell_6t
Xbit_r204_c151 bl_151 br_151 wl_204 vdd gnd cell_6t
Xbit_r205_c151 bl_151 br_151 wl_205 vdd gnd cell_6t
Xbit_r206_c151 bl_151 br_151 wl_206 vdd gnd cell_6t
Xbit_r207_c151 bl_151 br_151 wl_207 vdd gnd cell_6t
Xbit_r208_c151 bl_151 br_151 wl_208 vdd gnd cell_6t
Xbit_r209_c151 bl_151 br_151 wl_209 vdd gnd cell_6t
Xbit_r210_c151 bl_151 br_151 wl_210 vdd gnd cell_6t
Xbit_r211_c151 bl_151 br_151 wl_211 vdd gnd cell_6t
Xbit_r212_c151 bl_151 br_151 wl_212 vdd gnd cell_6t
Xbit_r213_c151 bl_151 br_151 wl_213 vdd gnd cell_6t
Xbit_r214_c151 bl_151 br_151 wl_214 vdd gnd cell_6t
Xbit_r215_c151 bl_151 br_151 wl_215 vdd gnd cell_6t
Xbit_r216_c151 bl_151 br_151 wl_216 vdd gnd cell_6t
Xbit_r217_c151 bl_151 br_151 wl_217 vdd gnd cell_6t
Xbit_r218_c151 bl_151 br_151 wl_218 vdd gnd cell_6t
Xbit_r219_c151 bl_151 br_151 wl_219 vdd gnd cell_6t
Xbit_r220_c151 bl_151 br_151 wl_220 vdd gnd cell_6t
Xbit_r221_c151 bl_151 br_151 wl_221 vdd gnd cell_6t
Xbit_r222_c151 bl_151 br_151 wl_222 vdd gnd cell_6t
Xbit_r223_c151 bl_151 br_151 wl_223 vdd gnd cell_6t
Xbit_r224_c151 bl_151 br_151 wl_224 vdd gnd cell_6t
Xbit_r225_c151 bl_151 br_151 wl_225 vdd gnd cell_6t
Xbit_r226_c151 bl_151 br_151 wl_226 vdd gnd cell_6t
Xbit_r227_c151 bl_151 br_151 wl_227 vdd gnd cell_6t
Xbit_r228_c151 bl_151 br_151 wl_228 vdd gnd cell_6t
Xbit_r229_c151 bl_151 br_151 wl_229 vdd gnd cell_6t
Xbit_r230_c151 bl_151 br_151 wl_230 vdd gnd cell_6t
Xbit_r231_c151 bl_151 br_151 wl_231 vdd gnd cell_6t
Xbit_r232_c151 bl_151 br_151 wl_232 vdd gnd cell_6t
Xbit_r233_c151 bl_151 br_151 wl_233 vdd gnd cell_6t
Xbit_r234_c151 bl_151 br_151 wl_234 vdd gnd cell_6t
Xbit_r235_c151 bl_151 br_151 wl_235 vdd gnd cell_6t
Xbit_r236_c151 bl_151 br_151 wl_236 vdd gnd cell_6t
Xbit_r237_c151 bl_151 br_151 wl_237 vdd gnd cell_6t
Xbit_r238_c151 bl_151 br_151 wl_238 vdd gnd cell_6t
Xbit_r239_c151 bl_151 br_151 wl_239 vdd gnd cell_6t
Xbit_r240_c151 bl_151 br_151 wl_240 vdd gnd cell_6t
Xbit_r241_c151 bl_151 br_151 wl_241 vdd gnd cell_6t
Xbit_r242_c151 bl_151 br_151 wl_242 vdd gnd cell_6t
Xbit_r243_c151 bl_151 br_151 wl_243 vdd gnd cell_6t
Xbit_r244_c151 bl_151 br_151 wl_244 vdd gnd cell_6t
Xbit_r245_c151 bl_151 br_151 wl_245 vdd gnd cell_6t
Xbit_r246_c151 bl_151 br_151 wl_246 vdd gnd cell_6t
Xbit_r247_c151 bl_151 br_151 wl_247 vdd gnd cell_6t
Xbit_r248_c151 bl_151 br_151 wl_248 vdd gnd cell_6t
Xbit_r249_c151 bl_151 br_151 wl_249 vdd gnd cell_6t
Xbit_r250_c151 bl_151 br_151 wl_250 vdd gnd cell_6t
Xbit_r251_c151 bl_151 br_151 wl_251 vdd gnd cell_6t
Xbit_r252_c151 bl_151 br_151 wl_252 vdd gnd cell_6t
Xbit_r253_c151 bl_151 br_151 wl_253 vdd gnd cell_6t
Xbit_r254_c151 bl_151 br_151 wl_254 vdd gnd cell_6t
Xbit_r255_c151 bl_151 br_151 wl_255 vdd gnd cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd cell_6t
Xbit_r1_c152 bl_152 br_152 wl_1 vdd gnd cell_6t
Xbit_r2_c152 bl_152 br_152 wl_2 vdd gnd cell_6t
Xbit_r3_c152 bl_152 br_152 wl_3 vdd gnd cell_6t
Xbit_r4_c152 bl_152 br_152 wl_4 vdd gnd cell_6t
Xbit_r5_c152 bl_152 br_152 wl_5 vdd gnd cell_6t
Xbit_r6_c152 bl_152 br_152 wl_6 vdd gnd cell_6t
Xbit_r7_c152 bl_152 br_152 wl_7 vdd gnd cell_6t
Xbit_r8_c152 bl_152 br_152 wl_8 vdd gnd cell_6t
Xbit_r9_c152 bl_152 br_152 wl_9 vdd gnd cell_6t
Xbit_r10_c152 bl_152 br_152 wl_10 vdd gnd cell_6t
Xbit_r11_c152 bl_152 br_152 wl_11 vdd gnd cell_6t
Xbit_r12_c152 bl_152 br_152 wl_12 vdd gnd cell_6t
Xbit_r13_c152 bl_152 br_152 wl_13 vdd gnd cell_6t
Xbit_r14_c152 bl_152 br_152 wl_14 vdd gnd cell_6t
Xbit_r15_c152 bl_152 br_152 wl_15 vdd gnd cell_6t
Xbit_r16_c152 bl_152 br_152 wl_16 vdd gnd cell_6t
Xbit_r17_c152 bl_152 br_152 wl_17 vdd gnd cell_6t
Xbit_r18_c152 bl_152 br_152 wl_18 vdd gnd cell_6t
Xbit_r19_c152 bl_152 br_152 wl_19 vdd gnd cell_6t
Xbit_r20_c152 bl_152 br_152 wl_20 vdd gnd cell_6t
Xbit_r21_c152 bl_152 br_152 wl_21 vdd gnd cell_6t
Xbit_r22_c152 bl_152 br_152 wl_22 vdd gnd cell_6t
Xbit_r23_c152 bl_152 br_152 wl_23 vdd gnd cell_6t
Xbit_r24_c152 bl_152 br_152 wl_24 vdd gnd cell_6t
Xbit_r25_c152 bl_152 br_152 wl_25 vdd gnd cell_6t
Xbit_r26_c152 bl_152 br_152 wl_26 vdd gnd cell_6t
Xbit_r27_c152 bl_152 br_152 wl_27 vdd gnd cell_6t
Xbit_r28_c152 bl_152 br_152 wl_28 vdd gnd cell_6t
Xbit_r29_c152 bl_152 br_152 wl_29 vdd gnd cell_6t
Xbit_r30_c152 bl_152 br_152 wl_30 vdd gnd cell_6t
Xbit_r31_c152 bl_152 br_152 wl_31 vdd gnd cell_6t
Xbit_r32_c152 bl_152 br_152 wl_32 vdd gnd cell_6t
Xbit_r33_c152 bl_152 br_152 wl_33 vdd gnd cell_6t
Xbit_r34_c152 bl_152 br_152 wl_34 vdd gnd cell_6t
Xbit_r35_c152 bl_152 br_152 wl_35 vdd gnd cell_6t
Xbit_r36_c152 bl_152 br_152 wl_36 vdd gnd cell_6t
Xbit_r37_c152 bl_152 br_152 wl_37 vdd gnd cell_6t
Xbit_r38_c152 bl_152 br_152 wl_38 vdd gnd cell_6t
Xbit_r39_c152 bl_152 br_152 wl_39 vdd gnd cell_6t
Xbit_r40_c152 bl_152 br_152 wl_40 vdd gnd cell_6t
Xbit_r41_c152 bl_152 br_152 wl_41 vdd gnd cell_6t
Xbit_r42_c152 bl_152 br_152 wl_42 vdd gnd cell_6t
Xbit_r43_c152 bl_152 br_152 wl_43 vdd gnd cell_6t
Xbit_r44_c152 bl_152 br_152 wl_44 vdd gnd cell_6t
Xbit_r45_c152 bl_152 br_152 wl_45 vdd gnd cell_6t
Xbit_r46_c152 bl_152 br_152 wl_46 vdd gnd cell_6t
Xbit_r47_c152 bl_152 br_152 wl_47 vdd gnd cell_6t
Xbit_r48_c152 bl_152 br_152 wl_48 vdd gnd cell_6t
Xbit_r49_c152 bl_152 br_152 wl_49 vdd gnd cell_6t
Xbit_r50_c152 bl_152 br_152 wl_50 vdd gnd cell_6t
Xbit_r51_c152 bl_152 br_152 wl_51 vdd gnd cell_6t
Xbit_r52_c152 bl_152 br_152 wl_52 vdd gnd cell_6t
Xbit_r53_c152 bl_152 br_152 wl_53 vdd gnd cell_6t
Xbit_r54_c152 bl_152 br_152 wl_54 vdd gnd cell_6t
Xbit_r55_c152 bl_152 br_152 wl_55 vdd gnd cell_6t
Xbit_r56_c152 bl_152 br_152 wl_56 vdd gnd cell_6t
Xbit_r57_c152 bl_152 br_152 wl_57 vdd gnd cell_6t
Xbit_r58_c152 bl_152 br_152 wl_58 vdd gnd cell_6t
Xbit_r59_c152 bl_152 br_152 wl_59 vdd gnd cell_6t
Xbit_r60_c152 bl_152 br_152 wl_60 vdd gnd cell_6t
Xbit_r61_c152 bl_152 br_152 wl_61 vdd gnd cell_6t
Xbit_r62_c152 bl_152 br_152 wl_62 vdd gnd cell_6t
Xbit_r63_c152 bl_152 br_152 wl_63 vdd gnd cell_6t
Xbit_r64_c152 bl_152 br_152 wl_64 vdd gnd cell_6t
Xbit_r65_c152 bl_152 br_152 wl_65 vdd gnd cell_6t
Xbit_r66_c152 bl_152 br_152 wl_66 vdd gnd cell_6t
Xbit_r67_c152 bl_152 br_152 wl_67 vdd gnd cell_6t
Xbit_r68_c152 bl_152 br_152 wl_68 vdd gnd cell_6t
Xbit_r69_c152 bl_152 br_152 wl_69 vdd gnd cell_6t
Xbit_r70_c152 bl_152 br_152 wl_70 vdd gnd cell_6t
Xbit_r71_c152 bl_152 br_152 wl_71 vdd gnd cell_6t
Xbit_r72_c152 bl_152 br_152 wl_72 vdd gnd cell_6t
Xbit_r73_c152 bl_152 br_152 wl_73 vdd gnd cell_6t
Xbit_r74_c152 bl_152 br_152 wl_74 vdd gnd cell_6t
Xbit_r75_c152 bl_152 br_152 wl_75 vdd gnd cell_6t
Xbit_r76_c152 bl_152 br_152 wl_76 vdd gnd cell_6t
Xbit_r77_c152 bl_152 br_152 wl_77 vdd gnd cell_6t
Xbit_r78_c152 bl_152 br_152 wl_78 vdd gnd cell_6t
Xbit_r79_c152 bl_152 br_152 wl_79 vdd gnd cell_6t
Xbit_r80_c152 bl_152 br_152 wl_80 vdd gnd cell_6t
Xbit_r81_c152 bl_152 br_152 wl_81 vdd gnd cell_6t
Xbit_r82_c152 bl_152 br_152 wl_82 vdd gnd cell_6t
Xbit_r83_c152 bl_152 br_152 wl_83 vdd gnd cell_6t
Xbit_r84_c152 bl_152 br_152 wl_84 vdd gnd cell_6t
Xbit_r85_c152 bl_152 br_152 wl_85 vdd gnd cell_6t
Xbit_r86_c152 bl_152 br_152 wl_86 vdd gnd cell_6t
Xbit_r87_c152 bl_152 br_152 wl_87 vdd gnd cell_6t
Xbit_r88_c152 bl_152 br_152 wl_88 vdd gnd cell_6t
Xbit_r89_c152 bl_152 br_152 wl_89 vdd gnd cell_6t
Xbit_r90_c152 bl_152 br_152 wl_90 vdd gnd cell_6t
Xbit_r91_c152 bl_152 br_152 wl_91 vdd gnd cell_6t
Xbit_r92_c152 bl_152 br_152 wl_92 vdd gnd cell_6t
Xbit_r93_c152 bl_152 br_152 wl_93 vdd gnd cell_6t
Xbit_r94_c152 bl_152 br_152 wl_94 vdd gnd cell_6t
Xbit_r95_c152 bl_152 br_152 wl_95 vdd gnd cell_6t
Xbit_r96_c152 bl_152 br_152 wl_96 vdd gnd cell_6t
Xbit_r97_c152 bl_152 br_152 wl_97 vdd gnd cell_6t
Xbit_r98_c152 bl_152 br_152 wl_98 vdd gnd cell_6t
Xbit_r99_c152 bl_152 br_152 wl_99 vdd gnd cell_6t
Xbit_r100_c152 bl_152 br_152 wl_100 vdd gnd cell_6t
Xbit_r101_c152 bl_152 br_152 wl_101 vdd gnd cell_6t
Xbit_r102_c152 bl_152 br_152 wl_102 vdd gnd cell_6t
Xbit_r103_c152 bl_152 br_152 wl_103 vdd gnd cell_6t
Xbit_r104_c152 bl_152 br_152 wl_104 vdd gnd cell_6t
Xbit_r105_c152 bl_152 br_152 wl_105 vdd gnd cell_6t
Xbit_r106_c152 bl_152 br_152 wl_106 vdd gnd cell_6t
Xbit_r107_c152 bl_152 br_152 wl_107 vdd gnd cell_6t
Xbit_r108_c152 bl_152 br_152 wl_108 vdd gnd cell_6t
Xbit_r109_c152 bl_152 br_152 wl_109 vdd gnd cell_6t
Xbit_r110_c152 bl_152 br_152 wl_110 vdd gnd cell_6t
Xbit_r111_c152 bl_152 br_152 wl_111 vdd gnd cell_6t
Xbit_r112_c152 bl_152 br_152 wl_112 vdd gnd cell_6t
Xbit_r113_c152 bl_152 br_152 wl_113 vdd gnd cell_6t
Xbit_r114_c152 bl_152 br_152 wl_114 vdd gnd cell_6t
Xbit_r115_c152 bl_152 br_152 wl_115 vdd gnd cell_6t
Xbit_r116_c152 bl_152 br_152 wl_116 vdd gnd cell_6t
Xbit_r117_c152 bl_152 br_152 wl_117 vdd gnd cell_6t
Xbit_r118_c152 bl_152 br_152 wl_118 vdd gnd cell_6t
Xbit_r119_c152 bl_152 br_152 wl_119 vdd gnd cell_6t
Xbit_r120_c152 bl_152 br_152 wl_120 vdd gnd cell_6t
Xbit_r121_c152 bl_152 br_152 wl_121 vdd gnd cell_6t
Xbit_r122_c152 bl_152 br_152 wl_122 vdd gnd cell_6t
Xbit_r123_c152 bl_152 br_152 wl_123 vdd gnd cell_6t
Xbit_r124_c152 bl_152 br_152 wl_124 vdd gnd cell_6t
Xbit_r125_c152 bl_152 br_152 wl_125 vdd gnd cell_6t
Xbit_r126_c152 bl_152 br_152 wl_126 vdd gnd cell_6t
Xbit_r127_c152 bl_152 br_152 wl_127 vdd gnd cell_6t
Xbit_r128_c152 bl_152 br_152 wl_128 vdd gnd cell_6t
Xbit_r129_c152 bl_152 br_152 wl_129 vdd gnd cell_6t
Xbit_r130_c152 bl_152 br_152 wl_130 vdd gnd cell_6t
Xbit_r131_c152 bl_152 br_152 wl_131 vdd gnd cell_6t
Xbit_r132_c152 bl_152 br_152 wl_132 vdd gnd cell_6t
Xbit_r133_c152 bl_152 br_152 wl_133 vdd gnd cell_6t
Xbit_r134_c152 bl_152 br_152 wl_134 vdd gnd cell_6t
Xbit_r135_c152 bl_152 br_152 wl_135 vdd gnd cell_6t
Xbit_r136_c152 bl_152 br_152 wl_136 vdd gnd cell_6t
Xbit_r137_c152 bl_152 br_152 wl_137 vdd gnd cell_6t
Xbit_r138_c152 bl_152 br_152 wl_138 vdd gnd cell_6t
Xbit_r139_c152 bl_152 br_152 wl_139 vdd gnd cell_6t
Xbit_r140_c152 bl_152 br_152 wl_140 vdd gnd cell_6t
Xbit_r141_c152 bl_152 br_152 wl_141 vdd gnd cell_6t
Xbit_r142_c152 bl_152 br_152 wl_142 vdd gnd cell_6t
Xbit_r143_c152 bl_152 br_152 wl_143 vdd gnd cell_6t
Xbit_r144_c152 bl_152 br_152 wl_144 vdd gnd cell_6t
Xbit_r145_c152 bl_152 br_152 wl_145 vdd gnd cell_6t
Xbit_r146_c152 bl_152 br_152 wl_146 vdd gnd cell_6t
Xbit_r147_c152 bl_152 br_152 wl_147 vdd gnd cell_6t
Xbit_r148_c152 bl_152 br_152 wl_148 vdd gnd cell_6t
Xbit_r149_c152 bl_152 br_152 wl_149 vdd gnd cell_6t
Xbit_r150_c152 bl_152 br_152 wl_150 vdd gnd cell_6t
Xbit_r151_c152 bl_152 br_152 wl_151 vdd gnd cell_6t
Xbit_r152_c152 bl_152 br_152 wl_152 vdd gnd cell_6t
Xbit_r153_c152 bl_152 br_152 wl_153 vdd gnd cell_6t
Xbit_r154_c152 bl_152 br_152 wl_154 vdd gnd cell_6t
Xbit_r155_c152 bl_152 br_152 wl_155 vdd gnd cell_6t
Xbit_r156_c152 bl_152 br_152 wl_156 vdd gnd cell_6t
Xbit_r157_c152 bl_152 br_152 wl_157 vdd gnd cell_6t
Xbit_r158_c152 bl_152 br_152 wl_158 vdd gnd cell_6t
Xbit_r159_c152 bl_152 br_152 wl_159 vdd gnd cell_6t
Xbit_r160_c152 bl_152 br_152 wl_160 vdd gnd cell_6t
Xbit_r161_c152 bl_152 br_152 wl_161 vdd gnd cell_6t
Xbit_r162_c152 bl_152 br_152 wl_162 vdd gnd cell_6t
Xbit_r163_c152 bl_152 br_152 wl_163 vdd gnd cell_6t
Xbit_r164_c152 bl_152 br_152 wl_164 vdd gnd cell_6t
Xbit_r165_c152 bl_152 br_152 wl_165 vdd gnd cell_6t
Xbit_r166_c152 bl_152 br_152 wl_166 vdd gnd cell_6t
Xbit_r167_c152 bl_152 br_152 wl_167 vdd gnd cell_6t
Xbit_r168_c152 bl_152 br_152 wl_168 vdd gnd cell_6t
Xbit_r169_c152 bl_152 br_152 wl_169 vdd gnd cell_6t
Xbit_r170_c152 bl_152 br_152 wl_170 vdd gnd cell_6t
Xbit_r171_c152 bl_152 br_152 wl_171 vdd gnd cell_6t
Xbit_r172_c152 bl_152 br_152 wl_172 vdd gnd cell_6t
Xbit_r173_c152 bl_152 br_152 wl_173 vdd gnd cell_6t
Xbit_r174_c152 bl_152 br_152 wl_174 vdd gnd cell_6t
Xbit_r175_c152 bl_152 br_152 wl_175 vdd gnd cell_6t
Xbit_r176_c152 bl_152 br_152 wl_176 vdd gnd cell_6t
Xbit_r177_c152 bl_152 br_152 wl_177 vdd gnd cell_6t
Xbit_r178_c152 bl_152 br_152 wl_178 vdd gnd cell_6t
Xbit_r179_c152 bl_152 br_152 wl_179 vdd gnd cell_6t
Xbit_r180_c152 bl_152 br_152 wl_180 vdd gnd cell_6t
Xbit_r181_c152 bl_152 br_152 wl_181 vdd gnd cell_6t
Xbit_r182_c152 bl_152 br_152 wl_182 vdd gnd cell_6t
Xbit_r183_c152 bl_152 br_152 wl_183 vdd gnd cell_6t
Xbit_r184_c152 bl_152 br_152 wl_184 vdd gnd cell_6t
Xbit_r185_c152 bl_152 br_152 wl_185 vdd gnd cell_6t
Xbit_r186_c152 bl_152 br_152 wl_186 vdd gnd cell_6t
Xbit_r187_c152 bl_152 br_152 wl_187 vdd gnd cell_6t
Xbit_r188_c152 bl_152 br_152 wl_188 vdd gnd cell_6t
Xbit_r189_c152 bl_152 br_152 wl_189 vdd gnd cell_6t
Xbit_r190_c152 bl_152 br_152 wl_190 vdd gnd cell_6t
Xbit_r191_c152 bl_152 br_152 wl_191 vdd gnd cell_6t
Xbit_r192_c152 bl_152 br_152 wl_192 vdd gnd cell_6t
Xbit_r193_c152 bl_152 br_152 wl_193 vdd gnd cell_6t
Xbit_r194_c152 bl_152 br_152 wl_194 vdd gnd cell_6t
Xbit_r195_c152 bl_152 br_152 wl_195 vdd gnd cell_6t
Xbit_r196_c152 bl_152 br_152 wl_196 vdd gnd cell_6t
Xbit_r197_c152 bl_152 br_152 wl_197 vdd gnd cell_6t
Xbit_r198_c152 bl_152 br_152 wl_198 vdd gnd cell_6t
Xbit_r199_c152 bl_152 br_152 wl_199 vdd gnd cell_6t
Xbit_r200_c152 bl_152 br_152 wl_200 vdd gnd cell_6t
Xbit_r201_c152 bl_152 br_152 wl_201 vdd gnd cell_6t
Xbit_r202_c152 bl_152 br_152 wl_202 vdd gnd cell_6t
Xbit_r203_c152 bl_152 br_152 wl_203 vdd gnd cell_6t
Xbit_r204_c152 bl_152 br_152 wl_204 vdd gnd cell_6t
Xbit_r205_c152 bl_152 br_152 wl_205 vdd gnd cell_6t
Xbit_r206_c152 bl_152 br_152 wl_206 vdd gnd cell_6t
Xbit_r207_c152 bl_152 br_152 wl_207 vdd gnd cell_6t
Xbit_r208_c152 bl_152 br_152 wl_208 vdd gnd cell_6t
Xbit_r209_c152 bl_152 br_152 wl_209 vdd gnd cell_6t
Xbit_r210_c152 bl_152 br_152 wl_210 vdd gnd cell_6t
Xbit_r211_c152 bl_152 br_152 wl_211 vdd gnd cell_6t
Xbit_r212_c152 bl_152 br_152 wl_212 vdd gnd cell_6t
Xbit_r213_c152 bl_152 br_152 wl_213 vdd gnd cell_6t
Xbit_r214_c152 bl_152 br_152 wl_214 vdd gnd cell_6t
Xbit_r215_c152 bl_152 br_152 wl_215 vdd gnd cell_6t
Xbit_r216_c152 bl_152 br_152 wl_216 vdd gnd cell_6t
Xbit_r217_c152 bl_152 br_152 wl_217 vdd gnd cell_6t
Xbit_r218_c152 bl_152 br_152 wl_218 vdd gnd cell_6t
Xbit_r219_c152 bl_152 br_152 wl_219 vdd gnd cell_6t
Xbit_r220_c152 bl_152 br_152 wl_220 vdd gnd cell_6t
Xbit_r221_c152 bl_152 br_152 wl_221 vdd gnd cell_6t
Xbit_r222_c152 bl_152 br_152 wl_222 vdd gnd cell_6t
Xbit_r223_c152 bl_152 br_152 wl_223 vdd gnd cell_6t
Xbit_r224_c152 bl_152 br_152 wl_224 vdd gnd cell_6t
Xbit_r225_c152 bl_152 br_152 wl_225 vdd gnd cell_6t
Xbit_r226_c152 bl_152 br_152 wl_226 vdd gnd cell_6t
Xbit_r227_c152 bl_152 br_152 wl_227 vdd gnd cell_6t
Xbit_r228_c152 bl_152 br_152 wl_228 vdd gnd cell_6t
Xbit_r229_c152 bl_152 br_152 wl_229 vdd gnd cell_6t
Xbit_r230_c152 bl_152 br_152 wl_230 vdd gnd cell_6t
Xbit_r231_c152 bl_152 br_152 wl_231 vdd gnd cell_6t
Xbit_r232_c152 bl_152 br_152 wl_232 vdd gnd cell_6t
Xbit_r233_c152 bl_152 br_152 wl_233 vdd gnd cell_6t
Xbit_r234_c152 bl_152 br_152 wl_234 vdd gnd cell_6t
Xbit_r235_c152 bl_152 br_152 wl_235 vdd gnd cell_6t
Xbit_r236_c152 bl_152 br_152 wl_236 vdd gnd cell_6t
Xbit_r237_c152 bl_152 br_152 wl_237 vdd gnd cell_6t
Xbit_r238_c152 bl_152 br_152 wl_238 vdd gnd cell_6t
Xbit_r239_c152 bl_152 br_152 wl_239 vdd gnd cell_6t
Xbit_r240_c152 bl_152 br_152 wl_240 vdd gnd cell_6t
Xbit_r241_c152 bl_152 br_152 wl_241 vdd gnd cell_6t
Xbit_r242_c152 bl_152 br_152 wl_242 vdd gnd cell_6t
Xbit_r243_c152 bl_152 br_152 wl_243 vdd gnd cell_6t
Xbit_r244_c152 bl_152 br_152 wl_244 vdd gnd cell_6t
Xbit_r245_c152 bl_152 br_152 wl_245 vdd gnd cell_6t
Xbit_r246_c152 bl_152 br_152 wl_246 vdd gnd cell_6t
Xbit_r247_c152 bl_152 br_152 wl_247 vdd gnd cell_6t
Xbit_r248_c152 bl_152 br_152 wl_248 vdd gnd cell_6t
Xbit_r249_c152 bl_152 br_152 wl_249 vdd gnd cell_6t
Xbit_r250_c152 bl_152 br_152 wl_250 vdd gnd cell_6t
Xbit_r251_c152 bl_152 br_152 wl_251 vdd gnd cell_6t
Xbit_r252_c152 bl_152 br_152 wl_252 vdd gnd cell_6t
Xbit_r253_c152 bl_152 br_152 wl_253 vdd gnd cell_6t
Xbit_r254_c152 bl_152 br_152 wl_254 vdd gnd cell_6t
Xbit_r255_c152 bl_152 br_152 wl_255 vdd gnd cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd cell_6t
Xbit_r1_c153 bl_153 br_153 wl_1 vdd gnd cell_6t
Xbit_r2_c153 bl_153 br_153 wl_2 vdd gnd cell_6t
Xbit_r3_c153 bl_153 br_153 wl_3 vdd gnd cell_6t
Xbit_r4_c153 bl_153 br_153 wl_4 vdd gnd cell_6t
Xbit_r5_c153 bl_153 br_153 wl_5 vdd gnd cell_6t
Xbit_r6_c153 bl_153 br_153 wl_6 vdd gnd cell_6t
Xbit_r7_c153 bl_153 br_153 wl_7 vdd gnd cell_6t
Xbit_r8_c153 bl_153 br_153 wl_8 vdd gnd cell_6t
Xbit_r9_c153 bl_153 br_153 wl_9 vdd gnd cell_6t
Xbit_r10_c153 bl_153 br_153 wl_10 vdd gnd cell_6t
Xbit_r11_c153 bl_153 br_153 wl_11 vdd gnd cell_6t
Xbit_r12_c153 bl_153 br_153 wl_12 vdd gnd cell_6t
Xbit_r13_c153 bl_153 br_153 wl_13 vdd gnd cell_6t
Xbit_r14_c153 bl_153 br_153 wl_14 vdd gnd cell_6t
Xbit_r15_c153 bl_153 br_153 wl_15 vdd gnd cell_6t
Xbit_r16_c153 bl_153 br_153 wl_16 vdd gnd cell_6t
Xbit_r17_c153 bl_153 br_153 wl_17 vdd gnd cell_6t
Xbit_r18_c153 bl_153 br_153 wl_18 vdd gnd cell_6t
Xbit_r19_c153 bl_153 br_153 wl_19 vdd gnd cell_6t
Xbit_r20_c153 bl_153 br_153 wl_20 vdd gnd cell_6t
Xbit_r21_c153 bl_153 br_153 wl_21 vdd gnd cell_6t
Xbit_r22_c153 bl_153 br_153 wl_22 vdd gnd cell_6t
Xbit_r23_c153 bl_153 br_153 wl_23 vdd gnd cell_6t
Xbit_r24_c153 bl_153 br_153 wl_24 vdd gnd cell_6t
Xbit_r25_c153 bl_153 br_153 wl_25 vdd gnd cell_6t
Xbit_r26_c153 bl_153 br_153 wl_26 vdd gnd cell_6t
Xbit_r27_c153 bl_153 br_153 wl_27 vdd gnd cell_6t
Xbit_r28_c153 bl_153 br_153 wl_28 vdd gnd cell_6t
Xbit_r29_c153 bl_153 br_153 wl_29 vdd gnd cell_6t
Xbit_r30_c153 bl_153 br_153 wl_30 vdd gnd cell_6t
Xbit_r31_c153 bl_153 br_153 wl_31 vdd gnd cell_6t
Xbit_r32_c153 bl_153 br_153 wl_32 vdd gnd cell_6t
Xbit_r33_c153 bl_153 br_153 wl_33 vdd gnd cell_6t
Xbit_r34_c153 bl_153 br_153 wl_34 vdd gnd cell_6t
Xbit_r35_c153 bl_153 br_153 wl_35 vdd gnd cell_6t
Xbit_r36_c153 bl_153 br_153 wl_36 vdd gnd cell_6t
Xbit_r37_c153 bl_153 br_153 wl_37 vdd gnd cell_6t
Xbit_r38_c153 bl_153 br_153 wl_38 vdd gnd cell_6t
Xbit_r39_c153 bl_153 br_153 wl_39 vdd gnd cell_6t
Xbit_r40_c153 bl_153 br_153 wl_40 vdd gnd cell_6t
Xbit_r41_c153 bl_153 br_153 wl_41 vdd gnd cell_6t
Xbit_r42_c153 bl_153 br_153 wl_42 vdd gnd cell_6t
Xbit_r43_c153 bl_153 br_153 wl_43 vdd gnd cell_6t
Xbit_r44_c153 bl_153 br_153 wl_44 vdd gnd cell_6t
Xbit_r45_c153 bl_153 br_153 wl_45 vdd gnd cell_6t
Xbit_r46_c153 bl_153 br_153 wl_46 vdd gnd cell_6t
Xbit_r47_c153 bl_153 br_153 wl_47 vdd gnd cell_6t
Xbit_r48_c153 bl_153 br_153 wl_48 vdd gnd cell_6t
Xbit_r49_c153 bl_153 br_153 wl_49 vdd gnd cell_6t
Xbit_r50_c153 bl_153 br_153 wl_50 vdd gnd cell_6t
Xbit_r51_c153 bl_153 br_153 wl_51 vdd gnd cell_6t
Xbit_r52_c153 bl_153 br_153 wl_52 vdd gnd cell_6t
Xbit_r53_c153 bl_153 br_153 wl_53 vdd gnd cell_6t
Xbit_r54_c153 bl_153 br_153 wl_54 vdd gnd cell_6t
Xbit_r55_c153 bl_153 br_153 wl_55 vdd gnd cell_6t
Xbit_r56_c153 bl_153 br_153 wl_56 vdd gnd cell_6t
Xbit_r57_c153 bl_153 br_153 wl_57 vdd gnd cell_6t
Xbit_r58_c153 bl_153 br_153 wl_58 vdd gnd cell_6t
Xbit_r59_c153 bl_153 br_153 wl_59 vdd gnd cell_6t
Xbit_r60_c153 bl_153 br_153 wl_60 vdd gnd cell_6t
Xbit_r61_c153 bl_153 br_153 wl_61 vdd gnd cell_6t
Xbit_r62_c153 bl_153 br_153 wl_62 vdd gnd cell_6t
Xbit_r63_c153 bl_153 br_153 wl_63 vdd gnd cell_6t
Xbit_r64_c153 bl_153 br_153 wl_64 vdd gnd cell_6t
Xbit_r65_c153 bl_153 br_153 wl_65 vdd gnd cell_6t
Xbit_r66_c153 bl_153 br_153 wl_66 vdd gnd cell_6t
Xbit_r67_c153 bl_153 br_153 wl_67 vdd gnd cell_6t
Xbit_r68_c153 bl_153 br_153 wl_68 vdd gnd cell_6t
Xbit_r69_c153 bl_153 br_153 wl_69 vdd gnd cell_6t
Xbit_r70_c153 bl_153 br_153 wl_70 vdd gnd cell_6t
Xbit_r71_c153 bl_153 br_153 wl_71 vdd gnd cell_6t
Xbit_r72_c153 bl_153 br_153 wl_72 vdd gnd cell_6t
Xbit_r73_c153 bl_153 br_153 wl_73 vdd gnd cell_6t
Xbit_r74_c153 bl_153 br_153 wl_74 vdd gnd cell_6t
Xbit_r75_c153 bl_153 br_153 wl_75 vdd gnd cell_6t
Xbit_r76_c153 bl_153 br_153 wl_76 vdd gnd cell_6t
Xbit_r77_c153 bl_153 br_153 wl_77 vdd gnd cell_6t
Xbit_r78_c153 bl_153 br_153 wl_78 vdd gnd cell_6t
Xbit_r79_c153 bl_153 br_153 wl_79 vdd gnd cell_6t
Xbit_r80_c153 bl_153 br_153 wl_80 vdd gnd cell_6t
Xbit_r81_c153 bl_153 br_153 wl_81 vdd gnd cell_6t
Xbit_r82_c153 bl_153 br_153 wl_82 vdd gnd cell_6t
Xbit_r83_c153 bl_153 br_153 wl_83 vdd gnd cell_6t
Xbit_r84_c153 bl_153 br_153 wl_84 vdd gnd cell_6t
Xbit_r85_c153 bl_153 br_153 wl_85 vdd gnd cell_6t
Xbit_r86_c153 bl_153 br_153 wl_86 vdd gnd cell_6t
Xbit_r87_c153 bl_153 br_153 wl_87 vdd gnd cell_6t
Xbit_r88_c153 bl_153 br_153 wl_88 vdd gnd cell_6t
Xbit_r89_c153 bl_153 br_153 wl_89 vdd gnd cell_6t
Xbit_r90_c153 bl_153 br_153 wl_90 vdd gnd cell_6t
Xbit_r91_c153 bl_153 br_153 wl_91 vdd gnd cell_6t
Xbit_r92_c153 bl_153 br_153 wl_92 vdd gnd cell_6t
Xbit_r93_c153 bl_153 br_153 wl_93 vdd gnd cell_6t
Xbit_r94_c153 bl_153 br_153 wl_94 vdd gnd cell_6t
Xbit_r95_c153 bl_153 br_153 wl_95 vdd gnd cell_6t
Xbit_r96_c153 bl_153 br_153 wl_96 vdd gnd cell_6t
Xbit_r97_c153 bl_153 br_153 wl_97 vdd gnd cell_6t
Xbit_r98_c153 bl_153 br_153 wl_98 vdd gnd cell_6t
Xbit_r99_c153 bl_153 br_153 wl_99 vdd gnd cell_6t
Xbit_r100_c153 bl_153 br_153 wl_100 vdd gnd cell_6t
Xbit_r101_c153 bl_153 br_153 wl_101 vdd gnd cell_6t
Xbit_r102_c153 bl_153 br_153 wl_102 vdd gnd cell_6t
Xbit_r103_c153 bl_153 br_153 wl_103 vdd gnd cell_6t
Xbit_r104_c153 bl_153 br_153 wl_104 vdd gnd cell_6t
Xbit_r105_c153 bl_153 br_153 wl_105 vdd gnd cell_6t
Xbit_r106_c153 bl_153 br_153 wl_106 vdd gnd cell_6t
Xbit_r107_c153 bl_153 br_153 wl_107 vdd gnd cell_6t
Xbit_r108_c153 bl_153 br_153 wl_108 vdd gnd cell_6t
Xbit_r109_c153 bl_153 br_153 wl_109 vdd gnd cell_6t
Xbit_r110_c153 bl_153 br_153 wl_110 vdd gnd cell_6t
Xbit_r111_c153 bl_153 br_153 wl_111 vdd gnd cell_6t
Xbit_r112_c153 bl_153 br_153 wl_112 vdd gnd cell_6t
Xbit_r113_c153 bl_153 br_153 wl_113 vdd gnd cell_6t
Xbit_r114_c153 bl_153 br_153 wl_114 vdd gnd cell_6t
Xbit_r115_c153 bl_153 br_153 wl_115 vdd gnd cell_6t
Xbit_r116_c153 bl_153 br_153 wl_116 vdd gnd cell_6t
Xbit_r117_c153 bl_153 br_153 wl_117 vdd gnd cell_6t
Xbit_r118_c153 bl_153 br_153 wl_118 vdd gnd cell_6t
Xbit_r119_c153 bl_153 br_153 wl_119 vdd gnd cell_6t
Xbit_r120_c153 bl_153 br_153 wl_120 vdd gnd cell_6t
Xbit_r121_c153 bl_153 br_153 wl_121 vdd gnd cell_6t
Xbit_r122_c153 bl_153 br_153 wl_122 vdd gnd cell_6t
Xbit_r123_c153 bl_153 br_153 wl_123 vdd gnd cell_6t
Xbit_r124_c153 bl_153 br_153 wl_124 vdd gnd cell_6t
Xbit_r125_c153 bl_153 br_153 wl_125 vdd gnd cell_6t
Xbit_r126_c153 bl_153 br_153 wl_126 vdd gnd cell_6t
Xbit_r127_c153 bl_153 br_153 wl_127 vdd gnd cell_6t
Xbit_r128_c153 bl_153 br_153 wl_128 vdd gnd cell_6t
Xbit_r129_c153 bl_153 br_153 wl_129 vdd gnd cell_6t
Xbit_r130_c153 bl_153 br_153 wl_130 vdd gnd cell_6t
Xbit_r131_c153 bl_153 br_153 wl_131 vdd gnd cell_6t
Xbit_r132_c153 bl_153 br_153 wl_132 vdd gnd cell_6t
Xbit_r133_c153 bl_153 br_153 wl_133 vdd gnd cell_6t
Xbit_r134_c153 bl_153 br_153 wl_134 vdd gnd cell_6t
Xbit_r135_c153 bl_153 br_153 wl_135 vdd gnd cell_6t
Xbit_r136_c153 bl_153 br_153 wl_136 vdd gnd cell_6t
Xbit_r137_c153 bl_153 br_153 wl_137 vdd gnd cell_6t
Xbit_r138_c153 bl_153 br_153 wl_138 vdd gnd cell_6t
Xbit_r139_c153 bl_153 br_153 wl_139 vdd gnd cell_6t
Xbit_r140_c153 bl_153 br_153 wl_140 vdd gnd cell_6t
Xbit_r141_c153 bl_153 br_153 wl_141 vdd gnd cell_6t
Xbit_r142_c153 bl_153 br_153 wl_142 vdd gnd cell_6t
Xbit_r143_c153 bl_153 br_153 wl_143 vdd gnd cell_6t
Xbit_r144_c153 bl_153 br_153 wl_144 vdd gnd cell_6t
Xbit_r145_c153 bl_153 br_153 wl_145 vdd gnd cell_6t
Xbit_r146_c153 bl_153 br_153 wl_146 vdd gnd cell_6t
Xbit_r147_c153 bl_153 br_153 wl_147 vdd gnd cell_6t
Xbit_r148_c153 bl_153 br_153 wl_148 vdd gnd cell_6t
Xbit_r149_c153 bl_153 br_153 wl_149 vdd gnd cell_6t
Xbit_r150_c153 bl_153 br_153 wl_150 vdd gnd cell_6t
Xbit_r151_c153 bl_153 br_153 wl_151 vdd gnd cell_6t
Xbit_r152_c153 bl_153 br_153 wl_152 vdd gnd cell_6t
Xbit_r153_c153 bl_153 br_153 wl_153 vdd gnd cell_6t
Xbit_r154_c153 bl_153 br_153 wl_154 vdd gnd cell_6t
Xbit_r155_c153 bl_153 br_153 wl_155 vdd gnd cell_6t
Xbit_r156_c153 bl_153 br_153 wl_156 vdd gnd cell_6t
Xbit_r157_c153 bl_153 br_153 wl_157 vdd gnd cell_6t
Xbit_r158_c153 bl_153 br_153 wl_158 vdd gnd cell_6t
Xbit_r159_c153 bl_153 br_153 wl_159 vdd gnd cell_6t
Xbit_r160_c153 bl_153 br_153 wl_160 vdd gnd cell_6t
Xbit_r161_c153 bl_153 br_153 wl_161 vdd gnd cell_6t
Xbit_r162_c153 bl_153 br_153 wl_162 vdd gnd cell_6t
Xbit_r163_c153 bl_153 br_153 wl_163 vdd gnd cell_6t
Xbit_r164_c153 bl_153 br_153 wl_164 vdd gnd cell_6t
Xbit_r165_c153 bl_153 br_153 wl_165 vdd gnd cell_6t
Xbit_r166_c153 bl_153 br_153 wl_166 vdd gnd cell_6t
Xbit_r167_c153 bl_153 br_153 wl_167 vdd gnd cell_6t
Xbit_r168_c153 bl_153 br_153 wl_168 vdd gnd cell_6t
Xbit_r169_c153 bl_153 br_153 wl_169 vdd gnd cell_6t
Xbit_r170_c153 bl_153 br_153 wl_170 vdd gnd cell_6t
Xbit_r171_c153 bl_153 br_153 wl_171 vdd gnd cell_6t
Xbit_r172_c153 bl_153 br_153 wl_172 vdd gnd cell_6t
Xbit_r173_c153 bl_153 br_153 wl_173 vdd gnd cell_6t
Xbit_r174_c153 bl_153 br_153 wl_174 vdd gnd cell_6t
Xbit_r175_c153 bl_153 br_153 wl_175 vdd gnd cell_6t
Xbit_r176_c153 bl_153 br_153 wl_176 vdd gnd cell_6t
Xbit_r177_c153 bl_153 br_153 wl_177 vdd gnd cell_6t
Xbit_r178_c153 bl_153 br_153 wl_178 vdd gnd cell_6t
Xbit_r179_c153 bl_153 br_153 wl_179 vdd gnd cell_6t
Xbit_r180_c153 bl_153 br_153 wl_180 vdd gnd cell_6t
Xbit_r181_c153 bl_153 br_153 wl_181 vdd gnd cell_6t
Xbit_r182_c153 bl_153 br_153 wl_182 vdd gnd cell_6t
Xbit_r183_c153 bl_153 br_153 wl_183 vdd gnd cell_6t
Xbit_r184_c153 bl_153 br_153 wl_184 vdd gnd cell_6t
Xbit_r185_c153 bl_153 br_153 wl_185 vdd gnd cell_6t
Xbit_r186_c153 bl_153 br_153 wl_186 vdd gnd cell_6t
Xbit_r187_c153 bl_153 br_153 wl_187 vdd gnd cell_6t
Xbit_r188_c153 bl_153 br_153 wl_188 vdd gnd cell_6t
Xbit_r189_c153 bl_153 br_153 wl_189 vdd gnd cell_6t
Xbit_r190_c153 bl_153 br_153 wl_190 vdd gnd cell_6t
Xbit_r191_c153 bl_153 br_153 wl_191 vdd gnd cell_6t
Xbit_r192_c153 bl_153 br_153 wl_192 vdd gnd cell_6t
Xbit_r193_c153 bl_153 br_153 wl_193 vdd gnd cell_6t
Xbit_r194_c153 bl_153 br_153 wl_194 vdd gnd cell_6t
Xbit_r195_c153 bl_153 br_153 wl_195 vdd gnd cell_6t
Xbit_r196_c153 bl_153 br_153 wl_196 vdd gnd cell_6t
Xbit_r197_c153 bl_153 br_153 wl_197 vdd gnd cell_6t
Xbit_r198_c153 bl_153 br_153 wl_198 vdd gnd cell_6t
Xbit_r199_c153 bl_153 br_153 wl_199 vdd gnd cell_6t
Xbit_r200_c153 bl_153 br_153 wl_200 vdd gnd cell_6t
Xbit_r201_c153 bl_153 br_153 wl_201 vdd gnd cell_6t
Xbit_r202_c153 bl_153 br_153 wl_202 vdd gnd cell_6t
Xbit_r203_c153 bl_153 br_153 wl_203 vdd gnd cell_6t
Xbit_r204_c153 bl_153 br_153 wl_204 vdd gnd cell_6t
Xbit_r205_c153 bl_153 br_153 wl_205 vdd gnd cell_6t
Xbit_r206_c153 bl_153 br_153 wl_206 vdd gnd cell_6t
Xbit_r207_c153 bl_153 br_153 wl_207 vdd gnd cell_6t
Xbit_r208_c153 bl_153 br_153 wl_208 vdd gnd cell_6t
Xbit_r209_c153 bl_153 br_153 wl_209 vdd gnd cell_6t
Xbit_r210_c153 bl_153 br_153 wl_210 vdd gnd cell_6t
Xbit_r211_c153 bl_153 br_153 wl_211 vdd gnd cell_6t
Xbit_r212_c153 bl_153 br_153 wl_212 vdd gnd cell_6t
Xbit_r213_c153 bl_153 br_153 wl_213 vdd gnd cell_6t
Xbit_r214_c153 bl_153 br_153 wl_214 vdd gnd cell_6t
Xbit_r215_c153 bl_153 br_153 wl_215 vdd gnd cell_6t
Xbit_r216_c153 bl_153 br_153 wl_216 vdd gnd cell_6t
Xbit_r217_c153 bl_153 br_153 wl_217 vdd gnd cell_6t
Xbit_r218_c153 bl_153 br_153 wl_218 vdd gnd cell_6t
Xbit_r219_c153 bl_153 br_153 wl_219 vdd gnd cell_6t
Xbit_r220_c153 bl_153 br_153 wl_220 vdd gnd cell_6t
Xbit_r221_c153 bl_153 br_153 wl_221 vdd gnd cell_6t
Xbit_r222_c153 bl_153 br_153 wl_222 vdd gnd cell_6t
Xbit_r223_c153 bl_153 br_153 wl_223 vdd gnd cell_6t
Xbit_r224_c153 bl_153 br_153 wl_224 vdd gnd cell_6t
Xbit_r225_c153 bl_153 br_153 wl_225 vdd gnd cell_6t
Xbit_r226_c153 bl_153 br_153 wl_226 vdd gnd cell_6t
Xbit_r227_c153 bl_153 br_153 wl_227 vdd gnd cell_6t
Xbit_r228_c153 bl_153 br_153 wl_228 vdd gnd cell_6t
Xbit_r229_c153 bl_153 br_153 wl_229 vdd gnd cell_6t
Xbit_r230_c153 bl_153 br_153 wl_230 vdd gnd cell_6t
Xbit_r231_c153 bl_153 br_153 wl_231 vdd gnd cell_6t
Xbit_r232_c153 bl_153 br_153 wl_232 vdd gnd cell_6t
Xbit_r233_c153 bl_153 br_153 wl_233 vdd gnd cell_6t
Xbit_r234_c153 bl_153 br_153 wl_234 vdd gnd cell_6t
Xbit_r235_c153 bl_153 br_153 wl_235 vdd gnd cell_6t
Xbit_r236_c153 bl_153 br_153 wl_236 vdd gnd cell_6t
Xbit_r237_c153 bl_153 br_153 wl_237 vdd gnd cell_6t
Xbit_r238_c153 bl_153 br_153 wl_238 vdd gnd cell_6t
Xbit_r239_c153 bl_153 br_153 wl_239 vdd gnd cell_6t
Xbit_r240_c153 bl_153 br_153 wl_240 vdd gnd cell_6t
Xbit_r241_c153 bl_153 br_153 wl_241 vdd gnd cell_6t
Xbit_r242_c153 bl_153 br_153 wl_242 vdd gnd cell_6t
Xbit_r243_c153 bl_153 br_153 wl_243 vdd gnd cell_6t
Xbit_r244_c153 bl_153 br_153 wl_244 vdd gnd cell_6t
Xbit_r245_c153 bl_153 br_153 wl_245 vdd gnd cell_6t
Xbit_r246_c153 bl_153 br_153 wl_246 vdd gnd cell_6t
Xbit_r247_c153 bl_153 br_153 wl_247 vdd gnd cell_6t
Xbit_r248_c153 bl_153 br_153 wl_248 vdd gnd cell_6t
Xbit_r249_c153 bl_153 br_153 wl_249 vdd gnd cell_6t
Xbit_r250_c153 bl_153 br_153 wl_250 vdd gnd cell_6t
Xbit_r251_c153 bl_153 br_153 wl_251 vdd gnd cell_6t
Xbit_r252_c153 bl_153 br_153 wl_252 vdd gnd cell_6t
Xbit_r253_c153 bl_153 br_153 wl_253 vdd gnd cell_6t
Xbit_r254_c153 bl_153 br_153 wl_254 vdd gnd cell_6t
Xbit_r255_c153 bl_153 br_153 wl_255 vdd gnd cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd cell_6t
Xbit_r1_c154 bl_154 br_154 wl_1 vdd gnd cell_6t
Xbit_r2_c154 bl_154 br_154 wl_2 vdd gnd cell_6t
Xbit_r3_c154 bl_154 br_154 wl_3 vdd gnd cell_6t
Xbit_r4_c154 bl_154 br_154 wl_4 vdd gnd cell_6t
Xbit_r5_c154 bl_154 br_154 wl_5 vdd gnd cell_6t
Xbit_r6_c154 bl_154 br_154 wl_6 vdd gnd cell_6t
Xbit_r7_c154 bl_154 br_154 wl_7 vdd gnd cell_6t
Xbit_r8_c154 bl_154 br_154 wl_8 vdd gnd cell_6t
Xbit_r9_c154 bl_154 br_154 wl_9 vdd gnd cell_6t
Xbit_r10_c154 bl_154 br_154 wl_10 vdd gnd cell_6t
Xbit_r11_c154 bl_154 br_154 wl_11 vdd gnd cell_6t
Xbit_r12_c154 bl_154 br_154 wl_12 vdd gnd cell_6t
Xbit_r13_c154 bl_154 br_154 wl_13 vdd gnd cell_6t
Xbit_r14_c154 bl_154 br_154 wl_14 vdd gnd cell_6t
Xbit_r15_c154 bl_154 br_154 wl_15 vdd gnd cell_6t
Xbit_r16_c154 bl_154 br_154 wl_16 vdd gnd cell_6t
Xbit_r17_c154 bl_154 br_154 wl_17 vdd gnd cell_6t
Xbit_r18_c154 bl_154 br_154 wl_18 vdd gnd cell_6t
Xbit_r19_c154 bl_154 br_154 wl_19 vdd gnd cell_6t
Xbit_r20_c154 bl_154 br_154 wl_20 vdd gnd cell_6t
Xbit_r21_c154 bl_154 br_154 wl_21 vdd gnd cell_6t
Xbit_r22_c154 bl_154 br_154 wl_22 vdd gnd cell_6t
Xbit_r23_c154 bl_154 br_154 wl_23 vdd gnd cell_6t
Xbit_r24_c154 bl_154 br_154 wl_24 vdd gnd cell_6t
Xbit_r25_c154 bl_154 br_154 wl_25 vdd gnd cell_6t
Xbit_r26_c154 bl_154 br_154 wl_26 vdd gnd cell_6t
Xbit_r27_c154 bl_154 br_154 wl_27 vdd gnd cell_6t
Xbit_r28_c154 bl_154 br_154 wl_28 vdd gnd cell_6t
Xbit_r29_c154 bl_154 br_154 wl_29 vdd gnd cell_6t
Xbit_r30_c154 bl_154 br_154 wl_30 vdd gnd cell_6t
Xbit_r31_c154 bl_154 br_154 wl_31 vdd gnd cell_6t
Xbit_r32_c154 bl_154 br_154 wl_32 vdd gnd cell_6t
Xbit_r33_c154 bl_154 br_154 wl_33 vdd gnd cell_6t
Xbit_r34_c154 bl_154 br_154 wl_34 vdd gnd cell_6t
Xbit_r35_c154 bl_154 br_154 wl_35 vdd gnd cell_6t
Xbit_r36_c154 bl_154 br_154 wl_36 vdd gnd cell_6t
Xbit_r37_c154 bl_154 br_154 wl_37 vdd gnd cell_6t
Xbit_r38_c154 bl_154 br_154 wl_38 vdd gnd cell_6t
Xbit_r39_c154 bl_154 br_154 wl_39 vdd gnd cell_6t
Xbit_r40_c154 bl_154 br_154 wl_40 vdd gnd cell_6t
Xbit_r41_c154 bl_154 br_154 wl_41 vdd gnd cell_6t
Xbit_r42_c154 bl_154 br_154 wl_42 vdd gnd cell_6t
Xbit_r43_c154 bl_154 br_154 wl_43 vdd gnd cell_6t
Xbit_r44_c154 bl_154 br_154 wl_44 vdd gnd cell_6t
Xbit_r45_c154 bl_154 br_154 wl_45 vdd gnd cell_6t
Xbit_r46_c154 bl_154 br_154 wl_46 vdd gnd cell_6t
Xbit_r47_c154 bl_154 br_154 wl_47 vdd gnd cell_6t
Xbit_r48_c154 bl_154 br_154 wl_48 vdd gnd cell_6t
Xbit_r49_c154 bl_154 br_154 wl_49 vdd gnd cell_6t
Xbit_r50_c154 bl_154 br_154 wl_50 vdd gnd cell_6t
Xbit_r51_c154 bl_154 br_154 wl_51 vdd gnd cell_6t
Xbit_r52_c154 bl_154 br_154 wl_52 vdd gnd cell_6t
Xbit_r53_c154 bl_154 br_154 wl_53 vdd gnd cell_6t
Xbit_r54_c154 bl_154 br_154 wl_54 vdd gnd cell_6t
Xbit_r55_c154 bl_154 br_154 wl_55 vdd gnd cell_6t
Xbit_r56_c154 bl_154 br_154 wl_56 vdd gnd cell_6t
Xbit_r57_c154 bl_154 br_154 wl_57 vdd gnd cell_6t
Xbit_r58_c154 bl_154 br_154 wl_58 vdd gnd cell_6t
Xbit_r59_c154 bl_154 br_154 wl_59 vdd gnd cell_6t
Xbit_r60_c154 bl_154 br_154 wl_60 vdd gnd cell_6t
Xbit_r61_c154 bl_154 br_154 wl_61 vdd gnd cell_6t
Xbit_r62_c154 bl_154 br_154 wl_62 vdd gnd cell_6t
Xbit_r63_c154 bl_154 br_154 wl_63 vdd gnd cell_6t
Xbit_r64_c154 bl_154 br_154 wl_64 vdd gnd cell_6t
Xbit_r65_c154 bl_154 br_154 wl_65 vdd gnd cell_6t
Xbit_r66_c154 bl_154 br_154 wl_66 vdd gnd cell_6t
Xbit_r67_c154 bl_154 br_154 wl_67 vdd gnd cell_6t
Xbit_r68_c154 bl_154 br_154 wl_68 vdd gnd cell_6t
Xbit_r69_c154 bl_154 br_154 wl_69 vdd gnd cell_6t
Xbit_r70_c154 bl_154 br_154 wl_70 vdd gnd cell_6t
Xbit_r71_c154 bl_154 br_154 wl_71 vdd gnd cell_6t
Xbit_r72_c154 bl_154 br_154 wl_72 vdd gnd cell_6t
Xbit_r73_c154 bl_154 br_154 wl_73 vdd gnd cell_6t
Xbit_r74_c154 bl_154 br_154 wl_74 vdd gnd cell_6t
Xbit_r75_c154 bl_154 br_154 wl_75 vdd gnd cell_6t
Xbit_r76_c154 bl_154 br_154 wl_76 vdd gnd cell_6t
Xbit_r77_c154 bl_154 br_154 wl_77 vdd gnd cell_6t
Xbit_r78_c154 bl_154 br_154 wl_78 vdd gnd cell_6t
Xbit_r79_c154 bl_154 br_154 wl_79 vdd gnd cell_6t
Xbit_r80_c154 bl_154 br_154 wl_80 vdd gnd cell_6t
Xbit_r81_c154 bl_154 br_154 wl_81 vdd gnd cell_6t
Xbit_r82_c154 bl_154 br_154 wl_82 vdd gnd cell_6t
Xbit_r83_c154 bl_154 br_154 wl_83 vdd gnd cell_6t
Xbit_r84_c154 bl_154 br_154 wl_84 vdd gnd cell_6t
Xbit_r85_c154 bl_154 br_154 wl_85 vdd gnd cell_6t
Xbit_r86_c154 bl_154 br_154 wl_86 vdd gnd cell_6t
Xbit_r87_c154 bl_154 br_154 wl_87 vdd gnd cell_6t
Xbit_r88_c154 bl_154 br_154 wl_88 vdd gnd cell_6t
Xbit_r89_c154 bl_154 br_154 wl_89 vdd gnd cell_6t
Xbit_r90_c154 bl_154 br_154 wl_90 vdd gnd cell_6t
Xbit_r91_c154 bl_154 br_154 wl_91 vdd gnd cell_6t
Xbit_r92_c154 bl_154 br_154 wl_92 vdd gnd cell_6t
Xbit_r93_c154 bl_154 br_154 wl_93 vdd gnd cell_6t
Xbit_r94_c154 bl_154 br_154 wl_94 vdd gnd cell_6t
Xbit_r95_c154 bl_154 br_154 wl_95 vdd gnd cell_6t
Xbit_r96_c154 bl_154 br_154 wl_96 vdd gnd cell_6t
Xbit_r97_c154 bl_154 br_154 wl_97 vdd gnd cell_6t
Xbit_r98_c154 bl_154 br_154 wl_98 vdd gnd cell_6t
Xbit_r99_c154 bl_154 br_154 wl_99 vdd gnd cell_6t
Xbit_r100_c154 bl_154 br_154 wl_100 vdd gnd cell_6t
Xbit_r101_c154 bl_154 br_154 wl_101 vdd gnd cell_6t
Xbit_r102_c154 bl_154 br_154 wl_102 vdd gnd cell_6t
Xbit_r103_c154 bl_154 br_154 wl_103 vdd gnd cell_6t
Xbit_r104_c154 bl_154 br_154 wl_104 vdd gnd cell_6t
Xbit_r105_c154 bl_154 br_154 wl_105 vdd gnd cell_6t
Xbit_r106_c154 bl_154 br_154 wl_106 vdd gnd cell_6t
Xbit_r107_c154 bl_154 br_154 wl_107 vdd gnd cell_6t
Xbit_r108_c154 bl_154 br_154 wl_108 vdd gnd cell_6t
Xbit_r109_c154 bl_154 br_154 wl_109 vdd gnd cell_6t
Xbit_r110_c154 bl_154 br_154 wl_110 vdd gnd cell_6t
Xbit_r111_c154 bl_154 br_154 wl_111 vdd gnd cell_6t
Xbit_r112_c154 bl_154 br_154 wl_112 vdd gnd cell_6t
Xbit_r113_c154 bl_154 br_154 wl_113 vdd gnd cell_6t
Xbit_r114_c154 bl_154 br_154 wl_114 vdd gnd cell_6t
Xbit_r115_c154 bl_154 br_154 wl_115 vdd gnd cell_6t
Xbit_r116_c154 bl_154 br_154 wl_116 vdd gnd cell_6t
Xbit_r117_c154 bl_154 br_154 wl_117 vdd gnd cell_6t
Xbit_r118_c154 bl_154 br_154 wl_118 vdd gnd cell_6t
Xbit_r119_c154 bl_154 br_154 wl_119 vdd gnd cell_6t
Xbit_r120_c154 bl_154 br_154 wl_120 vdd gnd cell_6t
Xbit_r121_c154 bl_154 br_154 wl_121 vdd gnd cell_6t
Xbit_r122_c154 bl_154 br_154 wl_122 vdd gnd cell_6t
Xbit_r123_c154 bl_154 br_154 wl_123 vdd gnd cell_6t
Xbit_r124_c154 bl_154 br_154 wl_124 vdd gnd cell_6t
Xbit_r125_c154 bl_154 br_154 wl_125 vdd gnd cell_6t
Xbit_r126_c154 bl_154 br_154 wl_126 vdd gnd cell_6t
Xbit_r127_c154 bl_154 br_154 wl_127 vdd gnd cell_6t
Xbit_r128_c154 bl_154 br_154 wl_128 vdd gnd cell_6t
Xbit_r129_c154 bl_154 br_154 wl_129 vdd gnd cell_6t
Xbit_r130_c154 bl_154 br_154 wl_130 vdd gnd cell_6t
Xbit_r131_c154 bl_154 br_154 wl_131 vdd gnd cell_6t
Xbit_r132_c154 bl_154 br_154 wl_132 vdd gnd cell_6t
Xbit_r133_c154 bl_154 br_154 wl_133 vdd gnd cell_6t
Xbit_r134_c154 bl_154 br_154 wl_134 vdd gnd cell_6t
Xbit_r135_c154 bl_154 br_154 wl_135 vdd gnd cell_6t
Xbit_r136_c154 bl_154 br_154 wl_136 vdd gnd cell_6t
Xbit_r137_c154 bl_154 br_154 wl_137 vdd gnd cell_6t
Xbit_r138_c154 bl_154 br_154 wl_138 vdd gnd cell_6t
Xbit_r139_c154 bl_154 br_154 wl_139 vdd gnd cell_6t
Xbit_r140_c154 bl_154 br_154 wl_140 vdd gnd cell_6t
Xbit_r141_c154 bl_154 br_154 wl_141 vdd gnd cell_6t
Xbit_r142_c154 bl_154 br_154 wl_142 vdd gnd cell_6t
Xbit_r143_c154 bl_154 br_154 wl_143 vdd gnd cell_6t
Xbit_r144_c154 bl_154 br_154 wl_144 vdd gnd cell_6t
Xbit_r145_c154 bl_154 br_154 wl_145 vdd gnd cell_6t
Xbit_r146_c154 bl_154 br_154 wl_146 vdd gnd cell_6t
Xbit_r147_c154 bl_154 br_154 wl_147 vdd gnd cell_6t
Xbit_r148_c154 bl_154 br_154 wl_148 vdd gnd cell_6t
Xbit_r149_c154 bl_154 br_154 wl_149 vdd gnd cell_6t
Xbit_r150_c154 bl_154 br_154 wl_150 vdd gnd cell_6t
Xbit_r151_c154 bl_154 br_154 wl_151 vdd gnd cell_6t
Xbit_r152_c154 bl_154 br_154 wl_152 vdd gnd cell_6t
Xbit_r153_c154 bl_154 br_154 wl_153 vdd gnd cell_6t
Xbit_r154_c154 bl_154 br_154 wl_154 vdd gnd cell_6t
Xbit_r155_c154 bl_154 br_154 wl_155 vdd gnd cell_6t
Xbit_r156_c154 bl_154 br_154 wl_156 vdd gnd cell_6t
Xbit_r157_c154 bl_154 br_154 wl_157 vdd gnd cell_6t
Xbit_r158_c154 bl_154 br_154 wl_158 vdd gnd cell_6t
Xbit_r159_c154 bl_154 br_154 wl_159 vdd gnd cell_6t
Xbit_r160_c154 bl_154 br_154 wl_160 vdd gnd cell_6t
Xbit_r161_c154 bl_154 br_154 wl_161 vdd gnd cell_6t
Xbit_r162_c154 bl_154 br_154 wl_162 vdd gnd cell_6t
Xbit_r163_c154 bl_154 br_154 wl_163 vdd gnd cell_6t
Xbit_r164_c154 bl_154 br_154 wl_164 vdd gnd cell_6t
Xbit_r165_c154 bl_154 br_154 wl_165 vdd gnd cell_6t
Xbit_r166_c154 bl_154 br_154 wl_166 vdd gnd cell_6t
Xbit_r167_c154 bl_154 br_154 wl_167 vdd gnd cell_6t
Xbit_r168_c154 bl_154 br_154 wl_168 vdd gnd cell_6t
Xbit_r169_c154 bl_154 br_154 wl_169 vdd gnd cell_6t
Xbit_r170_c154 bl_154 br_154 wl_170 vdd gnd cell_6t
Xbit_r171_c154 bl_154 br_154 wl_171 vdd gnd cell_6t
Xbit_r172_c154 bl_154 br_154 wl_172 vdd gnd cell_6t
Xbit_r173_c154 bl_154 br_154 wl_173 vdd gnd cell_6t
Xbit_r174_c154 bl_154 br_154 wl_174 vdd gnd cell_6t
Xbit_r175_c154 bl_154 br_154 wl_175 vdd gnd cell_6t
Xbit_r176_c154 bl_154 br_154 wl_176 vdd gnd cell_6t
Xbit_r177_c154 bl_154 br_154 wl_177 vdd gnd cell_6t
Xbit_r178_c154 bl_154 br_154 wl_178 vdd gnd cell_6t
Xbit_r179_c154 bl_154 br_154 wl_179 vdd gnd cell_6t
Xbit_r180_c154 bl_154 br_154 wl_180 vdd gnd cell_6t
Xbit_r181_c154 bl_154 br_154 wl_181 vdd gnd cell_6t
Xbit_r182_c154 bl_154 br_154 wl_182 vdd gnd cell_6t
Xbit_r183_c154 bl_154 br_154 wl_183 vdd gnd cell_6t
Xbit_r184_c154 bl_154 br_154 wl_184 vdd gnd cell_6t
Xbit_r185_c154 bl_154 br_154 wl_185 vdd gnd cell_6t
Xbit_r186_c154 bl_154 br_154 wl_186 vdd gnd cell_6t
Xbit_r187_c154 bl_154 br_154 wl_187 vdd gnd cell_6t
Xbit_r188_c154 bl_154 br_154 wl_188 vdd gnd cell_6t
Xbit_r189_c154 bl_154 br_154 wl_189 vdd gnd cell_6t
Xbit_r190_c154 bl_154 br_154 wl_190 vdd gnd cell_6t
Xbit_r191_c154 bl_154 br_154 wl_191 vdd gnd cell_6t
Xbit_r192_c154 bl_154 br_154 wl_192 vdd gnd cell_6t
Xbit_r193_c154 bl_154 br_154 wl_193 vdd gnd cell_6t
Xbit_r194_c154 bl_154 br_154 wl_194 vdd gnd cell_6t
Xbit_r195_c154 bl_154 br_154 wl_195 vdd gnd cell_6t
Xbit_r196_c154 bl_154 br_154 wl_196 vdd gnd cell_6t
Xbit_r197_c154 bl_154 br_154 wl_197 vdd gnd cell_6t
Xbit_r198_c154 bl_154 br_154 wl_198 vdd gnd cell_6t
Xbit_r199_c154 bl_154 br_154 wl_199 vdd gnd cell_6t
Xbit_r200_c154 bl_154 br_154 wl_200 vdd gnd cell_6t
Xbit_r201_c154 bl_154 br_154 wl_201 vdd gnd cell_6t
Xbit_r202_c154 bl_154 br_154 wl_202 vdd gnd cell_6t
Xbit_r203_c154 bl_154 br_154 wl_203 vdd gnd cell_6t
Xbit_r204_c154 bl_154 br_154 wl_204 vdd gnd cell_6t
Xbit_r205_c154 bl_154 br_154 wl_205 vdd gnd cell_6t
Xbit_r206_c154 bl_154 br_154 wl_206 vdd gnd cell_6t
Xbit_r207_c154 bl_154 br_154 wl_207 vdd gnd cell_6t
Xbit_r208_c154 bl_154 br_154 wl_208 vdd gnd cell_6t
Xbit_r209_c154 bl_154 br_154 wl_209 vdd gnd cell_6t
Xbit_r210_c154 bl_154 br_154 wl_210 vdd gnd cell_6t
Xbit_r211_c154 bl_154 br_154 wl_211 vdd gnd cell_6t
Xbit_r212_c154 bl_154 br_154 wl_212 vdd gnd cell_6t
Xbit_r213_c154 bl_154 br_154 wl_213 vdd gnd cell_6t
Xbit_r214_c154 bl_154 br_154 wl_214 vdd gnd cell_6t
Xbit_r215_c154 bl_154 br_154 wl_215 vdd gnd cell_6t
Xbit_r216_c154 bl_154 br_154 wl_216 vdd gnd cell_6t
Xbit_r217_c154 bl_154 br_154 wl_217 vdd gnd cell_6t
Xbit_r218_c154 bl_154 br_154 wl_218 vdd gnd cell_6t
Xbit_r219_c154 bl_154 br_154 wl_219 vdd gnd cell_6t
Xbit_r220_c154 bl_154 br_154 wl_220 vdd gnd cell_6t
Xbit_r221_c154 bl_154 br_154 wl_221 vdd gnd cell_6t
Xbit_r222_c154 bl_154 br_154 wl_222 vdd gnd cell_6t
Xbit_r223_c154 bl_154 br_154 wl_223 vdd gnd cell_6t
Xbit_r224_c154 bl_154 br_154 wl_224 vdd gnd cell_6t
Xbit_r225_c154 bl_154 br_154 wl_225 vdd gnd cell_6t
Xbit_r226_c154 bl_154 br_154 wl_226 vdd gnd cell_6t
Xbit_r227_c154 bl_154 br_154 wl_227 vdd gnd cell_6t
Xbit_r228_c154 bl_154 br_154 wl_228 vdd gnd cell_6t
Xbit_r229_c154 bl_154 br_154 wl_229 vdd gnd cell_6t
Xbit_r230_c154 bl_154 br_154 wl_230 vdd gnd cell_6t
Xbit_r231_c154 bl_154 br_154 wl_231 vdd gnd cell_6t
Xbit_r232_c154 bl_154 br_154 wl_232 vdd gnd cell_6t
Xbit_r233_c154 bl_154 br_154 wl_233 vdd gnd cell_6t
Xbit_r234_c154 bl_154 br_154 wl_234 vdd gnd cell_6t
Xbit_r235_c154 bl_154 br_154 wl_235 vdd gnd cell_6t
Xbit_r236_c154 bl_154 br_154 wl_236 vdd gnd cell_6t
Xbit_r237_c154 bl_154 br_154 wl_237 vdd gnd cell_6t
Xbit_r238_c154 bl_154 br_154 wl_238 vdd gnd cell_6t
Xbit_r239_c154 bl_154 br_154 wl_239 vdd gnd cell_6t
Xbit_r240_c154 bl_154 br_154 wl_240 vdd gnd cell_6t
Xbit_r241_c154 bl_154 br_154 wl_241 vdd gnd cell_6t
Xbit_r242_c154 bl_154 br_154 wl_242 vdd gnd cell_6t
Xbit_r243_c154 bl_154 br_154 wl_243 vdd gnd cell_6t
Xbit_r244_c154 bl_154 br_154 wl_244 vdd gnd cell_6t
Xbit_r245_c154 bl_154 br_154 wl_245 vdd gnd cell_6t
Xbit_r246_c154 bl_154 br_154 wl_246 vdd gnd cell_6t
Xbit_r247_c154 bl_154 br_154 wl_247 vdd gnd cell_6t
Xbit_r248_c154 bl_154 br_154 wl_248 vdd gnd cell_6t
Xbit_r249_c154 bl_154 br_154 wl_249 vdd gnd cell_6t
Xbit_r250_c154 bl_154 br_154 wl_250 vdd gnd cell_6t
Xbit_r251_c154 bl_154 br_154 wl_251 vdd gnd cell_6t
Xbit_r252_c154 bl_154 br_154 wl_252 vdd gnd cell_6t
Xbit_r253_c154 bl_154 br_154 wl_253 vdd gnd cell_6t
Xbit_r254_c154 bl_154 br_154 wl_254 vdd gnd cell_6t
Xbit_r255_c154 bl_154 br_154 wl_255 vdd gnd cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd cell_6t
Xbit_r1_c155 bl_155 br_155 wl_1 vdd gnd cell_6t
Xbit_r2_c155 bl_155 br_155 wl_2 vdd gnd cell_6t
Xbit_r3_c155 bl_155 br_155 wl_3 vdd gnd cell_6t
Xbit_r4_c155 bl_155 br_155 wl_4 vdd gnd cell_6t
Xbit_r5_c155 bl_155 br_155 wl_5 vdd gnd cell_6t
Xbit_r6_c155 bl_155 br_155 wl_6 vdd gnd cell_6t
Xbit_r7_c155 bl_155 br_155 wl_7 vdd gnd cell_6t
Xbit_r8_c155 bl_155 br_155 wl_8 vdd gnd cell_6t
Xbit_r9_c155 bl_155 br_155 wl_9 vdd gnd cell_6t
Xbit_r10_c155 bl_155 br_155 wl_10 vdd gnd cell_6t
Xbit_r11_c155 bl_155 br_155 wl_11 vdd gnd cell_6t
Xbit_r12_c155 bl_155 br_155 wl_12 vdd gnd cell_6t
Xbit_r13_c155 bl_155 br_155 wl_13 vdd gnd cell_6t
Xbit_r14_c155 bl_155 br_155 wl_14 vdd gnd cell_6t
Xbit_r15_c155 bl_155 br_155 wl_15 vdd gnd cell_6t
Xbit_r16_c155 bl_155 br_155 wl_16 vdd gnd cell_6t
Xbit_r17_c155 bl_155 br_155 wl_17 vdd gnd cell_6t
Xbit_r18_c155 bl_155 br_155 wl_18 vdd gnd cell_6t
Xbit_r19_c155 bl_155 br_155 wl_19 vdd gnd cell_6t
Xbit_r20_c155 bl_155 br_155 wl_20 vdd gnd cell_6t
Xbit_r21_c155 bl_155 br_155 wl_21 vdd gnd cell_6t
Xbit_r22_c155 bl_155 br_155 wl_22 vdd gnd cell_6t
Xbit_r23_c155 bl_155 br_155 wl_23 vdd gnd cell_6t
Xbit_r24_c155 bl_155 br_155 wl_24 vdd gnd cell_6t
Xbit_r25_c155 bl_155 br_155 wl_25 vdd gnd cell_6t
Xbit_r26_c155 bl_155 br_155 wl_26 vdd gnd cell_6t
Xbit_r27_c155 bl_155 br_155 wl_27 vdd gnd cell_6t
Xbit_r28_c155 bl_155 br_155 wl_28 vdd gnd cell_6t
Xbit_r29_c155 bl_155 br_155 wl_29 vdd gnd cell_6t
Xbit_r30_c155 bl_155 br_155 wl_30 vdd gnd cell_6t
Xbit_r31_c155 bl_155 br_155 wl_31 vdd gnd cell_6t
Xbit_r32_c155 bl_155 br_155 wl_32 vdd gnd cell_6t
Xbit_r33_c155 bl_155 br_155 wl_33 vdd gnd cell_6t
Xbit_r34_c155 bl_155 br_155 wl_34 vdd gnd cell_6t
Xbit_r35_c155 bl_155 br_155 wl_35 vdd gnd cell_6t
Xbit_r36_c155 bl_155 br_155 wl_36 vdd gnd cell_6t
Xbit_r37_c155 bl_155 br_155 wl_37 vdd gnd cell_6t
Xbit_r38_c155 bl_155 br_155 wl_38 vdd gnd cell_6t
Xbit_r39_c155 bl_155 br_155 wl_39 vdd gnd cell_6t
Xbit_r40_c155 bl_155 br_155 wl_40 vdd gnd cell_6t
Xbit_r41_c155 bl_155 br_155 wl_41 vdd gnd cell_6t
Xbit_r42_c155 bl_155 br_155 wl_42 vdd gnd cell_6t
Xbit_r43_c155 bl_155 br_155 wl_43 vdd gnd cell_6t
Xbit_r44_c155 bl_155 br_155 wl_44 vdd gnd cell_6t
Xbit_r45_c155 bl_155 br_155 wl_45 vdd gnd cell_6t
Xbit_r46_c155 bl_155 br_155 wl_46 vdd gnd cell_6t
Xbit_r47_c155 bl_155 br_155 wl_47 vdd gnd cell_6t
Xbit_r48_c155 bl_155 br_155 wl_48 vdd gnd cell_6t
Xbit_r49_c155 bl_155 br_155 wl_49 vdd gnd cell_6t
Xbit_r50_c155 bl_155 br_155 wl_50 vdd gnd cell_6t
Xbit_r51_c155 bl_155 br_155 wl_51 vdd gnd cell_6t
Xbit_r52_c155 bl_155 br_155 wl_52 vdd gnd cell_6t
Xbit_r53_c155 bl_155 br_155 wl_53 vdd gnd cell_6t
Xbit_r54_c155 bl_155 br_155 wl_54 vdd gnd cell_6t
Xbit_r55_c155 bl_155 br_155 wl_55 vdd gnd cell_6t
Xbit_r56_c155 bl_155 br_155 wl_56 vdd gnd cell_6t
Xbit_r57_c155 bl_155 br_155 wl_57 vdd gnd cell_6t
Xbit_r58_c155 bl_155 br_155 wl_58 vdd gnd cell_6t
Xbit_r59_c155 bl_155 br_155 wl_59 vdd gnd cell_6t
Xbit_r60_c155 bl_155 br_155 wl_60 vdd gnd cell_6t
Xbit_r61_c155 bl_155 br_155 wl_61 vdd gnd cell_6t
Xbit_r62_c155 bl_155 br_155 wl_62 vdd gnd cell_6t
Xbit_r63_c155 bl_155 br_155 wl_63 vdd gnd cell_6t
Xbit_r64_c155 bl_155 br_155 wl_64 vdd gnd cell_6t
Xbit_r65_c155 bl_155 br_155 wl_65 vdd gnd cell_6t
Xbit_r66_c155 bl_155 br_155 wl_66 vdd gnd cell_6t
Xbit_r67_c155 bl_155 br_155 wl_67 vdd gnd cell_6t
Xbit_r68_c155 bl_155 br_155 wl_68 vdd gnd cell_6t
Xbit_r69_c155 bl_155 br_155 wl_69 vdd gnd cell_6t
Xbit_r70_c155 bl_155 br_155 wl_70 vdd gnd cell_6t
Xbit_r71_c155 bl_155 br_155 wl_71 vdd gnd cell_6t
Xbit_r72_c155 bl_155 br_155 wl_72 vdd gnd cell_6t
Xbit_r73_c155 bl_155 br_155 wl_73 vdd gnd cell_6t
Xbit_r74_c155 bl_155 br_155 wl_74 vdd gnd cell_6t
Xbit_r75_c155 bl_155 br_155 wl_75 vdd gnd cell_6t
Xbit_r76_c155 bl_155 br_155 wl_76 vdd gnd cell_6t
Xbit_r77_c155 bl_155 br_155 wl_77 vdd gnd cell_6t
Xbit_r78_c155 bl_155 br_155 wl_78 vdd gnd cell_6t
Xbit_r79_c155 bl_155 br_155 wl_79 vdd gnd cell_6t
Xbit_r80_c155 bl_155 br_155 wl_80 vdd gnd cell_6t
Xbit_r81_c155 bl_155 br_155 wl_81 vdd gnd cell_6t
Xbit_r82_c155 bl_155 br_155 wl_82 vdd gnd cell_6t
Xbit_r83_c155 bl_155 br_155 wl_83 vdd gnd cell_6t
Xbit_r84_c155 bl_155 br_155 wl_84 vdd gnd cell_6t
Xbit_r85_c155 bl_155 br_155 wl_85 vdd gnd cell_6t
Xbit_r86_c155 bl_155 br_155 wl_86 vdd gnd cell_6t
Xbit_r87_c155 bl_155 br_155 wl_87 vdd gnd cell_6t
Xbit_r88_c155 bl_155 br_155 wl_88 vdd gnd cell_6t
Xbit_r89_c155 bl_155 br_155 wl_89 vdd gnd cell_6t
Xbit_r90_c155 bl_155 br_155 wl_90 vdd gnd cell_6t
Xbit_r91_c155 bl_155 br_155 wl_91 vdd gnd cell_6t
Xbit_r92_c155 bl_155 br_155 wl_92 vdd gnd cell_6t
Xbit_r93_c155 bl_155 br_155 wl_93 vdd gnd cell_6t
Xbit_r94_c155 bl_155 br_155 wl_94 vdd gnd cell_6t
Xbit_r95_c155 bl_155 br_155 wl_95 vdd gnd cell_6t
Xbit_r96_c155 bl_155 br_155 wl_96 vdd gnd cell_6t
Xbit_r97_c155 bl_155 br_155 wl_97 vdd gnd cell_6t
Xbit_r98_c155 bl_155 br_155 wl_98 vdd gnd cell_6t
Xbit_r99_c155 bl_155 br_155 wl_99 vdd gnd cell_6t
Xbit_r100_c155 bl_155 br_155 wl_100 vdd gnd cell_6t
Xbit_r101_c155 bl_155 br_155 wl_101 vdd gnd cell_6t
Xbit_r102_c155 bl_155 br_155 wl_102 vdd gnd cell_6t
Xbit_r103_c155 bl_155 br_155 wl_103 vdd gnd cell_6t
Xbit_r104_c155 bl_155 br_155 wl_104 vdd gnd cell_6t
Xbit_r105_c155 bl_155 br_155 wl_105 vdd gnd cell_6t
Xbit_r106_c155 bl_155 br_155 wl_106 vdd gnd cell_6t
Xbit_r107_c155 bl_155 br_155 wl_107 vdd gnd cell_6t
Xbit_r108_c155 bl_155 br_155 wl_108 vdd gnd cell_6t
Xbit_r109_c155 bl_155 br_155 wl_109 vdd gnd cell_6t
Xbit_r110_c155 bl_155 br_155 wl_110 vdd gnd cell_6t
Xbit_r111_c155 bl_155 br_155 wl_111 vdd gnd cell_6t
Xbit_r112_c155 bl_155 br_155 wl_112 vdd gnd cell_6t
Xbit_r113_c155 bl_155 br_155 wl_113 vdd gnd cell_6t
Xbit_r114_c155 bl_155 br_155 wl_114 vdd gnd cell_6t
Xbit_r115_c155 bl_155 br_155 wl_115 vdd gnd cell_6t
Xbit_r116_c155 bl_155 br_155 wl_116 vdd gnd cell_6t
Xbit_r117_c155 bl_155 br_155 wl_117 vdd gnd cell_6t
Xbit_r118_c155 bl_155 br_155 wl_118 vdd gnd cell_6t
Xbit_r119_c155 bl_155 br_155 wl_119 vdd gnd cell_6t
Xbit_r120_c155 bl_155 br_155 wl_120 vdd gnd cell_6t
Xbit_r121_c155 bl_155 br_155 wl_121 vdd gnd cell_6t
Xbit_r122_c155 bl_155 br_155 wl_122 vdd gnd cell_6t
Xbit_r123_c155 bl_155 br_155 wl_123 vdd gnd cell_6t
Xbit_r124_c155 bl_155 br_155 wl_124 vdd gnd cell_6t
Xbit_r125_c155 bl_155 br_155 wl_125 vdd gnd cell_6t
Xbit_r126_c155 bl_155 br_155 wl_126 vdd gnd cell_6t
Xbit_r127_c155 bl_155 br_155 wl_127 vdd gnd cell_6t
Xbit_r128_c155 bl_155 br_155 wl_128 vdd gnd cell_6t
Xbit_r129_c155 bl_155 br_155 wl_129 vdd gnd cell_6t
Xbit_r130_c155 bl_155 br_155 wl_130 vdd gnd cell_6t
Xbit_r131_c155 bl_155 br_155 wl_131 vdd gnd cell_6t
Xbit_r132_c155 bl_155 br_155 wl_132 vdd gnd cell_6t
Xbit_r133_c155 bl_155 br_155 wl_133 vdd gnd cell_6t
Xbit_r134_c155 bl_155 br_155 wl_134 vdd gnd cell_6t
Xbit_r135_c155 bl_155 br_155 wl_135 vdd gnd cell_6t
Xbit_r136_c155 bl_155 br_155 wl_136 vdd gnd cell_6t
Xbit_r137_c155 bl_155 br_155 wl_137 vdd gnd cell_6t
Xbit_r138_c155 bl_155 br_155 wl_138 vdd gnd cell_6t
Xbit_r139_c155 bl_155 br_155 wl_139 vdd gnd cell_6t
Xbit_r140_c155 bl_155 br_155 wl_140 vdd gnd cell_6t
Xbit_r141_c155 bl_155 br_155 wl_141 vdd gnd cell_6t
Xbit_r142_c155 bl_155 br_155 wl_142 vdd gnd cell_6t
Xbit_r143_c155 bl_155 br_155 wl_143 vdd gnd cell_6t
Xbit_r144_c155 bl_155 br_155 wl_144 vdd gnd cell_6t
Xbit_r145_c155 bl_155 br_155 wl_145 vdd gnd cell_6t
Xbit_r146_c155 bl_155 br_155 wl_146 vdd gnd cell_6t
Xbit_r147_c155 bl_155 br_155 wl_147 vdd gnd cell_6t
Xbit_r148_c155 bl_155 br_155 wl_148 vdd gnd cell_6t
Xbit_r149_c155 bl_155 br_155 wl_149 vdd gnd cell_6t
Xbit_r150_c155 bl_155 br_155 wl_150 vdd gnd cell_6t
Xbit_r151_c155 bl_155 br_155 wl_151 vdd gnd cell_6t
Xbit_r152_c155 bl_155 br_155 wl_152 vdd gnd cell_6t
Xbit_r153_c155 bl_155 br_155 wl_153 vdd gnd cell_6t
Xbit_r154_c155 bl_155 br_155 wl_154 vdd gnd cell_6t
Xbit_r155_c155 bl_155 br_155 wl_155 vdd gnd cell_6t
Xbit_r156_c155 bl_155 br_155 wl_156 vdd gnd cell_6t
Xbit_r157_c155 bl_155 br_155 wl_157 vdd gnd cell_6t
Xbit_r158_c155 bl_155 br_155 wl_158 vdd gnd cell_6t
Xbit_r159_c155 bl_155 br_155 wl_159 vdd gnd cell_6t
Xbit_r160_c155 bl_155 br_155 wl_160 vdd gnd cell_6t
Xbit_r161_c155 bl_155 br_155 wl_161 vdd gnd cell_6t
Xbit_r162_c155 bl_155 br_155 wl_162 vdd gnd cell_6t
Xbit_r163_c155 bl_155 br_155 wl_163 vdd gnd cell_6t
Xbit_r164_c155 bl_155 br_155 wl_164 vdd gnd cell_6t
Xbit_r165_c155 bl_155 br_155 wl_165 vdd gnd cell_6t
Xbit_r166_c155 bl_155 br_155 wl_166 vdd gnd cell_6t
Xbit_r167_c155 bl_155 br_155 wl_167 vdd gnd cell_6t
Xbit_r168_c155 bl_155 br_155 wl_168 vdd gnd cell_6t
Xbit_r169_c155 bl_155 br_155 wl_169 vdd gnd cell_6t
Xbit_r170_c155 bl_155 br_155 wl_170 vdd gnd cell_6t
Xbit_r171_c155 bl_155 br_155 wl_171 vdd gnd cell_6t
Xbit_r172_c155 bl_155 br_155 wl_172 vdd gnd cell_6t
Xbit_r173_c155 bl_155 br_155 wl_173 vdd gnd cell_6t
Xbit_r174_c155 bl_155 br_155 wl_174 vdd gnd cell_6t
Xbit_r175_c155 bl_155 br_155 wl_175 vdd gnd cell_6t
Xbit_r176_c155 bl_155 br_155 wl_176 vdd gnd cell_6t
Xbit_r177_c155 bl_155 br_155 wl_177 vdd gnd cell_6t
Xbit_r178_c155 bl_155 br_155 wl_178 vdd gnd cell_6t
Xbit_r179_c155 bl_155 br_155 wl_179 vdd gnd cell_6t
Xbit_r180_c155 bl_155 br_155 wl_180 vdd gnd cell_6t
Xbit_r181_c155 bl_155 br_155 wl_181 vdd gnd cell_6t
Xbit_r182_c155 bl_155 br_155 wl_182 vdd gnd cell_6t
Xbit_r183_c155 bl_155 br_155 wl_183 vdd gnd cell_6t
Xbit_r184_c155 bl_155 br_155 wl_184 vdd gnd cell_6t
Xbit_r185_c155 bl_155 br_155 wl_185 vdd gnd cell_6t
Xbit_r186_c155 bl_155 br_155 wl_186 vdd gnd cell_6t
Xbit_r187_c155 bl_155 br_155 wl_187 vdd gnd cell_6t
Xbit_r188_c155 bl_155 br_155 wl_188 vdd gnd cell_6t
Xbit_r189_c155 bl_155 br_155 wl_189 vdd gnd cell_6t
Xbit_r190_c155 bl_155 br_155 wl_190 vdd gnd cell_6t
Xbit_r191_c155 bl_155 br_155 wl_191 vdd gnd cell_6t
Xbit_r192_c155 bl_155 br_155 wl_192 vdd gnd cell_6t
Xbit_r193_c155 bl_155 br_155 wl_193 vdd gnd cell_6t
Xbit_r194_c155 bl_155 br_155 wl_194 vdd gnd cell_6t
Xbit_r195_c155 bl_155 br_155 wl_195 vdd gnd cell_6t
Xbit_r196_c155 bl_155 br_155 wl_196 vdd gnd cell_6t
Xbit_r197_c155 bl_155 br_155 wl_197 vdd gnd cell_6t
Xbit_r198_c155 bl_155 br_155 wl_198 vdd gnd cell_6t
Xbit_r199_c155 bl_155 br_155 wl_199 vdd gnd cell_6t
Xbit_r200_c155 bl_155 br_155 wl_200 vdd gnd cell_6t
Xbit_r201_c155 bl_155 br_155 wl_201 vdd gnd cell_6t
Xbit_r202_c155 bl_155 br_155 wl_202 vdd gnd cell_6t
Xbit_r203_c155 bl_155 br_155 wl_203 vdd gnd cell_6t
Xbit_r204_c155 bl_155 br_155 wl_204 vdd gnd cell_6t
Xbit_r205_c155 bl_155 br_155 wl_205 vdd gnd cell_6t
Xbit_r206_c155 bl_155 br_155 wl_206 vdd gnd cell_6t
Xbit_r207_c155 bl_155 br_155 wl_207 vdd gnd cell_6t
Xbit_r208_c155 bl_155 br_155 wl_208 vdd gnd cell_6t
Xbit_r209_c155 bl_155 br_155 wl_209 vdd gnd cell_6t
Xbit_r210_c155 bl_155 br_155 wl_210 vdd gnd cell_6t
Xbit_r211_c155 bl_155 br_155 wl_211 vdd gnd cell_6t
Xbit_r212_c155 bl_155 br_155 wl_212 vdd gnd cell_6t
Xbit_r213_c155 bl_155 br_155 wl_213 vdd gnd cell_6t
Xbit_r214_c155 bl_155 br_155 wl_214 vdd gnd cell_6t
Xbit_r215_c155 bl_155 br_155 wl_215 vdd gnd cell_6t
Xbit_r216_c155 bl_155 br_155 wl_216 vdd gnd cell_6t
Xbit_r217_c155 bl_155 br_155 wl_217 vdd gnd cell_6t
Xbit_r218_c155 bl_155 br_155 wl_218 vdd gnd cell_6t
Xbit_r219_c155 bl_155 br_155 wl_219 vdd gnd cell_6t
Xbit_r220_c155 bl_155 br_155 wl_220 vdd gnd cell_6t
Xbit_r221_c155 bl_155 br_155 wl_221 vdd gnd cell_6t
Xbit_r222_c155 bl_155 br_155 wl_222 vdd gnd cell_6t
Xbit_r223_c155 bl_155 br_155 wl_223 vdd gnd cell_6t
Xbit_r224_c155 bl_155 br_155 wl_224 vdd gnd cell_6t
Xbit_r225_c155 bl_155 br_155 wl_225 vdd gnd cell_6t
Xbit_r226_c155 bl_155 br_155 wl_226 vdd gnd cell_6t
Xbit_r227_c155 bl_155 br_155 wl_227 vdd gnd cell_6t
Xbit_r228_c155 bl_155 br_155 wl_228 vdd gnd cell_6t
Xbit_r229_c155 bl_155 br_155 wl_229 vdd gnd cell_6t
Xbit_r230_c155 bl_155 br_155 wl_230 vdd gnd cell_6t
Xbit_r231_c155 bl_155 br_155 wl_231 vdd gnd cell_6t
Xbit_r232_c155 bl_155 br_155 wl_232 vdd gnd cell_6t
Xbit_r233_c155 bl_155 br_155 wl_233 vdd gnd cell_6t
Xbit_r234_c155 bl_155 br_155 wl_234 vdd gnd cell_6t
Xbit_r235_c155 bl_155 br_155 wl_235 vdd gnd cell_6t
Xbit_r236_c155 bl_155 br_155 wl_236 vdd gnd cell_6t
Xbit_r237_c155 bl_155 br_155 wl_237 vdd gnd cell_6t
Xbit_r238_c155 bl_155 br_155 wl_238 vdd gnd cell_6t
Xbit_r239_c155 bl_155 br_155 wl_239 vdd gnd cell_6t
Xbit_r240_c155 bl_155 br_155 wl_240 vdd gnd cell_6t
Xbit_r241_c155 bl_155 br_155 wl_241 vdd gnd cell_6t
Xbit_r242_c155 bl_155 br_155 wl_242 vdd gnd cell_6t
Xbit_r243_c155 bl_155 br_155 wl_243 vdd gnd cell_6t
Xbit_r244_c155 bl_155 br_155 wl_244 vdd gnd cell_6t
Xbit_r245_c155 bl_155 br_155 wl_245 vdd gnd cell_6t
Xbit_r246_c155 bl_155 br_155 wl_246 vdd gnd cell_6t
Xbit_r247_c155 bl_155 br_155 wl_247 vdd gnd cell_6t
Xbit_r248_c155 bl_155 br_155 wl_248 vdd gnd cell_6t
Xbit_r249_c155 bl_155 br_155 wl_249 vdd gnd cell_6t
Xbit_r250_c155 bl_155 br_155 wl_250 vdd gnd cell_6t
Xbit_r251_c155 bl_155 br_155 wl_251 vdd gnd cell_6t
Xbit_r252_c155 bl_155 br_155 wl_252 vdd gnd cell_6t
Xbit_r253_c155 bl_155 br_155 wl_253 vdd gnd cell_6t
Xbit_r254_c155 bl_155 br_155 wl_254 vdd gnd cell_6t
Xbit_r255_c155 bl_155 br_155 wl_255 vdd gnd cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd cell_6t
Xbit_r1_c156 bl_156 br_156 wl_1 vdd gnd cell_6t
Xbit_r2_c156 bl_156 br_156 wl_2 vdd gnd cell_6t
Xbit_r3_c156 bl_156 br_156 wl_3 vdd gnd cell_6t
Xbit_r4_c156 bl_156 br_156 wl_4 vdd gnd cell_6t
Xbit_r5_c156 bl_156 br_156 wl_5 vdd gnd cell_6t
Xbit_r6_c156 bl_156 br_156 wl_6 vdd gnd cell_6t
Xbit_r7_c156 bl_156 br_156 wl_7 vdd gnd cell_6t
Xbit_r8_c156 bl_156 br_156 wl_8 vdd gnd cell_6t
Xbit_r9_c156 bl_156 br_156 wl_9 vdd gnd cell_6t
Xbit_r10_c156 bl_156 br_156 wl_10 vdd gnd cell_6t
Xbit_r11_c156 bl_156 br_156 wl_11 vdd gnd cell_6t
Xbit_r12_c156 bl_156 br_156 wl_12 vdd gnd cell_6t
Xbit_r13_c156 bl_156 br_156 wl_13 vdd gnd cell_6t
Xbit_r14_c156 bl_156 br_156 wl_14 vdd gnd cell_6t
Xbit_r15_c156 bl_156 br_156 wl_15 vdd gnd cell_6t
Xbit_r16_c156 bl_156 br_156 wl_16 vdd gnd cell_6t
Xbit_r17_c156 bl_156 br_156 wl_17 vdd gnd cell_6t
Xbit_r18_c156 bl_156 br_156 wl_18 vdd gnd cell_6t
Xbit_r19_c156 bl_156 br_156 wl_19 vdd gnd cell_6t
Xbit_r20_c156 bl_156 br_156 wl_20 vdd gnd cell_6t
Xbit_r21_c156 bl_156 br_156 wl_21 vdd gnd cell_6t
Xbit_r22_c156 bl_156 br_156 wl_22 vdd gnd cell_6t
Xbit_r23_c156 bl_156 br_156 wl_23 vdd gnd cell_6t
Xbit_r24_c156 bl_156 br_156 wl_24 vdd gnd cell_6t
Xbit_r25_c156 bl_156 br_156 wl_25 vdd gnd cell_6t
Xbit_r26_c156 bl_156 br_156 wl_26 vdd gnd cell_6t
Xbit_r27_c156 bl_156 br_156 wl_27 vdd gnd cell_6t
Xbit_r28_c156 bl_156 br_156 wl_28 vdd gnd cell_6t
Xbit_r29_c156 bl_156 br_156 wl_29 vdd gnd cell_6t
Xbit_r30_c156 bl_156 br_156 wl_30 vdd gnd cell_6t
Xbit_r31_c156 bl_156 br_156 wl_31 vdd gnd cell_6t
Xbit_r32_c156 bl_156 br_156 wl_32 vdd gnd cell_6t
Xbit_r33_c156 bl_156 br_156 wl_33 vdd gnd cell_6t
Xbit_r34_c156 bl_156 br_156 wl_34 vdd gnd cell_6t
Xbit_r35_c156 bl_156 br_156 wl_35 vdd gnd cell_6t
Xbit_r36_c156 bl_156 br_156 wl_36 vdd gnd cell_6t
Xbit_r37_c156 bl_156 br_156 wl_37 vdd gnd cell_6t
Xbit_r38_c156 bl_156 br_156 wl_38 vdd gnd cell_6t
Xbit_r39_c156 bl_156 br_156 wl_39 vdd gnd cell_6t
Xbit_r40_c156 bl_156 br_156 wl_40 vdd gnd cell_6t
Xbit_r41_c156 bl_156 br_156 wl_41 vdd gnd cell_6t
Xbit_r42_c156 bl_156 br_156 wl_42 vdd gnd cell_6t
Xbit_r43_c156 bl_156 br_156 wl_43 vdd gnd cell_6t
Xbit_r44_c156 bl_156 br_156 wl_44 vdd gnd cell_6t
Xbit_r45_c156 bl_156 br_156 wl_45 vdd gnd cell_6t
Xbit_r46_c156 bl_156 br_156 wl_46 vdd gnd cell_6t
Xbit_r47_c156 bl_156 br_156 wl_47 vdd gnd cell_6t
Xbit_r48_c156 bl_156 br_156 wl_48 vdd gnd cell_6t
Xbit_r49_c156 bl_156 br_156 wl_49 vdd gnd cell_6t
Xbit_r50_c156 bl_156 br_156 wl_50 vdd gnd cell_6t
Xbit_r51_c156 bl_156 br_156 wl_51 vdd gnd cell_6t
Xbit_r52_c156 bl_156 br_156 wl_52 vdd gnd cell_6t
Xbit_r53_c156 bl_156 br_156 wl_53 vdd gnd cell_6t
Xbit_r54_c156 bl_156 br_156 wl_54 vdd gnd cell_6t
Xbit_r55_c156 bl_156 br_156 wl_55 vdd gnd cell_6t
Xbit_r56_c156 bl_156 br_156 wl_56 vdd gnd cell_6t
Xbit_r57_c156 bl_156 br_156 wl_57 vdd gnd cell_6t
Xbit_r58_c156 bl_156 br_156 wl_58 vdd gnd cell_6t
Xbit_r59_c156 bl_156 br_156 wl_59 vdd gnd cell_6t
Xbit_r60_c156 bl_156 br_156 wl_60 vdd gnd cell_6t
Xbit_r61_c156 bl_156 br_156 wl_61 vdd gnd cell_6t
Xbit_r62_c156 bl_156 br_156 wl_62 vdd gnd cell_6t
Xbit_r63_c156 bl_156 br_156 wl_63 vdd gnd cell_6t
Xbit_r64_c156 bl_156 br_156 wl_64 vdd gnd cell_6t
Xbit_r65_c156 bl_156 br_156 wl_65 vdd gnd cell_6t
Xbit_r66_c156 bl_156 br_156 wl_66 vdd gnd cell_6t
Xbit_r67_c156 bl_156 br_156 wl_67 vdd gnd cell_6t
Xbit_r68_c156 bl_156 br_156 wl_68 vdd gnd cell_6t
Xbit_r69_c156 bl_156 br_156 wl_69 vdd gnd cell_6t
Xbit_r70_c156 bl_156 br_156 wl_70 vdd gnd cell_6t
Xbit_r71_c156 bl_156 br_156 wl_71 vdd gnd cell_6t
Xbit_r72_c156 bl_156 br_156 wl_72 vdd gnd cell_6t
Xbit_r73_c156 bl_156 br_156 wl_73 vdd gnd cell_6t
Xbit_r74_c156 bl_156 br_156 wl_74 vdd gnd cell_6t
Xbit_r75_c156 bl_156 br_156 wl_75 vdd gnd cell_6t
Xbit_r76_c156 bl_156 br_156 wl_76 vdd gnd cell_6t
Xbit_r77_c156 bl_156 br_156 wl_77 vdd gnd cell_6t
Xbit_r78_c156 bl_156 br_156 wl_78 vdd gnd cell_6t
Xbit_r79_c156 bl_156 br_156 wl_79 vdd gnd cell_6t
Xbit_r80_c156 bl_156 br_156 wl_80 vdd gnd cell_6t
Xbit_r81_c156 bl_156 br_156 wl_81 vdd gnd cell_6t
Xbit_r82_c156 bl_156 br_156 wl_82 vdd gnd cell_6t
Xbit_r83_c156 bl_156 br_156 wl_83 vdd gnd cell_6t
Xbit_r84_c156 bl_156 br_156 wl_84 vdd gnd cell_6t
Xbit_r85_c156 bl_156 br_156 wl_85 vdd gnd cell_6t
Xbit_r86_c156 bl_156 br_156 wl_86 vdd gnd cell_6t
Xbit_r87_c156 bl_156 br_156 wl_87 vdd gnd cell_6t
Xbit_r88_c156 bl_156 br_156 wl_88 vdd gnd cell_6t
Xbit_r89_c156 bl_156 br_156 wl_89 vdd gnd cell_6t
Xbit_r90_c156 bl_156 br_156 wl_90 vdd gnd cell_6t
Xbit_r91_c156 bl_156 br_156 wl_91 vdd gnd cell_6t
Xbit_r92_c156 bl_156 br_156 wl_92 vdd gnd cell_6t
Xbit_r93_c156 bl_156 br_156 wl_93 vdd gnd cell_6t
Xbit_r94_c156 bl_156 br_156 wl_94 vdd gnd cell_6t
Xbit_r95_c156 bl_156 br_156 wl_95 vdd gnd cell_6t
Xbit_r96_c156 bl_156 br_156 wl_96 vdd gnd cell_6t
Xbit_r97_c156 bl_156 br_156 wl_97 vdd gnd cell_6t
Xbit_r98_c156 bl_156 br_156 wl_98 vdd gnd cell_6t
Xbit_r99_c156 bl_156 br_156 wl_99 vdd gnd cell_6t
Xbit_r100_c156 bl_156 br_156 wl_100 vdd gnd cell_6t
Xbit_r101_c156 bl_156 br_156 wl_101 vdd gnd cell_6t
Xbit_r102_c156 bl_156 br_156 wl_102 vdd gnd cell_6t
Xbit_r103_c156 bl_156 br_156 wl_103 vdd gnd cell_6t
Xbit_r104_c156 bl_156 br_156 wl_104 vdd gnd cell_6t
Xbit_r105_c156 bl_156 br_156 wl_105 vdd gnd cell_6t
Xbit_r106_c156 bl_156 br_156 wl_106 vdd gnd cell_6t
Xbit_r107_c156 bl_156 br_156 wl_107 vdd gnd cell_6t
Xbit_r108_c156 bl_156 br_156 wl_108 vdd gnd cell_6t
Xbit_r109_c156 bl_156 br_156 wl_109 vdd gnd cell_6t
Xbit_r110_c156 bl_156 br_156 wl_110 vdd gnd cell_6t
Xbit_r111_c156 bl_156 br_156 wl_111 vdd gnd cell_6t
Xbit_r112_c156 bl_156 br_156 wl_112 vdd gnd cell_6t
Xbit_r113_c156 bl_156 br_156 wl_113 vdd gnd cell_6t
Xbit_r114_c156 bl_156 br_156 wl_114 vdd gnd cell_6t
Xbit_r115_c156 bl_156 br_156 wl_115 vdd gnd cell_6t
Xbit_r116_c156 bl_156 br_156 wl_116 vdd gnd cell_6t
Xbit_r117_c156 bl_156 br_156 wl_117 vdd gnd cell_6t
Xbit_r118_c156 bl_156 br_156 wl_118 vdd gnd cell_6t
Xbit_r119_c156 bl_156 br_156 wl_119 vdd gnd cell_6t
Xbit_r120_c156 bl_156 br_156 wl_120 vdd gnd cell_6t
Xbit_r121_c156 bl_156 br_156 wl_121 vdd gnd cell_6t
Xbit_r122_c156 bl_156 br_156 wl_122 vdd gnd cell_6t
Xbit_r123_c156 bl_156 br_156 wl_123 vdd gnd cell_6t
Xbit_r124_c156 bl_156 br_156 wl_124 vdd gnd cell_6t
Xbit_r125_c156 bl_156 br_156 wl_125 vdd gnd cell_6t
Xbit_r126_c156 bl_156 br_156 wl_126 vdd gnd cell_6t
Xbit_r127_c156 bl_156 br_156 wl_127 vdd gnd cell_6t
Xbit_r128_c156 bl_156 br_156 wl_128 vdd gnd cell_6t
Xbit_r129_c156 bl_156 br_156 wl_129 vdd gnd cell_6t
Xbit_r130_c156 bl_156 br_156 wl_130 vdd gnd cell_6t
Xbit_r131_c156 bl_156 br_156 wl_131 vdd gnd cell_6t
Xbit_r132_c156 bl_156 br_156 wl_132 vdd gnd cell_6t
Xbit_r133_c156 bl_156 br_156 wl_133 vdd gnd cell_6t
Xbit_r134_c156 bl_156 br_156 wl_134 vdd gnd cell_6t
Xbit_r135_c156 bl_156 br_156 wl_135 vdd gnd cell_6t
Xbit_r136_c156 bl_156 br_156 wl_136 vdd gnd cell_6t
Xbit_r137_c156 bl_156 br_156 wl_137 vdd gnd cell_6t
Xbit_r138_c156 bl_156 br_156 wl_138 vdd gnd cell_6t
Xbit_r139_c156 bl_156 br_156 wl_139 vdd gnd cell_6t
Xbit_r140_c156 bl_156 br_156 wl_140 vdd gnd cell_6t
Xbit_r141_c156 bl_156 br_156 wl_141 vdd gnd cell_6t
Xbit_r142_c156 bl_156 br_156 wl_142 vdd gnd cell_6t
Xbit_r143_c156 bl_156 br_156 wl_143 vdd gnd cell_6t
Xbit_r144_c156 bl_156 br_156 wl_144 vdd gnd cell_6t
Xbit_r145_c156 bl_156 br_156 wl_145 vdd gnd cell_6t
Xbit_r146_c156 bl_156 br_156 wl_146 vdd gnd cell_6t
Xbit_r147_c156 bl_156 br_156 wl_147 vdd gnd cell_6t
Xbit_r148_c156 bl_156 br_156 wl_148 vdd gnd cell_6t
Xbit_r149_c156 bl_156 br_156 wl_149 vdd gnd cell_6t
Xbit_r150_c156 bl_156 br_156 wl_150 vdd gnd cell_6t
Xbit_r151_c156 bl_156 br_156 wl_151 vdd gnd cell_6t
Xbit_r152_c156 bl_156 br_156 wl_152 vdd gnd cell_6t
Xbit_r153_c156 bl_156 br_156 wl_153 vdd gnd cell_6t
Xbit_r154_c156 bl_156 br_156 wl_154 vdd gnd cell_6t
Xbit_r155_c156 bl_156 br_156 wl_155 vdd gnd cell_6t
Xbit_r156_c156 bl_156 br_156 wl_156 vdd gnd cell_6t
Xbit_r157_c156 bl_156 br_156 wl_157 vdd gnd cell_6t
Xbit_r158_c156 bl_156 br_156 wl_158 vdd gnd cell_6t
Xbit_r159_c156 bl_156 br_156 wl_159 vdd gnd cell_6t
Xbit_r160_c156 bl_156 br_156 wl_160 vdd gnd cell_6t
Xbit_r161_c156 bl_156 br_156 wl_161 vdd gnd cell_6t
Xbit_r162_c156 bl_156 br_156 wl_162 vdd gnd cell_6t
Xbit_r163_c156 bl_156 br_156 wl_163 vdd gnd cell_6t
Xbit_r164_c156 bl_156 br_156 wl_164 vdd gnd cell_6t
Xbit_r165_c156 bl_156 br_156 wl_165 vdd gnd cell_6t
Xbit_r166_c156 bl_156 br_156 wl_166 vdd gnd cell_6t
Xbit_r167_c156 bl_156 br_156 wl_167 vdd gnd cell_6t
Xbit_r168_c156 bl_156 br_156 wl_168 vdd gnd cell_6t
Xbit_r169_c156 bl_156 br_156 wl_169 vdd gnd cell_6t
Xbit_r170_c156 bl_156 br_156 wl_170 vdd gnd cell_6t
Xbit_r171_c156 bl_156 br_156 wl_171 vdd gnd cell_6t
Xbit_r172_c156 bl_156 br_156 wl_172 vdd gnd cell_6t
Xbit_r173_c156 bl_156 br_156 wl_173 vdd gnd cell_6t
Xbit_r174_c156 bl_156 br_156 wl_174 vdd gnd cell_6t
Xbit_r175_c156 bl_156 br_156 wl_175 vdd gnd cell_6t
Xbit_r176_c156 bl_156 br_156 wl_176 vdd gnd cell_6t
Xbit_r177_c156 bl_156 br_156 wl_177 vdd gnd cell_6t
Xbit_r178_c156 bl_156 br_156 wl_178 vdd gnd cell_6t
Xbit_r179_c156 bl_156 br_156 wl_179 vdd gnd cell_6t
Xbit_r180_c156 bl_156 br_156 wl_180 vdd gnd cell_6t
Xbit_r181_c156 bl_156 br_156 wl_181 vdd gnd cell_6t
Xbit_r182_c156 bl_156 br_156 wl_182 vdd gnd cell_6t
Xbit_r183_c156 bl_156 br_156 wl_183 vdd gnd cell_6t
Xbit_r184_c156 bl_156 br_156 wl_184 vdd gnd cell_6t
Xbit_r185_c156 bl_156 br_156 wl_185 vdd gnd cell_6t
Xbit_r186_c156 bl_156 br_156 wl_186 vdd gnd cell_6t
Xbit_r187_c156 bl_156 br_156 wl_187 vdd gnd cell_6t
Xbit_r188_c156 bl_156 br_156 wl_188 vdd gnd cell_6t
Xbit_r189_c156 bl_156 br_156 wl_189 vdd gnd cell_6t
Xbit_r190_c156 bl_156 br_156 wl_190 vdd gnd cell_6t
Xbit_r191_c156 bl_156 br_156 wl_191 vdd gnd cell_6t
Xbit_r192_c156 bl_156 br_156 wl_192 vdd gnd cell_6t
Xbit_r193_c156 bl_156 br_156 wl_193 vdd gnd cell_6t
Xbit_r194_c156 bl_156 br_156 wl_194 vdd gnd cell_6t
Xbit_r195_c156 bl_156 br_156 wl_195 vdd gnd cell_6t
Xbit_r196_c156 bl_156 br_156 wl_196 vdd gnd cell_6t
Xbit_r197_c156 bl_156 br_156 wl_197 vdd gnd cell_6t
Xbit_r198_c156 bl_156 br_156 wl_198 vdd gnd cell_6t
Xbit_r199_c156 bl_156 br_156 wl_199 vdd gnd cell_6t
Xbit_r200_c156 bl_156 br_156 wl_200 vdd gnd cell_6t
Xbit_r201_c156 bl_156 br_156 wl_201 vdd gnd cell_6t
Xbit_r202_c156 bl_156 br_156 wl_202 vdd gnd cell_6t
Xbit_r203_c156 bl_156 br_156 wl_203 vdd gnd cell_6t
Xbit_r204_c156 bl_156 br_156 wl_204 vdd gnd cell_6t
Xbit_r205_c156 bl_156 br_156 wl_205 vdd gnd cell_6t
Xbit_r206_c156 bl_156 br_156 wl_206 vdd gnd cell_6t
Xbit_r207_c156 bl_156 br_156 wl_207 vdd gnd cell_6t
Xbit_r208_c156 bl_156 br_156 wl_208 vdd gnd cell_6t
Xbit_r209_c156 bl_156 br_156 wl_209 vdd gnd cell_6t
Xbit_r210_c156 bl_156 br_156 wl_210 vdd gnd cell_6t
Xbit_r211_c156 bl_156 br_156 wl_211 vdd gnd cell_6t
Xbit_r212_c156 bl_156 br_156 wl_212 vdd gnd cell_6t
Xbit_r213_c156 bl_156 br_156 wl_213 vdd gnd cell_6t
Xbit_r214_c156 bl_156 br_156 wl_214 vdd gnd cell_6t
Xbit_r215_c156 bl_156 br_156 wl_215 vdd gnd cell_6t
Xbit_r216_c156 bl_156 br_156 wl_216 vdd gnd cell_6t
Xbit_r217_c156 bl_156 br_156 wl_217 vdd gnd cell_6t
Xbit_r218_c156 bl_156 br_156 wl_218 vdd gnd cell_6t
Xbit_r219_c156 bl_156 br_156 wl_219 vdd gnd cell_6t
Xbit_r220_c156 bl_156 br_156 wl_220 vdd gnd cell_6t
Xbit_r221_c156 bl_156 br_156 wl_221 vdd gnd cell_6t
Xbit_r222_c156 bl_156 br_156 wl_222 vdd gnd cell_6t
Xbit_r223_c156 bl_156 br_156 wl_223 vdd gnd cell_6t
Xbit_r224_c156 bl_156 br_156 wl_224 vdd gnd cell_6t
Xbit_r225_c156 bl_156 br_156 wl_225 vdd gnd cell_6t
Xbit_r226_c156 bl_156 br_156 wl_226 vdd gnd cell_6t
Xbit_r227_c156 bl_156 br_156 wl_227 vdd gnd cell_6t
Xbit_r228_c156 bl_156 br_156 wl_228 vdd gnd cell_6t
Xbit_r229_c156 bl_156 br_156 wl_229 vdd gnd cell_6t
Xbit_r230_c156 bl_156 br_156 wl_230 vdd gnd cell_6t
Xbit_r231_c156 bl_156 br_156 wl_231 vdd gnd cell_6t
Xbit_r232_c156 bl_156 br_156 wl_232 vdd gnd cell_6t
Xbit_r233_c156 bl_156 br_156 wl_233 vdd gnd cell_6t
Xbit_r234_c156 bl_156 br_156 wl_234 vdd gnd cell_6t
Xbit_r235_c156 bl_156 br_156 wl_235 vdd gnd cell_6t
Xbit_r236_c156 bl_156 br_156 wl_236 vdd gnd cell_6t
Xbit_r237_c156 bl_156 br_156 wl_237 vdd gnd cell_6t
Xbit_r238_c156 bl_156 br_156 wl_238 vdd gnd cell_6t
Xbit_r239_c156 bl_156 br_156 wl_239 vdd gnd cell_6t
Xbit_r240_c156 bl_156 br_156 wl_240 vdd gnd cell_6t
Xbit_r241_c156 bl_156 br_156 wl_241 vdd gnd cell_6t
Xbit_r242_c156 bl_156 br_156 wl_242 vdd gnd cell_6t
Xbit_r243_c156 bl_156 br_156 wl_243 vdd gnd cell_6t
Xbit_r244_c156 bl_156 br_156 wl_244 vdd gnd cell_6t
Xbit_r245_c156 bl_156 br_156 wl_245 vdd gnd cell_6t
Xbit_r246_c156 bl_156 br_156 wl_246 vdd gnd cell_6t
Xbit_r247_c156 bl_156 br_156 wl_247 vdd gnd cell_6t
Xbit_r248_c156 bl_156 br_156 wl_248 vdd gnd cell_6t
Xbit_r249_c156 bl_156 br_156 wl_249 vdd gnd cell_6t
Xbit_r250_c156 bl_156 br_156 wl_250 vdd gnd cell_6t
Xbit_r251_c156 bl_156 br_156 wl_251 vdd gnd cell_6t
Xbit_r252_c156 bl_156 br_156 wl_252 vdd gnd cell_6t
Xbit_r253_c156 bl_156 br_156 wl_253 vdd gnd cell_6t
Xbit_r254_c156 bl_156 br_156 wl_254 vdd gnd cell_6t
Xbit_r255_c156 bl_156 br_156 wl_255 vdd gnd cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd cell_6t
Xbit_r1_c157 bl_157 br_157 wl_1 vdd gnd cell_6t
Xbit_r2_c157 bl_157 br_157 wl_2 vdd gnd cell_6t
Xbit_r3_c157 bl_157 br_157 wl_3 vdd gnd cell_6t
Xbit_r4_c157 bl_157 br_157 wl_4 vdd gnd cell_6t
Xbit_r5_c157 bl_157 br_157 wl_5 vdd gnd cell_6t
Xbit_r6_c157 bl_157 br_157 wl_6 vdd gnd cell_6t
Xbit_r7_c157 bl_157 br_157 wl_7 vdd gnd cell_6t
Xbit_r8_c157 bl_157 br_157 wl_8 vdd gnd cell_6t
Xbit_r9_c157 bl_157 br_157 wl_9 vdd gnd cell_6t
Xbit_r10_c157 bl_157 br_157 wl_10 vdd gnd cell_6t
Xbit_r11_c157 bl_157 br_157 wl_11 vdd gnd cell_6t
Xbit_r12_c157 bl_157 br_157 wl_12 vdd gnd cell_6t
Xbit_r13_c157 bl_157 br_157 wl_13 vdd gnd cell_6t
Xbit_r14_c157 bl_157 br_157 wl_14 vdd gnd cell_6t
Xbit_r15_c157 bl_157 br_157 wl_15 vdd gnd cell_6t
Xbit_r16_c157 bl_157 br_157 wl_16 vdd gnd cell_6t
Xbit_r17_c157 bl_157 br_157 wl_17 vdd gnd cell_6t
Xbit_r18_c157 bl_157 br_157 wl_18 vdd gnd cell_6t
Xbit_r19_c157 bl_157 br_157 wl_19 vdd gnd cell_6t
Xbit_r20_c157 bl_157 br_157 wl_20 vdd gnd cell_6t
Xbit_r21_c157 bl_157 br_157 wl_21 vdd gnd cell_6t
Xbit_r22_c157 bl_157 br_157 wl_22 vdd gnd cell_6t
Xbit_r23_c157 bl_157 br_157 wl_23 vdd gnd cell_6t
Xbit_r24_c157 bl_157 br_157 wl_24 vdd gnd cell_6t
Xbit_r25_c157 bl_157 br_157 wl_25 vdd gnd cell_6t
Xbit_r26_c157 bl_157 br_157 wl_26 vdd gnd cell_6t
Xbit_r27_c157 bl_157 br_157 wl_27 vdd gnd cell_6t
Xbit_r28_c157 bl_157 br_157 wl_28 vdd gnd cell_6t
Xbit_r29_c157 bl_157 br_157 wl_29 vdd gnd cell_6t
Xbit_r30_c157 bl_157 br_157 wl_30 vdd gnd cell_6t
Xbit_r31_c157 bl_157 br_157 wl_31 vdd gnd cell_6t
Xbit_r32_c157 bl_157 br_157 wl_32 vdd gnd cell_6t
Xbit_r33_c157 bl_157 br_157 wl_33 vdd gnd cell_6t
Xbit_r34_c157 bl_157 br_157 wl_34 vdd gnd cell_6t
Xbit_r35_c157 bl_157 br_157 wl_35 vdd gnd cell_6t
Xbit_r36_c157 bl_157 br_157 wl_36 vdd gnd cell_6t
Xbit_r37_c157 bl_157 br_157 wl_37 vdd gnd cell_6t
Xbit_r38_c157 bl_157 br_157 wl_38 vdd gnd cell_6t
Xbit_r39_c157 bl_157 br_157 wl_39 vdd gnd cell_6t
Xbit_r40_c157 bl_157 br_157 wl_40 vdd gnd cell_6t
Xbit_r41_c157 bl_157 br_157 wl_41 vdd gnd cell_6t
Xbit_r42_c157 bl_157 br_157 wl_42 vdd gnd cell_6t
Xbit_r43_c157 bl_157 br_157 wl_43 vdd gnd cell_6t
Xbit_r44_c157 bl_157 br_157 wl_44 vdd gnd cell_6t
Xbit_r45_c157 bl_157 br_157 wl_45 vdd gnd cell_6t
Xbit_r46_c157 bl_157 br_157 wl_46 vdd gnd cell_6t
Xbit_r47_c157 bl_157 br_157 wl_47 vdd gnd cell_6t
Xbit_r48_c157 bl_157 br_157 wl_48 vdd gnd cell_6t
Xbit_r49_c157 bl_157 br_157 wl_49 vdd gnd cell_6t
Xbit_r50_c157 bl_157 br_157 wl_50 vdd gnd cell_6t
Xbit_r51_c157 bl_157 br_157 wl_51 vdd gnd cell_6t
Xbit_r52_c157 bl_157 br_157 wl_52 vdd gnd cell_6t
Xbit_r53_c157 bl_157 br_157 wl_53 vdd gnd cell_6t
Xbit_r54_c157 bl_157 br_157 wl_54 vdd gnd cell_6t
Xbit_r55_c157 bl_157 br_157 wl_55 vdd gnd cell_6t
Xbit_r56_c157 bl_157 br_157 wl_56 vdd gnd cell_6t
Xbit_r57_c157 bl_157 br_157 wl_57 vdd gnd cell_6t
Xbit_r58_c157 bl_157 br_157 wl_58 vdd gnd cell_6t
Xbit_r59_c157 bl_157 br_157 wl_59 vdd gnd cell_6t
Xbit_r60_c157 bl_157 br_157 wl_60 vdd gnd cell_6t
Xbit_r61_c157 bl_157 br_157 wl_61 vdd gnd cell_6t
Xbit_r62_c157 bl_157 br_157 wl_62 vdd gnd cell_6t
Xbit_r63_c157 bl_157 br_157 wl_63 vdd gnd cell_6t
Xbit_r64_c157 bl_157 br_157 wl_64 vdd gnd cell_6t
Xbit_r65_c157 bl_157 br_157 wl_65 vdd gnd cell_6t
Xbit_r66_c157 bl_157 br_157 wl_66 vdd gnd cell_6t
Xbit_r67_c157 bl_157 br_157 wl_67 vdd gnd cell_6t
Xbit_r68_c157 bl_157 br_157 wl_68 vdd gnd cell_6t
Xbit_r69_c157 bl_157 br_157 wl_69 vdd gnd cell_6t
Xbit_r70_c157 bl_157 br_157 wl_70 vdd gnd cell_6t
Xbit_r71_c157 bl_157 br_157 wl_71 vdd gnd cell_6t
Xbit_r72_c157 bl_157 br_157 wl_72 vdd gnd cell_6t
Xbit_r73_c157 bl_157 br_157 wl_73 vdd gnd cell_6t
Xbit_r74_c157 bl_157 br_157 wl_74 vdd gnd cell_6t
Xbit_r75_c157 bl_157 br_157 wl_75 vdd gnd cell_6t
Xbit_r76_c157 bl_157 br_157 wl_76 vdd gnd cell_6t
Xbit_r77_c157 bl_157 br_157 wl_77 vdd gnd cell_6t
Xbit_r78_c157 bl_157 br_157 wl_78 vdd gnd cell_6t
Xbit_r79_c157 bl_157 br_157 wl_79 vdd gnd cell_6t
Xbit_r80_c157 bl_157 br_157 wl_80 vdd gnd cell_6t
Xbit_r81_c157 bl_157 br_157 wl_81 vdd gnd cell_6t
Xbit_r82_c157 bl_157 br_157 wl_82 vdd gnd cell_6t
Xbit_r83_c157 bl_157 br_157 wl_83 vdd gnd cell_6t
Xbit_r84_c157 bl_157 br_157 wl_84 vdd gnd cell_6t
Xbit_r85_c157 bl_157 br_157 wl_85 vdd gnd cell_6t
Xbit_r86_c157 bl_157 br_157 wl_86 vdd gnd cell_6t
Xbit_r87_c157 bl_157 br_157 wl_87 vdd gnd cell_6t
Xbit_r88_c157 bl_157 br_157 wl_88 vdd gnd cell_6t
Xbit_r89_c157 bl_157 br_157 wl_89 vdd gnd cell_6t
Xbit_r90_c157 bl_157 br_157 wl_90 vdd gnd cell_6t
Xbit_r91_c157 bl_157 br_157 wl_91 vdd gnd cell_6t
Xbit_r92_c157 bl_157 br_157 wl_92 vdd gnd cell_6t
Xbit_r93_c157 bl_157 br_157 wl_93 vdd gnd cell_6t
Xbit_r94_c157 bl_157 br_157 wl_94 vdd gnd cell_6t
Xbit_r95_c157 bl_157 br_157 wl_95 vdd gnd cell_6t
Xbit_r96_c157 bl_157 br_157 wl_96 vdd gnd cell_6t
Xbit_r97_c157 bl_157 br_157 wl_97 vdd gnd cell_6t
Xbit_r98_c157 bl_157 br_157 wl_98 vdd gnd cell_6t
Xbit_r99_c157 bl_157 br_157 wl_99 vdd gnd cell_6t
Xbit_r100_c157 bl_157 br_157 wl_100 vdd gnd cell_6t
Xbit_r101_c157 bl_157 br_157 wl_101 vdd gnd cell_6t
Xbit_r102_c157 bl_157 br_157 wl_102 vdd gnd cell_6t
Xbit_r103_c157 bl_157 br_157 wl_103 vdd gnd cell_6t
Xbit_r104_c157 bl_157 br_157 wl_104 vdd gnd cell_6t
Xbit_r105_c157 bl_157 br_157 wl_105 vdd gnd cell_6t
Xbit_r106_c157 bl_157 br_157 wl_106 vdd gnd cell_6t
Xbit_r107_c157 bl_157 br_157 wl_107 vdd gnd cell_6t
Xbit_r108_c157 bl_157 br_157 wl_108 vdd gnd cell_6t
Xbit_r109_c157 bl_157 br_157 wl_109 vdd gnd cell_6t
Xbit_r110_c157 bl_157 br_157 wl_110 vdd gnd cell_6t
Xbit_r111_c157 bl_157 br_157 wl_111 vdd gnd cell_6t
Xbit_r112_c157 bl_157 br_157 wl_112 vdd gnd cell_6t
Xbit_r113_c157 bl_157 br_157 wl_113 vdd gnd cell_6t
Xbit_r114_c157 bl_157 br_157 wl_114 vdd gnd cell_6t
Xbit_r115_c157 bl_157 br_157 wl_115 vdd gnd cell_6t
Xbit_r116_c157 bl_157 br_157 wl_116 vdd gnd cell_6t
Xbit_r117_c157 bl_157 br_157 wl_117 vdd gnd cell_6t
Xbit_r118_c157 bl_157 br_157 wl_118 vdd gnd cell_6t
Xbit_r119_c157 bl_157 br_157 wl_119 vdd gnd cell_6t
Xbit_r120_c157 bl_157 br_157 wl_120 vdd gnd cell_6t
Xbit_r121_c157 bl_157 br_157 wl_121 vdd gnd cell_6t
Xbit_r122_c157 bl_157 br_157 wl_122 vdd gnd cell_6t
Xbit_r123_c157 bl_157 br_157 wl_123 vdd gnd cell_6t
Xbit_r124_c157 bl_157 br_157 wl_124 vdd gnd cell_6t
Xbit_r125_c157 bl_157 br_157 wl_125 vdd gnd cell_6t
Xbit_r126_c157 bl_157 br_157 wl_126 vdd gnd cell_6t
Xbit_r127_c157 bl_157 br_157 wl_127 vdd gnd cell_6t
Xbit_r128_c157 bl_157 br_157 wl_128 vdd gnd cell_6t
Xbit_r129_c157 bl_157 br_157 wl_129 vdd gnd cell_6t
Xbit_r130_c157 bl_157 br_157 wl_130 vdd gnd cell_6t
Xbit_r131_c157 bl_157 br_157 wl_131 vdd gnd cell_6t
Xbit_r132_c157 bl_157 br_157 wl_132 vdd gnd cell_6t
Xbit_r133_c157 bl_157 br_157 wl_133 vdd gnd cell_6t
Xbit_r134_c157 bl_157 br_157 wl_134 vdd gnd cell_6t
Xbit_r135_c157 bl_157 br_157 wl_135 vdd gnd cell_6t
Xbit_r136_c157 bl_157 br_157 wl_136 vdd gnd cell_6t
Xbit_r137_c157 bl_157 br_157 wl_137 vdd gnd cell_6t
Xbit_r138_c157 bl_157 br_157 wl_138 vdd gnd cell_6t
Xbit_r139_c157 bl_157 br_157 wl_139 vdd gnd cell_6t
Xbit_r140_c157 bl_157 br_157 wl_140 vdd gnd cell_6t
Xbit_r141_c157 bl_157 br_157 wl_141 vdd gnd cell_6t
Xbit_r142_c157 bl_157 br_157 wl_142 vdd gnd cell_6t
Xbit_r143_c157 bl_157 br_157 wl_143 vdd gnd cell_6t
Xbit_r144_c157 bl_157 br_157 wl_144 vdd gnd cell_6t
Xbit_r145_c157 bl_157 br_157 wl_145 vdd gnd cell_6t
Xbit_r146_c157 bl_157 br_157 wl_146 vdd gnd cell_6t
Xbit_r147_c157 bl_157 br_157 wl_147 vdd gnd cell_6t
Xbit_r148_c157 bl_157 br_157 wl_148 vdd gnd cell_6t
Xbit_r149_c157 bl_157 br_157 wl_149 vdd gnd cell_6t
Xbit_r150_c157 bl_157 br_157 wl_150 vdd gnd cell_6t
Xbit_r151_c157 bl_157 br_157 wl_151 vdd gnd cell_6t
Xbit_r152_c157 bl_157 br_157 wl_152 vdd gnd cell_6t
Xbit_r153_c157 bl_157 br_157 wl_153 vdd gnd cell_6t
Xbit_r154_c157 bl_157 br_157 wl_154 vdd gnd cell_6t
Xbit_r155_c157 bl_157 br_157 wl_155 vdd gnd cell_6t
Xbit_r156_c157 bl_157 br_157 wl_156 vdd gnd cell_6t
Xbit_r157_c157 bl_157 br_157 wl_157 vdd gnd cell_6t
Xbit_r158_c157 bl_157 br_157 wl_158 vdd gnd cell_6t
Xbit_r159_c157 bl_157 br_157 wl_159 vdd gnd cell_6t
Xbit_r160_c157 bl_157 br_157 wl_160 vdd gnd cell_6t
Xbit_r161_c157 bl_157 br_157 wl_161 vdd gnd cell_6t
Xbit_r162_c157 bl_157 br_157 wl_162 vdd gnd cell_6t
Xbit_r163_c157 bl_157 br_157 wl_163 vdd gnd cell_6t
Xbit_r164_c157 bl_157 br_157 wl_164 vdd gnd cell_6t
Xbit_r165_c157 bl_157 br_157 wl_165 vdd gnd cell_6t
Xbit_r166_c157 bl_157 br_157 wl_166 vdd gnd cell_6t
Xbit_r167_c157 bl_157 br_157 wl_167 vdd gnd cell_6t
Xbit_r168_c157 bl_157 br_157 wl_168 vdd gnd cell_6t
Xbit_r169_c157 bl_157 br_157 wl_169 vdd gnd cell_6t
Xbit_r170_c157 bl_157 br_157 wl_170 vdd gnd cell_6t
Xbit_r171_c157 bl_157 br_157 wl_171 vdd gnd cell_6t
Xbit_r172_c157 bl_157 br_157 wl_172 vdd gnd cell_6t
Xbit_r173_c157 bl_157 br_157 wl_173 vdd gnd cell_6t
Xbit_r174_c157 bl_157 br_157 wl_174 vdd gnd cell_6t
Xbit_r175_c157 bl_157 br_157 wl_175 vdd gnd cell_6t
Xbit_r176_c157 bl_157 br_157 wl_176 vdd gnd cell_6t
Xbit_r177_c157 bl_157 br_157 wl_177 vdd gnd cell_6t
Xbit_r178_c157 bl_157 br_157 wl_178 vdd gnd cell_6t
Xbit_r179_c157 bl_157 br_157 wl_179 vdd gnd cell_6t
Xbit_r180_c157 bl_157 br_157 wl_180 vdd gnd cell_6t
Xbit_r181_c157 bl_157 br_157 wl_181 vdd gnd cell_6t
Xbit_r182_c157 bl_157 br_157 wl_182 vdd gnd cell_6t
Xbit_r183_c157 bl_157 br_157 wl_183 vdd gnd cell_6t
Xbit_r184_c157 bl_157 br_157 wl_184 vdd gnd cell_6t
Xbit_r185_c157 bl_157 br_157 wl_185 vdd gnd cell_6t
Xbit_r186_c157 bl_157 br_157 wl_186 vdd gnd cell_6t
Xbit_r187_c157 bl_157 br_157 wl_187 vdd gnd cell_6t
Xbit_r188_c157 bl_157 br_157 wl_188 vdd gnd cell_6t
Xbit_r189_c157 bl_157 br_157 wl_189 vdd gnd cell_6t
Xbit_r190_c157 bl_157 br_157 wl_190 vdd gnd cell_6t
Xbit_r191_c157 bl_157 br_157 wl_191 vdd gnd cell_6t
Xbit_r192_c157 bl_157 br_157 wl_192 vdd gnd cell_6t
Xbit_r193_c157 bl_157 br_157 wl_193 vdd gnd cell_6t
Xbit_r194_c157 bl_157 br_157 wl_194 vdd gnd cell_6t
Xbit_r195_c157 bl_157 br_157 wl_195 vdd gnd cell_6t
Xbit_r196_c157 bl_157 br_157 wl_196 vdd gnd cell_6t
Xbit_r197_c157 bl_157 br_157 wl_197 vdd gnd cell_6t
Xbit_r198_c157 bl_157 br_157 wl_198 vdd gnd cell_6t
Xbit_r199_c157 bl_157 br_157 wl_199 vdd gnd cell_6t
Xbit_r200_c157 bl_157 br_157 wl_200 vdd gnd cell_6t
Xbit_r201_c157 bl_157 br_157 wl_201 vdd gnd cell_6t
Xbit_r202_c157 bl_157 br_157 wl_202 vdd gnd cell_6t
Xbit_r203_c157 bl_157 br_157 wl_203 vdd gnd cell_6t
Xbit_r204_c157 bl_157 br_157 wl_204 vdd gnd cell_6t
Xbit_r205_c157 bl_157 br_157 wl_205 vdd gnd cell_6t
Xbit_r206_c157 bl_157 br_157 wl_206 vdd gnd cell_6t
Xbit_r207_c157 bl_157 br_157 wl_207 vdd gnd cell_6t
Xbit_r208_c157 bl_157 br_157 wl_208 vdd gnd cell_6t
Xbit_r209_c157 bl_157 br_157 wl_209 vdd gnd cell_6t
Xbit_r210_c157 bl_157 br_157 wl_210 vdd gnd cell_6t
Xbit_r211_c157 bl_157 br_157 wl_211 vdd gnd cell_6t
Xbit_r212_c157 bl_157 br_157 wl_212 vdd gnd cell_6t
Xbit_r213_c157 bl_157 br_157 wl_213 vdd gnd cell_6t
Xbit_r214_c157 bl_157 br_157 wl_214 vdd gnd cell_6t
Xbit_r215_c157 bl_157 br_157 wl_215 vdd gnd cell_6t
Xbit_r216_c157 bl_157 br_157 wl_216 vdd gnd cell_6t
Xbit_r217_c157 bl_157 br_157 wl_217 vdd gnd cell_6t
Xbit_r218_c157 bl_157 br_157 wl_218 vdd gnd cell_6t
Xbit_r219_c157 bl_157 br_157 wl_219 vdd gnd cell_6t
Xbit_r220_c157 bl_157 br_157 wl_220 vdd gnd cell_6t
Xbit_r221_c157 bl_157 br_157 wl_221 vdd gnd cell_6t
Xbit_r222_c157 bl_157 br_157 wl_222 vdd gnd cell_6t
Xbit_r223_c157 bl_157 br_157 wl_223 vdd gnd cell_6t
Xbit_r224_c157 bl_157 br_157 wl_224 vdd gnd cell_6t
Xbit_r225_c157 bl_157 br_157 wl_225 vdd gnd cell_6t
Xbit_r226_c157 bl_157 br_157 wl_226 vdd gnd cell_6t
Xbit_r227_c157 bl_157 br_157 wl_227 vdd gnd cell_6t
Xbit_r228_c157 bl_157 br_157 wl_228 vdd gnd cell_6t
Xbit_r229_c157 bl_157 br_157 wl_229 vdd gnd cell_6t
Xbit_r230_c157 bl_157 br_157 wl_230 vdd gnd cell_6t
Xbit_r231_c157 bl_157 br_157 wl_231 vdd gnd cell_6t
Xbit_r232_c157 bl_157 br_157 wl_232 vdd gnd cell_6t
Xbit_r233_c157 bl_157 br_157 wl_233 vdd gnd cell_6t
Xbit_r234_c157 bl_157 br_157 wl_234 vdd gnd cell_6t
Xbit_r235_c157 bl_157 br_157 wl_235 vdd gnd cell_6t
Xbit_r236_c157 bl_157 br_157 wl_236 vdd gnd cell_6t
Xbit_r237_c157 bl_157 br_157 wl_237 vdd gnd cell_6t
Xbit_r238_c157 bl_157 br_157 wl_238 vdd gnd cell_6t
Xbit_r239_c157 bl_157 br_157 wl_239 vdd gnd cell_6t
Xbit_r240_c157 bl_157 br_157 wl_240 vdd gnd cell_6t
Xbit_r241_c157 bl_157 br_157 wl_241 vdd gnd cell_6t
Xbit_r242_c157 bl_157 br_157 wl_242 vdd gnd cell_6t
Xbit_r243_c157 bl_157 br_157 wl_243 vdd gnd cell_6t
Xbit_r244_c157 bl_157 br_157 wl_244 vdd gnd cell_6t
Xbit_r245_c157 bl_157 br_157 wl_245 vdd gnd cell_6t
Xbit_r246_c157 bl_157 br_157 wl_246 vdd gnd cell_6t
Xbit_r247_c157 bl_157 br_157 wl_247 vdd gnd cell_6t
Xbit_r248_c157 bl_157 br_157 wl_248 vdd gnd cell_6t
Xbit_r249_c157 bl_157 br_157 wl_249 vdd gnd cell_6t
Xbit_r250_c157 bl_157 br_157 wl_250 vdd gnd cell_6t
Xbit_r251_c157 bl_157 br_157 wl_251 vdd gnd cell_6t
Xbit_r252_c157 bl_157 br_157 wl_252 vdd gnd cell_6t
Xbit_r253_c157 bl_157 br_157 wl_253 vdd gnd cell_6t
Xbit_r254_c157 bl_157 br_157 wl_254 vdd gnd cell_6t
Xbit_r255_c157 bl_157 br_157 wl_255 vdd gnd cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd cell_6t
Xbit_r1_c158 bl_158 br_158 wl_1 vdd gnd cell_6t
Xbit_r2_c158 bl_158 br_158 wl_2 vdd gnd cell_6t
Xbit_r3_c158 bl_158 br_158 wl_3 vdd gnd cell_6t
Xbit_r4_c158 bl_158 br_158 wl_4 vdd gnd cell_6t
Xbit_r5_c158 bl_158 br_158 wl_5 vdd gnd cell_6t
Xbit_r6_c158 bl_158 br_158 wl_6 vdd gnd cell_6t
Xbit_r7_c158 bl_158 br_158 wl_7 vdd gnd cell_6t
Xbit_r8_c158 bl_158 br_158 wl_8 vdd gnd cell_6t
Xbit_r9_c158 bl_158 br_158 wl_9 vdd gnd cell_6t
Xbit_r10_c158 bl_158 br_158 wl_10 vdd gnd cell_6t
Xbit_r11_c158 bl_158 br_158 wl_11 vdd gnd cell_6t
Xbit_r12_c158 bl_158 br_158 wl_12 vdd gnd cell_6t
Xbit_r13_c158 bl_158 br_158 wl_13 vdd gnd cell_6t
Xbit_r14_c158 bl_158 br_158 wl_14 vdd gnd cell_6t
Xbit_r15_c158 bl_158 br_158 wl_15 vdd gnd cell_6t
Xbit_r16_c158 bl_158 br_158 wl_16 vdd gnd cell_6t
Xbit_r17_c158 bl_158 br_158 wl_17 vdd gnd cell_6t
Xbit_r18_c158 bl_158 br_158 wl_18 vdd gnd cell_6t
Xbit_r19_c158 bl_158 br_158 wl_19 vdd gnd cell_6t
Xbit_r20_c158 bl_158 br_158 wl_20 vdd gnd cell_6t
Xbit_r21_c158 bl_158 br_158 wl_21 vdd gnd cell_6t
Xbit_r22_c158 bl_158 br_158 wl_22 vdd gnd cell_6t
Xbit_r23_c158 bl_158 br_158 wl_23 vdd gnd cell_6t
Xbit_r24_c158 bl_158 br_158 wl_24 vdd gnd cell_6t
Xbit_r25_c158 bl_158 br_158 wl_25 vdd gnd cell_6t
Xbit_r26_c158 bl_158 br_158 wl_26 vdd gnd cell_6t
Xbit_r27_c158 bl_158 br_158 wl_27 vdd gnd cell_6t
Xbit_r28_c158 bl_158 br_158 wl_28 vdd gnd cell_6t
Xbit_r29_c158 bl_158 br_158 wl_29 vdd gnd cell_6t
Xbit_r30_c158 bl_158 br_158 wl_30 vdd gnd cell_6t
Xbit_r31_c158 bl_158 br_158 wl_31 vdd gnd cell_6t
Xbit_r32_c158 bl_158 br_158 wl_32 vdd gnd cell_6t
Xbit_r33_c158 bl_158 br_158 wl_33 vdd gnd cell_6t
Xbit_r34_c158 bl_158 br_158 wl_34 vdd gnd cell_6t
Xbit_r35_c158 bl_158 br_158 wl_35 vdd gnd cell_6t
Xbit_r36_c158 bl_158 br_158 wl_36 vdd gnd cell_6t
Xbit_r37_c158 bl_158 br_158 wl_37 vdd gnd cell_6t
Xbit_r38_c158 bl_158 br_158 wl_38 vdd gnd cell_6t
Xbit_r39_c158 bl_158 br_158 wl_39 vdd gnd cell_6t
Xbit_r40_c158 bl_158 br_158 wl_40 vdd gnd cell_6t
Xbit_r41_c158 bl_158 br_158 wl_41 vdd gnd cell_6t
Xbit_r42_c158 bl_158 br_158 wl_42 vdd gnd cell_6t
Xbit_r43_c158 bl_158 br_158 wl_43 vdd gnd cell_6t
Xbit_r44_c158 bl_158 br_158 wl_44 vdd gnd cell_6t
Xbit_r45_c158 bl_158 br_158 wl_45 vdd gnd cell_6t
Xbit_r46_c158 bl_158 br_158 wl_46 vdd gnd cell_6t
Xbit_r47_c158 bl_158 br_158 wl_47 vdd gnd cell_6t
Xbit_r48_c158 bl_158 br_158 wl_48 vdd gnd cell_6t
Xbit_r49_c158 bl_158 br_158 wl_49 vdd gnd cell_6t
Xbit_r50_c158 bl_158 br_158 wl_50 vdd gnd cell_6t
Xbit_r51_c158 bl_158 br_158 wl_51 vdd gnd cell_6t
Xbit_r52_c158 bl_158 br_158 wl_52 vdd gnd cell_6t
Xbit_r53_c158 bl_158 br_158 wl_53 vdd gnd cell_6t
Xbit_r54_c158 bl_158 br_158 wl_54 vdd gnd cell_6t
Xbit_r55_c158 bl_158 br_158 wl_55 vdd gnd cell_6t
Xbit_r56_c158 bl_158 br_158 wl_56 vdd gnd cell_6t
Xbit_r57_c158 bl_158 br_158 wl_57 vdd gnd cell_6t
Xbit_r58_c158 bl_158 br_158 wl_58 vdd gnd cell_6t
Xbit_r59_c158 bl_158 br_158 wl_59 vdd gnd cell_6t
Xbit_r60_c158 bl_158 br_158 wl_60 vdd gnd cell_6t
Xbit_r61_c158 bl_158 br_158 wl_61 vdd gnd cell_6t
Xbit_r62_c158 bl_158 br_158 wl_62 vdd gnd cell_6t
Xbit_r63_c158 bl_158 br_158 wl_63 vdd gnd cell_6t
Xbit_r64_c158 bl_158 br_158 wl_64 vdd gnd cell_6t
Xbit_r65_c158 bl_158 br_158 wl_65 vdd gnd cell_6t
Xbit_r66_c158 bl_158 br_158 wl_66 vdd gnd cell_6t
Xbit_r67_c158 bl_158 br_158 wl_67 vdd gnd cell_6t
Xbit_r68_c158 bl_158 br_158 wl_68 vdd gnd cell_6t
Xbit_r69_c158 bl_158 br_158 wl_69 vdd gnd cell_6t
Xbit_r70_c158 bl_158 br_158 wl_70 vdd gnd cell_6t
Xbit_r71_c158 bl_158 br_158 wl_71 vdd gnd cell_6t
Xbit_r72_c158 bl_158 br_158 wl_72 vdd gnd cell_6t
Xbit_r73_c158 bl_158 br_158 wl_73 vdd gnd cell_6t
Xbit_r74_c158 bl_158 br_158 wl_74 vdd gnd cell_6t
Xbit_r75_c158 bl_158 br_158 wl_75 vdd gnd cell_6t
Xbit_r76_c158 bl_158 br_158 wl_76 vdd gnd cell_6t
Xbit_r77_c158 bl_158 br_158 wl_77 vdd gnd cell_6t
Xbit_r78_c158 bl_158 br_158 wl_78 vdd gnd cell_6t
Xbit_r79_c158 bl_158 br_158 wl_79 vdd gnd cell_6t
Xbit_r80_c158 bl_158 br_158 wl_80 vdd gnd cell_6t
Xbit_r81_c158 bl_158 br_158 wl_81 vdd gnd cell_6t
Xbit_r82_c158 bl_158 br_158 wl_82 vdd gnd cell_6t
Xbit_r83_c158 bl_158 br_158 wl_83 vdd gnd cell_6t
Xbit_r84_c158 bl_158 br_158 wl_84 vdd gnd cell_6t
Xbit_r85_c158 bl_158 br_158 wl_85 vdd gnd cell_6t
Xbit_r86_c158 bl_158 br_158 wl_86 vdd gnd cell_6t
Xbit_r87_c158 bl_158 br_158 wl_87 vdd gnd cell_6t
Xbit_r88_c158 bl_158 br_158 wl_88 vdd gnd cell_6t
Xbit_r89_c158 bl_158 br_158 wl_89 vdd gnd cell_6t
Xbit_r90_c158 bl_158 br_158 wl_90 vdd gnd cell_6t
Xbit_r91_c158 bl_158 br_158 wl_91 vdd gnd cell_6t
Xbit_r92_c158 bl_158 br_158 wl_92 vdd gnd cell_6t
Xbit_r93_c158 bl_158 br_158 wl_93 vdd gnd cell_6t
Xbit_r94_c158 bl_158 br_158 wl_94 vdd gnd cell_6t
Xbit_r95_c158 bl_158 br_158 wl_95 vdd gnd cell_6t
Xbit_r96_c158 bl_158 br_158 wl_96 vdd gnd cell_6t
Xbit_r97_c158 bl_158 br_158 wl_97 vdd gnd cell_6t
Xbit_r98_c158 bl_158 br_158 wl_98 vdd gnd cell_6t
Xbit_r99_c158 bl_158 br_158 wl_99 vdd gnd cell_6t
Xbit_r100_c158 bl_158 br_158 wl_100 vdd gnd cell_6t
Xbit_r101_c158 bl_158 br_158 wl_101 vdd gnd cell_6t
Xbit_r102_c158 bl_158 br_158 wl_102 vdd gnd cell_6t
Xbit_r103_c158 bl_158 br_158 wl_103 vdd gnd cell_6t
Xbit_r104_c158 bl_158 br_158 wl_104 vdd gnd cell_6t
Xbit_r105_c158 bl_158 br_158 wl_105 vdd gnd cell_6t
Xbit_r106_c158 bl_158 br_158 wl_106 vdd gnd cell_6t
Xbit_r107_c158 bl_158 br_158 wl_107 vdd gnd cell_6t
Xbit_r108_c158 bl_158 br_158 wl_108 vdd gnd cell_6t
Xbit_r109_c158 bl_158 br_158 wl_109 vdd gnd cell_6t
Xbit_r110_c158 bl_158 br_158 wl_110 vdd gnd cell_6t
Xbit_r111_c158 bl_158 br_158 wl_111 vdd gnd cell_6t
Xbit_r112_c158 bl_158 br_158 wl_112 vdd gnd cell_6t
Xbit_r113_c158 bl_158 br_158 wl_113 vdd gnd cell_6t
Xbit_r114_c158 bl_158 br_158 wl_114 vdd gnd cell_6t
Xbit_r115_c158 bl_158 br_158 wl_115 vdd gnd cell_6t
Xbit_r116_c158 bl_158 br_158 wl_116 vdd gnd cell_6t
Xbit_r117_c158 bl_158 br_158 wl_117 vdd gnd cell_6t
Xbit_r118_c158 bl_158 br_158 wl_118 vdd gnd cell_6t
Xbit_r119_c158 bl_158 br_158 wl_119 vdd gnd cell_6t
Xbit_r120_c158 bl_158 br_158 wl_120 vdd gnd cell_6t
Xbit_r121_c158 bl_158 br_158 wl_121 vdd gnd cell_6t
Xbit_r122_c158 bl_158 br_158 wl_122 vdd gnd cell_6t
Xbit_r123_c158 bl_158 br_158 wl_123 vdd gnd cell_6t
Xbit_r124_c158 bl_158 br_158 wl_124 vdd gnd cell_6t
Xbit_r125_c158 bl_158 br_158 wl_125 vdd gnd cell_6t
Xbit_r126_c158 bl_158 br_158 wl_126 vdd gnd cell_6t
Xbit_r127_c158 bl_158 br_158 wl_127 vdd gnd cell_6t
Xbit_r128_c158 bl_158 br_158 wl_128 vdd gnd cell_6t
Xbit_r129_c158 bl_158 br_158 wl_129 vdd gnd cell_6t
Xbit_r130_c158 bl_158 br_158 wl_130 vdd gnd cell_6t
Xbit_r131_c158 bl_158 br_158 wl_131 vdd gnd cell_6t
Xbit_r132_c158 bl_158 br_158 wl_132 vdd gnd cell_6t
Xbit_r133_c158 bl_158 br_158 wl_133 vdd gnd cell_6t
Xbit_r134_c158 bl_158 br_158 wl_134 vdd gnd cell_6t
Xbit_r135_c158 bl_158 br_158 wl_135 vdd gnd cell_6t
Xbit_r136_c158 bl_158 br_158 wl_136 vdd gnd cell_6t
Xbit_r137_c158 bl_158 br_158 wl_137 vdd gnd cell_6t
Xbit_r138_c158 bl_158 br_158 wl_138 vdd gnd cell_6t
Xbit_r139_c158 bl_158 br_158 wl_139 vdd gnd cell_6t
Xbit_r140_c158 bl_158 br_158 wl_140 vdd gnd cell_6t
Xbit_r141_c158 bl_158 br_158 wl_141 vdd gnd cell_6t
Xbit_r142_c158 bl_158 br_158 wl_142 vdd gnd cell_6t
Xbit_r143_c158 bl_158 br_158 wl_143 vdd gnd cell_6t
Xbit_r144_c158 bl_158 br_158 wl_144 vdd gnd cell_6t
Xbit_r145_c158 bl_158 br_158 wl_145 vdd gnd cell_6t
Xbit_r146_c158 bl_158 br_158 wl_146 vdd gnd cell_6t
Xbit_r147_c158 bl_158 br_158 wl_147 vdd gnd cell_6t
Xbit_r148_c158 bl_158 br_158 wl_148 vdd gnd cell_6t
Xbit_r149_c158 bl_158 br_158 wl_149 vdd gnd cell_6t
Xbit_r150_c158 bl_158 br_158 wl_150 vdd gnd cell_6t
Xbit_r151_c158 bl_158 br_158 wl_151 vdd gnd cell_6t
Xbit_r152_c158 bl_158 br_158 wl_152 vdd gnd cell_6t
Xbit_r153_c158 bl_158 br_158 wl_153 vdd gnd cell_6t
Xbit_r154_c158 bl_158 br_158 wl_154 vdd gnd cell_6t
Xbit_r155_c158 bl_158 br_158 wl_155 vdd gnd cell_6t
Xbit_r156_c158 bl_158 br_158 wl_156 vdd gnd cell_6t
Xbit_r157_c158 bl_158 br_158 wl_157 vdd gnd cell_6t
Xbit_r158_c158 bl_158 br_158 wl_158 vdd gnd cell_6t
Xbit_r159_c158 bl_158 br_158 wl_159 vdd gnd cell_6t
Xbit_r160_c158 bl_158 br_158 wl_160 vdd gnd cell_6t
Xbit_r161_c158 bl_158 br_158 wl_161 vdd gnd cell_6t
Xbit_r162_c158 bl_158 br_158 wl_162 vdd gnd cell_6t
Xbit_r163_c158 bl_158 br_158 wl_163 vdd gnd cell_6t
Xbit_r164_c158 bl_158 br_158 wl_164 vdd gnd cell_6t
Xbit_r165_c158 bl_158 br_158 wl_165 vdd gnd cell_6t
Xbit_r166_c158 bl_158 br_158 wl_166 vdd gnd cell_6t
Xbit_r167_c158 bl_158 br_158 wl_167 vdd gnd cell_6t
Xbit_r168_c158 bl_158 br_158 wl_168 vdd gnd cell_6t
Xbit_r169_c158 bl_158 br_158 wl_169 vdd gnd cell_6t
Xbit_r170_c158 bl_158 br_158 wl_170 vdd gnd cell_6t
Xbit_r171_c158 bl_158 br_158 wl_171 vdd gnd cell_6t
Xbit_r172_c158 bl_158 br_158 wl_172 vdd gnd cell_6t
Xbit_r173_c158 bl_158 br_158 wl_173 vdd gnd cell_6t
Xbit_r174_c158 bl_158 br_158 wl_174 vdd gnd cell_6t
Xbit_r175_c158 bl_158 br_158 wl_175 vdd gnd cell_6t
Xbit_r176_c158 bl_158 br_158 wl_176 vdd gnd cell_6t
Xbit_r177_c158 bl_158 br_158 wl_177 vdd gnd cell_6t
Xbit_r178_c158 bl_158 br_158 wl_178 vdd gnd cell_6t
Xbit_r179_c158 bl_158 br_158 wl_179 vdd gnd cell_6t
Xbit_r180_c158 bl_158 br_158 wl_180 vdd gnd cell_6t
Xbit_r181_c158 bl_158 br_158 wl_181 vdd gnd cell_6t
Xbit_r182_c158 bl_158 br_158 wl_182 vdd gnd cell_6t
Xbit_r183_c158 bl_158 br_158 wl_183 vdd gnd cell_6t
Xbit_r184_c158 bl_158 br_158 wl_184 vdd gnd cell_6t
Xbit_r185_c158 bl_158 br_158 wl_185 vdd gnd cell_6t
Xbit_r186_c158 bl_158 br_158 wl_186 vdd gnd cell_6t
Xbit_r187_c158 bl_158 br_158 wl_187 vdd gnd cell_6t
Xbit_r188_c158 bl_158 br_158 wl_188 vdd gnd cell_6t
Xbit_r189_c158 bl_158 br_158 wl_189 vdd gnd cell_6t
Xbit_r190_c158 bl_158 br_158 wl_190 vdd gnd cell_6t
Xbit_r191_c158 bl_158 br_158 wl_191 vdd gnd cell_6t
Xbit_r192_c158 bl_158 br_158 wl_192 vdd gnd cell_6t
Xbit_r193_c158 bl_158 br_158 wl_193 vdd gnd cell_6t
Xbit_r194_c158 bl_158 br_158 wl_194 vdd gnd cell_6t
Xbit_r195_c158 bl_158 br_158 wl_195 vdd gnd cell_6t
Xbit_r196_c158 bl_158 br_158 wl_196 vdd gnd cell_6t
Xbit_r197_c158 bl_158 br_158 wl_197 vdd gnd cell_6t
Xbit_r198_c158 bl_158 br_158 wl_198 vdd gnd cell_6t
Xbit_r199_c158 bl_158 br_158 wl_199 vdd gnd cell_6t
Xbit_r200_c158 bl_158 br_158 wl_200 vdd gnd cell_6t
Xbit_r201_c158 bl_158 br_158 wl_201 vdd gnd cell_6t
Xbit_r202_c158 bl_158 br_158 wl_202 vdd gnd cell_6t
Xbit_r203_c158 bl_158 br_158 wl_203 vdd gnd cell_6t
Xbit_r204_c158 bl_158 br_158 wl_204 vdd gnd cell_6t
Xbit_r205_c158 bl_158 br_158 wl_205 vdd gnd cell_6t
Xbit_r206_c158 bl_158 br_158 wl_206 vdd gnd cell_6t
Xbit_r207_c158 bl_158 br_158 wl_207 vdd gnd cell_6t
Xbit_r208_c158 bl_158 br_158 wl_208 vdd gnd cell_6t
Xbit_r209_c158 bl_158 br_158 wl_209 vdd gnd cell_6t
Xbit_r210_c158 bl_158 br_158 wl_210 vdd gnd cell_6t
Xbit_r211_c158 bl_158 br_158 wl_211 vdd gnd cell_6t
Xbit_r212_c158 bl_158 br_158 wl_212 vdd gnd cell_6t
Xbit_r213_c158 bl_158 br_158 wl_213 vdd gnd cell_6t
Xbit_r214_c158 bl_158 br_158 wl_214 vdd gnd cell_6t
Xbit_r215_c158 bl_158 br_158 wl_215 vdd gnd cell_6t
Xbit_r216_c158 bl_158 br_158 wl_216 vdd gnd cell_6t
Xbit_r217_c158 bl_158 br_158 wl_217 vdd gnd cell_6t
Xbit_r218_c158 bl_158 br_158 wl_218 vdd gnd cell_6t
Xbit_r219_c158 bl_158 br_158 wl_219 vdd gnd cell_6t
Xbit_r220_c158 bl_158 br_158 wl_220 vdd gnd cell_6t
Xbit_r221_c158 bl_158 br_158 wl_221 vdd gnd cell_6t
Xbit_r222_c158 bl_158 br_158 wl_222 vdd gnd cell_6t
Xbit_r223_c158 bl_158 br_158 wl_223 vdd gnd cell_6t
Xbit_r224_c158 bl_158 br_158 wl_224 vdd gnd cell_6t
Xbit_r225_c158 bl_158 br_158 wl_225 vdd gnd cell_6t
Xbit_r226_c158 bl_158 br_158 wl_226 vdd gnd cell_6t
Xbit_r227_c158 bl_158 br_158 wl_227 vdd gnd cell_6t
Xbit_r228_c158 bl_158 br_158 wl_228 vdd gnd cell_6t
Xbit_r229_c158 bl_158 br_158 wl_229 vdd gnd cell_6t
Xbit_r230_c158 bl_158 br_158 wl_230 vdd gnd cell_6t
Xbit_r231_c158 bl_158 br_158 wl_231 vdd gnd cell_6t
Xbit_r232_c158 bl_158 br_158 wl_232 vdd gnd cell_6t
Xbit_r233_c158 bl_158 br_158 wl_233 vdd gnd cell_6t
Xbit_r234_c158 bl_158 br_158 wl_234 vdd gnd cell_6t
Xbit_r235_c158 bl_158 br_158 wl_235 vdd gnd cell_6t
Xbit_r236_c158 bl_158 br_158 wl_236 vdd gnd cell_6t
Xbit_r237_c158 bl_158 br_158 wl_237 vdd gnd cell_6t
Xbit_r238_c158 bl_158 br_158 wl_238 vdd gnd cell_6t
Xbit_r239_c158 bl_158 br_158 wl_239 vdd gnd cell_6t
Xbit_r240_c158 bl_158 br_158 wl_240 vdd gnd cell_6t
Xbit_r241_c158 bl_158 br_158 wl_241 vdd gnd cell_6t
Xbit_r242_c158 bl_158 br_158 wl_242 vdd gnd cell_6t
Xbit_r243_c158 bl_158 br_158 wl_243 vdd gnd cell_6t
Xbit_r244_c158 bl_158 br_158 wl_244 vdd gnd cell_6t
Xbit_r245_c158 bl_158 br_158 wl_245 vdd gnd cell_6t
Xbit_r246_c158 bl_158 br_158 wl_246 vdd gnd cell_6t
Xbit_r247_c158 bl_158 br_158 wl_247 vdd gnd cell_6t
Xbit_r248_c158 bl_158 br_158 wl_248 vdd gnd cell_6t
Xbit_r249_c158 bl_158 br_158 wl_249 vdd gnd cell_6t
Xbit_r250_c158 bl_158 br_158 wl_250 vdd gnd cell_6t
Xbit_r251_c158 bl_158 br_158 wl_251 vdd gnd cell_6t
Xbit_r252_c158 bl_158 br_158 wl_252 vdd gnd cell_6t
Xbit_r253_c158 bl_158 br_158 wl_253 vdd gnd cell_6t
Xbit_r254_c158 bl_158 br_158 wl_254 vdd gnd cell_6t
Xbit_r255_c158 bl_158 br_158 wl_255 vdd gnd cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd cell_6t
Xbit_r1_c159 bl_159 br_159 wl_1 vdd gnd cell_6t
Xbit_r2_c159 bl_159 br_159 wl_2 vdd gnd cell_6t
Xbit_r3_c159 bl_159 br_159 wl_3 vdd gnd cell_6t
Xbit_r4_c159 bl_159 br_159 wl_4 vdd gnd cell_6t
Xbit_r5_c159 bl_159 br_159 wl_5 vdd gnd cell_6t
Xbit_r6_c159 bl_159 br_159 wl_6 vdd gnd cell_6t
Xbit_r7_c159 bl_159 br_159 wl_7 vdd gnd cell_6t
Xbit_r8_c159 bl_159 br_159 wl_8 vdd gnd cell_6t
Xbit_r9_c159 bl_159 br_159 wl_9 vdd gnd cell_6t
Xbit_r10_c159 bl_159 br_159 wl_10 vdd gnd cell_6t
Xbit_r11_c159 bl_159 br_159 wl_11 vdd gnd cell_6t
Xbit_r12_c159 bl_159 br_159 wl_12 vdd gnd cell_6t
Xbit_r13_c159 bl_159 br_159 wl_13 vdd gnd cell_6t
Xbit_r14_c159 bl_159 br_159 wl_14 vdd gnd cell_6t
Xbit_r15_c159 bl_159 br_159 wl_15 vdd gnd cell_6t
Xbit_r16_c159 bl_159 br_159 wl_16 vdd gnd cell_6t
Xbit_r17_c159 bl_159 br_159 wl_17 vdd gnd cell_6t
Xbit_r18_c159 bl_159 br_159 wl_18 vdd gnd cell_6t
Xbit_r19_c159 bl_159 br_159 wl_19 vdd gnd cell_6t
Xbit_r20_c159 bl_159 br_159 wl_20 vdd gnd cell_6t
Xbit_r21_c159 bl_159 br_159 wl_21 vdd gnd cell_6t
Xbit_r22_c159 bl_159 br_159 wl_22 vdd gnd cell_6t
Xbit_r23_c159 bl_159 br_159 wl_23 vdd gnd cell_6t
Xbit_r24_c159 bl_159 br_159 wl_24 vdd gnd cell_6t
Xbit_r25_c159 bl_159 br_159 wl_25 vdd gnd cell_6t
Xbit_r26_c159 bl_159 br_159 wl_26 vdd gnd cell_6t
Xbit_r27_c159 bl_159 br_159 wl_27 vdd gnd cell_6t
Xbit_r28_c159 bl_159 br_159 wl_28 vdd gnd cell_6t
Xbit_r29_c159 bl_159 br_159 wl_29 vdd gnd cell_6t
Xbit_r30_c159 bl_159 br_159 wl_30 vdd gnd cell_6t
Xbit_r31_c159 bl_159 br_159 wl_31 vdd gnd cell_6t
Xbit_r32_c159 bl_159 br_159 wl_32 vdd gnd cell_6t
Xbit_r33_c159 bl_159 br_159 wl_33 vdd gnd cell_6t
Xbit_r34_c159 bl_159 br_159 wl_34 vdd gnd cell_6t
Xbit_r35_c159 bl_159 br_159 wl_35 vdd gnd cell_6t
Xbit_r36_c159 bl_159 br_159 wl_36 vdd gnd cell_6t
Xbit_r37_c159 bl_159 br_159 wl_37 vdd gnd cell_6t
Xbit_r38_c159 bl_159 br_159 wl_38 vdd gnd cell_6t
Xbit_r39_c159 bl_159 br_159 wl_39 vdd gnd cell_6t
Xbit_r40_c159 bl_159 br_159 wl_40 vdd gnd cell_6t
Xbit_r41_c159 bl_159 br_159 wl_41 vdd gnd cell_6t
Xbit_r42_c159 bl_159 br_159 wl_42 vdd gnd cell_6t
Xbit_r43_c159 bl_159 br_159 wl_43 vdd gnd cell_6t
Xbit_r44_c159 bl_159 br_159 wl_44 vdd gnd cell_6t
Xbit_r45_c159 bl_159 br_159 wl_45 vdd gnd cell_6t
Xbit_r46_c159 bl_159 br_159 wl_46 vdd gnd cell_6t
Xbit_r47_c159 bl_159 br_159 wl_47 vdd gnd cell_6t
Xbit_r48_c159 bl_159 br_159 wl_48 vdd gnd cell_6t
Xbit_r49_c159 bl_159 br_159 wl_49 vdd gnd cell_6t
Xbit_r50_c159 bl_159 br_159 wl_50 vdd gnd cell_6t
Xbit_r51_c159 bl_159 br_159 wl_51 vdd gnd cell_6t
Xbit_r52_c159 bl_159 br_159 wl_52 vdd gnd cell_6t
Xbit_r53_c159 bl_159 br_159 wl_53 vdd gnd cell_6t
Xbit_r54_c159 bl_159 br_159 wl_54 vdd gnd cell_6t
Xbit_r55_c159 bl_159 br_159 wl_55 vdd gnd cell_6t
Xbit_r56_c159 bl_159 br_159 wl_56 vdd gnd cell_6t
Xbit_r57_c159 bl_159 br_159 wl_57 vdd gnd cell_6t
Xbit_r58_c159 bl_159 br_159 wl_58 vdd gnd cell_6t
Xbit_r59_c159 bl_159 br_159 wl_59 vdd gnd cell_6t
Xbit_r60_c159 bl_159 br_159 wl_60 vdd gnd cell_6t
Xbit_r61_c159 bl_159 br_159 wl_61 vdd gnd cell_6t
Xbit_r62_c159 bl_159 br_159 wl_62 vdd gnd cell_6t
Xbit_r63_c159 bl_159 br_159 wl_63 vdd gnd cell_6t
Xbit_r64_c159 bl_159 br_159 wl_64 vdd gnd cell_6t
Xbit_r65_c159 bl_159 br_159 wl_65 vdd gnd cell_6t
Xbit_r66_c159 bl_159 br_159 wl_66 vdd gnd cell_6t
Xbit_r67_c159 bl_159 br_159 wl_67 vdd gnd cell_6t
Xbit_r68_c159 bl_159 br_159 wl_68 vdd gnd cell_6t
Xbit_r69_c159 bl_159 br_159 wl_69 vdd gnd cell_6t
Xbit_r70_c159 bl_159 br_159 wl_70 vdd gnd cell_6t
Xbit_r71_c159 bl_159 br_159 wl_71 vdd gnd cell_6t
Xbit_r72_c159 bl_159 br_159 wl_72 vdd gnd cell_6t
Xbit_r73_c159 bl_159 br_159 wl_73 vdd gnd cell_6t
Xbit_r74_c159 bl_159 br_159 wl_74 vdd gnd cell_6t
Xbit_r75_c159 bl_159 br_159 wl_75 vdd gnd cell_6t
Xbit_r76_c159 bl_159 br_159 wl_76 vdd gnd cell_6t
Xbit_r77_c159 bl_159 br_159 wl_77 vdd gnd cell_6t
Xbit_r78_c159 bl_159 br_159 wl_78 vdd gnd cell_6t
Xbit_r79_c159 bl_159 br_159 wl_79 vdd gnd cell_6t
Xbit_r80_c159 bl_159 br_159 wl_80 vdd gnd cell_6t
Xbit_r81_c159 bl_159 br_159 wl_81 vdd gnd cell_6t
Xbit_r82_c159 bl_159 br_159 wl_82 vdd gnd cell_6t
Xbit_r83_c159 bl_159 br_159 wl_83 vdd gnd cell_6t
Xbit_r84_c159 bl_159 br_159 wl_84 vdd gnd cell_6t
Xbit_r85_c159 bl_159 br_159 wl_85 vdd gnd cell_6t
Xbit_r86_c159 bl_159 br_159 wl_86 vdd gnd cell_6t
Xbit_r87_c159 bl_159 br_159 wl_87 vdd gnd cell_6t
Xbit_r88_c159 bl_159 br_159 wl_88 vdd gnd cell_6t
Xbit_r89_c159 bl_159 br_159 wl_89 vdd gnd cell_6t
Xbit_r90_c159 bl_159 br_159 wl_90 vdd gnd cell_6t
Xbit_r91_c159 bl_159 br_159 wl_91 vdd gnd cell_6t
Xbit_r92_c159 bl_159 br_159 wl_92 vdd gnd cell_6t
Xbit_r93_c159 bl_159 br_159 wl_93 vdd gnd cell_6t
Xbit_r94_c159 bl_159 br_159 wl_94 vdd gnd cell_6t
Xbit_r95_c159 bl_159 br_159 wl_95 vdd gnd cell_6t
Xbit_r96_c159 bl_159 br_159 wl_96 vdd gnd cell_6t
Xbit_r97_c159 bl_159 br_159 wl_97 vdd gnd cell_6t
Xbit_r98_c159 bl_159 br_159 wl_98 vdd gnd cell_6t
Xbit_r99_c159 bl_159 br_159 wl_99 vdd gnd cell_6t
Xbit_r100_c159 bl_159 br_159 wl_100 vdd gnd cell_6t
Xbit_r101_c159 bl_159 br_159 wl_101 vdd gnd cell_6t
Xbit_r102_c159 bl_159 br_159 wl_102 vdd gnd cell_6t
Xbit_r103_c159 bl_159 br_159 wl_103 vdd gnd cell_6t
Xbit_r104_c159 bl_159 br_159 wl_104 vdd gnd cell_6t
Xbit_r105_c159 bl_159 br_159 wl_105 vdd gnd cell_6t
Xbit_r106_c159 bl_159 br_159 wl_106 vdd gnd cell_6t
Xbit_r107_c159 bl_159 br_159 wl_107 vdd gnd cell_6t
Xbit_r108_c159 bl_159 br_159 wl_108 vdd gnd cell_6t
Xbit_r109_c159 bl_159 br_159 wl_109 vdd gnd cell_6t
Xbit_r110_c159 bl_159 br_159 wl_110 vdd gnd cell_6t
Xbit_r111_c159 bl_159 br_159 wl_111 vdd gnd cell_6t
Xbit_r112_c159 bl_159 br_159 wl_112 vdd gnd cell_6t
Xbit_r113_c159 bl_159 br_159 wl_113 vdd gnd cell_6t
Xbit_r114_c159 bl_159 br_159 wl_114 vdd gnd cell_6t
Xbit_r115_c159 bl_159 br_159 wl_115 vdd gnd cell_6t
Xbit_r116_c159 bl_159 br_159 wl_116 vdd gnd cell_6t
Xbit_r117_c159 bl_159 br_159 wl_117 vdd gnd cell_6t
Xbit_r118_c159 bl_159 br_159 wl_118 vdd gnd cell_6t
Xbit_r119_c159 bl_159 br_159 wl_119 vdd gnd cell_6t
Xbit_r120_c159 bl_159 br_159 wl_120 vdd gnd cell_6t
Xbit_r121_c159 bl_159 br_159 wl_121 vdd gnd cell_6t
Xbit_r122_c159 bl_159 br_159 wl_122 vdd gnd cell_6t
Xbit_r123_c159 bl_159 br_159 wl_123 vdd gnd cell_6t
Xbit_r124_c159 bl_159 br_159 wl_124 vdd gnd cell_6t
Xbit_r125_c159 bl_159 br_159 wl_125 vdd gnd cell_6t
Xbit_r126_c159 bl_159 br_159 wl_126 vdd gnd cell_6t
Xbit_r127_c159 bl_159 br_159 wl_127 vdd gnd cell_6t
Xbit_r128_c159 bl_159 br_159 wl_128 vdd gnd cell_6t
Xbit_r129_c159 bl_159 br_159 wl_129 vdd gnd cell_6t
Xbit_r130_c159 bl_159 br_159 wl_130 vdd gnd cell_6t
Xbit_r131_c159 bl_159 br_159 wl_131 vdd gnd cell_6t
Xbit_r132_c159 bl_159 br_159 wl_132 vdd gnd cell_6t
Xbit_r133_c159 bl_159 br_159 wl_133 vdd gnd cell_6t
Xbit_r134_c159 bl_159 br_159 wl_134 vdd gnd cell_6t
Xbit_r135_c159 bl_159 br_159 wl_135 vdd gnd cell_6t
Xbit_r136_c159 bl_159 br_159 wl_136 vdd gnd cell_6t
Xbit_r137_c159 bl_159 br_159 wl_137 vdd gnd cell_6t
Xbit_r138_c159 bl_159 br_159 wl_138 vdd gnd cell_6t
Xbit_r139_c159 bl_159 br_159 wl_139 vdd gnd cell_6t
Xbit_r140_c159 bl_159 br_159 wl_140 vdd gnd cell_6t
Xbit_r141_c159 bl_159 br_159 wl_141 vdd gnd cell_6t
Xbit_r142_c159 bl_159 br_159 wl_142 vdd gnd cell_6t
Xbit_r143_c159 bl_159 br_159 wl_143 vdd gnd cell_6t
Xbit_r144_c159 bl_159 br_159 wl_144 vdd gnd cell_6t
Xbit_r145_c159 bl_159 br_159 wl_145 vdd gnd cell_6t
Xbit_r146_c159 bl_159 br_159 wl_146 vdd gnd cell_6t
Xbit_r147_c159 bl_159 br_159 wl_147 vdd gnd cell_6t
Xbit_r148_c159 bl_159 br_159 wl_148 vdd gnd cell_6t
Xbit_r149_c159 bl_159 br_159 wl_149 vdd gnd cell_6t
Xbit_r150_c159 bl_159 br_159 wl_150 vdd gnd cell_6t
Xbit_r151_c159 bl_159 br_159 wl_151 vdd gnd cell_6t
Xbit_r152_c159 bl_159 br_159 wl_152 vdd gnd cell_6t
Xbit_r153_c159 bl_159 br_159 wl_153 vdd gnd cell_6t
Xbit_r154_c159 bl_159 br_159 wl_154 vdd gnd cell_6t
Xbit_r155_c159 bl_159 br_159 wl_155 vdd gnd cell_6t
Xbit_r156_c159 bl_159 br_159 wl_156 vdd gnd cell_6t
Xbit_r157_c159 bl_159 br_159 wl_157 vdd gnd cell_6t
Xbit_r158_c159 bl_159 br_159 wl_158 vdd gnd cell_6t
Xbit_r159_c159 bl_159 br_159 wl_159 vdd gnd cell_6t
Xbit_r160_c159 bl_159 br_159 wl_160 vdd gnd cell_6t
Xbit_r161_c159 bl_159 br_159 wl_161 vdd gnd cell_6t
Xbit_r162_c159 bl_159 br_159 wl_162 vdd gnd cell_6t
Xbit_r163_c159 bl_159 br_159 wl_163 vdd gnd cell_6t
Xbit_r164_c159 bl_159 br_159 wl_164 vdd gnd cell_6t
Xbit_r165_c159 bl_159 br_159 wl_165 vdd gnd cell_6t
Xbit_r166_c159 bl_159 br_159 wl_166 vdd gnd cell_6t
Xbit_r167_c159 bl_159 br_159 wl_167 vdd gnd cell_6t
Xbit_r168_c159 bl_159 br_159 wl_168 vdd gnd cell_6t
Xbit_r169_c159 bl_159 br_159 wl_169 vdd gnd cell_6t
Xbit_r170_c159 bl_159 br_159 wl_170 vdd gnd cell_6t
Xbit_r171_c159 bl_159 br_159 wl_171 vdd gnd cell_6t
Xbit_r172_c159 bl_159 br_159 wl_172 vdd gnd cell_6t
Xbit_r173_c159 bl_159 br_159 wl_173 vdd gnd cell_6t
Xbit_r174_c159 bl_159 br_159 wl_174 vdd gnd cell_6t
Xbit_r175_c159 bl_159 br_159 wl_175 vdd gnd cell_6t
Xbit_r176_c159 bl_159 br_159 wl_176 vdd gnd cell_6t
Xbit_r177_c159 bl_159 br_159 wl_177 vdd gnd cell_6t
Xbit_r178_c159 bl_159 br_159 wl_178 vdd gnd cell_6t
Xbit_r179_c159 bl_159 br_159 wl_179 vdd gnd cell_6t
Xbit_r180_c159 bl_159 br_159 wl_180 vdd gnd cell_6t
Xbit_r181_c159 bl_159 br_159 wl_181 vdd gnd cell_6t
Xbit_r182_c159 bl_159 br_159 wl_182 vdd gnd cell_6t
Xbit_r183_c159 bl_159 br_159 wl_183 vdd gnd cell_6t
Xbit_r184_c159 bl_159 br_159 wl_184 vdd gnd cell_6t
Xbit_r185_c159 bl_159 br_159 wl_185 vdd gnd cell_6t
Xbit_r186_c159 bl_159 br_159 wl_186 vdd gnd cell_6t
Xbit_r187_c159 bl_159 br_159 wl_187 vdd gnd cell_6t
Xbit_r188_c159 bl_159 br_159 wl_188 vdd gnd cell_6t
Xbit_r189_c159 bl_159 br_159 wl_189 vdd gnd cell_6t
Xbit_r190_c159 bl_159 br_159 wl_190 vdd gnd cell_6t
Xbit_r191_c159 bl_159 br_159 wl_191 vdd gnd cell_6t
Xbit_r192_c159 bl_159 br_159 wl_192 vdd gnd cell_6t
Xbit_r193_c159 bl_159 br_159 wl_193 vdd gnd cell_6t
Xbit_r194_c159 bl_159 br_159 wl_194 vdd gnd cell_6t
Xbit_r195_c159 bl_159 br_159 wl_195 vdd gnd cell_6t
Xbit_r196_c159 bl_159 br_159 wl_196 vdd gnd cell_6t
Xbit_r197_c159 bl_159 br_159 wl_197 vdd gnd cell_6t
Xbit_r198_c159 bl_159 br_159 wl_198 vdd gnd cell_6t
Xbit_r199_c159 bl_159 br_159 wl_199 vdd gnd cell_6t
Xbit_r200_c159 bl_159 br_159 wl_200 vdd gnd cell_6t
Xbit_r201_c159 bl_159 br_159 wl_201 vdd gnd cell_6t
Xbit_r202_c159 bl_159 br_159 wl_202 vdd gnd cell_6t
Xbit_r203_c159 bl_159 br_159 wl_203 vdd gnd cell_6t
Xbit_r204_c159 bl_159 br_159 wl_204 vdd gnd cell_6t
Xbit_r205_c159 bl_159 br_159 wl_205 vdd gnd cell_6t
Xbit_r206_c159 bl_159 br_159 wl_206 vdd gnd cell_6t
Xbit_r207_c159 bl_159 br_159 wl_207 vdd gnd cell_6t
Xbit_r208_c159 bl_159 br_159 wl_208 vdd gnd cell_6t
Xbit_r209_c159 bl_159 br_159 wl_209 vdd gnd cell_6t
Xbit_r210_c159 bl_159 br_159 wl_210 vdd gnd cell_6t
Xbit_r211_c159 bl_159 br_159 wl_211 vdd gnd cell_6t
Xbit_r212_c159 bl_159 br_159 wl_212 vdd gnd cell_6t
Xbit_r213_c159 bl_159 br_159 wl_213 vdd gnd cell_6t
Xbit_r214_c159 bl_159 br_159 wl_214 vdd gnd cell_6t
Xbit_r215_c159 bl_159 br_159 wl_215 vdd gnd cell_6t
Xbit_r216_c159 bl_159 br_159 wl_216 vdd gnd cell_6t
Xbit_r217_c159 bl_159 br_159 wl_217 vdd gnd cell_6t
Xbit_r218_c159 bl_159 br_159 wl_218 vdd gnd cell_6t
Xbit_r219_c159 bl_159 br_159 wl_219 vdd gnd cell_6t
Xbit_r220_c159 bl_159 br_159 wl_220 vdd gnd cell_6t
Xbit_r221_c159 bl_159 br_159 wl_221 vdd gnd cell_6t
Xbit_r222_c159 bl_159 br_159 wl_222 vdd gnd cell_6t
Xbit_r223_c159 bl_159 br_159 wl_223 vdd gnd cell_6t
Xbit_r224_c159 bl_159 br_159 wl_224 vdd gnd cell_6t
Xbit_r225_c159 bl_159 br_159 wl_225 vdd gnd cell_6t
Xbit_r226_c159 bl_159 br_159 wl_226 vdd gnd cell_6t
Xbit_r227_c159 bl_159 br_159 wl_227 vdd gnd cell_6t
Xbit_r228_c159 bl_159 br_159 wl_228 vdd gnd cell_6t
Xbit_r229_c159 bl_159 br_159 wl_229 vdd gnd cell_6t
Xbit_r230_c159 bl_159 br_159 wl_230 vdd gnd cell_6t
Xbit_r231_c159 bl_159 br_159 wl_231 vdd gnd cell_6t
Xbit_r232_c159 bl_159 br_159 wl_232 vdd gnd cell_6t
Xbit_r233_c159 bl_159 br_159 wl_233 vdd gnd cell_6t
Xbit_r234_c159 bl_159 br_159 wl_234 vdd gnd cell_6t
Xbit_r235_c159 bl_159 br_159 wl_235 vdd gnd cell_6t
Xbit_r236_c159 bl_159 br_159 wl_236 vdd gnd cell_6t
Xbit_r237_c159 bl_159 br_159 wl_237 vdd gnd cell_6t
Xbit_r238_c159 bl_159 br_159 wl_238 vdd gnd cell_6t
Xbit_r239_c159 bl_159 br_159 wl_239 vdd gnd cell_6t
Xbit_r240_c159 bl_159 br_159 wl_240 vdd gnd cell_6t
Xbit_r241_c159 bl_159 br_159 wl_241 vdd gnd cell_6t
Xbit_r242_c159 bl_159 br_159 wl_242 vdd gnd cell_6t
Xbit_r243_c159 bl_159 br_159 wl_243 vdd gnd cell_6t
Xbit_r244_c159 bl_159 br_159 wl_244 vdd gnd cell_6t
Xbit_r245_c159 bl_159 br_159 wl_245 vdd gnd cell_6t
Xbit_r246_c159 bl_159 br_159 wl_246 vdd gnd cell_6t
Xbit_r247_c159 bl_159 br_159 wl_247 vdd gnd cell_6t
Xbit_r248_c159 bl_159 br_159 wl_248 vdd gnd cell_6t
Xbit_r249_c159 bl_159 br_159 wl_249 vdd gnd cell_6t
Xbit_r250_c159 bl_159 br_159 wl_250 vdd gnd cell_6t
Xbit_r251_c159 bl_159 br_159 wl_251 vdd gnd cell_6t
Xbit_r252_c159 bl_159 br_159 wl_252 vdd gnd cell_6t
Xbit_r253_c159 bl_159 br_159 wl_253 vdd gnd cell_6t
Xbit_r254_c159 bl_159 br_159 wl_254 vdd gnd cell_6t
Xbit_r255_c159 bl_159 br_159 wl_255 vdd gnd cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd cell_6t
Xbit_r1_c160 bl_160 br_160 wl_1 vdd gnd cell_6t
Xbit_r2_c160 bl_160 br_160 wl_2 vdd gnd cell_6t
Xbit_r3_c160 bl_160 br_160 wl_3 vdd gnd cell_6t
Xbit_r4_c160 bl_160 br_160 wl_4 vdd gnd cell_6t
Xbit_r5_c160 bl_160 br_160 wl_5 vdd gnd cell_6t
Xbit_r6_c160 bl_160 br_160 wl_6 vdd gnd cell_6t
Xbit_r7_c160 bl_160 br_160 wl_7 vdd gnd cell_6t
Xbit_r8_c160 bl_160 br_160 wl_8 vdd gnd cell_6t
Xbit_r9_c160 bl_160 br_160 wl_9 vdd gnd cell_6t
Xbit_r10_c160 bl_160 br_160 wl_10 vdd gnd cell_6t
Xbit_r11_c160 bl_160 br_160 wl_11 vdd gnd cell_6t
Xbit_r12_c160 bl_160 br_160 wl_12 vdd gnd cell_6t
Xbit_r13_c160 bl_160 br_160 wl_13 vdd gnd cell_6t
Xbit_r14_c160 bl_160 br_160 wl_14 vdd gnd cell_6t
Xbit_r15_c160 bl_160 br_160 wl_15 vdd gnd cell_6t
Xbit_r16_c160 bl_160 br_160 wl_16 vdd gnd cell_6t
Xbit_r17_c160 bl_160 br_160 wl_17 vdd gnd cell_6t
Xbit_r18_c160 bl_160 br_160 wl_18 vdd gnd cell_6t
Xbit_r19_c160 bl_160 br_160 wl_19 vdd gnd cell_6t
Xbit_r20_c160 bl_160 br_160 wl_20 vdd gnd cell_6t
Xbit_r21_c160 bl_160 br_160 wl_21 vdd gnd cell_6t
Xbit_r22_c160 bl_160 br_160 wl_22 vdd gnd cell_6t
Xbit_r23_c160 bl_160 br_160 wl_23 vdd gnd cell_6t
Xbit_r24_c160 bl_160 br_160 wl_24 vdd gnd cell_6t
Xbit_r25_c160 bl_160 br_160 wl_25 vdd gnd cell_6t
Xbit_r26_c160 bl_160 br_160 wl_26 vdd gnd cell_6t
Xbit_r27_c160 bl_160 br_160 wl_27 vdd gnd cell_6t
Xbit_r28_c160 bl_160 br_160 wl_28 vdd gnd cell_6t
Xbit_r29_c160 bl_160 br_160 wl_29 vdd gnd cell_6t
Xbit_r30_c160 bl_160 br_160 wl_30 vdd gnd cell_6t
Xbit_r31_c160 bl_160 br_160 wl_31 vdd gnd cell_6t
Xbit_r32_c160 bl_160 br_160 wl_32 vdd gnd cell_6t
Xbit_r33_c160 bl_160 br_160 wl_33 vdd gnd cell_6t
Xbit_r34_c160 bl_160 br_160 wl_34 vdd gnd cell_6t
Xbit_r35_c160 bl_160 br_160 wl_35 vdd gnd cell_6t
Xbit_r36_c160 bl_160 br_160 wl_36 vdd gnd cell_6t
Xbit_r37_c160 bl_160 br_160 wl_37 vdd gnd cell_6t
Xbit_r38_c160 bl_160 br_160 wl_38 vdd gnd cell_6t
Xbit_r39_c160 bl_160 br_160 wl_39 vdd gnd cell_6t
Xbit_r40_c160 bl_160 br_160 wl_40 vdd gnd cell_6t
Xbit_r41_c160 bl_160 br_160 wl_41 vdd gnd cell_6t
Xbit_r42_c160 bl_160 br_160 wl_42 vdd gnd cell_6t
Xbit_r43_c160 bl_160 br_160 wl_43 vdd gnd cell_6t
Xbit_r44_c160 bl_160 br_160 wl_44 vdd gnd cell_6t
Xbit_r45_c160 bl_160 br_160 wl_45 vdd gnd cell_6t
Xbit_r46_c160 bl_160 br_160 wl_46 vdd gnd cell_6t
Xbit_r47_c160 bl_160 br_160 wl_47 vdd gnd cell_6t
Xbit_r48_c160 bl_160 br_160 wl_48 vdd gnd cell_6t
Xbit_r49_c160 bl_160 br_160 wl_49 vdd gnd cell_6t
Xbit_r50_c160 bl_160 br_160 wl_50 vdd gnd cell_6t
Xbit_r51_c160 bl_160 br_160 wl_51 vdd gnd cell_6t
Xbit_r52_c160 bl_160 br_160 wl_52 vdd gnd cell_6t
Xbit_r53_c160 bl_160 br_160 wl_53 vdd gnd cell_6t
Xbit_r54_c160 bl_160 br_160 wl_54 vdd gnd cell_6t
Xbit_r55_c160 bl_160 br_160 wl_55 vdd gnd cell_6t
Xbit_r56_c160 bl_160 br_160 wl_56 vdd gnd cell_6t
Xbit_r57_c160 bl_160 br_160 wl_57 vdd gnd cell_6t
Xbit_r58_c160 bl_160 br_160 wl_58 vdd gnd cell_6t
Xbit_r59_c160 bl_160 br_160 wl_59 vdd gnd cell_6t
Xbit_r60_c160 bl_160 br_160 wl_60 vdd gnd cell_6t
Xbit_r61_c160 bl_160 br_160 wl_61 vdd gnd cell_6t
Xbit_r62_c160 bl_160 br_160 wl_62 vdd gnd cell_6t
Xbit_r63_c160 bl_160 br_160 wl_63 vdd gnd cell_6t
Xbit_r64_c160 bl_160 br_160 wl_64 vdd gnd cell_6t
Xbit_r65_c160 bl_160 br_160 wl_65 vdd gnd cell_6t
Xbit_r66_c160 bl_160 br_160 wl_66 vdd gnd cell_6t
Xbit_r67_c160 bl_160 br_160 wl_67 vdd gnd cell_6t
Xbit_r68_c160 bl_160 br_160 wl_68 vdd gnd cell_6t
Xbit_r69_c160 bl_160 br_160 wl_69 vdd gnd cell_6t
Xbit_r70_c160 bl_160 br_160 wl_70 vdd gnd cell_6t
Xbit_r71_c160 bl_160 br_160 wl_71 vdd gnd cell_6t
Xbit_r72_c160 bl_160 br_160 wl_72 vdd gnd cell_6t
Xbit_r73_c160 bl_160 br_160 wl_73 vdd gnd cell_6t
Xbit_r74_c160 bl_160 br_160 wl_74 vdd gnd cell_6t
Xbit_r75_c160 bl_160 br_160 wl_75 vdd gnd cell_6t
Xbit_r76_c160 bl_160 br_160 wl_76 vdd gnd cell_6t
Xbit_r77_c160 bl_160 br_160 wl_77 vdd gnd cell_6t
Xbit_r78_c160 bl_160 br_160 wl_78 vdd gnd cell_6t
Xbit_r79_c160 bl_160 br_160 wl_79 vdd gnd cell_6t
Xbit_r80_c160 bl_160 br_160 wl_80 vdd gnd cell_6t
Xbit_r81_c160 bl_160 br_160 wl_81 vdd gnd cell_6t
Xbit_r82_c160 bl_160 br_160 wl_82 vdd gnd cell_6t
Xbit_r83_c160 bl_160 br_160 wl_83 vdd gnd cell_6t
Xbit_r84_c160 bl_160 br_160 wl_84 vdd gnd cell_6t
Xbit_r85_c160 bl_160 br_160 wl_85 vdd gnd cell_6t
Xbit_r86_c160 bl_160 br_160 wl_86 vdd gnd cell_6t
Xbit_r87_c160 bl_160 br_160 wl_87 vdd gnd cell_6t
Xbit_r88_c160 bl_160 br_160 wl_88 vdd gnd cell_6t
Xbit_r89_c160 bl_160 br_160 wl_89 vdd gnd cell_6t
Xbit_r90_c160 bl_160 br_160 wl_90 vdd gnd cell_6t
Xbit_r91_c160 bl_160 br_160 wl_91 vdd gnd cell_6t
Xbit_r92_c160 bl_160 br_160 wl_92 vdd gnd cell_6t
Xbit_r93_c160 bl_160 br_160 wl_93 vdd gnd cell_6t
Xbit_r94_c160 bl_160 br_160 wl_94 vdd gnd cell_6t
Xbit_r95_c160 bl_160 br_160 wl_95 vdd gnd cell_6t
Xbit_r96_c160 bl_160 br_160 wl_96 vdd gnd cell_6t
Xbit_r97_c160 bl_160 br_160 wl_97 vdd gnd cell_6t
Xbit_r98_c160 bl_160 br_160 wl_98 vdd gnd cell_6t
Xbit_r99_c160 bl_160 br_160 wl_99 vdd gnd cell_6t
Xbit_r100_c160 bl_160 br_160 wl_100 vdd gnd cell_6t
Xbit_r101_c160 bl_160 br_160 wl_101 vdd gnd cell_6t
Xbit_r102_c160 bl_160 br_160 wl_102 vdd gnd cell_6t
Xbit_r103_c160 bl_160 br_160 wl_103 vdd gnd cell_6t
Xbit_r104_c160 bl_160 br_160 wl_104 vdd gnd cell_6t
Xbit_r105_c160 bl_160 br_160 wl_105 vdd gnd cell_6t
Xbit_r106_c160 bl_160 br_160 wl_106 vdd gnd cell_6t
Xbit_r107_c160 bl_160 br_160 wl_107 vdd gnd cell_6t
Xbit_r108_c160 bl_160 br_160 wl_108 vdd gnd cell_6t
Xbit_r109_c160 bl_160 br_160 wl_109 vdd gnd cell_6t
Xbit_r110_c160 bl_160 br_160 wl_110 vdd gnd cell_6t
Xbit_r111_c160 bl_160 br_160 wl_111 vdd gnd cell_6t
Xbit_r112_c160 bl_160 br_160 wl_112 vdd gnd cell_6t
Xbit_r113_c160 bl_160 br_160 wl_113 vdd gnd cell_6t
Xbit_r114_c160 bl_160 br_160 wl_114 vdd gnd cell_6t
Xbit_r115_c160 bl_160 br_160 wl_115 vdd gnd cell_6t
Xbit_r116_c160 bl_160 br_160 wl_116 vdd gnd cell_6t
Xbit_r117_c160 bl_160 br_160 wl_117 vdd gnd cell_6t
Xbit_r118_c160 bl_160 br_160 wl_118 vdd gnd cell_6t
Xbit_r119_c160 bl_160 br_160 wl_119 vdd gnd cell_6t
Xbit_r120_c160 bl_160 br_160 wl_120 vdd gnd cell_6t
Xbit_r121_c160 bl_160 br_160 wl_121 vdd gnd cell_6t
Xbit_r122_c160 bl_160 br_160 wl_122 vdd gnd cell_6t
Xbit_r123_c160 bl_160 br_160 wl_123 vdd gnd cell_6t
Xbit_r124_c160 bl_160 br_160 wl_124 vdd gnd cell_6t
Xbit_r125_c160 bl_160 br_160 wl_125 vdd gnd cell_6t
Xbit_r126_c160 bl_160 br_160 wl_126 vdd gnd cell_6t
Xbit_r127_c160 bl_160 br_160 wl_127 vdd gnd cell_6t
Xbit_r128_c160 bl_160 br_160 wl_128 vdd gnd cell_6t
Xbit_r129_c160 bl_160 br_160 wl_129 vdd gnd cell_6t
Xbit_r130_c160 bl_160 br_160 wl_130 vdd gnd cell_6t
Xbit_r131_c160 bl_160 br_160 wl_131 vdd gnd cell_6t
Xbit_r132_c160 bl_160 br_160 wl_132 vdd gnd cell_6t
Xbit_r133_c160 bl_160 br_160 wl_133 vdd gnd cell_6t
Xbit_r134_c160 bl_160 br_160 wl_134 vdd gnd cell_6t
Xbit_r135_c160 bl_160 br_160 wl_135 vdd gnd cell_6t
Xbit_r136_c160 bl_160 br_160 wl_136 vdd gnd cell_6t
Xbit_r137_c160 bl_160 br_160 wl_137 vdd gnd cell_6t
Xbit_r138_c160 bl_160 br_160 wl_138 vdd gnd cell_6t
Xbit_r139_c160 bl_160 br_160 wl_139 vdd gnd cell_6t
Xbit_r140_c160 bl_160 br_160 wl_140 vdd gnd cell_6t
Xbit_r141_c160 bl_160 br_160 wl_141 vdd gnd cell_6t
Xbit_r142_c160 bl_160 br_160 wl_142 vdd gnd cell_6t
Xbit_r143_c160 bl_160 br_160 wl_143 vdd gnd cell_6t
Xbit_r144_c160 bl_160 br_160 wl_144 vdd gnd cell_6t
Xbit_r145_c160 bl_160 br_160 wl_145 vdd gnd cell_6t
Xbit_r146_c160 bl_160 br_160 wl_146 vdd gnd cell_6t
Xbit_r147_c160 bl_160 br_160 wl_147 vdd gnd cell_6t
Xbit_r148_c160 bl_160 br_160 wl_148 vdd gnd cell_6t
Xbit_r149_c160 bl_160 br_160 wl_149 vdd gnd cell_6t
Xbit_r150_c160 bl_160 br_160 wl_150 vdd gnd cell_6t
Xbit_r151_c160 bl_160 br_160 wl_151 vdd gnd cell_6t
Xbit_r152_c160 bl_160 br_160 wl_152 vdd gnd cell_6t
Xbit_r153_c160 bl_160 br_160 wl_153 vdd gnd cell_6t
Xbit_r154_c160 bl_160 br_160 wl_154 vdd gnd cell_6t
Xbit_r155_c160 bl_160 br_160 wl_155 vdd gnd cell_6t
Xbit_r156_c160 bl_160 br_160 wl_156 vdd gnd cell_6t
Xbit_r157_c160 bl_160 br_160 wl_157 vdd gnd cell_6t
Xbit_r158_c160 bl_160 br_160 wl_158 vdd gnd cell_6t
Xbit_r159_c160 bl_160 br_160 wl_159 vdd gnd cell_6t
Xbit_r160_c160 bl_160 br_160 wl_160 vdd gnd cell_6t
Xbit_r161_c160 bl_160 br_160 wl_161 vdd gnd cell_6t
Xbit_r162_c160 bl_160 br_160 wl_162 vdd gnd cell_6t
Xbit_r163_c160 bl_160 br_160 wl_163 vdd gnd cell_6t
Xbit_r164_c160 bl_160 br_160 wl_164 vdd gnd cell_6t
Xbit_r165_c160 bl_160 br_160 wl_165 vdd gnd cell_6t
Xbit_r166_c160 bl_160 br_160 wl_166 vdd gnd cell_6t
Xbit_r167_c160 bl_160 br_160 wl_167 vdd gnd cell_6t
Xbit_r168_c160 bl_160 br_160 wl_168 vdd gnd cell_6t
Xbit_r169_c160 bl_160 br_160 wl_169 vdd gnd cell_6t
Xbit_r170_c160 bl_160 br_160 wl_170 vdd gnd cell_6t
Xbit_r171_c160 bl_160 br_160 wl_171 vdd gnd cell_6t
Xbit_r172_c160 bl_160 br_160 wl_172 vdd gnd cell_6t
Xbit_r173_c160 bl_160 br_160 wl_173 vdd gnd cell_6t
Xbit_r174_c160 bl_160 br_160 wl_174 vdd gnd cell_6t
Xbit_r175_c160 bl_160 br_160 wl_175 vdd gnd cell_6t
Xbit_r176_c160 bl_160 br_160 wl_176 vdd gnd cell_6t
Xbit_r177_c160 bl_160 br_160 wl_177 vdd gnd cell_6t
Xbit_r178_c160 bl_160 br_160 wl_178 vdd gnd cell_6t
Xbit_r179_c160 bl_160 br_160 wl_179 vdd gnd cell_6t
Xbit_r180_c160 bl_160 br_160 wl_180 vdd gnd cell_6t
Xbit_r181_c160 bl_160 br_160 wl_181 vdd gnd cell_6t
Xbit_r182_c160 bl_160 br_160 wl_182 vdd gnd cell_6t
Xbit_r183_c160 bl_160 br_160 wl_183 vdd gnd cell_6t
Xbit_r184_c160 bl_160 br_160 wl_184 vdd gnd cell_6t
Xbit_r185_c160 bl_160 br_160 wl_185 vdd gnd cell_6t
Xbit_r186_c160 bl_160 br_160 wl_186 vdd gnd cell_6t
Xbit_r187_c160 bl_160 br_160 wl_187 vdd gnd cell_6t
Xbit_r188_c160 bl_160 br_160 wl_188 vdd gnd cell_6t
Xbit_r189_c160 bl_160 br_160 wl_189 vdd gnd cell_6t
Xbit_r190_c160 bl_160 br_160 wl_190 vdd gnd cell_6t
Xbit_r191_c160 bl_160 br_160 wl_191 vdd gnd cell_6t
Xbit_r192_c160 bl_160 br_160 wl_192 vdd gnd cell_6t
Xbit_r193_c160 bl_160 br_160 wl_193 vdd gnd cell_6t
Xbit_r194_c160 bl_160 br_160 wl_194 vdd gnd cell_6t
Xbit_r195_c160 bl_160 br_160 wl_195 vdd gnd cell_6t
Xbit_r196_c160 bl_160 br_160 wl_196 vdd gnd cell_6t
Xbit_r197_c160 bl_160 br_160 wl_197 vdd gnd cell_6t
Xbit_r198_c160 bl_160 br_160 wl_198 vdd gnd cell_6t
Xbit_r199_c160 bl_160 br_160 wl_199 vdd gnd cell_6t
Xbit_r200_c160 bl_160 br_160 wl_200 vdd gnd cell_6t
Xbit_r201_c160 bl_160 br_160 wl_201 vdd gnd cell_6t
Xbit_r202_c160 bl_160 br_160 wl_202 vdd gnd cell_6t
Xbit_r203_c160 bl_160 br_160 wl_203 vdd gnd cell_6t
Xbit_r204_c160 bl_160 br_160 wl_204 vdd gnd cell_6t
Xbit_r205_c160 bl_160 br_160 wl_205 vdd gnd cell_6t
Xbit_r206_c160 bl_160 br_160 wl_206 vdd gnd cell_6t
Xbit_r207_c160 bl_160 br_160 wl_207 vdd gnd cell_6t
Xbit_r208_c160 bl_160 br_160 wl_208 vdd gnd cell_6t
Xbit_r209_c160 bl_160 br_160 wl_209 vdd gnd cell_6t
Xbit_r210_c160 bl_160 br_160 wl_210 vdd gnd cell_6t
Xbit_r211_c160 bl_160 br_160 wl_211 vdd gnd cell_6t
Xbit_r212_c160 bl_160 br_160 wl_212 vdd gnd cell_6t
Xbit_r213_c160 bl_160 br_160 wl_213 vdd gnd cell_6t
Xbit_r214_c160 bl_160 br_160 wl_214 vdd gnd cell_6t
Xbit_r215_c160 bl_160 br_160 wl_215 vdd gnd cell_6t
Xbit_r216_c160 bl_160 br_160 wl_216 vdd gnd cell_6t
Xbit_r217_c160 bl_160 br_160 wl_217 vdd gnd cell_6t
Xbit_r218_c160 bl_160 br_160 wl_218 vdd gnd cell_6t
Xbit_r219_c160 bl_160 br_160 wl_219 vdd gnd cell_6t
Xbit_r220_c160 bl_160 br_160 wl_220 vdd gnd cell_6t
Xbit_r221_c160 bl_160 br_160 wl_221 vdd gnd cell_6t
Xbit_r222_c160 bl_160 br_160 wl_222 vdd gnd cell_6t
Xbit_r223_c160 bl_160 br_160 wl_223 vdd gnd cell_6t
Xbit_r224_c160 bl_160 br_160 wl_224 vdd gnd cell_6t
Xbit_r225_c160 bl_160 br_160 wl_225 vdd gnd cell_6t
Xbit_r226_c160 bl_160 br_160 wl_226 vdd gnd cell_6t
Xbit_r227_c160 bl_160 br_160 wl_227 vdd gnd cell_6t
Xbit_r228_c160 bl_160 br_160 wl_228 vdd gnd cell_6t
Xbit_r229_c160 bl_160 br_160 wl_229 vdd gnd cell_6t
Xbit_r230_c160 bl_160 br_160 wl_230 vdd gnd cell_6t
Xbit_r231_c160 bl_160 br_160 wl_231 vdd gnd cell_6t
Xbit_r232_c160 bl_160 br_160 wl_232 vdd gnd cell_6t
Xbit_r233_c160 bl_160 br_160 wl_233 vdd gnd cell_6t
Xbit_r234_c160 bl_160 br_160 wl_234 vdd gnd cell_6t
Xbit_r235_c160 bl_160 br_160 wl_235 vdd gnd cell_6t
Xbit_r236_c160 bl_160 br_160 wl_236 vdd gnd cell_6t
Xbit_r237_c160 bl_160 br_160 wl_237 vdd gnd cell_6t
Xbit_r238_c160 bl_160 br_160 wl_238 vdd gnd cell_6t
Xbit_r239_c160 bl_160 br_160 wl_239 vdd gnd cell_6t
Xbit_r240_c160 bl_160 br_160 wl_240 vdd gnd cell_6t
Xbit_r241_c160 bl_160 br_160 wl_241 vdd gnd cell_6t
Xbit_r242_c160 bl_160 br_160 wl_242 vdd gnd cell_6t
Xbit_r243_c160 bl_160 br_160 wl_243 vdd gnd cell_6t
Xbit_r244_c160 bl_160 br_160 wl_244 vdd gnd cell_6t
Xbit_r245_c160 bl_160 br_160 wl_245 vdd gnd cell_6t
Xbit_r246_c160 bl_160 br_160 wl_246 vdd gnd cell_6t
Xbit_r247_c160 bl_160 br_160 wl_247 vdd gnd cell_6t
Xbit_r248_c160 bl_160 br_160 wl_248 vdd gnd cell_6t
Xbit_r249_c160 bl_160 br_160 wl_249 vdd gnd cell_6t
Xbit_r250_c160 bl_160 br_160 wl_250 vdd gnd cell_6t
Xbit_r251_c160 bl_160 br_160 wl_251 vdd gnd cell_6t
Xbit_r252_c160 bl_160 br_160 wl_252 vdd gnd cell_6t
Xbit_r253_c160 bl_160 br_160 wl_253 vdd gnd cell_6t
Xbit_r254_c160 bl_160 br_160 wl_254 vdd gnd cell_6t
Xbit_r255_c160 bl_160 br_160 wl_255 vdd gnd cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd cell_6t
Xbit_r1_c161 bl_161 br_161 wl_1 vdd gnd cell_6t
Xbit_r2_c161 bl_161 br_161 wl_2 vdd gnd cell_6t
Xbit_r3_c161 bl_161 br_161 wl_3 vdd gnd cell_6t
Xbit_r4_c161 bl_161 br_161 wl_4 vdd gnd cell_6t
Xbit_r5_c161 bl_161 br_161 wl_5 vdd gnd cell_6t
Xbit_r6_c161 bl_161 br_161 wl_6 vdd gnd cell_6t
Xbit_r7_c161 bl_161 br_161 wl_7 vdd gnd cell_6t
Xbit_r8_c161 bl_161 br_161 wl_8 vdd gnd cell_6t
Xbit_r9_c161 bl_161 br_161 wl_9 vdd gnd cell_6t
Xbit_r10_c161 bl_161 br_161 wl_10 vdd gnd cell_6t
Xbit_r11_c161 bl_161 br_161 wl_11 vdd gnd cell_6t
Xbit_r12_c161 bl_161 br_161 wl_12 vdd gnd cell_6t
Xbit_r13_c161 bl_161 br_161 wl_13 vdd gnd cell_6t
Xbit_r14_c161 bl_161 br_161 wl_14 vdd gnd cell_6t
Xbit_r15_c161 bl_161 br_161 wl_15 vdd gnd cell_6t
Xbit_r16_c161 bl_161 br_161 wl_16 vdd gnd cell_6t
Xbit_r17_c161 bl_161 br_161 wl_17 vdd gnd cell_6t
Xbit_r18_c161 bl_161 br_161 wl_18 vdd gnd cell_6t
Xbit_r19_c161 bl_161 br_161 wl_19 vdd gnd cell_6t
Xbit_r20_c161 bl_161 br_161 wl_20 vdd gnd cell_6t
Xbit_r21_c161 bl_161 br_161 wl_21 vdd gnd cell_6t
Xbit_r22_c161 bl_161 br_161 wl_22 vdd gnd cell_6t
Xbit_r23_c161 bl_161 br_161 wl_23 vdd gnd cell_6t
Xbit_r24_c161 bl_161 br_161 wl_24 vdd gnd cell_6t
Xbit_r25_c161 bl_161 br_161 wl_25 vdd gnd cell_6t
Xbit_r26_c161 bl_161 br_161 wl_26 vdd gnd cell_6t
Xbit_r27_c161 bl_161 br_161 wl_27 vdd gnd cell_6t
Xbit_r28_c161 bl_161 br_161 wl_28 vdd gnd cell_6t
Xbit_r29_c161 bl_161 br_161 wl_29 vdd gnd cell_6t
Xbit_r30_c161 bl_161 br_161 wl_30 vdd gnd cell_6t
Xbit_r31_c161 bl_161 br_161 wl_31 vdd gnd cell_6t
Xbit_r32_c161 bl_161 br_161 wl_32 vdd gnd cell_6t
Xbit_r33_c161 bl_161 br_161 wl_33 vdd gnd cell_6t
Xbit_r34_c161 bl_161 br_161 wl_34 vdd gnd cell_6t
Xbit_r35_c161 bl_161 br_161 wl_35 vdd gnd cell_6t
Xbit_r36_c161 bl_161 br_161 wl_36 vdd gnd cell_6t
Xbit_r37_c161 bl_161 br_161 wl_37 vdd gnd cell_6t
Xbit_r38_c161 bl_161 br_161 wl_38 vdd gnd cell_6t
Xbit_r39_c161 bl_161 br_161 wl_39 vdd gnd cell_6t
Xbit_r40_c161 bl_161 br_161 wl_40 vdd gnd cell_6t
Xbit_r41_c161 bl_161 br_161 wl_41 vdd gnd cell_6t
Xbit_r42_c161 bl_161 br_161 wl_42 vdd gnd cell_6t
Xbit_r43_c161 bl_161 br_161 wl_43 vdd gnd cell_6t
Xbit_r44_c161 bl_161 br_161 wl_44 vdd gnd cell_6t
Xbit_r45_c161 bl_161 br_161 wl_45 vdd gnd cell_6t
Xbit_r46_c161 bl_161 br_161 wl_46 vdd gnd cell_6t
Xbit_r47_c161 bl_161 br_161 wl_47 vdd gnd cell_6t
Xbit_r48_c161 bl_161 br_161 wl_48 vdd gnd cell_6t
Xbit_r49_c161 bl_161 br_161 wl_49 vdd gnd cell_6t
Xbit_r50_c161 bl_161 br_161 wl_50 vdd gnd cell_6t
Xbit_r51_c161 bl_161 br_161 wl_51 vdd gnd cell_6t
Xbit_r52_c161 bl_161 br_161 wl_52 vdd gnd cell_6t
Xbit_r53_c161 bl_161 br_161 wl_53 vdd gnd cell_6t
Xbit_r54_c161 bl_161 br_161 wl_54 vdd gnd cell_6t
Xbit_r55_c161 bl_161 br_161 wl_55 vdd gnd cell_6t
Xbit_r56_c161 bl_161 br_161 wl_56 vdd gnd cell_6t
Xbit_r57_c161 bl_161 br_161 wl_57 vdd gnd cell_6t
Xbit_r58_c161 bl_161 br_161 wl_58 vdd gnd cell_6t
Xbit_r59_c161 bl_161 br_161 wl_59 vdd gnd cell_6t
Xbit_r60_c161 bl_161 br_161 wl_60 vdd gnd cell_6t
Xbit_r61_c161 bl_161 br_161 wl_61 vdd gnd cell_6t
Xbit_r62_c161 bl_161 br_161 wl_62 vdd gnd cell_6t
Xbit_r63_c161 bl_161 br_161 wl_63 vdd gnd cell_6t
Xbit_r64_c161 bl_161 br_161 wl_64 vdd gnd cell_6t
Xbit_r65_c161 bl_161 br_161 wl_65 vdd gnd cell_6t
Xbit_r66_c161 bl_161 br_161 wl_66 vdd gnd cell_6t
Xbit_r67_c161 bl_161 br_161 wl_67 vdd gnd cell_6t
Xbit_r68_c161 bl_161 br_161 wl_68 vdd gnd cell_6t
Xbit_r69_c161 bl_161 br_161 wl_69 vdd gnd cell_6t
Xbit_r70_c161 bl_161 br_161 wl_70 vdd gnd cell_6t
Xbit_r71_c161 bl_161 br_161 wl_71 vdd gnd cell_6t
Xbit_r72_c161 bl_161 br_161 wl_72 vdd gnd cell_6t
Xbit_r73_c161 bl_161 br_161 wl_73 vdd gnd cell_6t
Xbit_r74_c161 bl_161 br_161 wl_74 vdd gnd cell_6t
Xbit_r75_c161 bl_161 br_161 wl_75 vdd gnd cell_6t
Xbit_r76_c161 bl_161 br_161 wl_76 vdd gnd cell_6t
Xbit_r77_c161 bl_161 br_161 wl_77 vdd gnd cell_6t
Xbit_r78_c161 bl_161 br_161 wl_78 vdd gnd cell_6t
Xbit_r79_c161 bl_161 br_161 wl_79 vdd gnd cell_6t
Xbit_r80_c161 bl_161 br_161 wl_80 vdd gnd cell_6t
Xbit_r81_c161 bl_161 br_161 wl_81 vdd gnd cell_6t
Xbit_r82_c161 bl_161 br_161 wl_82 vdd gnd cell_6t
Xbit_r83_c161 bl_161 br_161 wl_83 vdd gnd cell_6t
Xbit_r84_c161 bl_161 br_161 wl_84 vdd gnd cell_6t
Xbit_r85_c161 bl_161 br_161 wl_85 vdd gnd cell_6t
Xbit_r86_c161 bl_161 br_161 wl_86 vdd gnd cell_6t
Xbit_r87_c161 bl_161 br_161 wl_87 vdd gnd cell_6t
Xbit_r88_c161 bl_161 br_161 wl_88 vdd gnd cell_6t
Xbit_r89_c161 bl_161 br_161 wl_89 vdd gnd cell_6t
Xbit_r90_c161 bl_161 br_161 wl_90 vdd gnd cell_6t
Xbit_r91_c161 bl_161 br_161 wl_91 vdd gnd cell_6t
Xbit_r92_c161 bl_161 br_161 wl_92 vdd gnd cell_6t
Xbit_r93_c161 bl_161 br_161 wl_93 vdd gnd cell_6t
Xbit_r94_c161 bl_161 br_161 wl_94 vdd gnd cell_6t
Xbit_r95_c161 bl_161 br_161 wl_95 vdd gnd cell_6t
Xbit_r96_c161 bl_161 br_161 wl_96 vdd gnd cell_6t
Xbit_r97_c161 bl_161 br_161 wl_97 vdd gnd cell_6t
Xbit_r98_c161 bl_161 br_161 wl_98 vdd gnd cell_6t
Xbit_r99_c161 bl_161 br_161 wl_99 vdd gnd cell_6t
Xbit_r100_c161 bl_161 br_161 wl_100 vdd gnd cell_6t
Xbit_r101_c161 bl_161 br_161 wl_101 vdd gnd cell_6t
Xbit_r102_c161 bl_161 br_161 wl_102 vdd gnd cell_6t
Xbit_r103_c161 bl_161 br_161 wl_103 vdd gnd cell_6t
Xbit_r104_c161 bl_161 br_161 wl_104 vdd gnd cell_6t
Xbit_r105_c161 bl_161 br_161 wl_105 vdd gnd cell_6t
Xbit_r106_c161 bl_161 br_161 wl_106 vdd gnd cell_6t
Xbit_r107_c161 bl_161 br_161 wl_107 vdd gnd cell_6t
Xbit_r108_c161 bl_161 br_161 wl_108 vdd gnd cell_6t
Xbit_r109_c161 bl_161 br_161 wl_109 vdd gnd cell_6t
Xbit_r110_c161 bl_161 br_161 wl_110 vdd gnd cell_6t
Xbit_r111_c161 bl_161 br_161 wl_111 vdd gnd cell_6t
Xbit_r112_c161 bl_161 br_161 wl_112 vdd gnd cell_6t
Xbit_r113_c161 bl_161 br_161 wl_113 vdd gnd cell_6t
Xbit_r114_c161 bl_161 br_161 wl_114 vdd gnd cell_6t
Xbit_r115_c161 bl_161 br_161 wl_115 vdd gnd cell_6t
Xbit_r116_c161 bl_161 br_161 wl_116 vdd gnd cell_6t
Xbit_r117_c161 bl_161 br_161 wl_117 vdd gnd cell_6t
Xbit_r118_c161 bl_161 br_161 wl_118 vdd gnd cell_6t
Xbit_r119_c161 bl_161 br_161 wl_119 vdd gnd cell_6t
Xbit_r120_c161 bl_161 br_161 wl_120 vdd gnd cell_6t
Xbit_r121_c161 bl_161 br_161 wl_121 vdd gnd cell_6t
Xbit_r122_c161 bl_161 br_161 wl_122 vdd gnd cell_6t
Xbit_r123_c161 bl_161 br_161 wl_123 vdd gnd cell_6t
Xbit_r124_c161 bl_161 br_161 wl_124 vdd gnd cell_6t
Xbit_r125_c161 bl_161 br_161 wl_125 vdd gnd cell_6t
Xbit_r126_c161 bl_161 br_161 wl_126 vdd gnd cell_6t
Xbit_r127_c161 bl_161 br_161 wl_127 vdd gnd cell_6t
Xbit_r128_c161 bl_161 br_161 wl_128 vdd gnd cell_6t
Xbit_r129_c161 bl_161 br_161 wl_129 vdd gnd cell_6t
Xbit_r130_c161 bl_161 br_161 wl_130 vdd gnd cell_6t
Xbit_r131_c161 bl_161 br_161 wl_131 vdd gnd cell_6t
Xbit_r132_c161 bl_161 br_161 wl_132 vdd gnd cell_6t
Xbit_r133_c161 bl_161 br_161 wl_133 vdd gnd cell_6t
Xbit_r134_c161 bl_161 br_161 wl_134 vdd gnd cell_6t
Xbit_r135_c161 bl_161 br_161 wl_135 vdd gnd cell_6t
Xbit_r136_c161 bl_161 br_161 wl_136 vdd gnd cell_6t
Xbit_r137_c161 bl_161 br_161 wl_137 vdd gnd cell_6t
Xbit_r138_c161 bl_161 br_161 wl_138 vdd gnd cell_6t
Xbit_r139_c161 bl_161 br_161 wl_139 vdd gnd cell_6t
Xbit_r140_c161 bl_161 br_161 wl_140 vdd gnd cell_6t
Xbit_r141_c161 bl_161 br_161 wl_141 vdd gnd cell_6t
Xbit_r142_c161 bl_161 br_161 wl_142 vdd gnd cell_6t
Xbit_r143_c161 bl_161 br_161 wl_143 vdd gnd cell_6t
Xbit_r144_c161 bl_161 br_161 wl_144 vdd gnd cell_6t
Xbit_r145_c161 bl_161 br_161 wl_145 vdd gnd cell_6t
Xbit_r146_c161 bl_161 br_161 wl_146 vdd gnd cell_6t
Xbit_r147_c161 bl_161 br_161 wl_147 vdd gnd cell_6t
Xbit_r148_c161 bl_161 br_161 wl_148 vdd gnd cell_6t
Xbit_r149_c161 bl_161 br_161 wl_149 vdd gnd cell_6t
Xbit_r150_c161 bl_161 br_161 wl_150 vdd gnd cell_6t
Xbit_r151_c161 bl_161 br_161 wl_151 vdd gnd cell_6t
Xbit_r152_c161 bl_161 br_161 wl_152 vdd gnd cell_6t
Xbit_r153_c161 bl_161 br_161 wl_153 vdd gnd cell_6t
Xbit_r154_c161 bl_161 br_161 wl_154 vdd gnd cell_6t
Xbit_r155_c161 bl_161 br_161 wl_155 vdd gnd cell_6t
Xbit_r156_c161 bl_161 br_161 wl_156 vdd gnd cell_6t
Xbit_r157_c161 bl_161 br_161 wl_157 vdd gnd cell_6t
Xbit_r158_c161 bl_161 br_161 wl_158 vdd gnd cell_6t
Xbit_r159_c161 bl_161 br_161 wl_159 vdd gnd cell_6t
Xbit_r160_c161 bl_161 br_161 wl_160 vdd gnd cell_6t
Xbit_r161_c161 bl_161 br_161 wl_161 vdd gnd cell_6t
Xbit_r162_c161 bl_161 br_161 wl_162 vdd gnd cell_6t
Xbit_r163_c161 bl_161 br_161 wl_163 vdd gnd cell_6t
Xbit_r164_c161 bl_161 br_161 wl_164 vdd gnd cell_6t
Xbit_r165_c161 bl_161 br_161 wl_165 vdd gnd cell_6t
Xbit_r166_c161 bl_161 br_161 wl_166 vdd gnd cell_6t
Xbit_r167_c161 bl_161 br_161 wl_167 vdd gnd cell_6t
Xbit_r168_c161 bl_161 br_161 wl_168 vdd gnd cell_6t
Xbit_r169_c161 bl_161 br_161 wl_169 vdd gnd cell_6t
Xbit_r170_c161 bl_161 br_161 wl_170 vdd gnd cell_6t
Xbit_r171_c161 bl_161 br_161 wl_171 vdd gnd cell_6t
Xbit_r172_c161 bl_161 br_161 wl_172 vdd gnd cell_6t
Xbit_r173_c161 bl_161 br_161 wl_173 vdd gnd cell_6t
Xbit_r174_c161 bl_161 br_161 wl_174 vdd gnd cell_6t
Xbit_r175_c161 bl_161 br_161 wl_175 vdd gnd cell_6t
Xbit_r176_c161 bl_161 br_161 wl_176 vdd gnd cell_6t
Xbit_r177_c161 bl_161 br_161 wl_177 vdd gnd cell_6t
Xbit_r178_c161 bl_161 br_161 wl_178 vdd gnd cell_6t
Xbit_r179_c161 bl_161 br_161 wl_179 vdd gnd cell_6t
Xbit_r180_c161 bl_161 br_161 wl_180 vdd gnd cell_6t
Xbit_r181_c161 bl_161 br_161 wl_181 vdd gnd cell_6t
Xbit_r182_c161 bl_161 br_161 wl_182 vdd gnd cell_6t
Xbit_r183_c161 bl_161 br_161 wl_183 vdd gnd cell_6t
Xbit_r184_c161 bl_161 br_161 wl_184 vdd gnd cell_6t
Xbit_r185_c161 bl_161 br_161 wl_185 vdd gnd cell_6t
Xbit_r186_c161 bl_161 br_161 wl_186 vdd gnd cell_6t
Xbit_r187_c161 bl_161 br_161 wl_187 vdd gnd cell_6t
Xbit_r188_c161 bl_161 br_161 wl_188 vdd gnd cell_6t
Xbit_r189_c161 bl_161 br_161 wl_189 vdd gnd cell_6t
Xbit_r190_c161 bl_161 br_161 wl_190 vdd gnd cell_6t
Xbit_r191_c161 bl_161 br_161 wl_191 vdd gnd cell_6t
Xbit_r192_c161 bl_161 br_161 wl_192 vdd gnd cell_6t
Xbit_r193_c161 bl_161 br_161 wl_193 vdd gnd cell_6t
Xbit_r194_c161 bl_161 br_161 wl_194 vdd gnd cell_6t
Xbit_r195_c161 bl_161 br_161 wl_195 vdd gnd cell_6t
Xbit_r196_c161 bl_161 br_161 wl_196 vdd gnd cell_6t
Xbit_r197_c161 bl_161 br_161 wl_197 vdd gnd cell_6t
Xbit_r198_c161 bl_161 br_161 wl_198 vdd gnd cell_6t
Xbit_r199_c161 bl_161 br_161 wl_199 vdd gnd cell_6t
Xbit_r200_c161 bl_161 br_161 wl_200 vdd gnd cell_6t
Xbit_r201_c161 bl_161 br_161 wl_201 vdd gnd cell_6t
Xbit_r202_c161 bl_161 br_161 wl_202 vdd gnd cell_6t
Xbit_r203_c161 bl_161 br_161 wl_203 vdd gnd cell_6t
Xbit_r204_c161 bl_161 br_161 wl_204 vdd gnd cell_6t
Xbit_r205_c161 bl_161 br_161 wl_205 vdd gnd cell_6t
Xbit_r206_c161 bl_161 br_161 wl_206 vdd gnd cell_6t
Xbit_r207_c161 bl_161 br_161 wl_207 vdd gnd cell_6t
Xbit_r208_c161 bl_161 br_161 wl_208 vdd gnd cell_6t
Xbit_r209_c161 bl_161 br_161 wl_209 vdd gnd cell_6t
Xbit_r210_c161 bl_161 br_161 wl_210 vdd gnd cell_6t
Xbit_r211_c161 bl_161 br_161 wl_211 vdd gnd cell_6t
Xbit_r212_c161 bl_161 br_161 wl_212 vdd gnd cell_6t
Xbit_r213_c161 bl_161 br_161 wl_213 vdd gnd cell_6t
Xbit_r214_c161 bl_161 br_161 wl_214 vdd gnd cell_6t
Xbit_r215_c161 bl_161 br_161 wl_215 vdd gnd cell_6t
Xbit_r216_c161 bl_161 br_161 wl_216 vdd gnd cell_6t
Xbit_r217_c161 bl_161 br_161 wl_217 vdd gnd cell_6t
Xbit_r218_c161 bl_161 br_161 wl_218 vdd gnd cell_6t
Xbit_r219_c161 bl_161 br_161 wl_219 vdd gnd cell_6t
Xbit_r220_c161 bl_161 br_161 wl_220 vdd gnd cell_6t
Xbit_r221_c161 bl_161 br_161 wl_221 vdd gnd cell_6t
Xbit_r222_c161 bl_161 br_161 wl_222 vdd gnd cell_6t
Xbit_r223_c161 bl_161 br_161 wl_223 vdd gnd cell_6t
Xbit_r224_c161 bl_161 br_161 wl_224 vdd gnd cell_6t
Xbit_r225_c161 bl_161 br_161 wl_225 vdd gnd cell_6t
Xbit_r226_c161 bl_161 br_161 wl_226 vdd gnd cell_6t
Xbit_r227_c161 bl_161 br_161 wl_227 vdd gnd cell_6t
Xbit_r228_c161 bl_161 br_161 wl_228 vdd gnd cell_6t
Xbit_r229_c161 bl_161 br_161 wl_229 vdd gnd cell_6t
Xbit_r230_c161 bl_161 br_161 wl_230 vdd gnd cell_6t
Xbit_r231_c161 bl_161 br_161 wl_231 vdd gnd cell_6t
Xbit_r232_c161 bl_161 br_161 wl_232 vdd gnd cell_6t
Xbit_r233_c161 bl_161 br_161 wl_233 vdd gnd cell_6t
Xbit_r234_c161 bl_161 br_161 wl_234 vdd gnd cell_6t
Xbit_r235_c161 bl_161 br_161 wl_235 vdd gnd cell_6t
Xbit_r236_c161 bl_161 br_161 wl_236 vdd gnd cell_6t
Xbit_r237_c161 bl_161 br_161 wl_237 vdd gnd cell_6t
Xbit_r238_c161 bl_161 br_161 wl_238 vdd gnd cell_6t
Xbit_r239_c161 bl_161 br_161 wl_239 vdd gnd cell_6t
Xbit_r240_c161 bl_161 br_161 wl_240 vdd gnd cell_6t
Xbit_r241_c161 bl_161 br_161 wl_241 vdd gnd cell_6t
Xbit_r242_c161 bl_161 br_161 wl_242 vdd gnd cell_6t
Xbit_r243_c161 bl_161 br_161 wl_243 vdd gnd cell_6t
Xbit_r244_c161 bl_161 br_161 wl_244 vdd gnd cell_6t
Xbit_r245_c161 bl_161 br_161 wl_245 vdd gnd cell_6t
Xbit_r246_c161 bl_161 br_161 wl_246 vdd gnd cell_6t
Xbit_r247_c161 bl_161 br_161 wl_247 vdd gnd cell_6t
Xbit_r248_c161 bl_161 br_161 wl_248 vdd gnd cell_6t
Xbit_r249_c161 bl_161 br_161 wl_249 vdd gnd cell_6t
Xbit_r250_c161 bl_161 br_161 wl_250 vdd gnd cell_6t
Xbit_r251_c161 bl_161 br_161 wl_251 vdd gnd cell_6t
Xbit_r252_c161 bl_161 br_161 wl_252 vdd gnd cell_6t
Xbit_r253_c161 bl_161 br_161 wl_253 vdd gnd cell_6t
Xbit_r254_c161 bl_161 br_161 wl_254 vdd gnd cell_6t
Xbit_r255_c161 bl_161 br_161 wl_255 vdd gnd cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd cell_6t
Xbit_r1_c162 bl_162 br_162 wl_1 vdd gnd cell_6t
Xbit_r2_c162 bl_162 br_162 wl_2 vdd gnd cell_6t
Xbit_r3_c162 bl_162 br_162 wl_3 vdd gnd cell_6t
Xbit_r4_c162 bl_162 br_162 wl_4 vdd gnd cell_6t
Xbit_r5_c162 bl_162 br_162 wl_5 vdd gnd cell_6t
Xbit_r6_c162 bl_162 br_162 wl_6 vdd gnd cell_6t
Xbit_r7_c162 bl_162 br_162 wl_7 vdd gnd cell_6t
Xbit_r8_c162 bl_162 br_162 wl_8 vdd gnd cell_6t
Xbit_r9_c162 bl_162 br_162 wl_9 vdd gnd cell_6t
Xbit_r10_c162 bl_162 br_162 wl_10 vdd gnd cell_6t
Xbit_r11_c162 bl_162 br_162 wl_11 vdd gnd cell_6t
Xbit_r12_c162 bl_162 br_162 wl_12 vdd gnd cell_6t
Xbit_r13_c162 bl_162 br_162 wl_13 vdd gnd cell_6t
Xbit_r14_c162 bl_162 br_162 wl_14 vdd gnd cell_6t
Xbit_r15_c162 bl_162 br_162 wl_15 vdd gnd cell_6t
Xbit_r16_c162 bl_162 br_162 wl_16 vdd gnd cell_6t
Xbit_r17_c162 bl_162 br_162 wl_17 vdd gnd cell_6t
Xbit_r18_c162 bl_162 br_162 wl_18 vdd gnd cell_6t
Xbit_r19_c162 bl_162 br_162 wl_19 vdd gnd cell_6t
Xbit_r20_c162 bl_162 br_162 wl_20 vdd gnd cell_6t
Xbit_r21_c162 bl_162 br_162 wl_21 vdd gnd cell_6t
Xbit_r22_c162 bl_162 br_162 wl_22 vdd gnd cell_6t
Xbit_r23_c162 bl_162 br_162 wl_23 vdd gnd cell_6t
Xbit_r24_c162 bl_162 br_162 wl_24 vdd gnd cell_6t
Xbit_r25_c162 bl_162 br_162 wl_25 vdd gnd cell_6t
Xbit_r26_c162 bl_162 br_162 wl_26 vdd gnd cell_6t
Xbit_r27_c162 bl_162 br_162 wl_27 vdd gnd cell_6t
Xbit_r28_c162 bl_162 br_162 wl_28 vdd gnd cell_6t
Xbit_r29_c162 bl_162 br_162 wl_29 vdd gnd cell_6t
Xbit_r30_c162 bl_162 br_162 wl_30 vdd gnd cell_6t
Xbit_r31_c162 bl_162 br_162 wl_31 vdd gnd cell_6t
Xbit_r32_c162 bl_162 br_162 wl_32 vdd gnd cell_6t
Xbit_r33_c162 bl_162 br_162 wl_33 vdd gnd cell_6t
Xbit_r34_c162 bl_162 br_162 wl_34 vdd gnd cell_6t
Xbit_r35_c162 bl_162 br_162 wl_35 vdd gnd cell_6t
Xbit_r36_c162 bl_162 br_162 wl_36 vdd gnd cell_6t
Xbit_r37_c162 bl_162 br_162 wl_37 vdd gnd cell_6t
Xbit_r38_c162 bl_162 br_162 wl_38 vdd gnd cell_6t
Xbit_r39_c162 bl_162 br_162 wl_39 vdd gnd cell_6t
Xbit_r40_c162 bl_162 br_162 wl_40 vdd gnd cell_6t
Xbit_r41_c162 bl_162 br_162 wl_41 vdd gnd cell_6t
Xbit_r42_c162 bl_162 br_162 wl_42 vdd gnd cell_6t
Xbit_r43_c162 bl_162 br_162 wl_43 vdd gnd cell_6t
Xbit_r44_c162 bl_162 br_162 wl_44 vdd gnd cell_6t
Xbit_r45_c162 bl_162 br_162 wl_45 vdd gnd cell_6t
Xbit_r46_c162 bl_162 br_162 wl_46 vdd gnd cell_6t
Xbit_r47_c162 bl_162 br_162 wl_47 vdd gnd cell_6t
Xbit_r48_c162 bl_162 br_162 wl_48 vdd gnd cell_6t
Xbit_r49_c162 bl_162 br_162 wl_49 vdd gnd cell_6t
Xbit_r50_c162 bl_162 br_162 wl_50 vdd gnd cell_6t
Xbit_r51_c162 bl_162 br_162 wl_51 vdd gnd cell_6t
Xbit_r52_c162 bl_162 br_162 wl_52 vdd gnd cell_6t
Xbit_r53_c162 bl_162 br_162 wl_53 vdd gnd cell_6t
Xbit_r54_c162 bl_162 br_162 wl_54 vdd gnd cell_6t
Xbit_r55_c162 bl_162 br_162 wl_55 vdd gnd cell_6t
Xbit_r56_c162 bl_162 br_162 wl_56 vdd gnd cell_6t
Xbit_r57_c162 bl_162 br_162 wl_57 vdd gnd cell_6t
Xbit_r58_c162 bl_162 br_162 wl_58 vdd gnd cell_6t
Xbit_r59_c162 bl_162 br_162 wl_59 vdd gnd cell_6t
Xbit_r60_c162 bl_162 br_162 wl_60 vdd gnd cell_6t
Xbit_r61_c162 bl_162 br_162 wl_61 vdd gnd cell_6t
Xbit_r62_c162 bl_162 br_162 wl_62 vdd gnd cell_6t
Xbit_r63_c162 bl_162 br_162 wl_63 vdd gnd cell_6t
Xbit_r64_c162 bl_162 br_162 wl_64 vdd gnd cell_6t
Xbit_r65_c162 bl_162 br_162 wl_65 vdd gnd cell_6t
Xbit_r66_c162 bl_162 br_162 wl_66 vdd gnd cell_6t
Xbit_r67_c162 bl_162 br_162 wl_67 vdd gnd cell_6t
Xbit_r68_c162 bl_162 br_162 wl_68 vdd gnd cell_6t
Xbit_r69_c162 bl_162 br_162 wl_69 vdd gnd cell_6t
Xbit_r70_c162 bl_162 br_162 wl_70 vdd gnd cell_6t
Xbit_r71_c162 bl_162 br_162 wl_71 vdd gnd cell_6t
Xbit_r72_c162 bl_162 br_162 wl_72 vdd gnd cell_6t
Xbit_r73_c162 bl_162 br_162 wl_73 vdd gnd cell_6t
Xbit_r74_c162 bl_162 br_162 wl_74 vdd gnd cell_6t
Xbit_r75_c162 bl_162 br_162 wl_75 vdd gnd cell_6t
Xbit_r76_c162 bl_162 br_162 wl_76 vdd gnd cell_6t
Xbit_r77_c162 bl_162 br_162 wl_77 vdd gnd cell_6t
Xbit_r78_c162 bl_162 br_162 wl_78 vdd gnd cell_6t
Xbit_r79_c162 bl_162 br_162 wl_79 vdd gnd cell_6t
Xbit_r80_c162 bl_162 br_162 wl_80 vdd gnd cell_6t
Xbit_r81_c162 bl_162 br_162 wl_81 vdd gnd cell_6t
Xbit_r82_c162 bl_162 br_162 wl_82 vdd gnd cell_6t
Xbit_r83_c162 bl_162 br_162 wl_83 vdd gnd cell_6t
Xbit_r84_c162 bl_162 br_162 wl_84 vdd gnd cell_6t
Xbit_r85_c162 bl_162 br_162 wl_85 vdd gnd cell_6t
Xbit_r86_c162 bl_162 br_162 wl_86 vdd gnd cell_6t
Xbit_r87_c162 bl_162 br_162 wl_87 vdd gnd cell_6t
Xbit_r88_c162 bl_162 br_162 wl_88 vdd gnd cell_6t
Xbit_r89_c162 bl_162 br_162 wl_89 vdd gnd cell_6t
Xbit_r90_c162 bl_162 br_162 wl_90 vdd gnd cell_6t
Xbit_r91_c162 bl_162 br_162 wl_91 vdd gnd cell_6t
Xbit_r92_c162 bl_162 br_162 wl_92 vdd gnd cell_6t
Xbit_r93_c162 bl_162 br_162 wl_93 vdd gnd cell_6t
Xbit_r94_c162 bl_162 br_162 wl_94 vdd gnd cell_6t
Xbit_r95_c162 bl_162 br_162 wl_95 vdd gnd cell_6t
Xbit_r96_c162 bl_162 br_162 wl_96 vdd gnd cell_6t
Xbit_r97_c162 bl_162 br_162 wl_97 vdd gnd cell_6t
Xbit_r98_c162 bl_162 br_162 wl_98 vdd gnd cell_6t
Xbit_r99_c162 bl_162 br_162 wl_99 vdd gnd cell_6t
Xbit_r100_c162 bl_162 br_162 wl_100 vdd gnd cell_6t
Xbit_r101_c162 bl_162 br_162 wl_101 vdd gnd cell_6t
Xbit_r102_c162 bl_162 br_162 wl_102 vdd gnd cell_6t
Xbit_r103_c162 bl_162 br_162 wl_103 vdd gnd cell_6t
Xbit_r104_c162 bl_162 br_162 wl_104 vdd gnd cell_6t
Xbit_r105_c162 bl_162 br_162 wl_105 vdd gnd cell_6t
Xbit_r106_c162 bl_162 br_162 wl_106 vdd gnd cell_6t
Xbit_r107_c162 bl_162 br_162 wl_107 vdd gnd cell_6t
Xbit_r108_c162 bl_162 br_162 wl_108 vdd gnd cell_6t
Xbit_r109_c162 bl_162 br_162 wl_109 vdd gnd cell_6t
Xbit_r110_c162 bl_162 br_162 wl_110 vdd gnd cell_6t
Xbit_r111_c162 bl_162 br_162 wl_111 vdd gnd cell_6t
Xbit_r112_c162 bl_162 br_162 wl_112 vdd gnd cell_6t
Xbit_r113_c162 bl_162 br_162 wl_113 vdd gnd cell_6t
Xbit_r114_c162 bl_162 br_162 wl_114 vdd gnd cell_6t
Xbit_r115_c162 bl_162 br_162 wl_115 vdd gnd cell_6t
Xbit_r116_c162 bl_162 br_162 wl_116 vdd gnd cell_6t
Xbit_r117_c162 bl_162 br_162 wl_117 vdd gnd cell_6t
Xbit_r118_c162 bl_162 br_162 wl_118 vdd gnd cell_6t
Xbit_r119_c162 bl_162 br_162 wl_119 vdd gnd cell_6t
Xbit_r120_c162 bl_162 br_162 wl_120 vdd gnd cell_6t
Xbit_r121_c162 bl_162 br_162 wl_121 vdd gnd cell_6t
Xbit_r122_c162 bl_162 br_162 wl_122 vdd gnd cell_6t
Xbit_r123_c162 bl_162 br_162 wl_123 vdd gnd cell_6t
Xbit_r124_c162 bl_162 br_162 wl_124 vdd gnd cell_6t
Xbit_r125_c162 bl_162 br_162 wl_125 vdd gnd cell_6t
Xbit_r126_c162 bl_162 br_162 wl_126 vdd gnd cell_6t
Xbit_r127_c162 bl_162 br_162 wl_127 vdd gnd cell_6t
Xbit_r128_c162 bl_162 br_162 wl_128 vdd gnd cell_6t
Xbit_r129_c162 bl_162 br_162 wl_129 vdd gnd cell_6t
Xbit_r130_c162 bl_162 br_162 wl_130 vdd gnd cell_6t
Xbit_r131_c162 bl_162 br_162 wl_131 vdd gnd cell_6t
Xbit_r132_c162 bl_162 br_162 wl_132 vdd gnd cell_6t
Xbit_r133_c162 bl_162 br_162 wl_133 vdd gnd cell_6t
Xbit_r134_c162 bl_162 br_162 wl_134 vdd gnd cell_6t
Xbit_r135_c162 bl_162 br_162 wl_135 vdd gnd cell_6t
Xbit_r136_c162 bl_162 br_162 wl_136 vdd gnd cell_6t
Xbit_r137_c162 bl_162 br_162 wl_137 vdd gnd cell_6t
Xbit_r138_c162 bl_162 br_162 wl_138 vdd gnd cell_6t
Xbit_r139_c162 bl_162 br_162 wl_139 vdd gnd cell_6t
Xbit_r140_c162 bl_162 br_162 wl_140 vdd gnd cell_6t
Xbit_r141_c162 bl_162 br_162 wl_141 vdd gnd cell_6t
Xbit_r142_c162 bl_162 br_162 wl_142 vdd gnd cell_6t
Xbit_r143_c162 bl_162 br_162 wl_143 vdd gnd cell_6t
Xbit_r144_c162 bl_162 br_162 wl_144 vdd gnd cell_6t
Xbit_r145_c162 bl_162 br_162 wl_145 vdd gnd cell_6t
Xbit_r146_c162 bl_162 br_162 wl_146 vdd gnd cell_6t
Xbit_r147_c162 bl_162 br_162 wl_147 vdd gnd cell_6t
Xbit_r148_c162 bl_162 br_162 wl_148 vdd gnd cell_6t
Xbit_r149_c162 bl_162 br_162 wl_149 vdd gnd cell_6t
Xbit_r150_c162 bl_162 br_162 wl_150 vdd gnd cell_6t
Xbit_r151_c162 bl_162 br_162 wl_151 vdd gnd cell_6t
Xbit_r152_c162 bl_162 br_162 wl_152 vdd gnd cell_6t
Xbit_r153_c162 bl_162 br_162 wl_153 vdd gnd cell_6t
Xbit_r154_c162 bl_162 br_162 wl_154 vdd gnd cell_6t
Xbit_r155_c162 bl_162 br_162 wl_155 vdd gnd cell_6t
Xbit_r156_c162 bl_162 br_162 wl_156 vdd gnd cell_6t
Xbit_r157_c162 bl_162 br_162 wl_157 vdd gnd cell_6t
Xbit_r158_c162 bl_162 br_162 wl_158 vdd gnd cell_6t
Xbit_r159_c162 bl_162 br_162 wl_159 vdd gnd cell_6t
Xbit_r160_c162 bl_162 br_162 wl_160 vdd gnd cell_6t
Xbit_r161_c162 bl_162 br_162 wl_161 vdd gnd cell_6t
Xbit_r162_c162 bl_162 br_162 wl_162 vdd gnd cell_6t
Xbit_r163_c162 bl_162 br_162 wl_163 vdd gnd cell_6t
Xbit_r164_c162 bl_162 br_162 wl_164 vdd gnd cell_6t
Xbit_r165_c162 bl_162 br_162 wl_165 vdd gnd cell_6t
Xbit_r166_c162 bl_162 br_162 wl_166 vdd gnd cell_6t
Xbit_r167_c162 bl_162 br_162 wl_167 vdd gnd cell_6t
Xbit_r168_c162 bl_162 br_162 wl_168 vdd gnd cell_6t
Xbit_r169_c162 bl_162 br_162 wl_169 vdd gnd cell_6t
Xbit_r170_c162 bl_162 br_162 wl_170 vdd gnd cell_6t
Xbit_r171_c162 bl_162 br_162 wl_171 vdd gnd cell_6t
Xbit_r172_c162 bl_162 br_162 wl_172 vdd gnd cell_6t
Xbit_r173_c162 bl_162 br_162 wl_173 vdd gnd cell_6t
Xbit_r174_c162 bl_162 br_162 wl_174 vdd gnd cell_6t
Xbit_r175_c162 bl_162 br_162 wl_175 vdd gnd cell_6t
Xbit_r176_c162 bl_162 br_162 wl_176 vdd gnd cell_6t
Xbit_r177_c162 bl_162 br_162 wl_177 vdd gnd cell_6t
Xbit_r178_c162 bl_162 br_162 wl_178 vdd gnd cell_6t
Xbit_r179_c162 bl_162 br_162 wl_179 vdd gnd cell_6t
Xbit_r180_c162 bl_162 br_162 wl_180 vdd gnd cell_6t
Xbit_r181_c162 bl_162 br_162 wl_181 vdd gnd cell_6t
Xbit_r182_c162 bl_162 br_162 wl_182 vdd gnd cell_6t
Xbit_r183_c162 bl_162 br_162 wl_183 vdd gnd cell_6t
Xbit_r184_c162 bl_162 br_162 wl_184 vdd gnd cell_6t
Xbit_r185_c162 bl_162 br_162 wl_185 vdd gnd cell_6t
Xbit_r186_c162 bl_162 br_162 wl_186 vdd gnd cell_6t
Xbit_r187_c162 bl_162 br_162 wl_187 vdd gnd cell_6t
Xbit_r188_c162 bl_162 br_162 wl_188 vdd gnd cell_6t
Xbit_r189_c162 bl_162 br_162 wl_189 vdd gnd cell_6t
Xbit_r190_c162 bl_162 br_162 wl_190 vdd gnd cell_6t
Xbit_r191_c162 bl_162 br_162 wl_191 vdd gnd cell_6t
Xbit_r192_c162 bl_162 br_162 wl_192 vdd gnd cell_6t
Xbit_r193_c162 bl_162 br_162 wl_193 vdd gnd cell_6t
Xbit_r194_c162 bl_162 br_162 wl_194 vdd gnd cell_6t
Xbit_r195_c162 bl_162 br_162 wl_195 vdd gnd cell_6t
Xbit_r196_c162 bl_162 br_162 wl_196 vdd gnd cell_6t
Xbit_r197_c162 bl_162 br_162 wl_197 vdd gnd cell_6t
Xbit_r198_c162 bl_162 br_162 wl_198 vdd gnd cell_6t
Xbit_r199_c162 bl_162 br_162 wl_199 vdd gnd cell_6t
Xbit_r200_c162 bl_162 br_162 wl_200 vdd gnd cell_6t
Xbit_r201_c162 bl_162 br_162 wl_201 vdd gnd cell_6t
Xbit_r202_c162 bl_162 br_162 wl_202 vdd gnd cell_6t
Xbit_r203_c162 bl_162 br_162 wl_203 vdd gnd cell_6t
Xbit_r204_c162 bl_162 br_162 wl_204 vdd gnd cell_6t
Xbit_r205_c162 bl_162 br_162 wl_205 vdd gnd cell_6t
Xbit_r206_c162 bl_162 br_162 wl_206 vdd gnd cell_6t
Xbit_r207_c162 bl_162 br_162 wl_207 vdd gnd cell_6t
Xbit_r208_c162 bl_162 br_162 wl_208 vdd gnd cell_6t
Xbit_r209_c162 bl_162 br_162 wl_209 vdd gnd cell_6t
Xbit_r210_c162 bl_162 br_162 wl_210 vdd gnd cell_6t
Xbit_r211_c162 bl_162 br_162 wl_211 vdd gnd cell_6t
Xbit_r212_c162 bl_162 br_162 wl_212 vdd gnd cell_6t
Xbit_r213_c162 bl_162 br_162 wl_213 vdd gnd cell_6t
Xbit_r214_c162 bl_162 br_162 wl_214 vdd gnd cell_6t
Xbit_r215_c162 bl_162 br_162 wl_215 vdd gnd cell_6t
Xbit_r216_c162 bl_162 br_162 wl_216 vdd gnd cell_6t
Xbit_r217_c162 bl_162 br_162 wl_217 vdd gnd cell_6t
Xbit_r218_c162 bl_162 br_162 wl_218 vdd gnd cell_6t
Xbit_r219_c162 bl_162 br_162 wl_219 vdd gnd cell_6t
Xbit_r220_c162 bl_162 br_162 wl_220 vdd gnd cell_6t
Xbit_r221_c162 bl_162 br_162 wl_221 vdd gnd cell_6t
Xbit_r222_c162 bl_162 br_162 wl_222 vdd gnd cell_6t
Xbit_r223_c162 bl_162 br_162 wl_223 vdd gnd cell_6t
Xbit_r224_c162 bl_162 br_162 wl_224 vdd gnd cell_6t
Xbit_r225_c162 bl_162 br_162 wl_225 vdd gnd cell_6t
Xbit_r226_c162 bl_162 br_162 wl_226 vdd gnd cell_6t
Xbit_r227_c162 bl_162 br_162 wl_227 vdd gnd cell_6t
Xbit_r228_c162 bl_162 br_162 wl_228 vdd gnd cell_6t
Xbit_r229_c162 bl_162 br_162 wl_229 vdd gnd cell_6t
Xbit_r230_c162 bl_162 br_162 wl_230 vdd gnd cell_6t
Xbit_r231_c162 bl_162 br_162 wl_231 vdd gnd cell_6t
Xbit_r232_c162 bl_162 br_162 wl_232 vdd gnd cell_6t
Xbit_r233_c162 bl_162 br_162 wl_233 vdd gnd cell_6t
Xbit_r234_c162 bl_162 br_162 wl_234 vdd gnd cell_6t
Xbit_r235_c162 bl_162 br_162 wl_235 vdd gnd cell_6t
Xbit_r236_c162 bl_162 br_162 wl_236 vdd gnd cell_6t
Xbit_r237_c162 bl_162 br_162 wl_237 vdd gnd cell_6t
Xbit_r238_c162 bl_162 br_162 wl_238 vdd gnd cell_6t
Xbit_r239_c162 bl_162 br_162 wl_239 vdd gnd cell_6t
Xbit_r240_c162 bl_162 br_162 wl_240 vdd gnd cell_6t
Xbit_r241_c162 bl_162 br_162 wl_241 vdd gnd cell_6t
Xbit_r242_c162 bl_162 br_162 wl_242 vdd gnd cell_6t
Xbit_r243_c162 bl_162 br_162 wl_243 vdd gnd cell_6t
Xbit_r244_c162 bl_162 br_162 wl_244 vdd gnd cell_6t
Xbit_r245_c162 bl_162 br_162 wl_245 vdd gnd cell_6t
Xbit_r246_c162 bl_162 br_162 wl_246 vdd gnd cell_6t
Xbit_r247_c162 bl_162 br_162 wl_247 vdd gnd cell_6t
Xbit_r248_c162 bl_162 br_162 wl_248 vdd gnd cell_6t
Xbit_r249_c162 bl_162 br_162 wl_249 vdd gnd cell_6t
Xbit_r250_c162 bl_162 br_162 wl_250 vdd gnd cell_6t
Xbit_r251_c162 bl_162 br_162 wl_251 vdd gnd cell_6t
Xbit_r252_c162 bl_162 br_162 wl_252 vdd gnd cell_6t
Xbit_r253_c162 bl_162 br_162 wl_253 vdd gnd cell_6t
Xbit_r254_c162 bl_162 br_162 wl_254 vdd gnd cell_6t
Xbit_r255_c162 bl_162 br_162 wl_255 vdd gnd cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd cell_6t
Xbit_r1_c163 bl_163 br_163 wl_1 vdd gnd cell_6t
Xbit_r2_c163 bl_163 br_163 wl_2 vdd gnd cell_6t
Xbit_r3_c163 bl_163 br_163 wl_3 vdd gnd cell_6t
Xbit_r4_c163 bl_163 br_163 wl_4 vdd gnd cell_6t
Xbit_r5_c163 bl_163 br_163 wl_5 vdd gnd cell_6t
Xbit_r6_c163 bl_163 br_163 wl_6 vdd gnd cell_6t
Xbit_r7_c163 bl_163 br_163 wl_7 vdd gnd cell_6t
Xbit_r8_c163 bl_163 br_163 wl_8 vdd gnd cell_6t
Xbit_r9_c163 bl_163 br_163 wl_9 vdd gnd cell_6t
Xbit_r10_c163 bl_163 br_163 wl_10 vdd gnd cell_6t
Xbit_r11_c163 bl_163 br_163 wl_11 vdd gnd cell_6t
Xbit_r12_c163 bl_163 br_163 wl_12 vdd gnd cell_6t
Xbit_r13_c163 bl_163 br_163 wl_13 vdd gnd cell_6t
Xbit_r14_c163 bl_163 br_163 wl_14 vdd gnd cell_6t
Xbit_r15_c163 bl_163 br_163 wl_15 vdd gnd cell_6t
Xbit_r16_c163 bl_163 br_163 wl_16 vdd gnd cell_6t
Xbit_r17_c163 bl_163 br_163 wl_17 vdd gnd cell_6t
Xbit_r18_c163 bl_163 br_163 wl_18 vdd gnd cell_6t
Xbit_r19_c163 bl_163 br_163 wl_19 vdd gnd cell_6t
Xbit_r20_c163 bl_163 br_163 wl_20 vdd gnd cell_6t
Xbit_r21_c163 bl_163 br_163 wl_21 vdd gnd cell_6t
Xbit_r22_c163 bl_163 br_163 wl_22 vdd gnd cell_6t
Xbit_r23_c163 bl_163 br_163 wl_23 vdd gnd cell_6t
Xbit_r24_c163 bl_163 br_163 wl_24 vdd gnd cell_6t
Xbit_r25_c163 bl_163 br_163 wl_25 vdd gnd cell_6t
Xbit_r26_c163 bl_163 br_163 wl_26 vdd gnd cell_6t
Xbit_r27_c163 bl_163 br_163 wl_27 vdd gnd cell_6t
Xbit_r28_c163 bl_163 br_163 wl_28 vdd gnd cell_6t
Xbit_r29_c163 bl_163 br_163 wl_29 vdd gnd cell_6t
Xbit_r30_c163 bl_163 br_163 wl_30 vdd gnd cell_6t
Xbit_r31_c163 bl_163 br_163 wl_31 vdd gnd cell_6t
Xbit_r32_c163 bl_163 br_163 wl_32 vdd gnd cell_6t
Xbit_r33_c163 bl_163 br_163 wl_33 vdd gnd cell_6t
Xbit_r34_c163 bl_163 br_163 wl_34 vdd gnd cell_6t
Xbit_r35_c163 bl_163 br_163 wl_35 vdd gnd cell_6t
Xbit_r36_c163 bl_163 br_163 wl_36 vdd gnd cell_6t
Xbit_r37_c163 bl_163 br_163 wl_37 vdd gnd cell_6t
Xbit_r38_c163 bl_163 br_163 wl_38 vdd gnd cell_6t
Xbit_r39_c163 bl_163 br_163 wl_39 vdd gnd cell_6t
Xbit_r40_c163 bl_163 br_163 wl_40 vdd gnd cell_6t
Xbit_r41_c163 bl_163 br_163 wl_41 vdd gnd cell_6t
Xbit_r42_c163 bl_163 br_163 wl_42 vdd gnd cell_6t
Xbit_r43_c163 bl_163 br_163 wl_43 vdd gnd cell_6t
Xbit_r44_c163 bl_163 br_163 wl_44 vdd gnd cell_6t
Xbit_r45_c163 bl_163 br_163 wl_45 vdd gnd cell_6t
Xbit_r46_c163 bl_163 br_163 wl_46 vdd gnd cell_6t
Xbit_r47_c163 bl_163 br_163 wl_47 vdd gnd cell_6t
Xbit_r48_c163 bl_163 br_163 wl_48 vdd gnd cell_6t
Xbit_r49_c163 bl_163 br_163 wl_49 vdd gnd cell_6t
Xbit_r50_c163 bl_163 br_163 wl_50 vdd gnd cell_6t
Xbit_r51_c163 bl_163 br_163 wl_51 vdd gnd cell_6t
Xbit_r52_c163 bl_163 br_163 wl_52 vdd gnd cell_6t
Xbit_r53_c163 bl_163 br_163 wl_53 vdd gnd cell_6t
Xbit_r54_c163 bl_163 br_163 wl_54 vdd gnd cell_6t
Xbit_r55_c163 bl_163 br_163 wl_55 vdd gnd cell_6t
Xbit_r56_c163 bl_163 br_163 wl_56 vdd gnd cell_6t
Xbit_r57_c163 bl_163 br_163 wl_57 vdd gnd cell_6t
Xbit_r58_c163 bl_163 br_163 wl_58 vdd gnd cell_6t
Xbit_r59_c163 bl_163 br_163 wl_59 vdd gnd cell_6t
Xbit_r60_c163 bl_163 br_163 wl_60 vdd gnd cell_6t
Xbit_r61_c163 bl_163 br_163 wl_61 vdd gnd cell_6t
Xbit_r62_c163 bl_163 br_163 wl_62 vdd gnd cell_6t
Xbit_r63_c163 bl_163 br_163 wl_63 vdd gnd cell_6t
Xbit_r64_c163 bl_163 br_163 wl_64 vdd gnd cell_6t
Xbit_r65_c163 bl_163 br_163 wl_65 vdd gnd cell_6t
Xbit_r66_c163 bl_163 br_163 wl_66 vdd gnd cell_6t
Xbit_r67_c163 bl_163 br_163 wl_67 vdd gnd cell_6t
Xbit_r68_c163 bl_163 br_163 wl_68 vdd gnd cell_6t
Xbit_r69_c163 bl_163 br_163 wl_69 vdd gnd cell_6t
Xbit_r70_c163 bl_163 br_163 wl_70 vdd gnd cell_6t
Xbit_r71_c163 bl_163 br_163 wl_71 vdd gnd cell_6t
Xbit_r72_c163 bl_163 br_163 wl_72 vdd gnd cell_6t
Xbit_r73_c163 bl_163 br_163 wl_73 vdd gnd cell_6t
Xbit_r74_c163 bl_163 br_163 wl_74 vdd gnd cell_6t
Xbit_r75_c163 bl_163 br_163 wl_75 vdd gnd cell_6t
Xbit_r76_c163 bl_163 br_163 wl_76 vdd gnd cell_6t
Xbit_r77_c163 bl_163 br_163 wl_77 vdd gnd cell_6t
Xbit_r78_c163 bl_163 br_163 wl_78 vdd gnd cell_6t
Xbit_r79_c163 bl_163 br_163 wl_79 vdd gnd cell_6t
Xbit_r80_c163 bl_163 br_163 wl_80 vdd gnd cell_6t
Xbit_r81_c163 bl_163 br_163 wl_81 vdd gnd cell_6t
Xbit_r82_c163 bl_163 br_163 wl_82 vdd gnd cell_6t
Xbit_r83_c163 bl_163 br_163 wl_83 vdd gnd cell_6t
Xbit_r84_c163 bl_163 br_163 wl_84 vdd gnd cell_6t
Xbit_r85_c163 bl_163 br_163 wl_85 vdd gnd cell_6t
Xbit_r86_c163 bl_163 br_163 wl_86 vdd gnd cell_6t
Xbit_r87_c163 bl_163 br_163 wl_87 vdd gnd cell_6t
Xbit_r88_c163 bl_163 br_163 wl_88 vdd gnd cell_6t
Xbit_r89_c163 bl_163 br_163 wl_89 vdd gnd cell_6t
Xbit_r90_c163 bl_163 br_163 wl_90 vdd gnd cell_6t
Xbit_r91_c163 bl_163 br_163 wl_91 vdd gnd cell_6t
Xbit_r92_c163 bl_163 br_163 wl_92 vdd gnd cell_6t
Xbit_r93_c163 bl_163 br_163 wl_93 vdd gnd cell_6t
Xbit_r94_c163 bl_163 br_163 wl_94 vdd gnd cell_6t
Xbit_r95_c163 bl_163 br_163 wl_95 vdd gnd cell_6t
Xbit_r96_c163 bl_163 br_163 wl_96 vdd gnd cell_6t
Xbit_r97_c163 bl_163 br_163 wl_97 vdd gnd cell_6t
Xbit_r98_c163 bl_163 br_163 wl_98 vdd gnd cell_6t
Xbit_r99_c163 bl_163 br_163 wl_99 vdd gnd cell_6t
Xbit_r100_c163 bl_163 br_163 wl_100 vdd gnd cell_6t
Xbit_r101_c163 bl_163 br_163 wl_101 vdd gnd cell_6t
Xbit_r102_c163 bl_163 br_163 wl_102 vdd gnd cell_6t
Xbit_r103_c163 bl_163 br_163 wl_103 vdd gnd cell_6t
Xbit_r104_c163 bl_163 br_163 wl_104 vdd gnd cell_6t
Xbit_r105_c163 bl_163 br_163 wl_105 vdd gnd cell_6t
Xbit_r106_c163 bl_163 br_163 wl_106 vdd gnd cell_6t
Xbit_r107_c163 bl_163 br_163 wl_107 vdd gnd cell_6t
Xbit_r108_c163 bl_163 br_163 wl_108 vdd gnd cell_6t
Xbit_r109_c163 bl_163 br_163 wl_109 vdd gnd cell_6t
Xbit_r110_c163 bl_163 br_163 wl_110 vdd gnd cell_6t
Xbit_r111_c163 bl_163 br_163 wl_111 vdd gnd cell_6t
Xbit_r112_c163 bl_163 br_163 wl_112 vdd gnd cell_6t
Xbit_r113_c163 bl_163 br_163 wl_113 vdd gnd cell_6t
Xbit_r114_c163 bl_163 br_163 wl_114 vdd gnd cell_6t
Xbit_r115_c163 bl_163 br_163 wl_115 vdd gnd cell_6t
Xbit_r116_c163 bl_163 br_163 wl_116 vdd gnd cell_6t
Xbit_r117_c163 bl_163 br_163 wl_117 vdd gnd cell_6t
Xbit_r118_c163 bl_163 br_163 wl_118 vdd gnd cell_6t
Xbit_r119_c163 bl_163 br_163 wl_119 vdd gnd cell_6t
Xbit_r120_c163 bl_163 br_163 wl_120 vdd gnd cell_6t
Xbit_r121_c163 bl_163 br_163 wl_121 vdd gnd cell_6t
Xbit_r122_c163 bl_163 br_163 wl_122 vdd gnd cell_6t
Xbit_r123_c163 bl_163 br_163 wl_123 vdd gnd cell_6t
Xbit_r124_c163 bl_163 br_163 wl_124 vdd gnd cell_6t
Xbit_r125_c163 bl_163 br_163 wl_125 vdd gnd cell_6t
Xbit_r126_c163 bl_163 br_163 wl_126 vdd gnd cell_6t
Xbit_r127_c163 bl_163 br_163 wl_127 vdd gnd cell_6t
Xbit_r128_c163 bl_163 br_163 wl_128 vdd gnd cell_6t
Xbit_r129_c163 bl_163 br_163 wl_129 vdd gnd cell_6t
Xbit_r130_c163 bl_163 br_163 wl_130 vdd gnd cell_6t
Xbit_r131_c163 bl_163 br_163 wl_131 vdd gnd cell_6t
Xbit_r132_c163 bl_163 br_163 wl_132 vdd gnd cell_6t
Xbit_r133_c163 bl_163 br_163 wl_133 vdd gnd cell_6t
Xbit_r134_c163 bl_163 br_163 wl_134 vdd gnd cell_6t
Xbit_r135_c163 bl_163 br_163 wl_135 vdd gnd cell_6t
Xbit_r136_c163 bl_163 br_163 wl_136 vdd gnd cell_6t
Xbit_r137_c163 bl_163 br_163 wl_137 vdd gnd cell_6t
Xbit_r138_c163 bl_163 br_163 wl_138 vdd gnd cell_6t
Xbit_r139_c163 bl_163 br_163 wl_139 vdd gnd cell_6t
Xbit_r140_c163 bl_163 br_163 wl_140 vdd gnd cell_6t
Xbit_r141_c163 bl_163 br_163 wl_141 vdd gnd cell_6t
Xbit_r142_c163 bl_163 br_163 wl_142 vdd gnd cell_6t
Xbit_r143_c163 bl_163 br_163 wl_143 vdd gnd cell_6t
Xbit_r144_c163 bl_163 br_163 wl_144 vdd gnd cell_6t
Xbit_r145_c163 bl_163 br_163 wl_145 vdd gnd cell_6t
Xbit_r146_c163 bl_163 br_163 wl_146 vdd gnd cell_6t
Xbit_r147_c163 bl_163 br_163 wl_147 vdd gnd cell_6t
Xbit_r148_c163 bl_163 br_163 wl_148 vdd gnd cell_6t
Xbit_r149_c163 bl_163 br_163 wl_149 vdd gnd cell_6t
Xbit_r150_c163 bl_163 br_163 wl_150 vdd gnd cell_6t
Xbit_r151_c163 bl_163 br_163 wl_151 vdd gnd cell_6t
Xbit_r152_c163 bl_163 br_163 wl_152 vdd gnd cell_6t
Xbit_r153_c163 bl_163 br_163 wl_153 vdd gnd cell_6t
Xbit_r154_c163 bl_163 br_163 wl_154 vdd gnd cell_6t
Xbit_r155_c163 bl_163 br_163 wl_155 vdd gnd cell_6t
Xbit_r156_c163 bl_163 br_163 wl_156 vdd gnd cell_6t
Xbit_r157_c163 bl_163 br_163 wl_157 vdd gnd cell_6t
Xbit_r158_c163 bl_163 br_163 wl_158 vdd gnd cell_6t
Xbit_r159_c163 bl_163 br_163 wl_159 vdd gnd cell_6t
Xbit_r160_c163 bl_163 br_163 wl_160 vdd gnd cell_6t
Xbit_r161_c163 bl_163 br_163 wl_161 vdd gnd cell_6t
Xbit_r162_c163 bl_163 br_163 wl_162 vdd gnd cell_6t
Xbit_r163_c163 bl_163 br_163 wl_163 vdd gnd cell_6t
Xbit_r164_c163 bl_163 br_163 wl_164 vdd gnd cell_6t
Xbit_r165_c163 bl_163 br_163 wl_165 vdd gnd cell_6t
Xbit_r166_c163 bl_163 br_163 wl_166 vdd gnd cell_6t
Xbit_r167_c163 bl_163 br_163 wl_167 vdd gnd cell_6t
Xbit_r168_c163 bl_163 br_163 wl_168 vdd gnd cell_6t
Xbit_r169_c163 bl_163 br_163 wl_169 vdd gnd cell_6t
Xbit_r170_c163 bl_163 br_163 wl_170 vdd gnd cell_6t
Xbit_r171_c163 bl_163 br_163 wl_171 vdd gnd cell_6t
Xbit_r172_c163 bl_163 br_163 wl_172 vdd gnd cell_6t
Xbit_r173_c163 bl_163 br_163 wl_173 vdd gnd cell_6t
Xbit_r174_c163 bl_163 br_163 wl_174 vdd gnd cell_6t
Xbit_r175_c163 bl_163 br_163 wl_175 vdd gnd cell_6t
Xbit_r176_c163 bl_163 br_163 wl_176 vdd gnd cell_6t
Xbit_r177_c163 bl_163 br_163 wl_177 vdd gnd cell_6t
Xbit_r178_c163 bl_163 br_163 wl_178 vdd gnd cell_6t
Xbit_r179_c163 bl_163 br_163 wl_179 vdd gnd cell_6t
Xbit_r180_c163 bl_163 br_163 wl_180 vdd gnd cell_6t
Xbit_r181_c163 bl_163 br_163 wl_181 vdd gnd cell_6t
Xbit_r182_c163 bl_163 br_163 wl_182 vdd gnd cell_6t
Xbit_r183_c163 bl_163 br_163 wl_183 vdd gnd cell_6t
Xbit_r184_c163 bl_163 br_163 wl_184 vdd gnd cell_6t
Xbit_r185_c163 bl_163 br_163 wl_185 vdd gnd cell_6t
Xbit_r186_c163 bl_163 br_163 wl_186 vdd gnd cell_6t
Xbit_r187_c163 bl_163 br_163 wl_187 vdd gnd cell_6t
Xbit_r188_c163 bl_163 br_163 wl_188 vdd gnd cell_6t
Xbit_r189_c163 bl_163 br_163 wl_189 vdd gnd cell_6t
Xbit_r190_c163 bl_163 br_163 wl_190 vdd gnd cell_6t
Xbit_r191_c163 bl_163 br_163 wl_191 vdd gnd cell_6t
Xbit_r192_c163 bl_163 br_163 wl_192 vdd gnd cell_6t
Xbit_r193_c163 bl_163 br_163 wl_193 vdd gnd cell_6t
Xbit_r194_c163 bl_163 br_163 wl_194 vdd gnd cell_6t
Xbit_r195_c163 bl_163 br_163 wl_195 vdd gnd cell_6t
Xbit_r196_c163 bl_163 br_163 wl_196 vdd gnd cell_6t
Xbit_r197_c163 bl_163 br_163 wl_197 vdd gnd cell_6t
Xbit_r198_c163 bl_163 br_163 wl_198 vdd gnd cell_6t
Xbit_r199_c163 bl_163 br_163 wl_199 vdd gnd cell_6t
Xbit_r200_c163 bl_163 br_163 wl_200 vdd gnd cell_6t
Xbit_r201_c163 bl_163 br_163 wl_201 vdd gnd cell_6t
Xbit_r202_c163 bl_163 br_163 wl_202 vdd gnd cell_6t
Xbit_r203_c163 bl_163 br_163 wl_203 vdd gnd cell_6t
Xbit_r204_c163 bl_163 br_163 wl_204 vdd gnd cell_6t
Xbit_r205_c163 bl_163 br_163 wl_205 vdd gnd cell_6t
Xbit_r206_c163 bl_163 br_163 wl_206 vdd gnd cell_6t
Xbit_r207_c163 bl_163 br_163 wl_207 vdd gnd cell_6t
Xbit_r208_c163 bl_163 br_163 wl_208 vdd gnd cell_6t
Xbit_r209_c163 bl_163 br_163 wl_209 vdd gnd cell_6t
Xbit_r210_c163 bl_163 br_163 wl_210 vdd gnd cell_6t
Xbit_r211_c163 bl_163 br_163 wl_211 vdd gnd cell_6t
Xbit_r212_c163 bl_163 br_163 wl_212 vdd gnd cell_6t
Xbit_r213_c163 bl_163 br_163 wl_213 vdd gnd cell_6t
Xbit_r214_c163 bl_163 br_163 wl_214 vdd gnd cell_6t
Xbit_r215_c163 bl_163 br_163 wl_215 vdd gnd cell_6t
Xbit_r216_c163 bl_163 br_163 wl_216 vdd gnd cell_6t
Xbit_r217_c163 bl_163 br_163 wl_217 vdd gnd cell_6t
Xbit_r218_c163 bl_163 br_163 wl_218 vdd gnd cell_6t
Xbit_r219_c163 bl_163 br_163 wl_219 vdd gnd cell_6t
Xbit_r220_c163 bl_163 br_163 wl_220 vdd gnd cell_6t
Xbit_r221_c163 bl_163 br_163 wl_221 vdd gnd cell_6t
Xbit_r222_c163 bl_163 br_163 wl_222 vdd gnd cell_6t
Xbit_r223_c163 bl_163 br_163 wl_223 vdd gnd cell_6t
Xbit_r224_c163 bl_163 br_163 wl_224 vdd gnd cell_6t
Xbit_r225_c163 bl_163 br_163 wl_225 vdd gnd cell_6t
Xbit_r226_c163 bl_163 br_163 wl_226 vdd gnd cell_6t
Xbit_r227_c163 bl_163 br_163 wl_227 vdd gnd cell_6t
Xbit_r228_c163 bl_163 br_163 wl_228 vdd gnd cell_6t
Xbit_r229_c163 bl_163 br_163 wl_229 vdd gnd cell_6t
Xbit_r230_c163 bl_163 br_163 wl_230 vdd gnd cell_6t
Xbit_r231_c163 bl_163 br_163 wl_231 vdd gnd cell_6t
Xbit_r232_c163 bl_163 br_163 wl_232 vdd gnd cell_6t
Xbit_r233_c163 bl_163 br_163 wl_233 vdd gnd cell_6t
Xbit_r234_c163 bl_163 br_163 wl_234 vdd gnd cell_6t
Xbit_r235_c163 bl_163 br_163 wl_235 vdd gnd cell_6t
Xbit_r236_c163 bl_163 br_163 wl_236 vdd gnd cell_6t
Xbit_r237_c163 bl_163 br_163 wl_237 vdd gnd cell_6t
Xbit_r238_c163 bl_163 br_163 wl_238 vdd gnd cell_6t
Xbit_r239_c163 bl_163 br_163 wl_239 vdd gnd cell_6t
Xbit_r240_c163 bl_163 br_163 wl_240 vdd gnd cell_6t
Xbit_r241_c163 bl_163 br_163 wl_241 vdd gnd cell_6t
Xbit_r242_c163 bl_163 br_163 wl_242 vdd gnd cell_6t
Xbit_r243_c163 bl_163 br_163 wl_243 vdd gnd cell_6t
Xbit_r244_c163 bl_163 br_163 wl_244 vdd gnd cell_6t
Xbit_r245_c163 bl_163 br_163 wl_245 vdd gnd cell_6t
Xbit_r246_c163 bl_163 br_163 wl_246 vdd gnd cell_6t
Xbit_r247_c163 bl_163 br_163 wl_247 vdd gnd cell_6t
Xbit_r248_c163 bl_163 br_163 wl_248 vdd gnd cell_6t
Xbit_r249_c163 bl_163 br_163 wl_249 vdd gnd cell_6t
Xbit_r250_c163 bl_163 br_163 wl_250 vdd gnd cell_6t
Xbit_r251_c163 bl_163 br_163 wl_251 vdd gnd cell_6t
Xbit_r252_c163 bl_163 br_163 wl_252 vdd gnd cell_6t
Xbit_r253_c163 bl_163 br_163 wl_253 vdd gnd cell_6t
Xbit_r254_c163 bl_163 br_163 wl_254 vdd gnd cell_6t
Xbit_r255_c163 bl_163 br_163 wl_255 vdd gnd cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd cell_6t
Xbit_r1_c164 bl_164 br_164 wl_1 vdd gnd cell_6t
Xbit_r2_c164 bl_164 br_164 wl_2 vdd gnd cell_6t
Xbit_r3_c164 bl_164 br_164 wl_3 vdd gnd cell_6t
Xbit_r4_c164 bl_164 br_164 wl_4 vdd gnd cell_6t
Xbit_r5_c164 bl_164 br_164 wl_5 vdd gnd cell_6t
Xbit_r6_c164 bl_164 br_164 wl_6 vdd gnd cell_6t
Xbit_r7_c164 bl_164 br_164 wl_7 vdd gnd cell_6t
Xbit_r8_c164 bl_164 br_164 wl_8 vdd gnd cell_6t
Xbit_r9_c164 bl_164 br_164 wl_9 vdd gnd cell_6t
Xbit_r10_c164 bl_164 br_164 wl_10 vdd gnd cell_6t
Xbit_r11_c164 bl_164 br_164 wl_11 vdd gnd cell_6t
Xbit_r12_c164 bl_164 br_164 wl_12 vdd gnd cell_6t
Xbit_r13_c164 bl_164 br_164 wl_13 vdd gnd cell_6t
Xbit_r14_c164 bl_164 br_164 wl_14 vdd gnd cell_6t
Xbit_r15_c164 bl_164 br_164 wl_15 vdd gnd cell_6t
Xbit_r16_c164 bl_164 br_164 wl_16 vdd gnd cell_6t
Xbit_r17_c164 bl_164 br_164 wl_17 vdd gnd cell_6t
Xbit_r18_c164 bl_164 br_164 wl_18 vdd gnd cell_6t
Xbit_r19_c164 bl_164 br_164 wl_19 vdd gnd cell_6t
Xbit_r20_c164 bl_164 br_164 wl_20 vdd gnd cell_6t
Xbit_r21_c164 bl_164 br_164 wl_21 vdd gnd cell_6t
Xbit_r22_c164 bl_164 br_164 wl_22 vdd gnd cell_6t
Xbit_r23_c164 bl_164 br_164 wl_23 vdd gnd cell_6t
Xbit_r24_c164 bl_164 br_164 wl_24 vdd gnd cell_6t
Xbit_r25_c164 bl_164 br_164 wl_25 vdd gnd cell_6t
Xbit_r26_c164 bl_164 br_164 wl_26 vdd gnd cell_6t
Xbit_r27_c164 bl_164 br_164 wl_27 vdd gnd cell_6t
Xbit_r28_c164 bl_164 br_164 wl_28 vdd gnd cell_6t
Xbit_r29_c164 bl_164 br_164 wl_29 vdd gnd cell_6t
Xbit_r30_c164 bl_164 br_164 wl_30 vdd gnd cell_6t
Xbit_r31_c164 bl_164 br_164 wl_31 vdd gnd cell_6t
Xbit_r32_c164 bl_164 br_164 wl_32 vdd gnd cell_6t
Xbit_r33_c164 bl_164 br_164 wl_33 vdd gnd cell_6t
Xbit_r34_c164 bl_164 br_164 wl_34 vdd gnd cell_6t
Xbit_r35_c164 bl_164 br_164 wl_35 vdd gnd cell_6t
Xbit_r36_c164 bl_164 br_164 wl_36 vdd gnd cell_6t
Xbit_r37_c164 bl_164 br_164 wl_37 vdd gnd cell_6t
Xbit_r38_c164 bl_164 br_164 wl_38 vdd gnd cell_6t
Xbit_r39_c164 bl_164 br_164 wl_39 vdd gnd cell_6t
Xbit_r40_c164 bl_164 br_164 wl_40 vdd gnd cell_6t
Xbit_r41_c164 bl_164 br_164 wl_41 vdd gnd cell_6t
Xbit_r42_c164 bl_164 br_164 wl_42 vdd gnd cell_6t
Xbit_r43_c164 bl_164 br_164 wl_43 vdd gnd cell_6t
Xbit_r44_c164 bl_164 br_164 wl_44 vdd gnd cell_6t
Xbit_r45_c164 bl_164 br_164 wl_45 vdd gnd cell_6t
Xbit_r46_c164 bl_164 br_164 wl_46 vdd gnd cell_6t
Xbit_r47_c164 bl_164 br_164 wl_47 vdd gnd cell_6t
Xbit_r48_c164 bl_164 br_164 wl_48 vdd gnd cell_6t
Xbit_r49_c164 bl_164 br_164 wl_49 vdd gnd cell_6t
Xbit_r50_c164 bl_164 br_164 wl_50 vdd gnd cell_6t
Xbit_r51_c164 bl_164 br_164 wl_51 vdd gnd cell_6t
Xbit_r52_c164 bl_164 br_164 wl_52 vdd gnd cell_6t
Xbit_r53_c164 bl_164 br_164 wl_53 vdd gnd cell_6t
Xbit_r54_c164 bl_164 br_164 wl_54 vdd gnd cell_6t
Xbit_r55_c164 bl_164 br_164 wl_55 vdd gnd cell_6t
Xbit_r56_c164 bl_164 br_164 wl_56 vdd gnd cell_6t
Xbit_r57_c164 bl_164 br_164 wl_57 vdd gnd cell_6t
Xbit_r58_c164 bl_164 br_164 wl_58 vdd gnd cell_6t
Xbit_r59_c164 bl_164 br_164 wl_59 vdd gnd cell_6t
Xbit_r60_c164 bl_164 br_164 wl_60 vdd gnd cell_6t
Xbit_r61_c164 bl_164 br_164 wl_61 vdd gnd cell_6t
Xbit_r62_c164 bl_164 br_164 wl_62 vdd gnd cell_6t
Xbit_r63_c164 bl_164 br_164 wl_63 vdd gnd cell_6t
Xbit_r64_c164 bl_164 br_164 wl_64 vdd gnd cell_6t
Xbit_r65_c164 bl_164 br_164 wl_65 vdd gnd cell_6t
Xbit_r66_c164 bl_164 br_164 wl_66 vdd gnd cell_6t
Xbit_r67_c164 bl_164 br_164 wl_67 vdd gnd cell_6t
Xbit_r68_c164 bl_164 br_164 wl_68 vdd gnd cell_6t
Xbit_r69_c164 bl_164 br_164 wl_69 vdd gnd cell_6t
Xbit_r70_c164 bl_164 br_164 wl_70 vdd gnd cell_6t
Xbit_r71_c164 bl_164 br_164 wl_71 vdd gnd cell_6t
Xbit_r72_c164 bl_164 br_164 wl_72 vdd gnd cell_6t
Xbit_r73_c164 bl_164 br_164 wl_73 vdd gnd cell_6t
Xbit_r74_c164 bl_164 br_164 wl_74 vdd gnd cell_6t
Xbit_r75_c164 bl_164 br_164 wl_75 vdd gnd cell_6t
Xbit_r76_c164 bl_164 br_164 wl_76 vdd gnd cell_6t
Xbit_r77_c164 bl_164 br_164 wl_77 vdd gnd cell_6t
Xbit_r78_c164 bl_164 br_164 wl_78 vdd gnd cell_6t
Xbit_r79_c164 bl_164 br_164 wl_79 vdd gnd cell_6t
Xbit_r80_c164 bl_164 br_164 wl_80 vdd gnd cell_6t
Xbit_r81_c164 bl_164 br_164 wl_81 vdd gnd cell_6t
Xbit_r82_c164 bl_164 br_164 wl_82 vdd gnd cell_6t
Xbit_r83_c164 bl_164 br_164 wl_83 vdd gnd cell_6t
Xbit_r84_c164 bl_164 br_164 wl_84 vdd gnd cell_6t
Xbit_r85_c164 bl_164 br_164 wl_85 vdd gnd cell_6t
Xbit_r86_c164 bl_164 br_164 wl_86 vdd gnd cell_6t
Xbit_r87_c164 bl_164 br_164 wl_87 vdd gnd cell_6t
Xbit_r88_c164 bl_164 br_164 wl_88 vdd gnd cell_6t
Xbit_r89_c164 bl_164 br_164 wl_89 vdd gnd cell_6t
Xbit_r90_c164 bl_164 br_164 wl_90 vdd gnd cell_6t
Xbit_r91_c164 bl_164 br_164 wl_91 vdd gnd cell_6t
Xbit_r92_c164 bl_164 br_164 wl_92 vdd gnd cell_6t
Xbit_r93_c164 bl_164 br_164 wl_93 vdd gnd cell_6t
Xbit_r94_c164 bl_164 br_164 wl_94 vdd gnd cell_6t
Xbit_r95_c164 bl_164 br_164 wl_95 vdd gnd cell_6t
Xbit_r96_c164 bl_164 br_164 wl_96 vdd gnd cell_6t
Xbit_r97_c164 bl_164 br_164 wl_97 vdd gnd cell_6t
Xbit_r98_c164 bl_164 br_164 wl_98 vdd gnd cell_6t
Xbit_r99_c164 bl_164 br_164 wl_99 vdd gnd cell_6t
Xbit_r100_c164 bl_164 br_164 wl_100 vdd gnd cell_6t
Xbit_r101_c164 bl_164 br_164 wl_101 vdd gnd cell_6t
Xbit_r102_c164 bl_164 br_164 wl_102 vdd gnd cell_6t
Xbit_r103_c164 bl_164 br_164 wl_103 vdd gnd cell_6t
Xbit_r104_c164 bl_164 br_164 wl_104 vdd gnd cell_6t
Xbit_r105_c164 bl_164 br_164 wl_105 vdd gnd cell_6t
Xbit_r106_c164 bl_164 br_164 wl_106 vdd gnd cell_6t
Xbit_r107_c164 bl_164 br_164 wl_107 vdd gnd cell_6t
Xbit_r108_c164 bl_164 br_164 wl_108 vdd gnd cell_6t
Xbit_r109_c164 bl_164 br_164 wl_109 vdd gnd cell_6t
Xbit_r110_c164 bl_164 br_164 wl_110 vdd gnd cell_6t
Xbit_r111_c164 bl_164 br_164 wl_111 vdd gnd cell_6t
Xbit_r112_c164 bl_164 br_164 wl_112 vdd gnd cell_6t
Xbit_r113_c164 bl_164 br_164 wl_113 vdd gnd cell_6t
Xbit_r114_c164 bl_164 br_164 wl_114 vdd gnd cell_6t
Xbit_r115_c164 bl_164 br_164 wl_115 vdd gnd cell_6t
Xbit_r116_c164 bl_164 br_164 wl_116 vdd gnd cell_6t
Xbit_r117_c164 bl_164 br_164 wl_117 vdd gnd cell_6t
Xbit_r118_c164 bl_164 br_164 wl_118 vdd gnd cell_6t
Xbit_r119_c164 bl_164 br_164 wl_119 vdd gnd cell_6t
Xbit_r120_c164 bl_164 br_164 wl_120 vdd gnd cell_6t
Xbit_r121_c164 bl_164 br_164 wl_121 vdd gnd cell_6t
Xbit_r122_c164 bl_164 br_164 wl_122 vdd gnd cell_6t
Xbit_r123_c164 bl_164 br_164 wl_123 vdd gnd cell_6t
Xbit_r124_c164 bl_164 br_164 wl_124 vdd gnd cell_6t
Xbit_r125_c164 bl_164 br_164 wl_125 vdd gnd cell_6t
Xbit_r126_c164 bl_164 br_164 wl_126 vdd gnd cell_6t
Xbit_r127_c164 bl_164 br_164 wl_127 vdd gnd cell_6t
Xbit_r128_c164 bl_164 br_164 wl_128 vdd gnd cell_6t
Xbit_r129_c164 bl_164 br_164 wl_129 vdd gnd cell_6t
Xbit_r130_c164 bl_164 br_164 wl_130 vdd gnd cell_6t
Xbit_r131_c164 bl_164 br_164 wl_131 vdd gnd cell_6t
Xbit_r132_c164 bl_164 br_164 wl_132 vdd gnd cell_6t
Xbit_r133_c164 bl_164 br_164 wl_133 vdd gnd cell_6t
Xbit_r134_c164 bl_164 br_164 wl_134 vdd gnd cell_6t
Xbit_r135_c164 bl_164 br_164 wl_135 vdd gnd cell_6t
Xbit_r136_c164 bl_164 br_164 wl_136 vdd gnd cell_6t
Xbit_r137_c164 bl_164 br_164 wl_137 vdd gnd cell_6t
Xbit_r138_c164 bl_164 br_164 wl_138 vdd gnd cell_6t
Xbit_r139_c164 bl_164 br_164 wl_139 vdd gnd cell_6t
Xbit_r140_c164 bl_164 br_164 wl_140 vdd gnd cell_6t
Xbit_r141_c164 bl_164 br_164 wl_141 vdd gnd cell_6t
Xbit_r142_c164 bl_164 br_164 wl_142 vdd gnd cell_6t
Xbit_r143_c164 bl_164 br_164 wl_143 vdd gnd cell_6t
Xbit_r144_c164 bl_164 br_164 wl_144 vdd gnd cell_6t
Xbit_r145_c164 bl_164 br_164 wl_145 vdd gnd cell_6t
Xbit_r146_c164 bl_164 br_164 wl_146 vdd gnd cell_6t
Xbit_r147_c164 bl_164 br_164 wl_147 vdd gnd cell_6t
Xbit_r148_c164 bl_164 br_164 wl_148 vdd gnd cell_6t
Xbit_r149_c164 bl_164 br_164 wl_149 vdd gnd cell_6t
Xbit_r150_c164 bl_164 br_164 wl_150 vdd gnd cell_6t
Xbit_r151_c164 bl_164 br_164 wl_151 vdd gnd cell_6t
Xbit_r152_c164 bl_164 br_164 wl_152 vdd gnd cell_6t
Xbit_r153_c164 bl_164 br_164 wl_153 vdd gnd cell_6t
Xbit_r154_c164 bl_164 br_164 wl_154 vdd gnd cell_6t
Xbit_r155_c164 bl_164 br_164 wl_155 vdd gnd cell_6t
Xbit_r156_c164 bl_164 br_164 wl_156 vdd gnd cell_6t
Xbit_r157_c164 bl_164 br_164 wl_157 vdd gnd cell_6t
Xbit_r158_c164 bl_164 br_164 wl_158 vdd gnd cell_6t
Xbit_r159_c164 bl_164 br_164 wl_159 vdd gnd cell_6t
Xbit_r160_c164 bl_164 br_164 wl_160 vdd gnd cell_6t
Xbit_r161_c164 bl_164 br_164 wl_161 vdd gnd cell_6t
Xbit_r162_c164 bl_164 br_164 wl_162 vdd gnd cell_6t
Xbit_r163_c164 bl_164 br_164 wl_163 vdd gnd cell_6t
Xbit_r164_c164 bl_164 br_164 wl_164 vdd gnd cell_6t
Xbit_r165_c164 bl_164 br_164 wl_165 vdd gnd cell_6t
Xbit_r166_c164 bl_164 br_164 wl_166 vdd gnd cell_6t
Xbit_r167_c164 bl_164 br_164 wl_167 vdd gnd cell_6t
Xbit_r168_c164 bl_164 br_164 wl_168 vdd gnd cell_6t
Xbit_r169_c164 bl_164 br_164 wl_169 vdd gnd cell_6t
Xbit_r170_c164 bl_164 br_164 wl_170 vdd gnd cell_6t
Xbit_r171_c164 bl_164 br_164 wl_171 vdd gnd cell_6t
Xbit_r172_c164 bl_164 br_164 wl_172 vdd gnd cell_6t
Xbit_r173_c164 bl_164 br_164 wl_173 vdd gnd cell_6t
Xbit_r174_c164 bl_164 br_164 wl_174 vdd gnd cell_6t
Xbit_r175_c164 bl_164 br_164 wl_175 vdd gnd cell_6t
Xbit_r176_c164 bl_164 br_164 wl_176 vdd gnd cell_6t
Xbit_r177_c164 bl_164 br_164 wl_177 vdd gnd cell_6t
Xbit_r178_c164 bl_164 br_164 wl_178 vdd gnd cell_6t
Xbit_r179_c164 bl_164 br_164 wl_179 vdd gnd cell_6t
Xbit_r180_c164 bl_164 br_164 wl_180 vdd gnd cell_6t
Xbit_r181_c164 bl_164 br_164 wl_181 vdd gnd cell_6t
Xbit_r182_c164 bl_164 br_164 wl_182 vdd gnd cell_6t
Xbit_r183_c164 bl_164 br_164 wl_183 vdd gnd cell_6t
Xbit_r184_c164 bl_164 br_164 wl_184 vdd gnd cell_6t
Xbit_r185_c164 bl_164 br_164 wl_185 vdd gnd cell_6t
Xbit_r186_c164 bl_164 br_164 wl_186 vdd gnd cell_6t
Xbit_r187_c164 bl_164 br_164 wl_187 vdd gnd cell_6t
Xbit_r188_c164 bl_164 br_164 wl_188 vdd gnd cell_6t
Xbit_r189_c164 bl_164 br_164 wl_189 vdd gnd cell_6t
Xbit_r190_c164 bl_164 br_164 wl_190 vdd gnd cell_6t
Xbit_r191_c164 bl_164 br_164 wl_191 vdd gnd cell_6t
Xbit_r192_c164 bl_164 br_164 wl_192 vdd gnd cell_6t
Xbit_r193_c164 bl_164 br_164 wl_193 vdd gnd cell_6t
Xbit_r194_c164 bl_164 br_164 wl_194 vdd gnd cell_6t
Xbit_r195_c164 bl_164 br_164 wl_195 vdd gnd cell_6t
Xbit_r196_c164 bl_164 br_164 wl_196 vdd gnd cell_6t
Xbit_r197_c164 bl_164 br_164 wl_197 vdd gnd cell_6t
Xbit_r198_c164 bl_164 br_164 wl_198 vdd gnd cell_6t
Xbit_r199_c164 bl_164 br_164 wl_199 vdd gnd cell_6t
Xbit_r200_c164 bl_164 br_164 wl_200 vdd gnd cell_6t
Xbit_r201_c164 bl_164 br_164 wl_201 vdd gnd cell_6t
Xbit_r202_c164 bl_164 br_164 wl_202 vdd gnd cell_6t
Xbit_r203_c164 bl_164 br_164 wl_203 vdd gnd cell_6t
Xbit_r204_c164 bl_164 br_164 wl_204 vdd gnd cell_6t
Xbit_r205_c164 bl_164 br_164 wl_205 vdd gnd cell_6t
Xbit_r206_c164 bl_164 br_164 wl_206 vdd gnd cell_6t
Xbit_r207_c164 bl_164 br_164 wl_207 vdd gnd cell_6t
Xbit_r208_c164 bl_164 br_164 wl_208 vdd gnd cell_6t
Xbit_r209_c164 bl_164 br_164 wl_209 vdd gnd cell_6t
Xbit_r210_c164 bl_164 br_164 wl_210 vdd gnd cell_6t
Xbit_r211_c164 bl_164 br_164 wl_211 vdd gnd cell_6t
Xbit_r212_c164 bl_164 br_164 wl_212 vdd gnd cell_6t
Xbit_r213_c164 bl_164 br_164 wl_213 vdd gnd cell_6t
Xbit_r214_c164 bl_164 br_164 wl_214 vdd gnd cell_6t
Xbit_r215_c164 bl_164 br_164 wl_215 vdd gnd cell_6t
Xbit_r216_c164 bl_164 br_164 wl_216 vdd gnd cell_6t
Xbit_r217_c164 bl_164 br_164 wl_217 vdd gnd cell_6t
Xbit_r218_c164 bl_164 br_164 wl_218 vdd gnd cell_6t
Xbit_r219_c164 bl_164 br_164 wl_219 vdd gnd cell_6t
Xbit_r220_c164 bl_164 br_164 wl_220 vdd gnd cell_6t
Xbit_r221_c164 bl_164 br_164 wl_221 vdd gnd cell_6t
Xbit_r222_c164 bl_164 br_164 wl_222 vdd gnd cell_6t
Xbit_r223_c164 bl_164 br_164 wl_223 vdd gnd cell_6t
Xbit_r224_c164 bl_164 br_164 wl_224 vdd gnd cell_6t
Xbit_r225_c164 bl_164 br_164 wl_225 vdd gnd cell_6t
Xbit_r226_c164 bl_164 br_164 wl_226 vdd gnd cell_6t
Xbit_r227_c164 bl_164 br_164 wl_227 vdd gnd cell_6t
Xbit_r228_c164 bl_164 br_164 wl_228 vdd gnd cell_6t
Xbit_r229_c164 bl_164 br_164 wl_229 vdd gnd cell_6t
Xbit_r230_c164 bl_164 br_164 wl_230 vdd gnd cell_6t
Xbit_r231_c164 bl_164 br_164 wl_231 vdd gnd cell_6t
Xbit_r232_c164 bl_164 br_164 wl_232 vdd gnd cell_6t
Xbit_r233_c164 bl_164 br_164 wl_233 vdd gnd cell_6t
Xbit_r234_c164 bl_164 br_164 wl_234 vdd gnd cell_6t
Xbit_r235_c164 bl_164 br_164 wl_235 vdd gnd cell_6t
Xbit_r236_c164 bl_164 br_164 wl_236 vdd gnd cell_6t
Xbit_r237_c164 bl_164 br_164 wl_237 vdd gnd cell_6t
Xbit_r238_c164 bl_164 br_164 wl_238 vdd gnd cell_6t
Xbit_r239_c164 bl_164 br_164 wl_239 vdd gnd cell_6t
Xbit_r240_c164 bl_164 br_164 wl_240 vdd gnd cell_6t
Xbit_r241_c164 bl_164 br_164 wl_241 vdd gnd cell_6t
Xbit_r242_c164 bl_164 br_164 wl_242 vdd gnd cell_6t
Xbit_r243_c164 bl_164 br_164 wl_243 vdd gnd cell_6t
Xbit_r244_c164 bl_164 br_164 wl_244 vdd gnd cell_6t
Xbit_r245_c164 bl_164 br_164 wl_245 vdd gnd cell_6t
Xbit_r246_c164 bl_164 br_164 wl_246 vdd gnd cell_6t
Xbit_r247_c164 bl_164 br_164 wl_247 vdd gnd cell_6t
Xbit_r248_c164 bl_164 br_164 wl_248 vdd gnd cell_6t
Xbit_r249_c164 bl_164 br_164 wl_249 vdd gnd cell_6t
Xbit_r250_c164 bl_164 br_164 wl_250 vdd gnd cell_6t
Xbit_r251_c164 bl_164 br_164 wl_251 vdd gnd cell_6t
Xbit_r252_c164 bl_164 br_164 wl_252 vdd gnd cell_6t
Xbit_r253_c164 bl_164 br_164 wl_253 vdd gnd cell_6t
Xbit_r254_c164 bl_164 br_164 wl_254 vdd gnd cell_6t
Xbit_r255_c164 bl_164 br_164 wl_255 vdd gnd cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd cell_6t
Xbit_r1_c165 bl_165 br_165 wl_1 vdd gnd cell_6t
Xbit_r2_c165 bl_165 br_165 wl_2 vdd gnd cell_6t
Xbit_r3_c165 bl_165 br_165 wl_3 vdd gnd cell_6t
Xbit_r4_c165 bl_165 br_165 wl_4 vdd gnd cell_6t
Xbit_r5_c165 bl_165 br_165 wl_5 vdd gnd cell_6t
Xbit_r6_c165 bl_165 br_165 wl_6 vdd gnd cell_6t
Xbit_r7_c165 bl_165 br_165 wl_7 vdd gnd cell_6t
Xbit_r8_c165 bl_165 br_165 wl_8 vdd gnd cell_6t
Xbit_r9_c165 bl_165 br_165 wl_9 vdd gnd cell_6t
Xbit_r10_c165 bl_165 br_165 wl_10 vdd gnd cell_6t
Xbit_r11_c165 bl_165 br_165 wl_11 vdd gnd cell_6t
Xbit_r12_c165 bl_165 br_165 wl_12 vdd gnd cell_6t
Xbit_r13_c165 bl_165 br_165 wl_13 vdd gnd cell_6t
Xbit_r14_c165 bl_165 br_165 wl_14 vdd gnd cell_6t
Xbit_r15_c165 bl_165 br_165 wl_15 vdd gnd cell_6t
Xbit_r16_c165 bl_165 br_165 wl_16 vdd gnd cell_6t
Xbit_r17_c165 bl_165 br_165 wl_17 vdd gnd cell_6t
Xbit_r18_c165 bl_165 br_165 wl_18 vdd gnd cell_6t
Xbit_r19_c165 bl_165 br_165 wl_19 vdd gnd cell_6t
Xbit_r20_c165 bl_165 br_165 wl_20 vdd gnd cell_6t
Xbit_r21_c165 bl_165 br_165 wl_21 vdd gnd cell_6t
Xbit_r22_c165 bl_165 br_165 wl_22 vdd gnd cell_6t
Xbit_r23_c165 bl_165 br_165 wl_23 vdd gnd cell_6t
Xbit_r24_c165 bl_165 br_165 wl_24 vdd gnd cell_6t
Xbit_r25_c165 bl_165 br_165 wl_25 vdd gnd cell_6t
Xbit_r26_c165 bl_165 br_165 wl_26 vdd gnd cell_6t
Xbit_r27_c165 bl_165 br_165 wl_27 vdd gnd cell_6t
Xbit_r28_c165 bl_165 br_165 wl_28 vdd gnd cell_6t
Xbit_r29_c165 bl_165 br_165 wl_29 vdd gnd cell_6t
Xbit_r30_c165 bl_165 br_165 wl_30 vdd gnd cell_6t
Xbit_r31_c165 bl_165 br_165 wl_31 vdd gnd cell_6t
Xbit_r32_c165 bl_165 br_165 wl_32 vdd gnd cell_6t
Xbit_r33_c165 bl_165 br_165 wl_33 vdd gnd cell_6t
Xbit_r34_c165 bl_165 br_165 wl_34 vdd gnd cell_6t
Xbit_r35_c165 bl_165 br_165 wl_35 vdd gnd cell_6t
Xbit_r36_c165 bl_165 br_165 wl_36 vdd gnd cell_6t
Xbit_r37_c165 bl_165 br_165 wl_37 vdd gnd cell_6t
Xbit_r38_c165 bl_165 br_165 wl_38 vdd gnd cell_6t
Xbit_r39_c165 bl_165 br_165 wl_39 vdd gnd cell_6t
Xbit_r40_c165 bl_165 br_165 wl_40 vdd gnd cell_6t
Xbit_r41_c165 bl_165 br_165 wl_41 vdd gnd cell_6t
Xbit_r42_c165 bl_165 br_165 wl_42 vdd gnd cell_6t
Xbit_r43_c165 bl_165 br_165 wl_43 vdd gnd cell_6t
Xbit_r44_c165 bl_165 br_165 wl_44 vdd gnd cell_6t
Xbit_r45_c165 bl_165 br_165 wl_45 vdd gnd cell_6t
Xbit_r46_c165 bl_165 br_165 wl_46 vdd gnd cell_6t
Xbit_r47_c165 bl_165 br_165 wl_47 vdd gnd cell_6t
Xbit_r48_c165 bl_165 br_165 wl_48 vdd gnd cell_6t
Xbit_r49_c165 bl_165 br_165 wl_49 vdd gnd cell_6t
Xbit_r50_c165 bl_165 br_165 wl_50 vdd gnd cell_6t
Xbit_r51_c165 bl_165 br_165 wl_51 vdd gnd cell_6t
Xbit_r52_c165 bl_165 br_165 wl_52 vdd gnd cell_6t
Xbit_r53_c165 bl_165 br_165 wl_53 vdd gnd cell_6t
Xbit_r54_c165 bl_165 br_165 wl_54 vdd gnd cell_6t
Xbit_r55_c165 bl_165 br_165 wl_55 vdd gnd cell_6t
Xbit_r56_c165 bl_165 br_165 wl_56 vdd gnd cell_6t
Xbit_r57_c165 bl_165 br_165 wl_57 vdd gnd cell_6t
Xbit_r58_c165 bl_165 br_165 wl_58 vdd gnd cell_6t
Xbit_r59_c165 bl_165 br_165 wl_59 vdd gnd cell_6t
Xbit_r60_c165 bl_165 br_165 wl_60 vdd gnd cell_6t
Xbit_r61_c165 bl_165 br_165 wl_61 vdd gnd cell_6t
Xbit_r62_c165 bl_165 br_165 wl_62 vdd gnd cell_6t
Xbit_r63_c165 bl_165 br_165 wl_63 vdd gnd cell_6t
Xbit_r64_c165 bl_165 br_165 wl_64 vdd gnd cell_6t
Xbit_r65_c165 bl_165 br_165 wl_65 vdd gnd cell_6t
Xbit_r66_c165 bl_165 br_165 wl_66 vdd gnd cell_6t
Xbit_r67_c165 bl_165 br_165 wl_67 vdd gnd cell_6t
Xbit_r68_c165 bl_165 br_165 wl_68 vdd gnd cell_6t
Xbit_r69_c165 bl_165 br_165 wl_69 vdd gnd cell_6t
Xbit_r70_c165 bl_165 br_165 wl_70 vdd gnd cell_6t
Xbit_r71_c165 bl_165 br_165 wl_71 vdd gnd cell_6t
Xbit_r72_c165 bl_165 br_165 wl_72 vdd gnd cell_6t
Xbit_r73_c165 bl_165 br_165 wl_73 vdd gnd cell_6t
Xbit_r74_c165 bl_165 br_165 wl_74 vdd gnd cell_6t
Xbit_r75_c165 bl_165 br_165 wl_75 vdd gnd cell_6t
Xbit_r76_c165 bl_165 br_165 wl_76 vdd gnd cell_6t
Xbit_r77_c165 bl_165 br_165 wl_77 vdd gnd cell_6t
Xbit_r78_c165 bl_165 br_165 wl_78 vdd gnd cell_6t
Xbit_r79_c165 bl_165 br_165 wl_79 vdd gnd cell_6t
Xbit_r80_c165 bl_165 br_165 wl_80 vdd gnd cell_6t
Xbit_r81_c165 bl_165 br_165 wl_81 vdd gnd cell_6t
Xbit_r82_c165 bl_165 br_165 wl_82 vdd gnd cell_6t
Xbit_r83_c165 bl_165 br_165 wl_83 vdd gnd cell_6t
Xbit_r84_c165 bl_165 br_165 wl_84 vdd gnd cell_6t
Xbit_r85_c165 bl_165 br_165 wl_85 vdd gnd cell_6t
Xbit_r86_c165 bl_165 br_165 wl_86 vdd gnd cell_6t
Xbit_r87_c165 bl_165 br_165 wl_87 vdd gnd cell_6t
Xbit_r88_c165 bl_165 br_165 wl_88 vdd gnd cell_6t
Xbit_r89_c165 bl_165 br_165 wl_89 vdd gnd cell_6t
Xbit_r90_c165 bl_165 br_165 wl_90 vdd gnd cell_6t
Xbit_r91_c165 bl_165 br_165 wl_91 vdd gnd cell_6t
Xbit_r92_c165 bl_165 br_165 wl_92 vdd gnd cell_6t
Xbit_r93_c165 bl_165 br_165 wl_93 vdd gnd cell_6t
Xbit_r94_c165 bl_165 br_165 wl_94 vdd gnd cell_6t
Xbit_r95_c165 bl_165 br_165 wl_95 vdd gnd cell_6t
Xbit_r96_c165 bl_165 br_165 wl_96 vdd gnd cell_6t
Xbit_r97_c165 bl_165 br_165 wl_97 vdd gnd cell_6t
Xbit_r98_c165 bl_165 br_165 wl_98 vdd gnd cell_6t
Xbit_r99_c165 bl_165 br_165 wl_99 vdd gnd cell_6t
Xbit_r100_c165 bl_165 br_165 wl_100 vdd gnd cell_6t
Xbit_r101_c165 bl_165 br_165 wl_101 vdd gnd cell_6t
Xbit_r102_c165 bl_165 br_165 wl_102 vdd gnd cell_6t
Xbit_r103_c165 bl_165 br_165 wl_103 vdd gnd cell_6t
Xbit_r104_c165 bl_165 br_165 wl_104 vdd gnd cell_6t
Xbit_r105_c165 bl_165 br_165 wl_105 vdd gnd cell_6t
Xbit_r106_c165 bl_165 br_165 wl_106 vdd gnd cell_6t
Xbit_r107_c165 bl_165 br_165 wl_107 vdd gnd cell_6t
Xbit_r108_c165 bl_165 br_165 wl_108 vdd gnd cell_6t
Xbit_r109_c165 bl_165 br_165 wl_109 vdd gnd cell_6t
Xbit_r110_c165 bl_165 br_165 wl_110 vdd gnd cell_6t
Xbit_r111_c165 bl_165 br_165 wl_111 vdd gnd cell_6t
Xbit_r112_c165 bl_165 br_165 wl_112 vdd gnd cell_6t
Xbit_r113_c165 bl_165 br_165 wl_113 vdd gnd cell_6t
Xbit_r114_c165 bl_165 br_165 wl_114 vdd gnd cell_6t
Xbit_r115_c165 bl_165 br_165 wl_115 vdd gnd cell_6t
Xbit_r116_c165 bl_165 br_165 wl_116 vdd gnd cell_6t
Xbit_r117_c165 bl_165 br_165 wl_117 vdd gnd cell_6t
Xbit_r118_c165 bl_165 br_165 wl_118 vdd gnd cell_6t
Xbit_r119_c165 bl_165 br_165 wl_119 vdd gnd cell_6t
Xbit_r120_c165 bl_165 br_165 wl_120 vdd gnd cell_6t
Xbit_r121_c165 bl_165 br_165 wl_121 vdd gnd cell_6t
Xbit_r122_c165 bl_165 br_165 wl_122 vdd gnd cell_6t
Xbit_r123_c165 bl_165 br_165 wl_123 vdd gnd cell_6t
Xbit_r124_c165 bl_165 br_165 wl_124 vdd gnd cell_6t
Xbit_r125_c165 bl_165 br_165 wl_125 vdd gnd cell_6t
Xbit_r126_c165 bl_165 br_165 wl_126 vdd gnd cell_6t
Xbit_r127_c165 bl_165 br_165 wl_127 vdd gnd cell_6t
Xbit_r128_c165 bl_165 br_165 wl_128 vdd gnd cell_6t
Xbit_r129_c165 bl_165 br_165 wl_129 vdd gnd cell_6t
Xbit_r130_c165 bl_165 br_165 wl_130 vdd gnd cell_6t
Xbit_r131_c165 bl_165 br_165 wl_131 vdd gnd cell_6t
Xbit_r132_c165 bl_165 br_165 wl_132 vdd gnd cell_6t
Xbit_r133_c165 bl_165 br_165 wl_133 vdd gnd cell_6t
Xbit_r134_c165 bl_165 br_165 wl_134 vdd gnd cell_6t
Xbit_r135_c165 bl_165 br_165 wl_135 vdd gnd cell_6t
Xbit_r136_c165 bl_165 br_165 wl_136 vdd gnd cell_6t
Xbit_r137_c165 bl_165 br_165 wl_137 vdd gnd cell_6t
Xbit_r138_c165 bl_165 br_165 wl_138 vdd gnd cell_6t
Xbit_r139_c165 bl_165 br_165 wl_139 vdd gnd cell_6t
Xbit_r140_c165 bl_165 br_165 wl_140 vdd gnd cell_6t
Xbit_r141_c165 bl_165 br_165 wl_141 vdd gnd cell_6t
Xbit_r142_c165 bl_165 br_165 wl_142 vdd gnd cell_6t
Xbit_r143_c165 bl_165 br_165 wl_143 vdd gnd cell_6t
Xbit_r144_c165 bl_165 br_165 wl_144 vdd gnd cell_6t
Xbit_r145_c165 bl_165 br_165 wl_145 vdd gnd cell_6t
Xbit_r146_c165 bl_165 br_165 wl_146 vdd gnd cell_6t
Xbit_r147_c165 bl_165 br_165 wl_147 vdd gnd cell_6t
Xbit_r148_c165 bl_165 br_165 wl_148 vdd gnd cell_6t
Xbit_r149_c165 bl_165 br_165 wl_149 vdd gnd cell_6t
Xbit_r150_c165 bl_165 br_165 wl_150 vdd gnd cell_6t
Xbit_r151_c165 bl_165 br_165 wl_151 vdd gnd cell_6t
Xbit_r152_c165 bl_165 br_165 wl_152 vdd gnd cell_6t
Xbit_r153_c165 bl_165 br_165 wl_153 vdd gnd cell_6t
Xbit_r154_c165 bl_165 br_165 wl_154 vdd gnd cell_6t
Xbit_r155_c165 bl_165 br_165 wl_155 vdd gnd cell_6t
Xbit_r156_c165 bl_165 br_165 wl_156 vdd gnd cell_6t
Xbit_r157_c165 bl_165 br_165 wl_157 vdd gnd cell_6t
Xbit_r158_c165 bl_165 br_165 wl_158 vdd gnd cell_6t
Xbit_r159_c165 bl_165 br_165 wl_159 vdd gnd cell_6t
Xbit_r160_c165 bl_165 br_165 wl_160 vdd gnd cell_6t
Xbit_r161_c165 bl_165 br_165 wl_161 vdd gnd cell_6t
Xbit_r162_c165 bl_165 br_165 wl_162 vdd gnd cell_6t
Xbit_r163_c165 bl_165 br_165 wl_163 vdd gnd cell_6t
Xbit_r164_c165 bl_165 br_165 wl_164 vdd gnd cell_6t
Xbit_r165_c165 bl_165 br_165 wl_165 vdd gnd cell_6t
Xbit_r166_c165 bl_165 br_165 wl_166 vdd gnd cell_6t
Xbit_r167_c165 bl_165 br_165 wl_167 vdd gnd cell_6t
Xbit_r168_c165 bl_165 br_165 wl_168 vdd gnd cell_6t
Xbit_r169_c165 bl_165 br_165 wl_169 vdd gnd cell_6t
Xbit_r170_c165 bl_165 br_165 wl_170 vdd gnd cell_6t
Xbit_r171_c165 bl_165 br_165 wl_171 vdd gnd cell_6t
Xbit_r172_c165 bl_165 br_165 wl_172 vdd gnd cell_6t
Xbit_r173_c165 bl_165 br_165 wl_173 vdd gnd cell_6t
Xbit_r174_c165 bl_165 br_165 wl_174 vdd gnd cell_6t
Xbit_r175_c165 bl_165 br_165 wl_175 vdd gnd cell_6t
Xbit_r176_c165 bl_165 br_165 wl_176 vdd gnd cell_6t
Xbit_r177_c165 bl_165 br_165 wl_177 vdd gnd cell_6t
Xbit_r178_c165 bl_165 br_165 wl_178 vdd gnd cell_6t
Xbit_r179_c165 bl_165 br_165 wl_179 vdd gnd cell_6t
Xbit_r180_c165 bl_165 br_165 wl_180 vdd gnd cell_6t
Xbit_r181_c165 bl_165 br_165 wl_181 vdd gnd cell_6t
Xbit_r182_c165 bl_165 br_165 wl_182 vdd gnd cell_6t
Xbit_r183_c165 bl_165 br_165 wl_183 vdd gnd cell_6t
Xbit_r184_c165 bl_165 br_165 wl_184 vdd gnd cell_6t
Xbit_r185_c165 bl_165 br_165 wl_185 vdd gnd cell_6t
Xbit_r186_c165 bl_165 br_165 wl_186 vdd gnd cell_6t
Xbit_r187_c165 bl_165 br_165 wl_187 vdd gnd cell_6t
Xbit_r188_c165 bl_165 br_165 wl_188 vdd gnd cell_6t
Xbit_r189_c165 bl_165 br_165 wl_189 vdd gnd cell_6t
Xbit_r190_c165 bl_165 br_165 wl_190 vdd gnd cell_6t
Xbit_r191_c165 bl_165 br_165 wl_191 vdd gnd cell_6t
Xbit_r192_c165 bl_165 br_165 wl_192 vdd gnd cell_6t
Xbit_r193_c165 bl_165 br_165 wl_193 vdd gnd cell_6t
Xbit_r194_c165 bl_165 br_165 wl_194 vdd gnd cell_6t
Xbit_r195_c165 bl_165 br_165 wl_195 vdd gnd cell_6t
Xbit_r196_c165 bl_165 br_165 wl_196 vdd gnd cell_6t
Xbit_r197_c165 bl_165 br_165 wl_197 vdd gnd cell_6t
Xbit_r198_c165 bl_165 br_165 wl_198 vdd gnd cell_6t
Xbit_r199_c165 bl_165 br_165 wl_199 vdd gnd cell_6t
Xbit_r200_c165 bl_165 br_165 wl_200 vdd gnd cell_6t
Xbit_r201_c165 bl_165 br_165 wl_201 vdd gnd cell_6t
Xbit_r202_c165 bl_165 br_165 wl_202 vdd gnd cell_6t
Xbit_r203_c165 bl_165 br_165 wl_203 vdd gnd cell_6t
Xbit_r204_c165 bl_165 br_165 wl_204 vdd gnd cell_6t
Xbit_r205_c165 bl_165 br_165 wl_205 vdd gnd cell_6t
Xbit_r206_c165 bl_165 br_165 wl_206 vdd gnd cell_6t
Xbit_r207_c165 bl_165 br_165 wl_207 vdd gnd cell_6t
Xbit_r208_c165 bl_165 br_165 wl_208 vdd gnd cell_6t
Xbit_r209_c165 bl_165 br_165 wl_209 vdd gnd cell_6t
Xbit_r210_c165 bl_165 br_165 wl_210 vdd gnd cell_6t
Xbit_r211_c165 bl_165 br_165 wl_211 vdd gnd cell_6t
Xbit_r212_c165 bl_165 br_165 wl_212 vdd gnd cell_6t
Xbit_r213_c165 bl_165 br_165 wl_213 vdd gnd cell_6t
Xbit_r214_c165 bl_165 br_165 wl_214 vdd gnd cell_6t
Xbit_r215_c165 bl_165 br_165 wl_215 vdd gnd cell_6t
Xbit_r216_c165 bl_165 br_165 wl_216 vdd gnd cell_6t
Xbit_r217_c165 bl_165 br_165 wl_217 vdd gnd cell_6t
Xbit_r218_c165 bl_165 br_165 wl_218 vdd gnd cell_6t
Xbit_r219_c165 bl_165 br_165 wl_219 vdd gnd cell_6t
Xbit_r220_c165 bl_165 br_165 wl_220 vdd gnd cell_6t
Xbit_r221_c165 bl_165 br_165 wl_221 vdd gnd cell_6t
Xbit_r222_c165 bl_165 br_165 wl_222 vdd gnd cell_6t
Xbit_r223_c165 bl_165 br_165 wl_223 vdd gnd cell_6t
Xbit_r224_c165 bl_165 br_165 wl_224 vdd gnd cell_6t
Xbit_r225_c165 bl_165 br_165 wl_225 vdd gnd cell_6t
Xbit_r226_c165 bl_165 br_165 wl_226 vdd gnd cell_6t
Xbit_r227_c165 bl_165 br_165 wl_227 vdd gnd cell_6t
Xbit_r228_c165 bl_165 br_165 wl_228 vdd gnd cell_6t
Xbit_r229_c165 bl_165 br_165 wl_229 vdd gnd cell_6t
Xbit_r230_c165 bl_165 br_165 wl_230 vdd gnd cell_6t
Xbit_r231_c165 bl_165 br_165 wl_231 vdd gnd cell_6t
Xbit_r232_c165 bl_165 br_165 wl_232 vdd gnd cell_6t
Xbit_r233_c165 bl_165 br_165 wl_233 vdd gnd cell_6t
Xbit_r234_c165 bl_165 br_165 wl_234 vdd gnd cell_6t
Xbit_r235_c165 bl_165 br_165 wl_235 vdd gnd cell_6t
Xbit_r236_c165 bl_165 br_165 wl_236 vdd gnd cell_6t
Xbit_r237_c165 bl_165 br_165 wl_237 vdd gnd cell_6t
Xbit_r238_c165 bl_165 br_165 wl_238 vdd gnd cell_6t
Xbit_r239_c165 bl_165 br_165 wl_239 vdd gnd cell_6t
Xbit_r240_c165 bl_165 br_165 wl_240 vdd gnd cell_6t
Xbit_r241_c165 bl_165 br_165 wl_241 vdd gnd cell_6t
Xbit_r242_c165 bl_165 br_165 wl_242 vdd gnd cell_6t
Xbit_r243_c165 bl_165 br_165 wl_243 vdd gnd cell_6t
Xbit_r244_c165 bl_165 br_165 wl_244 vdd gnd cell_6t
Xbit_r245_c165 bl_165 br_165 wl_245 vdd gnd cell_6t
Xbit_r246_c165 bl_165 br_165 wl_246 vdd gnd cell_6t
Xbit_r247_c165 bl_165 br_165 wl_247 vdd gnd cell_6t
Xbit_r248_c165 bl_165 br_165 wl_248 vdd gnd cell_6t
Xbit_r249_c165 bl_165 br_165 wl_249 vdd gnd cell_6t
Xbit_r250_c165 bl_165 br_165 wl_250 vdd gnd cell_6t
Xbit_r251_c165 bl_165 br_165 wl_251 vdd gnd cell_6t
Xbit_r252_c165 bl_165 br_165 wl_252 vdd gnd cell_6t
Xbit_r253_c165 bl_165 br_165 wl_253 vdd gnd cell_6t
Xbit_r254_c165 bl_165 br_165 wl_254 vdd gnd cell_6t
Xbit_r255_c165 bl_165 br_165 wl_255 vdd gnd cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd cell_6t
Xbit_r1_c166 bl_166 br_166 wl_1 vdd gnd cell_6t
Xbit_r2_c166 bl_166 br_166 wl_2 vdd gnd cell_6t
Xbit_r3_c166 bl_166 br_166 wl_3 vdd gnd cell_6t
Xbit_r4_c166 bl_166 br_166 wl_4 vdd gnd cell_6t
Xbit_r5_c166 bl_166 br_166 wl_5 vdd gnd cell_6t
Xbit_r6_c166 bl_166 br_166 wl_6 vdd gnd cell_6t
Xbit_r7_c166 bl_166 br_166 wl_7 vdd gnd cell_6t
Xbit_r8_c166 bl_166 br_166 wl_8 vdd gnd cell_6t
Xbit_r9_c166 bl_166 br_166 wl_9 vdd gnd cell_6t
Xbit_r10_c166 bl_166 br_166 wl_10 vdd gnd cell_6t
Xbit_r11_c166 bl_166 br_166 wl_11 vdd gnd cell_6t
Xbit_r12_c166 bl_166 br_166 wl_12 vdd gnd cell_6t
Xbit_r13_c166 bl_166 br_166 wl_13 vdd gnd cell_6t
Xbit_r14_c166 bl_166 br_166 wl_14 vdd gnd cell_6t
Xbit_r15_c166 bl_166 br_166 wl_15 vdd gnd cell_6t
Xbit_r16_c166 bl_166 br_166 wl_16 vdd gnd cell_6t
Xbit_r17_c166 bl_166 br_166 wl_17 vdd gnd cell_6t
Xbit_r18_c166 bl_166 br_166 wl_18 vdd gnd cell_6t
Xbit_r19_c166 bl_166 br_166 wl_19 vdd gnd cell_6t
Xbit_r20_c166 bl_166 br_166 wl_20 vdd gnd cell_6t
Xbit_r21_c166 bl_166 br_166 wl_21 vdd gnd cell_6t
Xbit_r22_c166 bl_166 br_166 wl_22 vdd gnd cell_6t
Xbit_r23_c166 bl_166 br_166 wl_23 vdd gnd cell_6t
Xbit_r24_c166 bl_166 br_166 wl_24 vdd gnd cell_6t
Xbit_r25_c166 bl_166 br_166 wl_25 vdd gnd cell_6t
Xbit_r26_c166 bl_166 br_166 wl_26 vdd gnd cell_6t
Xbit_r27_c166 bl_166 br_166 wl_27 vdd gnd cell_6t
Xbit_r28_c166 bl_166 br_166 wl_28 vdd gnd cell_6t
Xbit_r29_c166 bl_166 br_166 wl_29 vdd gnd cell_6t
Xbit_r30_c166 bl_166 br_166 wl_30 vdd gnd cell_6t
Xbit_r31_c166 bl_166 br_166 wl_31 vdd gnd cell_6t
Xbit_r32_c166 bl_166 br_166 wl_32 vdd gnd cell_6t
Xbit_r33_c166 bl_166 br_166 wl_33 vdd gnd cell_6t
Xbit_r34_c166 bl_166 br_166 wl_34 vdd gnd cell_6t
Xbit_r35_c166 bl_166 br_166 wl_35 vdd gnd cell_6t
Xbit_r36_c166 bl_166 br_166 wl_36 vdd gnd cell_6t
Xbit_r37_c166 bl_166 br_166 wl_37 vdd gnd cell_6t
Xbit_r38_c166 bl_166 br_166 wl_38 vdd gnd cell_6t
Xbit_r39_c166 bl_166 br_166 wl_39 vdd gnd cell_6t
Xbit_r40_c166 bl_166 br_166 wl_40 vdd gnd cell_6t
Xbit_r41_c166 bl_166 br_166 wl_41 vdd gnd cell_6t
Xbit_r42_c166 bl_166 br_166 wl_42 vdd gnd cell_6t
Xbit_r43_c166 bl_166 br_166 wl_43 vdd gnd cell_6t
Xbit_r44_c166 bl_166 br_166 wl_44 vdd gnd cell_6t
Xbit_r45_c166 bl_166 br_166 wl_45 vdd gnd cell_6t
Xbit_r46_c166 bl_166 br_166 wl_46 vdd gnd cell_6t
Xbit_r47_c166 bl_166 br_166 wl_47 vdd gnd cell_6t
Xbit_r48_c166 bl_166 br_166 wl_48 vdd gnd cell_6t
Xbit_r49_c166 bl_166 br_166 wl_49 vdd gnd cell_6t
Xbit_r50_c166 bl_166 br_166 wl_50 vdd gnd cell_6t
Xbit_r51_c166 bl_166 br_166 wl_51 vdd gnd cell_6t
Xbit_r52_c166 bl_166 br_166 wl_52 vdd gnd cell_6t
Xbit_r53_c166 bl_166 br_166 wl_53 vdd gnd cell_6t
Xbit_r54_c166 bl_166 br_166 wl_54 vdd gnd cell_6t
Xbit_r55_c166 bl_166 br_166 wl_55 vdd gnd cell_6t
Xbit_r56_c166 bl_166 br_166 wl_56 vdd gnd cell_6t
Xbit_r57_c166 bl_166 br_166 wl_57 vdd gnd cell_6t
Xbit_r58_c166 bl_166 br_166 wl_58 vdd gnd cell_6t
Xbit_r59_c166 bl_166 br_166 wl_59 vdd gnd cell_6t
Xbit_r60_c166 bl_166 br_166 wl_60 vdd gnd cell_6t
Xbit_r61_c166 bl_166 br_166 wl_61 vdd gnd cell_6t
Xbit_r62_c166 bl_166 br_166 wl_62 vdd gnd cell_6t
Xbit_r63_c166 bl_166 br_166 wl_63 vdd gnd cell_6t
Xbit_r64_c166 bl_166 br_166 wl_64 vdd gnd cell_6t
Xbit_r65_c166 bl_166 br_166 wl_65 vdd gnd cell_6t
Xbit_r66_c166 bl_166 br_166 wl_66 vdd gnd cell_6t
Xbit_r67_c166 bl_166 br_166 wl_67 vdd gnd cell_6t
Xbit_r68_c166 bl_166 br_166 wl_68 vdd gnd cell_6t
Xbit_r69_c166 bl_166 br_166 wl_69 vdd gnd cell_6t
Xbit_r70_c166 bl_166 br_166 wl_70 vdd gnd cell_6t
Xbit_r71_c166 bl_166 br_166 wl_71 vdd gnd cell_6t
Xbit_r72_c166 bl_166 br_166 wl_72 vdd gnd cell_6t
Xbit_r73_c166 bl_166 br_166 wl_73 vdd gnd cell_6t
Xbit_r74_c166 bl_166 br_166 wl_74 vdd gnd cell_6t
Xbit_r75_c166 bl_166 br_166 wl_75 vdd gnd cell_6t
Xbit_r76_c166 bl_166 br_166 wl_76 vdd gnd cell_6t
Xbit_r77_c166 bl_166 br_166 wl_77 vdd gnd cell_6t
Xbit_r78_c166 bl_166 br_166 wl_78 vdd gnd cell_6t
Xbit_r79_c166 bl_166 br_166 wl_79 vdd gnd cell_6t
Xbit_r80_c166 bl_166 br_166 wl_80 vdd gnd cell_6t
Xbit_r81_c166 bl_166 br_166 wl_81 vdd gnd cell_6t
Xbit_r82_c166 bl_166 br_166 wl_82 vdd gnd cell_6t
Xbit_r83_c166 bl_166 br_166 wl_83 vdd gnd cell_6t
Xbit_r84_c166 bl_166 br_166 wl_84 vdd gnd cell_6t
Xbit_r85_c166 bl_166 br_166 wl_85 vdd gnd cell_6t
Xbit_r86_c166 bl_166 br_166 wl_86 vdd gnd cell_6t
Xbit_r87_c166 bl_166 br_166 wl_87 vdd gnd cell_6t
Xbit_r88_c166 bl_166 br_166 wl_88 vdd gnd cell_6t
Xbit_r89_c166 bl_166 br_166 wl_89 vdd gnd cell_6t
Xbit_r90_c166 bl_166 br_166 wl_90 vdd gnd cell_6t
Xbit_r91_c166 bl_166 br_166 wl_91 vdd gnd cell_6t
Xbit_r92_c166 bl_166 br_166 wl_92 vdd gnd cell_6t
Xbit_r93_c166 bl_166 br_166 wl_93 vdd gnd cell_6t
Xbit_r94_c166 bl_166 br_166 wl_94 vdd gnd cell_6t
Xbit_r95_c166 bl_166 br_166 wl_95 vdd gnd cell_6t
Xbit_r96_c166 bl_166 br_166 wl_96 vdd gnd cell_6t
Xbit_r97_c166 bl_166 br_166 wl_97 vdd gnd cell_6t
Xbit_r98_c166 bl_166 br_166 wl_98 vdd gnd cell_6t
Xbit_r99_c166 bl_166 br_166 wl_99 vdd gnd cell_6t
Xbit_r100_c166 bl_166 br_166 wl_100 vdd gnd cell_6t
Xbit_r101_c166 bl_166 br_166 wl_101 vdd gnd cell_6t
Xbit_r102_c166 bl_166 br_166 wl_102 vdd gnd cell_6t
Xbit_r103_c166 bl_166 br_166 wl_103 vdd gnd cell_6t
Xbit_r104_c166 bl_166 br_166 wl_104 vdd gnd cell_6t
Xbit_r105_c166 bl_166 br_166 wl_105 vdd gnd cell_6t
Xbit_r106_c166 bl_166 br_166 wl_106 vdd gnd cell_6t
Xbit_r107_c166 bl_166 br_166 wl_107 vdd gnd cell_6t
Xbit_r108_c166 bl_166 br_166 wl_108 vdd gnd cell_6t
Xbit_r109_c166 bl_166 br_166 wl_109 vdd gnd cell_6t
Xbit_r110_c166 bl_166 br_166 wl_110 vdd gnd cell_6t
Xbit_r111_c166 bl_166 br_166 wl_111 vdd gnd cell_6t
Xbit_r112_c166 bl_166 br_166 wl_112 vdd gnd cell_6t
Xbit_r113_c166 bl_166 br_166 wl_113 vdd gnd cell_6t
Xbit_r114_c166 bl_166 br_166 wl_114 vdd gnd cell_6t
Xbit_r115_c166 bl_166 br_166 wl_115 vdd gnd cell_6t
Xbit_r116_c166 bl_166 br_166 wl_116 vdd gnd cell_6t
Xbit_r117_c166 bl_166 br_166 wl_117 vdd gnd cell_6t
Xbit_r118_c166 bl_166 br_166 wl_118 vdd gnd cell_6t
Xbit_r119_c166 bl_166 br_166 wl_119 vdd gnd cell_6t
Xbit_r120_c166 bl_166 br_166 wl_120 vdd gnd cell_6t
Xbit_r121_c166 bl_166 br_166 wl_121 vdd gnd cell_6t
Xbit_r122_c166 bl_166 br_166 wl_122 vdd gnd cell_6t
Xbit_r123_c166 bl_166 br_166 wl_123 vdd gnd cell_6t
Xbit_r124_c166 bl_166 br_166 wl_124 vdd gnd cell_6t
Xbit_r125_c166 bl_166 br_166 wl_125 vdd gnd cell_6t
Xbit_r126_c166 bl_166 br_166 wl_126 vdd gnd cell_6t
Xbit_r127_c166 bl_166 br_166 wl_127 vdd gnd cell_6t
Xbit_r128_c166 bl_166 br_166 wl_128 vdd gnd cell_6t
Xbit_r129_c166 bl_166 br_166 wl_129 vdd gnd cell_6t
Xbit_r130_c166 bl_166 br_166 wl_130 vdd gnd cell_6t
Xbit_r131_c166 bl_166 br_166 wl_131 vdd gnd cell_6t
Xbit_r132_c166 bl_166 br_166 wl_132 vdd gnd cell_6t
Xbit_r133_c166 bl_166 br_166 wl_133 vdd gnd cell_6t
Xbit_r134_c166 bl_166 br_166 wl_134 vdd gnd cell_6t
Xbit_r135_c166 bl_166 br_166 wl_135 vdd gnd cell_6t
Xbit_r136_c166 bl_166 br_166 wl_136 vdd gnd cell_6t
Xbit_r137_c166 bl_166 br_166 wl_137 vdd gnd cell_6t
Xbit_r138_c166 bl_166 br_166 wl_138 vdd gnd cell_6t
Xbit_r139_c166 bl_166 br_166 wl_139 vdd gnd cell_6t
Xbit_r140_c166 bl_166 br_166 wl_140 vdd gnd cell_6t
Xbit_r141_c166 bl_166 br_166 wl_141 vdd gnd cell_6t
Xbit_r142_c166 bl_166 br_166 wl_142 vdd gnd cell_6t
Xbit_r143_c166 bl_166 br_166 wl_143 vdd gnd cell_6t
Xbit_r144_c166 bl_166 br_166 wl_144 vdd gnd cell_6t
Xbit_r145_c166 bl_166 br_166 wl_145 vdd gnd cell_6t
Xbit_r146_c166 bl_166 br_166 wl_146 vdd gnd cell_6t
Xbit_r147_c166 bl_166 br_166 wl_147 vdd gnd cell_6t
Xbit_r148_c166 bl_166 br_166 wl_148 vdd gnd cell_6t
Xbit_r149_c166 bl_166 br_166 wl_149 vdd gnd cell_6t
Xbit_r150_c166 bl_166 br_166 wl_150 vdd gnd cell_6t
Xbit_r151_c166 bl_166 br_166 wl_151 vdd gnd cell_6t
Xbit_r152_c166 bl_166 br_166 wl_152 vdd gnd cell_6t
Xbit_r153_c166 bl_166 br_166 wl_153 vdd gnd cell_6t
Xbit_r154_c166 bl_166 br_166 wl_154 vdd gnd cell_6t
Xbit_r155_c166 bl_166 br_166 wl_155 vdd gnd cell_6t
Xbit_r156_c166 bl_166 br_166 wl_156 vdd gnd cell_6t
Xbit_r157_c166 bl_166 br_166 wl_157 vdd gnd cell_6t
Xbit_r158_c166 bl_166 br_166 wl_158 vdd gnd cell_6t
Xbit_r159_c166 bl_166 br_166 wl_159 vdd gnd cell_6t
Xbit_r160_c166 bl_166 br_166 wl_160 vdd gnd cell_6t
Xbit_r161_c166 bl_166 br_166 wl_161 vdd gnd cell_6t
Xbit_r162_c166 bl_166 br_166 wl_162 vdd gnd cell_6t
Xbit_r163_c166 bl_166 br_166 wl_163 vdd gnd cell_6t
Xbit_r164_c166 bl_166 br_166 wl_164 vdd gnd cell_6t
Xbit_r165_c166 bl_166 br_166 wl_165 vdd gnd cell_6t
Xbit_r166_c166 bl_166 br_166 wl_166 vdd gnd cell_6t
Xbit_r167_c166 bl_166 br_166 wl_167 vdd gnd cell_6t
Xbit_r168_c166 bl_166 br_166 wl_168 vdd gnd cell_6t
Xbit_r169_c166 bl_166 br_166 wl_169 vdd gnd cell_6t
Xbit_r170_c166 bl_166 br_166 wl_170 vdd gnd cell_6t
Xbit_r171_c166 bl_166 br_166 wl_171 vdd gnd cell_6t
Xbit_r172_c166 bl_166 br_166 wl_172 vdd gnd cell_6t
Xbit_r173_c166 bl_166 br_166 wl_173 vdd gnd cell_6t
Xbit_r174_c166 bl_166 br_166 wl_174 vdd gnd cell_6t
Xbit_r175_c166 bl_166 br_166 wl_175 vdd gnd cell_6t
Xbit_r176_c166 bl_166 br_166 wl_176 vdd gnd cell_6t
Xbit_r177_c166 bl_166 br_166 wl_177 vdd gnd cell_6t
Xbit_r178_c166 bl_166 br_166 wl_178 vdd gnd cell_6t
Xbit_r179_c166 bl_166 br_166 wl_179 vdd gnd cell_6t
Xbit_r180_c166 bl_166 br_166 wl_180 vdd gnd cell_6t
Xbit_r181_c166 bl_166 br_166 wl_181 vdd gnd cell_6t
Xbit_r182_c166 bl_166 br_166 wl_182 vdd gnd cell_6t
Xbit_r183_c166 bl_166 br_166 wl_183 vdd gnd cell_6t
Xbit_r184_c166 bl_166 br_166 wl_184 vdd gnd cell_6t
Xbit_r185_c166 bl_166 br_166 wl_185 vdd gnd cell_6t
Xbit_r186_c166 bl_166 br_166 wl_186 vdd gnd cell_6t
Xbit_r187_c166 bl_166 br_166 wl_187 vdd gnd cell_6t
Xbit_r188_c166 bl_166 br_166 wl_188 vdd gnd cell_6t
Xbit_r189_c166 bl_166 br_166 wl_189 vdd gnd cell_6t
Xbit_r190_c166 bl_166 br_166 wl_190 vdd gnd cell_6t
Xbit_r191_c166 bl_166 br_166 wl_191 vdd gnd cell_6t
Xbit_r192_c166 bl_166 br_166 wl_192 vdd gnd cell_6t
Xbit_r193_c166 bl_166 br_166 wl_193 vdd gnd cell_6t
Xbit_r194_c166 bl_166 br_166 wl_194 vdd gnd cell_6t
Xbit_r195_c166 bl_166 br_166 wl_195 vdd gnd cell_6t
Xbit_r196_c166 bl_166 br_166 wl_196 vdd gnd cell_6t
Xbit_r197_c166 bl_166 br_166 wl_197 vdd gnd cell_6t
Xbit_r198_c166 bl_166 br_166 wl_198 vdd gnd cell_6t
Xbit_r199_c166 bl_166 br_166 wl_199 vdd gnd cell_6t
Xbit_r200_c166 bl_166 br_166 wl_200 vdd gnd cell_6t
Xbit_r201_c166 bl_166 br_166 wl_201 vdd gnd cell_6t
Xbit_r202_c166 bl_166 br_166 wl_202 vdd gnd cell_6t
Xbit_r203_c166 bl_166 br_166 wl_203 vdd gnd cell_6t
Xbit_r204_c166 bl_166 br_166 wl_204 vdd gnd cell_6t
Xbit_r205_c166 bl_166 br_166 wl_205 vdd gnd cell_6t
Xbit_r206_c166 bl_166 br_166 wl_206 vdd gnd cell_6t
Xbit_r207_c166 bl_166 br_166 wl_207 vdd gnd cell_6t
Xbit_r208_c166 bl_166 br_166 wl_208 vdd gnd cell_6t
Xbit_r209_c166 bl_166 br_166 wl_209 vdd gnd cell_6t
Xbit_r210_c166 bl_166 br_166 wl_210 vdd gnd cell_6t
Xbit_r211_c166 bl_166 br_166 wl_211 vdd gnd cell_6t
Xbit_r212_c166 bl_166 br_166 wl_212 vdd gnd cell_6t
Xbit_r213_c166 bl_166 br_166 wl_213 vdd gnd cell_6t
Xbit_r214_c166 bl_166 br_166 wl_214 vdd gnd cell_6t
Xbit_r215_c166 bl_166 br_166 wl_215 vdd gnd cell_6t
Xbit_r216_c166 bl_166 br_166 wl_216 vdd gnd cell_6t
Xbit_r217_c166 bl_166 br_166 wl_217 vdd gnd cell_6t
Xbit_r218_c166 bl_166 br_166 wl_218 vdd gnd cell_6t
Xbit_r219_c166 bl_166 br_166 wl_219 vdd gnd cell_6t
Xbit_r220_c166 bl_166 br_166 wl_220 vdd gnd cell_6t
Xbit_r221_c166 bl_166 br_166 wl_221 vdd gnd cell_6t
Xbit_r222_c166 bl_166 br_166 wl_222 vdd gnd cell_6t
Xbit_r223_c166 bl_166 br_166 wl_223 vdd gnd cell_6t
Xbit_r224_c166 bl_166 br_166 wl_224 vdd gnd cell_6t
Xbit_r225_c166 bl_166 br_166 wl_225 vdd gnd cell_6t
Xbit_r226_c166 bl_166 br_166 wl_226 vdd gnd cell_6t
Xbit_r227_c166 bl_166 br_166 wl_227 vdd gnd cell_6t
Xbit_r228_c166 bl_166 br_166 wl_228 vdd gnd cell_6t
Xbit_r229_c166 bl_166 br_166 wl_229 vdd gnd cell_6t
Xbit_r230_c166 bl_166 br_166 wl_230 vdd gnd cell_6t
Xbit_r231_c166 bl_166 br_166 wl_231 vdd gnd cell_6t
Xbit_r232_c166 bl_166 br_166 wl_232 vdd gnd cell_6t
Xbit_r233_c166 bl_166 br_166 wl_233 vdd gnd cell_6t
Xbit_r234_c166 bl_166 br_166 wl_234 vdd gnd cell_6t
Xbit_r235_c166 bl_166 br_166 wl_235 vdd gnd cell_6t
Xbit_r236_c166 bl_166 br_166 wl_236 vdd gnd cell_6t
Xbit_r237_c166 bl_166 br_166 wl_237 vdd gnd cell_6t
Xbit_r238_c166 bl_166 br_166 wl_238 vdd gnd cell_6t
Xbit_r239_c166 bl_166 br_166 wl_239 vdd gnd cell_6t
Xbit_r240_c166 bl_166 br_166 wl_240 vdd gnd cell_6t
Xbit_r241_c166 bl_166 br_166 wl_241 vdd gnd cell_6t
Xbit_r242_c166 bl_166 br_166 wl_242 vdd gnd cell_6t
Xbit_r243_c166 bl_166 br_166 wl_243 vdd gnd cell_6t
Xbit_r244_c166 bl_166 br_166 wl_244 vdd gnd cell_6t
Xbit_r245_c166 bl_166 br_166 wl_245 vdd gnd cell_6t
Xbit_r246_c166 bl_166 br_166 wl_246 vdd gnd cell_6t
Xbit_r247_c166 bl_166 br_166 wl_247 vdd gnd cell_6t
Xbit_r248_c166 bl_166 br_166 wl_248 vdd gnd cell_6t
Xbit_r249_c166 bl_166 br_166 wl_249 vdd gnd cell_6t
Xbit_r250_c166 bl_166 br_166 wl_250 vdd gnd cell_6t
Xbit_r251_c166 bl_166 br_166 wl_251 vdd gnd cell_6t
Xbit_r252_c166 bl_166 br_166 wl_252 vdd gnd cell_6t
Xbit_r253_c166 bl_166 br_166 wl_253 vdd gnd cell_6t
Xbit_r254_c166 bl_166 br_166 wl_254 vdd gnd cell_6t
Xbit_r255_c166 bl_166 br_166 wl_255 vdd gnd cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd cell_6t
Xbit_r1_c167 bl_167 br_167 wl_1 vdd gnd cell_6t
Xbit_r2_c167 bl_167 br_167 wl_2 vdd gnd cell_6t
Xbit_r3_c167 bl_167 br_167 wl_3 vdd gnd cell_6t
Xbit_r4_c167 bl_167 br_167 wl_4 vdd gnd cell_6t
Xbit_r5_c167 bl_167 br_167 wl_5 vdd gnd cell_6t
Xbit_r6_c167 bl_167 br_167 wl_6 vdd gnd cell_6t
Xbit_r7_c167 bl_167 br_167 wl_7 vdd gnd cell_6t
Xbit_r8_c167 bl_167 br_167 wl_8 vdd gnd cell_6t
Xbit_r9_c167 bl_167 br_167 wl_9 vdd gnd cell_6t
Xbit_r10_c167 bl_167 br_167 wl_10 vdd gnd cell_6t
Xbit_r11_c167 bl_167 br_167 wl_11 vdd gnd cell_6t
Xbit_r12_c167 bl_167 br_167 wl_12 vdd gnd cell_6t
Xbit_r13_c167 bl_167 br_167 wl_13 vdd gnd cell_6t
Xbit_r14_c167 bl_167 br_167 wl_14 vdd gnd cell_6t
Xbit_r15_c167 bl_167 br_167 wl_15 vdd gnd cell_6t
Xbit_r16_c167 bl_167 br_167 wl_16 vdd gnd cell_6t
Xbit_r17_c167 bl_167 br_167 wl_17 vdd gnd cell_6t
Xbit_r18_c167 bl_167 br_167 wl_18 vdd gnd cell_6t
Xbit_r19_c167 bl_167 br_167 wl_19 vdd gnd cell_6t
Xbit_r20_c167 bl_167 br_167 wl_20 vdd gnd cell_6t
Xbit_r21_c167 bl_167 br_167 wl_21 vdd gnd cell_6t
Xbit_r22_c167 bl_167 br_167 wl_22 vdd gnd cell_6t
Xbit_r23_c167 bl_167 br_167 wl_23 vdd gnd cell_6t
Xbit_r24_c167 bl_167 br_167 wl_24 vdd gnd cell_6t
Xbit_r25_c167 bl_167 br_167 wl_25 vdd gnd cell_6t
Xbit_r26_c167 bl_167 br_167 wl_26 vdd gnd cell_6t
Xbit_r27_c167 bl_167 br_167 wl_27 vdd gnd cell_6t
Xbit_r28_c167 bl_167 br_167 wl_28 vdd gnd cell_6t
Xbit_r29_c167 bl_167 br_167 wl_29 vdd gnd cell_6t
Xbit_r30_c167 bl_167 br_167 wl_30 vdd gnd cell_6t
Xbit_r31_c167 bl_167 br_167 wl_31 vdd gnd cell_6t
Xbit_r32_c167 bl_167 br_167 wl_32 vdd gnd cell_6t
Xbit_r33_c167 bl_167 br_167 wl_33 vdd gnd cell_6t
Xbit_r34_c167 bl_167 br_167 wl_34 vdd gnd cell_6t
Xbit_r35_c167 bl_167 br_167 wl_35 vdd gnd cell_6t
Xbit_r36_c167 bl_167 br_167 wl_36 vdd gnd cell_6t
Xbit_r37_c167 bl_167 br_167 wl_37 vdd gnd cell_6t
Xbit_r38_c167 bl_167 br_167 wl_38 vdd gnd cell_6t
Xbit_r39_c167 bl_167 br_167 wl_39 vdd gnd cell_6t
Xbit_r40_c167 bl_167 br_167 wl_40 vdd gnd cell_6t
Xbit_r41_c167 bl_167 br_167 wl_41 vdd gnd cell_6t
Xbit_r42_c167 bl_167 br_167 wl_42 vdd gnd cell_6t
Xbit_r43_c167 bl_167 br_167 wl_43 vdd gnd cell_6t
Xbit_r44_c167 bl_167 br_167 wl_44 vdd gnd cell_6t
Xbit_r45_c167 bl_167 br_167 wl_45 vdd gnd cell_6t
Xbit_r46_c167 bl_167 br_167 wl_46 vdd gnd cell_6t
Xbit_r47_c167 bl_167 br_167 wl_47 vdd gnd cell_6t
Xbit_r48_c167 bl_167 br_167 wl_48 vdd gnd cell_6t
Xbit_r49_c167 bl_167 br_167 wl_49 vdd gnd cell_6t
Xbit_r50_c167 bl_167 br_167 wl_50 vdd gnd cell_6t
Xbit_r51_c167 bl_167 br_167 wl_51 vdd gnd cell_6t
Xbit_r52_c167 bl_167 br_167 wl_52 vdd gnd cell_6t
Xbit_r53_c167 bl_167 br_167 wl_53 vdd gnd cell_6t
Xbit_r54_c167 bl_167 br_167 wl_54 vdd gnd cell_6t
Xbit_r55_c167 bl_167 br_167 wl_55 vdd gnd cell_6t
Xbit_r56_c167 bl_167 br_167 wl_56 vdd gnd cell_6t
Xbit_r57_c167 bl_167 br_167 wl_57 vdd gnd cell_6t
Xbit_r58_c167 bl_167 br_167 wl_58 vdd gnd cell_6t
Xbit_r59_c167 bl_167 br_167 wl_59 vdd gnd cell_6t
Xbit_r60_c167 bl_167 br_167 wl_60 vdd gnd cell_6t
Xbit_r61_c167 bl_167 br_167 wl_61 vdd gnd cell_6t
Xbit_r62_c167 bl_167 br_167 wl_62 vdd gnd cell_6t
Xbit_r63_c167 bl_167 br_167 wl_63 vdd gnd cell_6t
Xbit_r64_c167 bl_167 br_167 wl_64 vdd gnd cell_6t
Xbit_r65_c167 bl_167 br_167 wl_65 vdd gnd cell_6t
Xbit_r66_c167 bl_167 br_167 wl_66 vdd gnd cell_6t
Xbit_r67_c167 bl_167 br_167 wl_67 vdd gnd cell_6t
Xbit_r68_c167 bl_167 br_167 wl_68 vdd gnd cell_6t
Xbit_r69_c167 bl_167 br_167 wl_69 vdd gnd cell_6t
Xbit_r70_c167 bl_167 br_167 wl_70 vdd gnd cell_6t
Xbit_r71_c167 bl_167 br_167 wl_71 vdd gnd cell_6t
Xbit_r72_c167 bl_167 br_167 wl_72 vdd gnd cell_6t
Xbit_r73_c167 bl_167 br_167 wl_73 vdd gnd cell_6t
Xbit_r74_c167 bl_167 br_167 wl_74 vdd gnd cell_6t
Xbit_r75_c167 bl_167 br_167 wl_75 vdd gnd cell_6t
Xbit_r76_c167 bl_167 br_167 wl_76 vdd gnd cell_6t
Xbit_r77_c167 bl_167 br_167 wl_77 vdd gnd cell_6t
Xbit_r78_c167 bl_167 br_167 wl_78 vdd gnd cell_6t
Xbit_r79_c167 bl_167 br_167 wl_79 vdd gnd cell_6t
Xbit_r80_c167 bl_167 br_167 wl_80 vdd gnd cell_6t
Xbit_r81_c167 bl_167 br_167 wl_81 vdd gnd cell_6t
Xbit_r82_c167 bl_167 br_167 wl_82 vdd gnd cell_6t
Xbit_r83_c167 bl_167 br_167 wl_83 vdd gnd cell_6t
Xbit_r84_c167 bl_167 br_167 wl_84 vdd gnd cell_6t
Xbit_r85_c167 bl_167 br_167 wl_85 vdd gnd cell_6t
Xbit_r86_c167 bl_167 br_167 wl_86 vdd gnd cell_6t
Xbit_r87_c167 bl_167 br_167 wl_87 vdd gnd cell_6t
Xbit_r88_c167 bl_167 br_167 wl_88 vdd gnd cell_6t
Xbit_r89_c167 bl_167 br_167 wl_89 vdd gnd cell_6t
Xbit_r90_c167 bl_167 br_167 wl_90 vdd gnd cell_6t
Xbit_r91_c167 bl_167 br_167 wl_91 vdd gnd cell_6t
Xbit_r92_c167 bl_167 br_167 wl_92 vdd gnd cell_6t
Xbit_r93_c167 bl_167 br_167 wl_93 vdd gnd cell_6t
Xbit_r94_c167 bl_167 br_167 wl_94 vdd gnd cell_6t
Xbit_r95_c167 bl_167 br_167 wl_95 vdd gnd cell_6t
Xbit_r96_c167 bl_167 br_167 wl_96 vdd gnd cell_6t
Xbit_r97_c167 bl_167 br_167 wl_97 vdd gnd cell_6t
Xbit_r98_c167 bl_167 br_167 wl_98 vdd gnd cell_6t
Xbit_r99_c167 bl_167 br_167 wl_99 vdd gnd cell_6t
Xbit_r100_c167 bl_167 br_167 wl_100 vdd gnd cell_6t
Xbit_r101_c167 bl_167 br_167 wl_101 vdd gnd cell_6t
Xbit_r102_c167 bl_167 br_167 wl_102 vdd gnd cell_6t
Xbit_r103_c167 bl_167 br_167 wl_103 vdd gnd cell_6t
Xbit_r104_c167 bl_167 br_167 wl_104 vdd gnd cell_6t
Xbit_r105_c167 bl_167 br_167 wl_105 vdd gnd cell_6t
Xbit_r106_c167 bl_167 br_167 wl_106 vdd gnd cell_6t
Xbit_r107_c167 bl_167 br_167 wl_107 vdd gnd cell_6t
Xbit_r108_c167 bl_167 br_167 wl_108 vdd gnd cell_6t
Xbit_r109_c167 bl_167 br_167 wl_109 vdd gnd cell_6t
Xbit_r110_c167 bl_167 br_167 wl_110 vdd gnd cell_6t
Xbit_r111_c167 bl_167 br_167 wl_111 vdd gnd cell_6t
Xbit_r112_c167 bl_167 br_167 wl_112 vdd gnd cell_6t
Xbit_r113_c167 bl_167 br_167 wl_113 vdd gnd cell_6t
Xbit_r114_c167 bl_167 br_167 wl_114 vdd gnd cell_6t
Xbit_r115_c167 bl_167 br_167 wl_115 vdd gnd cell_6t
Xbit_r116_c167 bl_167 br_167 wl_116 vdd gnd cell_6t
Xbit_r117_c167 bl_167 br_167 wl_117 vdd gnd cell_6t
Xbit_r118_c167 bl_167 br_167 wl_118 vdd gnd cell_6t
Xbit_r119_c167 bl_167 br_167 wl_119 vdd gnd cell_6t
Xbit_r120_c167 bl_167 br_167 wl_120 vdd gnd cell_6t
Xbit_r121_c167 bl_167 br_167 wl_121 vdd gnd cell_6t
Xbit_r122_c167 bl_167 br_167 wl_122 vdd gnd cell_6t
Xbit_r123_c167 bl_167 br_167 wl_123 vdd gnd cell_6t
Xbit_r124_c167 bl_167 br_167 wl_124 vdd gnd cell_6t
Xbit_r125_c167 bl_167 br_167 wl_125 vdd gnd cell_6t
Xbit_r126_c167 bl_167 br_167 wl_126 vdd gnd cell_6t
Xbit_r127_c167 bl_167 br_167 wl_127 vdd gnd cell_6t
Xbit_r128_c167 bl_167 br_167 wl_128 vdd gnd cell_6t
Xbit_r129_c167 bl_167 br_167 wl_129 vdd gnd cell_6t
Xbit_r130_c167 bl_167 br_167 wl_130 vdd gnd cell_6t
Xbit_r131_c167 bl_167 br_167 wl_131 vdd gnd cell_6t
Xbit_r132_c167 bl_167 br_167 wl_132 vdd gnd cell_6t
Xbit_r133_c167 bl_167 br_167 wl_133 vdd gnd cell_6t
Xbit_r134_c167 bl_167 br_167 wl_134 vdd gnd cell_6t
Xbit_r135_c167 bl_167 br_167 wl_135 vdd gnd cell_6t
Xbit_r136_c167 bl_167 br_167 wl_136 vdd gnd cell_6t
Xbit_r137_c167 bl_167 br_167 wl_137 vdd gnd cell_6t
Xbit_r138_c167 bl_167 br_167 wl_138 vdd gnd cell_6t
Xbit_r139_c167 bl_167 br_167 wl_139 vdd gnd cell_6t
Xbit_r140_c167 bl_167 br_167 wl_140 vdd gnd cell_6t
Xbit_r141_c167 bl_167 br_167 wl_141 vdd gnd cell_6t
Xbit_r142_c167 bl_167 br_167 wl_142 vdd gnd cell_6t
Xbit_r143_c167 bl_167 br_167 wl_143 vdd gnd cell_6t
Xbit_r144_c167 bl_167 br_167 wl_144 vdd gnd cell_6t
Xbit_r145_c167 bl_167 br_167 wl_145 vdd gnd cell_6t
Xbit_r146_c167 bl_167 br_167 wl_146 vdd gnd cell_6t
Xbit_r147_c167 bl_167 br_167 wl_147 vdd gnd cell_6t
Xbit_r148_c167 bl_167 br_167 wl_148 vdd gnd cell_6t
Xbit_r149_c167 bl_167 br_167 wl_149 vdd gnd cell_6t
Xbit_r150_c167 bl_167 br_167 wl_150 vdd gnd cell_6t
Xbit_r151_c167 bl_167 br_167 wl_151 vdd gnd cell_6t
Xbit_r152_c167 bl_167 br_167 wl_152 vdd gnd cell_6t
Xbit_r153_c167 bl_167 br_167 wl_153 vdd gnd cell_6t
Xbit_r154_c167 bl_167 br_167 wl_154 vdd gnd cell_6t
Xbit_r155_c167 bl_167 br_167 wl_155 vdd gnd cell_6t
Xbit_r156_c167 bl_167 br_167 wl_156 vdd gnd cell_6t
Xbit_r157_c167 bl_167 br_167 wl_157 vdd gnd cell_6t
Xbit_r158_c167 bl_167 br_167 wl_158 vdd gnd cell_6t
Xbit_r159_c167 bl_167 br_167 wl_159 vdd gnd cell_6t
Xbit_r160_c167 bl_167 br_167 wl_160 vdd gnd cell_6t
Xbit_r161_c167 bl_167 br_167 wl_161 vdd gnd cell_6t
Xbit_r162_c167 bl_167 br_167 wl_162 vdd gnd cell_6t
Xbit_r163_c167 bl_167 br_167 wl_163 vdd gnd cell_6t
Xbit_r164_c167 bl_167 br_167 wl_164 vdd gnd cell_6t
Xbit_r165_c167 bl_167 br_167 wl_165 vdd gnd cell_6t
Xbit_r166_c167 bl_167 br_167 wl_166 vdd gnd cell_6t
Xbit_r167_c167 bl_167 br_167 wl_167 vdd gnd cell_6t
Xbit_r168_c167 bl_167 br_167 wl_168 vdd gnd cell_6t
Xbit_r169_c167 bl_167 br_167 wl_169 vdd gnd cell_6t
Xbit_r170_c167 bl_167 br_167 wl_170 vdd gnd cell_6t
Xbit_r171_c167 bl_167 br_167 wl_171 vdd gnd cell_6t
Xbit_r172_c167 bl_167 br_167 wl_172 vdd gnd cell_6t
Xbit_r173_c167 bl_167 br_167 wl_173 vdd gnd cell_6t
Xbit_r174_c167 bl_167 br_167 wl_174 vdd gnd cell_6t
Xbit_r175_c167 bl_167 br_167 wl_175 vdd gnd cell_6t
Xbit_r176_c167 bl_167 br_167 wl_176 vdd gnd cell_6t
Xbit_r177_c167 bl_167 br_167 wl_177 vdd gnd cell_6t
Xbit_r178_c167 bl_167 br_167 wl_178 vdd gnd cell_6t
Xbit_r179_c167 bl_167 br_167 wl_179 vdd gnd cell_6t
Xbit_r180_c167 bl_167 br_167 wl_180 vdd gnd cell_6t
Xbit_r181_c167 bl_167 br_167 wl_181 vdd gnd cell_6t
Xbit_r182_c167 bl_167 br_167 wl_182 vdd gnd cell_6t
Xbit_r183_c167 bl_167 br_167 wl_183 vdd gnd cell_6t
Xbit_r184_c167 bl_167 br_167 wl_184 vdd gnd cell_6t
Xbit_r185_c167 bl_167 br_167 wl_185 vdd gnd cell_6t
Xbit_r186_c167 bl_167 br_167 wl_186 vdd gnd cell_6t
Xbit_r187_c167 bl_167 br_167 wl_187 vdd gnd cell_6t
Xbit_r188_c167 bl_167 br_167 wl_188 vdd gnd cell_6t
Xbit_r189_c167 bl_167 br_167 wl_189 vdd gnd cell_6t
Xbit_r190_c167 bl_167 br_167 wl_190 vdd gnd cell_6t
Xbit_r191_c167 bl_167 br_167 wl_191 vdd gnd cell_6t
Xbit_r192_c167 bl_167 br_167 wl_192 vdd gnd cell_6t
Xbit_r193_c167 bl_167 br_167 wl_193 vdd gnd cell_6t
Xbit_r194_c167 bl_167 br_167 wl_194 vdd gnd cell_6t
Xbit_r195_c167 bl_167 br_167 wl_195 vdd gnd cell_6t
Xbit_r196_c167 bl_167 br_167 wl_196 vdd gnd cell_6t
Xbit_r197_c167 bl_167 br_167 wl_197 vdd gnd cell_6t
Xbit_r198_c167 bl_167 br_167 wl_198 vdd gnd cell_6t
Xbit_r199_c167 bl_167 br_167 wl_199 vdd gnd cell_6t
Xbit_r200_c167 bl_167 br_167 wl_200 vdd gnd cell_6t
Xbit_r201_c167 bl_167 br_167 wl_201 vdd gnd cell_6t
Xbit_r202_c167 bl_167 br_167 wl_202 vdd gnd cell_6t
Xbit_r203_c167 bl_167 br_167 wl_203 vdd gnd cell_6t
Xbit_r204_c167 bl_167 br_167 wl_204 vdd gnd cell_6t
Xbit_r205_c167 bl_167 br_167 wl_205 vdd gnd cell_6t
Xbit_r206_c167 bl_167 br_167 wl_206 vdd gnd cell_6t
Xbit_r207_c167 bl_167 br_167 wl_207 vdd gnd cell_6t
Xbit_r208_c167 bl_167 br_167 wl_208 vdd gnd cell_6t
Xbit_r209_c167 bl_167 br_167 wl_209 vdd gnd cell_6t
Xbit_r210_c167 bl_167 br_167 wl_210 vdd gnd cell_6t
Xbit_r211_c167 bl_167 br_167 wl_211 vdd gnd cell_6t
Xbit_r212_c167 bl_167 br_167 wl_212 vdd gnd cell_6t
Xbit_r213_c167 bl_167 br_167 wl_213 vdd gnd cell_6t
Xbit_r214_c167 bl_167 br_167 wl_214 vdd gnd cell_6t
Xbit_r215_c167 bl_167 br_167 wl_215 vdd gnd cell_6t
Xbit_r216_c167 bl_167 br_167 wl_216 vdd gnd cell_6t
Xbit_r217_c167 bl_167 br_167 wl_217 vdd gnd cell_6t
Xbit_r218_c167 bl_167 br_167 wl_218 vdd gnd cell_6t
Xbit_r219_c167 bl_167 br_167 wl_219 vdd gnd cell_6t
Xbit_r220_c167 bl_167 br_167 wl_220 vdd gnd cell_6t
Xbit_r221_c167 bl_167 br_167 wl_221 vdd gnd cell_6t
Xbit_r222_c167 bl_167 br_167 wl_222 vdd gnd cell_6t
Xbit_r223_c167 bl_167 br_167 wl_223 vdd gnd cell_6t
Xbit_r224_c167 bl_167 br_167 wl_224 vdd gnd cell_6t
Xbit_r225_c167 bl_167 br_167 wl_225 vdd gnd cell_6t
Xbit_r226_c167 bl_167 br_167 wl_226 vdd gnd cell_6t
Xbit_r227_c167 bl_167 br_167 wl_227 vdd gnd cell_6t
Xbit_r228_c167 bl_167 br_167 wl_228 vdd gnd cell_6t
Xbit_r229_c167 bl_167 br_167 wl_229 vdd gnd cell_6t
Xbit_r230_c167 bl_167 br_167 wl_230 vdd gnd cell_6t
Xbit_r231_c167 bl_167 br_167 wl_231 vdd gnd cell_6t
Xbit_r232_c167 bl_167 br_167 wl_232 vdd gnd cell_6t
Xbit_r233_c167 bl_167 br_167 wl_233 vdd gnd cell_6t
Xbit_r234_c167 bl_167 br_167 wl_234 vdd gnd cell_6t
Xbit_r235_c167 bl_167 br_167 wl_235 vdd gnd cell_6t
Xbit_r236_c167 bl_167 br_167 wl_236 vdd gnd cell_6t
Xbit_r237_c167 bl_167 br_167 wl_237 vdd gnd cell_6t
Xbit_r238_c167 bl_167 br_167 wl_238 vdd gnd cell_6t
Xbit_r239_c167 bl_167 br_167 wl_239 vdd gnd cell_6t
Xbit_r240_c167 bl_167 br_167 wl_240 vdd gnd cell_6t
Xbit_r241_c167 bl_167 br_167 wl_241 vdd gnd cell_6t
Xbit_r242_c167 bl_167 br_167 wl_242 vdd gnd cell_6t
Xbit_r243_c167 bl_167 br_167 wl_243 vdd gnd cell_6t
Xbit_r244_c167 bl_167 br_167 wl_244 vdd gnd cell_6t
Xbit_r245_c167 bl_167 br_167 wl_245 vdd gnd cell_6t
Xbit_r246_c167 bl_167 br_167 wl_246 vdd gnd cell_6t
Xbit_r247_c167 bl_167 br_167 wl_247 vdd gnd cell_6t
Xbit_r248_c167 bl_167 br_167 wl_248 vdd gnd cell_6t
Xbit_r249_c167 bl_167 br_167 wl_249 vdd gnd cell_6t
Xbit_r250_c167 bl_167 br_167 wl_250 vdd gnd cell_6t
Xbit_r251_c167 bl_167 br_167 wl_251 vdd gnd cell_6t
Xbit_r252_c167 bl_167 br_167 wl_252 vdd gnd cell_6t
Xbit_r253_c167 bl_167 br_167 wl_253 vdd gnd cell_6t
Xbit_r254_c167 bl_167 br_167 wl_254 vdd gnd cell_6t
Xbit_r255_c167 bl_167 br_167 wl_255 vdd gnd cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd cell_6t
Xbit_r1_c168 bl_168 br_168 wl_1 vdd gnd cell_6t
Xbit_r2_c168 bl_168 br_168 wl_2 vdd gnd cell_6t
Xbit_r3_c168 bl_168 br_168 wl_3 vdd gnd cell_6t
Xbit_r4_c168 bl_168 br_168 wl_4 vdd gnd cell_6t
Xbit_r5_c168 bl_168 br_168 wl_5 vdd gnd cell_6t
Xbit_r6_c168 bl_168 br_168 wl_6 vdd gnd cell_6t
Xbit_r7_c168 bl_168 br_168 wl_7 vdd gnd cell_6t
Xbit_r8_c168 bl_168 br_168 wl_8 vdd gnd cell_6t
Xbit_r9_c168 bl_168 br_168 wl_9 vdd gnd cell_6t
Xbit_r10_c168 bl_168 br_168 wl_10 vdd gnd cell_6t
Xbit_r11_c168 bl_168 br_168 wl_11 vdd gnd cell_6t
Xbit_r12_c168 bl_168 br_168 wl_12 vdd gnd cell_6t
Xbit_r13_c168 bl_168 br_168 wl_13 vdd gnd cell_6t
Xbit_r14_c168 bl_168 br_168 wl_14 vdd gnd cell_6t
Xbit_r15_c168 bl_168 br_168 wl_15 vdd gnd cell_6t
Xbit_r16_c168 bl_168 br_168 wl_16 vdd gnd cell_6t
Xbit_r17_c168 bl_168 br_168 wl_17 vdd gnd cell_6t
Xbit_r18_c168 bl_168 br_168 wl_18 vdd gnd cell_6t
Xbit_r19_c168 bl_168 br_168 wl_19 vdd gnd cell_6t
Xbit_r20_c168 bl_168 br_168 wl_20 vdd gnd cell_6t
Xbit_r21_c168 bl_168 br_168 wl_21 vdd gnd cell_6t
Xbit_r22_c168 bl_168 br_168 wl_22 vdd gnd cell_6t
Xbit_r23_c168 bl_168 br_168 wl_23 vdd gnd cell_6t
Xbit_r24_c168 bl_168 br_168 wl_24 vdd gnd cell_6t
Xbit_r25_c168 bl_168 br_168 wl_25 vdd gnd cell_6t
Xbit_r26_c168 bl_168 br_168 wl_26 vdd gnd cell_6t
Xbit_r27_c168 bl_168 br_168 wl_27 vdd gnd cell_6t
Xbit_r28_c168 bl_168 br_168 wl_28 vdd gnd cell_6t
Xbit_r29_c168 bl_168 br_168 wl_29 vdd gnd cell_6t
Xbit_r30_c168 bl_168 br_168 wl_30 vdd gnd cell_6t
Xbit_r31_c168 bl_168 br_168 wl_31 vdd gnd cell_6t
Xbit_r32_c168 bl_168 br_168 wl_32 vdd gnd cell_6t
Xbit_r33_c168 bl_168 br_168 wl_33 vdd gnd cell_6t
Xbit_r34_c168 bl_168 br_168 wl_34 vdd gnd cell_6t
Xbit_r35_c168 bl_168 br_168 wl_35 vdd gnd cell_6t
Xbit_r36_c168 bl_168 br_168 wl_36 vdd gnd cell_6t
Xbit_r37_c168 bl_168 br_168 wl_37 vdd gnd cell_6t
Xbit_r38_c168 bl_168 br_168 wl_38 vdd gnd cell_6t
Xbit_r39_c168 bl_168 br_168 wl_39 vdd gnd cell_6t
Xbit_r40_c168 bl_168 br_168 wl_40 vdd gnd cell_6t
Xbit_r41_c168 bl_168 br_168 wl_41 vdd gnd cell_6t
Xbit_r42_c168 bl_168 br_168 wl_42 vdd gnd cell_6t
Xbit_r43_c168 bl_168 br_168 wl_43 vdd gnd cell_6t
Xbit_r44_c168 bl_168 br_168 wl_44 vdd gnd cell_6t
Xbit_r45_c168 bl_168 br_168 wl_45 vdd gnd cell_6t
Xbit_r46_c168 bl_168 br_168 wl_46 vdd gnd cell_6t
Xbit_r47_c168 bl_168 br_168 wl_47 vdd gnd cell_6t
Xbit_r48_c168 bl_168 br_168 wl_48 vdd gnd cell_6t
Xbit_r49_c168 bl_168 br_168 wl_49 vdd gnd cell_6t
Xbit_r50_c168 bl_168 br_168 wl_50 vdd gnd cell_6t
Xbit_r51_c168 bl_168 br_168 wl_51 vdd gnd cell_6t
Xbit_r52_c168 bl_168 br_168 wl_52 vdd gnd cell_6t
Xbit_r53_c168 bl_168 br_168 wl_53 vdd gnd cell_6t
Xbit_r54_c168 bl_168 br_168 wl_54 vdd gnd cell_6t
Xbit_r55_c168 bl_168 br_168 wl_55 vdd gnd cell_6t
Xbit_r56_c168 bl_168 br_168 wl_56 vdd gnd cell_6t
Xbit_r57_c168 bl_168 br_168 wl_57 vdd gnd cell_6t
Xbit_r58_c168 bl_168 br_168 wl_58 vdd gnd cell_6t
Xbit_r59_c168 bl_168 br_168 wl_59 vdd gnd cell_6t
Xbit_r60_c168 bl_168 br_168 wl_60 vdd gnd cell_6t
Xbit_r61_c168 bl_168 br_168 wl_61 vdd gnd cell_6t
Xbit_r62_c168 bl_168 br_168 wl_62 vdd gnd cell_6t
Xbit_r63_c168 bl_168 br_168 wl_63 vdd gnd cell_6t
Xbit_r64_c168 bl_168 br_168 wl_64 vdd gnd cell_6t
Xbit_r65_c168 bl_168 br_168 wl_65 vdd gnd cell_6t
Xbit_r66_c168 bl_168 br_168 wl_66 vdd gnd cell_6t
Xbit_r67_c168 bl_168 br_168 wl_67 vdd gnd cell_6t
Xbit_r68_c168 bl_168 br_168 wl_68 vdd gnd cell_6t
Xbit_r69_c168 bl_168 br_168 wl_69 vdd gnd cell_6t
Xbit_r70_c168 bl_168 br_168 wl_70 vdd gnd cell_6t
Xbit_r71_c168 bl_168 br_168 wl_71 vdd gnd cell_6t
Xbit_r72_c168 bl_168 br_168 wl_72 vdd gnd cell_6t
Xbit_r73_c168 bl_168 br_168 wl_73 vdd gnd cell_6t
Xbit_r74_c168 bl_168 br_168 wl_74 vdd gnd cell_6t
Xbit_r75_c168 bl_168 br_168 wl_75 vdd gnd cell_6t
Xbit_r76_c168 bl_168 br_168 wl_76 vdd gnd cell_6t
Xbit_r77_c168 bl_168 br_168 wl_77 vdd gnd cell_6t
Xbit_r78_c168 bl_168 br_168 wl_78 vdd gnd cell_6t
Xbit_r79_c168 bl_168 br_168 wl_79 vdd gnd cell_6t
Xbit_r80_c168 bl_168 br_168 wl_80 vdd gnd cell_6t
Xbit_r81_c168 bl_168 br_168 wl_81 vdd gnd cell_6t
Xbit_r82_c168 bl_168 br_168 wl_82 vdd gnd cell_6t
Xbit_r83_c168 bl_168 br_168 wl_83 vdd gnd cell_6t
Xbit_r84_c168 bl_168 br_168 wl_84 vdd gnd cell_6t
Xbit_r85_c168 bl_168 br_168 wl_85 vdd gnd cell_6t
Xbit_r86_c168 bl_168 br_168 wl_86 vdd gnd cell_6t
Xbit_r87_c168 bl_168 br_168 wl_87 vdd gnd cell_6t
Xbit_r88_c168 bl_168 br_168 wl_88 vdd gnd cell_6t
Xbit_r89_c168 bl_168 br_168 wl_89 vdd gnd cell_6t
Xbit_r90_c168 bl_168 br_168 wl_90 vdd gnd cell_6t
Xbit_r91_c168 bl_168 br_168 wl_91 vdd gnd cell_6t
Xbit_r92_c168 bl_168 br_168 wl_92 vdd gnd cell_6t
Xbit_r93_c168 bl_168 br_168 wl_93 vdd gnd cell_6t
Xbit_r94_c168 bl_168 br_168 wl_94 vdd gnd cell_6t
Xbit_r95_c168 bl_168 br_168 wl_95 vdd gnd cell_6t
Xbit_r96_c168 bl_168 br_168 wl_96 vdd gnd cell_6t
Xbit_r97_c168 bl_168 br_168 wl_97 vdd gnd cell_6t
Xbit_r98_c168 bl_168 br_168 wl_98 vdd gnd cell_6t
Xbit_r99_c168 bl_168 br_168 wl_99 vdd gnd cell_6t
Xbit_r100_c168 bl_168 br_168 wl_100 vdd gnd cell_6t
Xbit_r101_c168 bl_168 br_168 wl_101 vdd gnd cell_6t
Xbit_r102_c168 bl_168 br_168 wl_102 vdd gnd cell_6t
Xbit_r103_c168 bl_168 br_168 wl_103 vdd gnd cell_6t
Xbit_r104_c168 bl_168 br_168 wl_104 vdd gnd cell_6t
Xbit_r105_c168 bl_168 br_168 wl_105 vdd gnd cell_6t
Xbit_r106_c168 bl_168 br_168 wl_106 vdd gnd cell_6t
Xbit_r107_c168 bl_168 br_168 wl_107 vdd gnd cell_6t
Xbit_r108_c168 bl_168 br_168 wl_108 vdd gnd cell_6t
Xbit_r109_c168 bl_168 br_168 wl_109 vdd gnd cell_6t
Xbit_r110_c168 bl_168 br_168 wl_110 vdd gnd cell_6t
Xbit_r111_c168 bl_168 br_168 wl_111 vdd gnd cell_6t
Xbit_r112_c168 bl_168 br_168 wl_112 vdd gnd cell_6t
Xbit_r113_c168 bl_168 br_168 wl_113 vdd gnd cell_6t
Xbit_r114_c168 bl_168 br_168 wl_114 vdd gnd cell_6t
Xbit_r115_c168 bl_168 br_168 wl_115 vdd gnd cell_6t
Xbit_r116_c168 bl_168 br_168 wl_116 vdd gnd cell_6t
Xbit_r117_c168 bl_168 br_168 wl_117 vdd gnd cell_6t
Xbit_r118_c168 bl_168 br_168 wl_118 vdd gnd cell_6t
Xbit_r119_c168 bl_168 br_168 wl_119 vdd gnd cell_6t
Xbit_r120_c168 bl_168 br_168 wl_120 vdd gnd cell_6t
Xbit_r121_c168 bl_168 br_168 wl_121 vdd gnd cell_6t
Xbit_r122_c168 bl_168 br_168 wl_122 vdd gnd cell_6t
Xbit_r123_c168 bl_168 br_168 wl_123 vdd gnd cell_6t
Xbit_r124_c168 bl_168 br_168 wl_124 vdd gnd cell_6t
Xbit_r125_c168 bl_168 br_168 wl_125 vdd gnd cell_6t
Xbit_r126_c168 bl_168 br_168 wl_126 vdd gnd cell_6t
Xbit_r127_c168 bl_168 br_168 wl_127 vdd gnd cell_6t
Xbit_r128_c168 bl_168 br_168 wl_128 vdd gnd cell_6t
Xbit_r129_c168 bl_168 br_168 wl_129 vdd gnd cell_6t
Xbit_r130_c168 bl_168 br_168 wl_130 vdd gnd cell_6t
Xbit_r131_c168 bl_168 br_168 wl_131 vdd gnd cell_6t
Xbit_r132_c168 bl_168 br_168 wl_132 vdd gnd cell_6t
Xbit_r133_c168 bl_168 br_168 wl_133 vdd gnd cell_6t
Xbit_r134_c168 bl_168 br_168 wl_134 vdd gnd cell_6t
Xbit_r135_c168 bl_168 br_168 wl_135 vdd gnd cell_6t
Xbit_r136_c168 bl_168 br_168 wl_136 vdd gnd cell_6t
Xbit_r137_c168 bl_168 br_168 wl_137 vdd gnd cell_6t
Xbit_r138_c168 bl_168 br_168 wl_138 vdd gnd cell_6t
Xbit_r139_c168 bl_168 br_168 wl_139 vdd gnd cell_6t
Xbit_r140_c168 bl_168 br_168 wl_140 vdd gnd cell_6t
Xbit_r141_c168 bl_168 br_168 wl_141 vdd gnd cell_6t
Xbit_r142_c168 bl_168 br_168 wl_142 vdd gnd cell_6t
Xbit_r143_c168 bl_168 br_168 wl_143 vdd gnd cell_6t
Xbit_r144_c168 bl_168 br_168 wl_144 vdd gnd cell_6t
Xbit_r145_c168 bl_168 br_168 wl_145 vdd gnd cell_6t
Xbit_r146_c168 bl_168 br_168 wl_146 vdd gnd cell_6t
Xbit_r147_c168 bl_168 br_168 wl_147 vdd gnd cell_6t
Xbit_r148_c168 bl_168 br_168 wl_148 vdd gnd cell_6t
Xbit_r149_c168 bl_168 br_168 wl_149 vdd gnd cell_6t
Xbit_r150_c168 bl_168 br_168 wl_150 vdd gnd cell_6t
Xbit_r151_c168 bl_168 br_168 wl_151 vdd gnd cell_6t
Xbit_r152_c168 bl_168 br_168 wl_152 vdd gnd cell_6t
Xbit_r153_c168 bl_168 br_168 wl_153 vdd gnd cell_6t
Xbit_r154_c168 bl_168 br_168 wl_154 vdd gnd cell_6t
Xbit_r155_c168 bl_168 br_168 wl_155 vdd gnd cell_6t
Xbit_r156_c168 bl_168 br_168 wl_156 vdd gnd cell_6t
Xbit_r157_c168 bl_168 br_168 wl_157 vdd gnd cell_6t
Xbit_r158_c168 bl_168 br_168 wl_158 vdd gnd cell_6t
Xbit_r159_c168 bl_168 br_168 wl_159 vdd gnd cell_6t
Xbit_r160_c168 bl_168 br_168 wl_160 vdd gnd cell_6t
Xbit_r161_c168 bl_168 br_168 wl_161 vdd gnd cell_6t
Xbit_r162_c168 bl_168 br_168 wl_162 vdd gnd cell_6t
Xbit_r163_c168 bl_168 br_168 wl_163 vdd gnd cell_6t
Xbit_r164_c168 bl_168 br_168 wl_164 vdd gnd cell_6t
Xbit_r165_c168 bl_168 br_168 wl_165 vdd gnd cell_6t
Xbit_r166_c168 bl_168 br_168 wl_166 vdd gnd cell_6t
Xbit_r167_c168 bl_168 br_168 wl_167 vdd gnd cell_6t
Xbit_r168_c168 bl_168 br_168 wl_168 vdd gnd cell_6t
Xbit_r169_c168 bl_168 br_168 wl_169 vdd gnd cell_6t
Xbit_r170_c168 bl_168 br_168 wl_170 vdd gnd cell_6t
Xbit_r171_c168 bl_168 br_168 wl_171 vdd gnd cell_6t
Xbit_r172_c168 bl_168 br_168 wl_172 vdd gnd cell_6t
Xbit_r173_c168 bl_168 br_168 wl_173 vdd gnd cell_6t
Xbit_r174_c168 bl_168 br_168 wl_174 vdd gnd cell_6t
Xbit_r175_c168 bl_168 br_168 wl_175 vdd gnd cell_6t
Xbit_r176_c168 bl_168 br_168 wl_176 vdd gnd cell_6t
Xbit_r177_c168 bl_168 br_168 wl_177 vdd gnd cell_6t
Xbit_r178_c168 bl_168 br_168 wl_178 vdd gnd cell_6t
Xbit_r179_c168 bl_168 br_168 wl_179 vdd gnd cell_6t
Xbit_r180_c168 bl_168 br_168 wl_180 vdd gnd cell_6t
Xbit_r181_c168 bl_168 br_168 wl_181 vdd gnd cell_6t
Xbit_r182_c168 bl_168 br_168 wl_182 vdd gnd cell_6t
Xbit_r183_c168 bl_168 br_168 wl_183 vdd gnd cell_6t
Xbit_r184_c168 bl_168 br_168 wl_184 vdd gnd cell_6t
Xbit_r185_c168 bl_168 br_168 wl_185 vdd gnd cell_6t
Xbit_r186_c168 bl_168 br_168 wl_186 vdd gnd cell_6t
Xbit_r187_c168 bl_168 br_168 wl_187 vdd gnd cell_6t
Xbit_r188_c168 bl_168 br_168 wl_188 vdd gnd cell_6t
Xbit_r189_c168 bl_168 br_168 wl_189 vdd gnd cell_6t
Xbit_r190_c168 bl_168 br_168 wl_190 vdd gnd cell_6t
Xbit_r191_c168 bl_168 br_168 wl_191 vdd gnd cell_6t
Xbit_r192_c168 bl_168 br_168 wl_192 vdd gnd cell_6t
Xbit_r193_c168 bl_168 br_168 wl_193 vdd gnd cell_6t
Xbit_r194_c168 bl_168 br_168 wl_194 vdd gnd cell_6t
Xbit_r195_c168 bl_168 br_168 wl_195 vdd gnd cell_6t
Xbit_r196_c168 bl_168 br_168 wl_196 vdd gnd cell_6t
Xbit_r197_c168 bl_168 br_168 wl_197 vdd gnd cell_6t
Xbit_r198_c168 bl_168 br_168 wl_198 vdd gnd cell_6t
Xbit_r199_c168 bl_168 br_168 wl_199 vdd gnd cell_6t
Xbit_r200_c168 bl_168 br_168 wl_200 vdd gnd cell_6t
Xbit_r201_c168 bl_168 br_168 wl_201 vdd gnd cell_6t
Xbit_r202_c168 bl_168 br_168 wl_202 vdd gnd cell_6t
Xbit_r203_c168 bl_168 br_168 wl_203 vdd gnd cell_6t
Xbit_r204_c168 bl_168 br_168 wl_204 vdd gnd cell_6t
Xbit_r205_c168 bl_168 br_168 wl_205 vdd gnd cell_6t
Xbit_r206_c168 bl_168 br_168 wl_206 vdd gnd cell_6t
Xbit_r207_c168 bl_168 br_168 wl_207 vdd gnd cell_6t
Xbit_r208_c168 bl_168 br_168 wl_208 vdd gnd cell_6t
Xbit_r209_c168 bl_168 br_168 wl_209 vdd gnd cell_6t
Xbit_r210_c168 bl_168 br_168 wl_210 vdd gnd cell_6t
Xbit_r211_c168 bl_168 br_168 wl_211 vdd gnd cell_6t
Xbit_r212_c168 bl_168 br_168 wl_212 vdd gnd cell_6t
Xbit_r213_c168 bl_168 br_168 wl_213 vdd gnd cell_6t
Xbit_r214_c168 bl_168 br_168 wl_214 vdd gnd cell_6t
Xbit_r215_c168 bl_168 br_168 wl_215 vdd gnd cell_6t
Xbit_r216_c168 bl_168 br_168 wl_216 vdd gnd cell_6t
Xbit_r217_c168 bl_168 br_168 wl_217 vdd gnd cell_6t
Xbit_r218_c168 bl_168 br_168 wl_218 vdd gnd cell_6t
Xbit_r219_c168 bl_168 br_168 wl_219 vdd gnd cell_6t
Xbit_r220_c168 bl_168 br_168 wl_220 vdd gnd cell_6t
Xbit_r221_c168 bl_168 br_168 wl_221 vdd gnd cell_6t
Xbit_r222_c168 bl_168 br_168 wl_222 vdd gnd cell_6t
Xbit_r223_c168 bl_168 br_168 wl_223 vdd gnd cell_6t
Xbit_r224_c168 bl_168 br_168 wl_224 vdd gnd cell_6t
Xbit_r225_c168 bl_168 br_168 wl_225 vdd gnd cell_6t
Xbit_r226_c168 bl_168 br_168 wl_226 vdd gnd cell_6t
Xbit_r227_c168 bl_168 br_168 wl_227 vdd gnd cell_6t
Xbit_r228_c168 bl_168 br_168 wl_228 vdd gnd cell_6t
Xbit_r229_c168 bl_168 br_168 wl_229 vdd gnd cell_6t
Xbit_r230_c168 bl_168 br_168 wl_230 vdd gnd cell_6t
Xbit_r231_c168 bl_168 br_168 wl_231 vdd gnd cell_6t
Xbit_r232_c168 bl_168 br_168 wl_232 vdd gnd cell_6t
Xbit_r233_c168 bl_168 br_168 wl_233 vdd gnd cell_6t
Xbit_r234_c168 bl_168 br_168 wl_234 vdd gnd cell_6t
Xbit_r235_c168 bl_168 br_168 wl_235 vdd gnd cell_6t
Xbit_r236_c168 bl_168 br_168 wl_236 vdd gnd cell_6t
Xbit_r237_c168 bl_168 br_168 wl_237 vdd gnd cell_6t
Xbit_r238_c168 bl_168 br_168 wl_238 vdd gnd cell_6t
Xbit_r239_c168 bl_168 br_168 wl_239 vdd gnd cell_6t
Xbit_r240_c168 bl_168 br_168 wl_240 vdd gnd cell_6t
Xbit_r241_c168 bl_168 br_168 wl_241 vdd gnd cell_6t
Xbit_r242_c168 bl_168 br_168 wl_242 vdd gnd cell_6t
Xbit_r243_c168 bl_168 br_168 wl_243 vdd gnd cell_6t
Xbit_r244_c168 bl_168 br_168 wl_244 vdd gnd cell_6t
Xbit_r245_c168 bl_168 br_168 wl_245 vdd gnd cell_6t
Xbit_r246_c168 bl_168 br_168 wl_246 vdd gnd cell_6t
Xbit_r247_c168 bl_168 br_168 wl_247 vdd gnd cell_6t
Xbit_r248_c168 bl_168 br_168 wl_248 vdd gnd cell_6t
Xbit_r249_c168 bl_168 br_168 wl_249 vdd gnd cell_6t
Xbit_r250_c168 bl_168 br_168 wl_250 vdd gnd cell_6t
Xbit_r251_c168 bl_168 br_168 wl_251 vdd gnd cell_6t
Xbit_r252_c168 bl_168 br_168 wl_252 vdd gnd cell_6t
Xbit_r253_c168 bl_168 br_168 wl_253 vdd gnd cell_6t
Xbit_r254_c168 bl_168 br_168 wl_254 vdd gnd cell_6t
Xbit_r255_c168 bl_168 br_168 wl_255 vdd gnd cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd cell_6t
Xbit_r1_c169 bl_169 br_169 wl_1 vdd gnd cell_6t
Xbit_r2_c169 bl_169 br_169 wl_2 vdd gnd cell_6t
Xbit_r3_c169 bl_169 br_169 wl_3 vdd gnd cell_6t
Xbit_r4_c169 bl_169 br_169 wl_4 vdd gnd cell_6t
Xbit_r5_c169 bl_169 br_169 wl_5 vdd gnd cell_6t
Xbit_r6_c169 bl_169 br_169 wl_6 vdd gnd cell_6t
Xbit_r7_c169 bl_169 br_169 wl_7 vdd gnd cell_6t
Xbit_r8_c169 bl_169 br_169 wl_8 vdd gnd cell_6t
Xbit_r9_c169 bl_169 br_169 wl_9 vdd gnd cell_6t
Xbit_r10_c169 bl_169 br_169 wl_10 vdd gnd cell_6t
Xbit_r11_c169 bl_169 br_169 wl_11 vdd gnd cell_6t
Xbit_r12_c169 bl_169 br_169 wl_12 vdd gnd cell_6t
Xbit_r13_c169 bl_169 br_169 wl_13 vdd gnd cell_6t
Xbit_r14_c169 bl_169 br_169 wl_14 vdd gnd cell_6t
Xbit_r15_c169 bl_169 br_169 wl_15 vdd gnd cell_6t
Xbit_r16_c169 bl_169 br_169 wl_16 vdd gnd cell_6t
Xbit_r17_c169 bl_169 br_169 wl_17 vdd gnd cell_6t
Xbit_r18_c169 bl_169 br_169 wl_18 vdd gnd cell_6t
Xbit_r19_c169 bl_169 br_169 wl_19 vdd gnd cell_6t
Xbit_r20_c169 bl_169 br_169 wl_20 vdd gnd cell_6t
Xbit_r21_c169 bl_169 br_169 wl_21 vdd gnd cell_6t
Xbit_r22_c169 bl_169 br_169 wl_22 vdd gnd cell_6t
Xbit_r23_c169 bl_169 br_169 wl_23 vdd gnd cell_6t
Xbit_r24_c169 bl_169 br_169 wl_24 vdd gnd cell_6t
Xbit_r25_c169 bl_169 br_169 wl_25 vdd gnd cell_6t
Xbit_r26_c169 bl_169 br_169 wl_26 vdd gnd cell_6t
Xbit_r27_c169 bl_169 br_169 wl_27 vdd gnd cell_6t
Xbit_r28_c169 bl_169 br_169 wl_28 vdd gnd cell_6t
Xbit_r29_c169 bl_169 br_169 wl_29 vdd gnd cell_6t
Xbit_r30_c169 bl_169 br_169 wl_30 vdd gnd cell_6t
Xbit_r31_c169 bl_169 br_169 wl_31 vdd gnd cell_6t
Xbit_r32_c169 bl_169 br_169 wl_32 vdd gnd cell_6t
Xbit_r33_c169 bl_169 br_169 wl_33 vdd gnd cell_6t
Xbit_r34_c169 bl_169 br_169 wl_34 vdd gnd cell_6t
Xbit_r35_c169 bl_169 br_169 wl_35 vdd gnd cell_6t
Xbit_r36_c169 bl_169 br_169 wl_36 vdd gnd cell_6t
Xbit_r37_c169 bl_169 br_169 wl_37 vdd gnd cell_6t
Xbit_r38_c169 bl_169 br_169 wl_38 vdd gnd cell_6t
Xbit_r39_c169 bl_169 br_169 wl_39 vdd gnd cell_6t
Xbit_r40_c169 bl_169 br_169 wl_40 vdd gnd cell_6t
Xbit_r41_c169 bl_169 br_169 wl_41 vdd gnd cell_6t
Xbit_r42_c169 bl_169 br_169 wl_42 vdd gnd cell_6t
Xbit_r43_c169 bl_169 br_169 wl_43 vdd gnd cell_6t
Xbit_r44_c169 bl_169 br_169 wl_44 vdd gnd cell_6t
Xbit_r45_c169 bl_169 br_169 wl_45 vdd gnd cell_6t
Xbit_r46_c169 bl_169 br_169 wl_46 vdd gnd cell_6t
Xbit_r47_c169 bl_169 br_169 wl_47 vdd gnd cell_6t
Xbit_r48_c169 bl_169 br_169 wl_48 vdd gnd cell_6t
Xbit_r49_c169 bl_169 br_169 wl_49 vdd gnd cell_6t
Xbit_r50_c169 bl_169 br_169 wl_50 vdd gnd cell_6t
Xbit_r51_c169 bl_169 br_169 wl_51 vdd gnd cell_6t
Xbit_r52_c169 bl_169 br_169 wl_52 vdd gnd cell_6t
Xbit_r53_c169 bl_169 br_169 wl_53 vdd gnd cell_6t
Xbit_r54_c169 bl_169 br_169 wl_54 vdd gnd cell_6t
Xbit_r55_c169 bl_169 br_169 wl_55 vdd gnd cell_6t
Xbit_r56_c169 bl_169 br_169 wl_56 vdd gnd cell_6t
Xbit_r57_c169 bl_169 br_169 wl_57 vdd gnd cell_6t
Xbit_r58_c169 bl_169 br_169 wl_58 vdd gnd cell_6t
Xbit_r59_c169 bl_169 br_169 wl_59 vdd gnd cell_6t
Xbit_r60_c169 bl_169 br_169 wl_60 vdd gnd cell_6t
Xbit_r61_c169 bl_169 br_169 wl_61 vdd gnd cell_6t
Xbit_r62_c169 bl_169 br_169 wl_62 vdd gnd cell_6t
Xbit_r63_c169 bl_169 br_169 wl_63 vdd gnd cell_6t
Xbit_r64_c169 bl_169 br_169 wl_64 vdd gnd cell_6t
Xbit_r65_c169 bl_169 br_169 wl_65 vdd gnd cell_6t
Xbit_r66_c169 bl_169 br_169 wl_66 vdd gnd cell_6t
Xbit_r67_c169 bl_169 br_169 wl_67 vdd gnd cell_6t
Xbit_r68_c169 bl_169 br_169 wl_68 vdd gnd cell_6t
Xbit_r69_c169 bl_169 br_169 wl_69 vdd gnd cell_6t
Xbit_r70_c169 bl_169 br_169 wl_70 vdd gnd cell_6t
Xbit_r71_c169 bl_169 br_169 wl_71 vdd gnd cell_6t
Xbit_r72_c169 bl_169 br_169 wl_72 vdd gnd cell_6t
Xbit_r73_c169 bl_169 br_169 wl_73 vdd gnd cell_6t
Xbit_r74_c169 bl_169 br_169 wl_74 vdd gnd cell_6t
Xbit_r75_c169 bl_169 br_169 wl_75 vdd gnd cell_6t
Xbit_r76_c169 bl_169 br_169 wl_76 vdd gnd cell_6t
Xbit_r77_c169 bl_169 br_169 wl_77 vdd gnd cell_6t
Xbit_r78_c169 bl_169 br_169 wl_78 vdd gnd cell_6t
Xbit_r79_c169 bl_169 br_169 wl_79 vdd gnd cell_6t
Xbit_r80_c169 bl_169 br_169 wl_80 vdd gnd cell_6t
Xbit_r81_c169 bl_169 br_169 wl_81 vdd gnd cell_6t
Xbit_r82_c169 bl_169 br_169 wl_82 vdd gnd cell_6t
Xbit_r83_c169 bl_169 br_169 wl_83 vdd gnd cell_6t
Xbit_r84_c169 bl_169 br_169 wl_84 vdd gnd cell_6t
Xbit_r85_c169 bl_169 br_169 wl_85 vdd gnd cell_6t
Xbit_r86_c169 bl_169 br_169 wl_86 vdd gnd cell_6t
Xbit_r87_c169 bl_169 br_169 wl_87 vdd gnd cell_6t
Xbit_r88_c169 bl_169 br_169 wl_88 vdd gnd cell_6t
Xbit_r89_c169 bl_169 br_169 wl_89 vdd gnd cell_6t
Xbit_r90_c169 bl_169 br_169 wl_90 vdd gnd cell_6t
Xbit_r91_c169 bl_169 br_169 wl_91 vdd gnd cell_6t
Xbit_r92_c169 bl_169 br_169 wl_92 vdd gnd cell_6t
Xbit_r93_c169 bl_169 br_169 wl_93 vdd gnd cell_6t
Xbit_r94_c169 bl_169 br_169 wl_94 vdd gnd cell_6t
Xbit_r95_c169 bl_169 br_169 wl_95 vdd gnd cell_6t
Xbit_r96_c169 bl_169 br_169 wl_96 vdd gnd cell_6t
Xbit_r97_c169 bl_169 br_169 wl_97 vdd gnd cell_6t
Xbit_r98_c169 bl_169 br_169 wl_98 vdd gnd cell_6t
Xbit_r99_c169 bl_169 br_169 wl_99 vdd gnd cell_6t
Xbit_r100_c169 bl_169 br_169 wl_100 vdd gnd cell_6t
Xbit_r101_c169 bl_169 br_169 wl_101 vdd gnd cell_6t
Xbit_r102_c169 bl_169 br_169 wl_102 vdd gnd cell_6t
Xbit_r103_c169 bl_169 br_169 wl_103 vdd gnd cell_6t
Xbit_r104_c169 bl_169 br_169 wl_104 vdd gnd cell_6t
Xbit_r105_c169 bl_169 br_169 wl_105 vdd gnd cell_6t
Xbit_r106_c169 bl_169 br_169 wl_106 vdd gnd cell_6t
Xbit_r107_c169 bl_169 br_169 wl_107 vdd gnd cell_6t
Xbit_r108_c169 bl_169 br_169 wl_108 vdd gnd cell_6t
Xbit_r109_c169 bl_169 br_169 wl_109 vdd gnd cell_6t
Xbit_r110_c169 bl_169 br_169 wl_110 vdd gnd cell_6t
Xbit_r111_c169 bl_169 br_169 wl_111 vdd gnd cell_6t
Xbit_r112_c169 bl_169 br_169 wl_112 vdd gnd cell_6t
Xbit_r113_c169 bl_169 br_169 wl_113 vdd gnd cell_6t
Xbit_r114_c169 bl_169 br_169 wl_114 vdd gnd cell_6t
Xbit_r115_c169 bl_169 br_169 wl_115 vdd gnd cell_6t
Xbit_r116_c169 bl_169 br_169 wl_116 vdd gnd cell_6t
Xbit_r117_c169 bl_169 br_169 wl_117 vdd gnd cell_6t
Xbit_r118_c169 bl_169 br_169 wl_118 vdd gnd cell_6t
Xbit_r119_c169 bl_169 br_169 wl_119 vdd gnd cell_6t
Xbit_r120_c169 bl_169 br_169 wl_120 vdd gnd cell_6t
Xbit_r121_c169 bl_169 br_169 wl_121 vdd gnd cell_6t
Xbit_r122_c169 bl_169 br_169 wl_122 vdd gnd cell_6t
Xbit_r123_c169 bl_169 br_169 wl_123 vdd gnd cell_6t
Xbit_r124_c169 bl_169 br_169 wl_124 vdd gnd cell_6t
Xbit_r125_c169 bl_169 br_169 wl_125 vdd gnd cell_6t
Xbit_r126_c169 bl_169 br_169 wl_126 vdd gnd cell_6t
Xbit_r127_c169 bl_169 br_169 wl_127 vdd gnd cell_6t
Xbit_r128_c169 bl_169 br_169 wl_128 vdd gnd cell_6t
Xbit_r129_c169 bl_169 br_169 wl_129 vdd gnd cell_6t
Xbit_r130_c169 bl_169 br_169 wl_130 vdd gnd cell_6t
Xbit_r131_c169 bl_169 br_169 wl_131 vdd gnd cell_6t
Xbit_r132_c169 bl_169 br_169 wl_132 vdd gnd cell_6t
Xbit_r133_c169 bl_169 br_169 wl_133 vdd gnd cell_6t
Xbit_r134_c169 bl_169 br_169 wl_134 vdd gnd cell_6t
Xbit_r135_c169 bl_169 br_169 wl_135 vdd gnd cell_6t
Xbit_r136_c169 bl_169 br_169 wl_136 vdd gnd cell_6t
Xbit_r137_c169 bl_169 br_169 wl_137 vdd gnd cell_6t
Xbit_r138_c169 bl_169 br_169 wl_138 vdd gnd cell_6t
Xbit_r139_c169 bl_169 br_169 wl_139 vdd gnd cell_6t
Xbit_r140_c169 bl_169 br_169 wl_140 vdd gnd cell_6t
Xbit_r141_c169 bl_169 br_169 wl_141 vdd gnd cell_6t
Xbit_r142_c169 bl_169 br_169 wl_142 vdd gnd cell_6t
Xbit_r143_c169 bl_169 br_169 wl_143 vdd gnd cell_6t
Xbit_r144_c169 bl_169 br_169 wl_144 vdd gnd cell_6t
Xbit_r145_c169 bl_169 br_169 wl_145 vdd gnd cell_6t
Xbit_r146_c169 bl_169 br_169 wl_146 vdd gnd cell_6t
Xbit_r147_c169 bl_169 br_169 wl_147 vdd gnd cell_6t
Xbit_r148_c169 bl_169 br_169 wl_148 vdd gnd cell_6t
Xbit_r149_c169 bl_169 br_169 wl_149 vdd gnd cell_6t
Xbit_r150_c169 bl_169 br_169 wl_150 vdd gnd cell_6t
Xbit_r151_c169 bl_169 br_169 wl_151 vdd gnd cell_6t
Xbit_r152_c169 bl_169 br_169 wl_152 vdd gnd cell_6t
Xbit_r153_c169 bl_169 br_169 wl_153 vdd gnd cell_6t
Xbit_r154_c169 bl_169 br_169 wl_154 vdd gnd cell_6t
Xbit_r155_c169 bl_169 br_169 wl_155 vdd gnd cell_6t
Xbit_r156_c169 bl_169 br_169 wl_156 vdd gnd cell_6t
Xbit_r157_c169 bl_169 br_169 wl_157 vdd gnd cell_6t
Xbit_r158_c169 bl_169 br_169 wl_158 vdd gnd cell_6t
Xbit_r159_c169 bl_169 br_169 wl_159 vdd gnd cell_6t
Xbit_r160_c169 bl_169 br_169 wl_160 vdd gnd cell_6t
Xbit_r161_c169 bl_169 br_169 wl_161 vdd gnd cell_6t
Xbit_r162_c169 bl_169 br_169 wl_162 vdd gnd cell_6t
Xbit_r163_c169 bl_169 br_169 wl_163 vdd gnd cell_6t
Xbit_r164_c169 bl_169 br_169 wl_164 vdd gnd cell_6t
Xbit_r165_c169 bl_169 br_169 wl_165 vdd gnd cell_6t
Xbit_r166_c169 bl_169 br_169 wl_166 vdd gnd cell_6t
Xbit_r167_c169 bl_169 br_169 wl_167 vdd gnd cell_6t
Xbit_r168_c169 bl_169 br_169 wl_168 vdd gnd cell_6t
Xbit_r169_c169 bl_169 br_169 wl_169 vdd gnd cell_6t
Xbit_r170_c169 bl_169 br_169 wl_170 vdd gnd cell_6t
Xbit_r171_c169 bl_169 br_169 wl_171 vdd gnd cell_6t
Xbit_r172_c169 bl_169 br_169 wl_172 vdd gnd cell_6t
Xbit_r173_c169 bl_169 br_169 wl_173 vdd gnd cell_6t
Xbit_r174_c169 bl_169 br_169 wl_174 vdd gnd cell_6t
Xbit_r175_c169 bl_169 br_169 wl_175 vdd gnd cell_6t
Xbit_r176_c169 bl_169 br_169 wl_176 vdd gnd cell_6t
Xbit_r177_c169 bl_169 br_169 wl_177 vdd gnd cell_6t
Xbit_r178_c169 bl_169 br_169 wl_178 vdd gnd cell_6t
Xbit_r179_c169 bl_169 br_169 wl_179 vdd gnd cell_6t
Xbit_r180_c169 bl_169 br_169 wl_180 vdd gnd cell_6t
Xbit_r181_c169 bl_169 br_169 wl_181 vdd gnd cell_6t
Xbit_r182_c169 bl_169 br_169 wl_182 vdd gnd cell_6t
Xbit_r183_c169 bl_169 br_169 wl_183 vdd gnd cell_6t
Xbit_r184_c169 bl_169 br_169 wl_184 vdd gnd cell_6t
Xbit_r185_c169 bl_169 br_169 wl_185 vdd gnd cell_6t
Xbit_r186_c169 bl_169 br_169 wl_186 vdd gnd cell_6t
Xbit_r187_c169 bl_169 br_169 wl_187 vdd gnd cell_6t
Xbit_r188_c169 bl_169 br_169 wl_188 vdd gnd cell_6t
Xbit_r189_c169 bl_169 br_169 wl_189 vdd gnd cell_6t
Xbit_r190_c169 bl_169 br_169 wl_190 vdd gnd cell_6t
Xbit_r191_c169 bl_169 br_169 wl_191 vdd gnd cell_6t
Xbit_r192_c169 bl_169 br_169 wl_192 vdd gnd cell_6t
Xbit_r193_c169 bl_169 br_169 wl_193 vdd gnd cell_6t
Xbit_r194_c169 bl_169 br_169 wl_194 vdd gnd cell_6t
Xbit_r195_c169 bl_169 br_169 wl_195 vdd gnd cell_6t
Xbit_r196_c169 bl_169 br_169 wl_196 vdd gnd cell_6t
Xbit_r197_c169 bl_169 br_169 wl_197 vdd gnd cell_6t
Xbit_r198_c169 bl_169 br_169 wl_198 vdd gnd cell_6t
Xbit_r199_c169 bl_169 br_169 wl_199 vdd gnd cell_6t
Xbit_r200_c169 bl_169 br_169 wl_200 vdd gnd cell_6t
Xbit_r201_c169 bl_169 br_169 wl_201 vdd gnd cell_6t
Xbit_r202_c169 bl_169 br_169 wl_202 vdd gnd cell_6t
Xbit_r203_c169 bl_169 br_169 wl_203 vdd gnd cell_6t
Xbit_r204_c169 bl_169 br_169 wl_204 vdd gnd cell_6t
Xbit_r205_c169 bl_169 br_169 wl_205 vdd gnd cell_6t
Xbit_r206_c169 bl_169 br_169 wl_206 vdd gnd cell_6t
Xbit_r207_c169 bl_169 br_169 wl_207 vdd gnd cell_6t
Xbit_r208_c169 bl_169 br_169 wl_208 vdd gnd cell_6t
Xbit_r209_c169 bl_169 br_169 wl_209 vdd gnd cell_6t
Xbit_r210_c169 bl_169 br_169 wl_210 vdd gnd cell_6t
Xbit_r211_c169 bl_169 br_169 wl_211 vdd gnd cell_6t
Xbit_r212_c169 bl_169 br_169 wl_212 vdd gnd cell_6t
Xbit_r213_c169 bl_169 br_169 wl_213 vdd gnd cell_6t
Xbit_r214_c169 bl_169 br_169 wl_214 vdd gnd cell_6t
Xbit_r215_c169 bl_169 br_169 wl_215 vdd gnd cell_6t
Xbit_r216_c169 bl_169 br_169 wl_216 vdd gnd cell_6t
Xbit_r217_c169 bl_169 br_169 wl_217 vdd gnd cell_6t
Xbit_r218_c169 bl_169 br_169 wl_218 vdd gnd cell_6t
Xbit_r219_c169 bl_169 br_169 wl_219 vdd gnd cell_6t
Xbit_r220_c169 bl_169 br_169 wl_220 vdd gnd cell_6t
Xbit_r221_c169 bl_169 br_169 wl_221 vdd gnd cell_6t
Xbit_r222_c169 bl_169 br_169 wl_222 vdd gnd cell_6t
Xbit_r223_c169 bl_169 br_169 wl_223 vdd gnd cell_6t
Xbit_r224_c169 bl_169 br_169 wl_224 vdd gnd cell_6t
Xbit_r225_c169 bl_169 br_169 wl_225 vdd gnd cell_6t
Xbit_r226_c169 bl_169 br_169 wl_226 vdd gnd cell_6t
Xbit_r227_c169 bl_169 br_169 wl_227 vdd gnd cell_6t
Xbit_r228_c169 bl_169 br_169 wl_228 vdd gnd cell_6t
Xbit_r229_c169 bl_169 br_169 wl_229 vdd gnd cell_6t
Xbit_r230_c169 bl_169 br_169 wl_230 vdd gnd cell_6t
Xbit_r231_c169 bl_169 br_169 wl_231 vdd gnd cell_6t
Xbit_r232_c169 bl_169 br_169 wl_232 vdd gnd cell_6t
Xbit_r233_c169 bl_169 br_169 wl_233 vdd gnd cell_6t
Xbit_r234_c169 bl_169 br_169 wl_234 vdd gnd cell_6t
Xbit_r235_c169 bl_169 br_169 wl_235 vdd gnd cell_6t
Xbit_r236_c169 bl_169 br_169 wl_236 vdd gnd cell_6t
Xbit_r237_c169 bl_169 br_169 wl_237 vdd gnd cell_6t
Xbit_r238_c169 bl_169 br_169 wl_238 vdd gnd cell_6t
Xbit_r239_c169 bl_169 br_169 wl_239 vdd gnd cell_6t
Xbit_r240_c169 bl_169 br_169 wl_240 vdd gnd cell_6t
Xbit_r241_c169 bl_169 br_169 wl_241 vdd gnd cell_6t
Xbit_r242_c169 bl_169 br_169 wl_242 vdd gnd cell_6t
Xbit_r243_c169 bl_169 br_169 wl_243 vdd gnd cell_6t
Xbit_r244_c169 bl_169 br_169 wl_244 vdd gnd cell_6t
Xbit_r245_c169 bl_169 br_169 wl_245 vdd gnd cell_6t
Xbit_r246_c169 bl_169 br_169 wl_246 vdd gnd cell_6t
Xbit_r247_c169 bl_169 br_169 wl_247 vdd gnd cell_6t
Xbit_r248_c169 bl_169 br_169 wl_248 vdd gnd cell_6t
Xbit_r249_c169 bl_169 br_169 wl_249 vdd gnd cell_6t
Xbit_r250_c169 bl_169 br_169 wl_250 vdd gnd cell_6t
Xbit_r251_c169 bl_169 br_169 wl_251 vdd gnd cell_6t
Xbit_r252_c169 bl_169 br_169 wl_252 vdd gnd cell_6t
Xbit_r253_c169 bl_169 br_169 wl_253 vdd gnd cell_6t
Xbit_r254_c169 bl_169 br_169 wl_254 vdd gnd cell_6t
Xbit_r255_c169 bl_169 br_169 wl_255 vdd gnd cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd cell_6t
Xbit_r1_c170 bl_170 br_170 wl_1 vdd gnd cell_6t
Xbit_r2_c170 bl_170 br_170 wl_2 vdd gnd cell_6t
Xbit_r3_c170 bl_170 br_170 wl_3 vdd gnd cell_6t
Xbit_r4_c170 bl_170 br_170 wl_4 vdd gnd cell_6t
Xbit_r5_c170 bl_170 br_170 wl_5 vdd gnd cell_6t
Xbit_r6_c170 bl_170 br_170 wl_6 vdd gnd cell_6t
Xbit_r7_c170 bl_170 br_170 wl_7 vdd gnd cell_6t
Xbit_r8_c170 bl_170 br_170 wl_8 vdd gnd cell_6t
Xbit_r9_c170 bl_170 br_170 wl_9 vdd gnd cell_6t
Xbit_r10_c170 bl_170 br_170 wl_10 vdd gnd cell_6t
Xbit_r11_c170 bl_170 br_170 wl_11 vdd gnd cell_6t
Xbit_r12_c170 bl_170 br_170 wl_12 vdd gnd cell_6t
Xbit_r13_c170 bl_170 br_170 wl_13 vdd gnd cell_6t
Xbit_r14_c170 bl_170 br_170 wl_14 vdd gnd cell_6t
Xbit_r15_c170 bl_170 br_170 wl_15 vdd gnd cell_6t
Xbit_r16_c170 bl_170 br_170 wl_16 vdd gnd cell_6t
Xbit_r17_c170 bl_170 br_170 wl_17 vdd gnd cell_6t
Xbit_r18_c170 bl_170 br_170 wl_18 vdd gnd cell_6t
Xbit_r19_c170 bl_170 br_170 wl_19 vdd gnd cell_6t
Xbit_r20_c170 bl_170 br_170 wl_20 vdd gnd cell_6t
Xbit_r21_c170 bl_170 br_170 wl_21 vdd gnd cell_6t
Xbit_r22_c170 bl_170 br_170 wl_22 vdd gnd cell_6t
Xbit_r23_c170 bl_170 br_170 wl_23 vdd gnd cell_6t
Xbit_r24_c170 bl_170 br_170 wl_24 vdd gnd cell_6t
Xbit_r25_c170 bl_170 br_170 wl_25 vdd gnd cell_6t
Xbit_r26_c170 bl_170 br_170 wl_26 vdd gnd cell_6t
Xbit_r27_c170 bl_170 br_170 wl_27 vdd gnd cell_6t
Xbit_r28_c170 bl_170 br_170 wl_28 vdd gnd cell_6t
Xbit_r29_c170 bl_170 br_170 wl_29 vdd gnd cell_6t
Xbit_r30_c170 bl_170 br_170 wl_30 vdd gnd cell_6t
Xbit_r31_c170 bl_170 br_170 wl_31 vdd gnd cell_6t
Xbit_r32_c170 bl_170 br_170 wl_32 vdd gnd cell_6t
Xbit_r33_c170 bl_170 br_170 wl_33 vdd gnd cell_6t
Xbit_r34_c170 bl_170 br_170 wl_34 vdd gnd cell_6t
Xbit_r35_c170 bl_170 br_170 wl_35 vdd gnd cell_6t
Xbit_r36_c170 bl_170 br_170 wl_36 vdd gnd cell_6t
Xbit_r37_c170 bl_170 br_170 wl_37 vdd gnd cell_6t
Xbit_r38_c170 bl_170 br_170 wl_38 vdd gnd cell_6t
Xbit_r39_c170 bl_170 br_170 wl_39 vdd gnd cell_6t
Xbit_r40_c170 bl_170 br_170 wl_40 vdd gnd cell_6t
Xbit_r41_c170 bl_170 br_170 wl_41 vdd gnd cell_6t
Xbit_r42_c170 bl_170 br_170 wl_42 vdd gnd cell_6t
Xbit_r43_c170 bl_170 br_170 wl_43 vdd gnd cell_6t
Xbit_r44_c170 bl_170 br_170 wl_44 vdd gnd cell_6t
Xbit_r45_c170 bl_170 br_170 wl_45 vdd gnd cell_6t
Xbit_r46_c170 bl_170 br_170 wl_46 vdd gnd cell_6t
Xbit_r47_c170 bl_170 br_170 wl_47 vdd gnd cell_6t
Xbit_r48_c170 bl_170 br_170 wl_48 vdd gnd cell_6t
Xbit_r49_c170 bl_170 br_170 wl_49 vdd gnd cell_6t
Xbit_r50_c170 bl_170 br_170 wl_50 vdd gnd cell_6t
Xbit_r51_c170 bl_170 br_170 wl_51 vdd gnd cell_6t
Xbit_r52_c170 bl_170 br_170 wl_52 vdd gnd cell_6t
Xbit_r53_c170 bl_170 br_170 wl_53 vdd gnd cell_6t
Xbit_r54_c170 bl_170 br_170 wl_54 vdd gnd cell_6t
Xbit_r55_c170 bl_170 br_170 wl_55 vdd gnd cell_6t
Xbit_r56_c170 bl_170 br_170 wl_56 vdd gnd cell_6t
Xbit_r57_c170 bl_170 br_170 wl_57 vdd gnd cell_6t
Xbit_r58_c170 bl_170 br_170 wl_58 vdd gnd cell_6t
Xbit_r59_c170 bl_170 br_170 wl_59 vdd gnd cell_6t
Xbit_r60_c170 bl_170 br_170 wl_60 vdd gnd cell_6t
Xbit_r61_c170 bl_170 br_170 wl_61 vdd gnd cell_6t
Xbit_r62_c170 bl_170 br_170 wl_62 vdd gnd cell_6t
Xbit_r63_c170 bl_170 br_170 wl_63 vdd gnd cell_6t
Xbit_r64_c170 bl_170 br_170 wl_64 vdd gnd cell_6t
Xbit_r65_c170 bl_170 br_170 wl_65 vdd gnd cell_6t
Xbit_r66_c170 bl_170 br_170 wl_66 vdd gnd cell_6t
Xbit_r67_c170 bl_170 br_170 wl_67 vdd gnd cell_6t
Xbit_r68_c170 bl_170 br_170 wl_68 vdd gnd cell_6t
Xbit_r69_c170 bl_170 br_170 wl_69 vdd gnd cell_6t
Xbit_r70_c170 bl_170 br_170 wl_70 vdd gnd cell_6t
Xbit_r71_c170 bl_170 br_170 wl_71 vdd gnd cell_6t
Xbit_r72_c170 bl_170 br_170 wl_72 vdd gnd cell_6t
Xbit_r73_c170 bl_170 br_170 wl_73 vdd gnd cell_6t
Xbit_r74_c170 bl_170 br_170 wl_74 vdd gnd cell_6t
Xbit_r75_c170 bl_170 br_170 wl_75 vdd gnd cell_6t
Xbit_r76_c170 bl_170 br_170 wl_76 vdd gnd cell_6t
Xbit_r77_c170 bl_170 br_170 wl_77 vdd gnd cell_6t
Xbit_r78_c170 bl_170 br_170 wl_78 vdd gnd cell_6t
Xbit_r79_c170 bl_170 br_170 wl_79 vdd gnd cell_6t
Xbit_r80_c170 bl_170 br_170 wl_80 vdd gnd cell_6t
Xbit_r81_c170 bl_170 br_170 wl_81 vdd gnd cell_6t
Xbit_r82_c170 bl_170 br_170 wl_82 vdd gnd cell_6t
Xbit_r83_c170 bl_170 br_170 wl_83 vdd gnd cell_6t
Xbit_r84_c170 bl_170 br_170 wl_84 vdd gnd cell_6t
Xbit_r85_c170 bl_170 br_170 wl_85 vdd gnd cell_6t
Xbit_r86_c170 bl_170 br_170 wl_86 vdd gnd cell_6t
Xbit_r87_c170 bl_170 br_170 wl_87 vdd gnd cell_6t
Xbit_r88_c170 bl_170 br_170 wl_88 vdd gnd cell_6t
Xbit_r89_c170 bl_170 br_170 wl_89 vdd gnd cell_6t
Xbit_r90_c170 bl_170 br_170 wl_90 vdd gnd cell_6t
Xbit_r91_c170 bl_170 br_170 wl_91 vdd gnd cell_6t
Xbit_r92_c170 bl_170 br_170 wl_92 vdd gnd cell_6t
Xbit_r93_c170 bl_170 br_170 wl_93 vdd gnd cell_6t
Xbit_r94_c170 bl_170 br_170 wl_94 vdd gnd cell_6t
Xbit_r95_c170 bl_170 br_170 wl_95 vdd gnd cell_6t
Xbit_r96_c170 bl_170 br_170 wl_96 vdd gnd cell_6t
Xbit_r97_c170 bl_170 br_170 wl_97 vdd gnd cell_6t
Xbit_r98_c170 bl_170 br_170 wl_98 vdd gnd cell_6t
Xbit_r99_c170 bl_170 br_170 wl_99 vdd gnd cell_6t
Xbit_r100_c170 bl_170 br_170 wl_100 vdd gnd cell_6t
Xbit_r101_c170 bl_170 br_170 wl_101 vdd gnd cell_6t
Xbit_r102_c170 bl_170 br_170 wl_102 vdd gnd cell_6t
Xbit_r103_c170 bl_170 br_170 wl_103 vdd gnd cell_6t
Xbit_r104_c170 bl_170 br_170 wl_104 vdd gnd cell_6t
Xbit_r105_c170 bl_170 br_170 wl_105 vdd gnd cell_6t
Xbit_r106_c170 bl_170 br_170 wl_106 vdd gnd cell_6t
Xbit_r107_c170 bl_170 br_170 wl_107 vdd gnd cell_6t
Xbit_r108_c170 bl_170 br_170 wl_108 vdd gnd cell_6t
Xbit_r109_c170 bl_170 br_170 wl_109 vdd gnd cell_6t
Xbit_r110_c170 bl_170 br_170 wl_110 vdd gnd cell_6t
Xbit_r111_c170 bl_170 br_170 wl_111 vdd gnd cell_6t
Xbit_r112_c170 bl_170 br_170 wl_112 vdd gnd cell_6t
Xbit_r113_c170 bl_170 br_170 wl_113 vdd gnd cell_6t
Xbit_r114_c170 bl_170 br_170 wl_114 vdd gnd cell_6t
Xbit_r115_c170 bl_170 br_170 wl_115 vdd gnd cell_6t
Xbit_r116_c170 bl_170 br_170 wl_116 vdd gnd cell_6t
Xbit_r117_c170 bl_170 br_170 wl_117 vdd gnd cell_6t
Xbit_r118_c170 bl_170 br_170 wl_118 vdd gnd cell_6t
Xbit_r119_c170 bl_170 br_170 wl_119 vdd gnd cell_6t
Xbit_r120_c170 bl_170 br_170 wl_120 vdd gnd cell_6t
Xbit_r121_c170 bl_170 br_170 wl_121 vdd gnd cell_6t
Xbit_r122_c170 bl_170 br_170 wl_122 vdd gnd cell_6t
Xbit_r123_c170 bl_170 br_170 wl_123 vdd gnd cell_6t
Xbit_r124_c170 bl_170 br_170 wl_124 vdd gnd cell_6t
Xbit_r125_c170 bl_170 br_170 wl_125 vdd gnd cell_6t
Xbit_r126_c170 bl_170 br_170 wl_126 vdd gnd cell_6t
Xbit_r127_c170 bl_170 br_170 wl_127 vdd gnd cell_6t
Xbit_r128_c170 bl_170 br_170 wl_128 vdd gnd cell_6t
Xbit_r129_c170 bl_170 br_170 wl_129 vdd gnd cell_6t
Xbit_r130_c170 bl_170 br_170 wl_130 vdd gnd cell_6t
Xbit_r131_c170 bl_170 br_170 wl_131 vdd gnd cell_6t
Xbit_r132_c170 bl_170 br_170 wl_132 vdd gnd cell_6t
Xbit_r133_c170 bl_170 br_170 wl_133 vdd gnd cell_6t
Xbit_r134_c170 bl_170 br_170 wl_134 vdd gnd cell_6t
Xbit_r135_c170 bl_170 br_170 wl_135 vdd gnd cell_6t
Xbit_r136_c170 bl_170 br_170 wl_136 vdd gnd cell_6t
Xbit_r137_c170 bl_170 br_170 wl_137 vdd gnd cell_6t
Xbit_r138_c170 bl_170 br_170 wl_138 vdd gnd cell_6t
Xbit_r139_c170 bl_170 br_170 wl_139 vdd gnd cell_6t
Xbit_r140_c170 bl_170 br_170 wl_140 vdd gnd cell_6t
Xbit_r141_c170 bl_170 br_170 wl_141 vdd gnd cell_6t
Xbit_r142_c170 bl_170 br_170 wl_142 vdd gnd cell_6t
Xbit_r143_c170 bl_170 br_170 wl_143 vdd gnd cell_6t
Xbit_r144_c170 bl_170 br_170 wl_144 vdd gnd cell_6t
Xbit_r145_c170 bl_170 br_170 wl_145 vdd gnd cell_6t
Xbit_r146_c170 bl_170 br_170 wl_146 vdd gnd cell_6t
Xbit_r147_c170 bl_170 br_170 wl_147 vdd gnd cell_6t
Xbit_r148_c170 bl_170 br_170 wl_148 vdd gnd cell_6t
Xbit_r149_c170 bl_170 br_170 wl_149 vdd gnd cell_6t
Xbit_r150_c170 bl_170 br_170 wl_150 vdd gnd cell_6t
Xbit_r151_c170 bl_170 br_170 wl_151 vdd gnd cell_6t
Xbit_r152_c170 bl_170 br_170 wl_152 vdd gnd cell_6t
Xbit_r153_c170 bl_170 br_170 wl_153 vdd gnd cell_6t
Xbit_r154_c170 bl_170 br_170 wl_154 vdd gnd cell_6t
Xbit_r155_c170 bl_170 br_170 wl_155 vdd gnd cell_6t
Xbit_r156_c170 bl_170 br_170 wl_156 vdd gnd cell_6t
Xbit_r157_c170 bl_170 br_170 wl_157 vdd gnd cell_6t
Xbit_r158_c170 bl_170 br_170 wl_158 vdd gnd cell_6t
Xbit_r159_c170 bl_170 br_170 wl_159 vdd gnd cell_6t
Xbit_r160_c170 bl_170 br_170 wl_160 vdd gnd cell_6t
Xbit_r161_c170 bl_170 br_170 wl_161 vdd gnd cell_6t
Xbit_r162_c170 bl_170 br_170 wl_162 vdd gnd cell_6t
Xbit_r163_c170 bl_170 br_170 wl_163 vdd gnd cell_6t
Xbit_r164_c170 bl_170 br_170 wl_164 vdd gnd cell_6t
Xbit_r165_c170 bl_170 br_170 wl_165 vdd gnd cell_6t
Xbit_r166_c170 bl_170 br_170 wl_166 vdd gnd cell_6t
Xbit_r167_c170 bl_170 br_170 wl_167 vdd gnd cell_6t
Xbit_r168_c170 bl_170 br_170 wl_168 vdd gnd cell_6t
Xbit_r169_c170 bl_170 br_170 wl_169 vdd gnd cell_6t
Xbit_r170_c170 bl_170 br_170 wl_170 vdd gnd cell_6t
Xbit_r171_c170 bl_170 br_170 wl_171 vdd gnd cell_6t
Xbit_r172_c170 bl_170 br_170 wl_172 vdd gnd cell_6t
Xbit_r173_c170 bl_170 br_170 wl_173 vdd gnd cell_6t
Xbit_r174_c170 bl_170 br_170 wl_174 vdd gnd cell_6t
Xbit_r175_c170 bl_170 br_170 wl_175 vdd gnd cell_6t
Xbit_r176_c170 bl_170 br_170 wl_176 vdd gnd cell_6t
Xbit_r177_c170 bl_170 br_170 wl_177 vdd gnd cell_6t
Xbit_r178_c170 bl_170 br_170 wl_178 vdd gnd cell_6t
Xbit_r179_c170 bl_170 br_170 wl_179 vdd gnd cell_6t
Xbit_r180_c170 bl_170 br_170 wl_180 vdd gnd cell_6t
Xbit_r181_c170 bl_170 br_170 wl_181 vdd gnd cell_6t
Xbit_r182_c170 bl_170 br_170 wl_182 vdd gnd cell_6t
Xbit_r183_c170 bl_170 br_170 wl_183 vdd gnd cell_6t
Xbit_r184_c170 bl_170 br_170 wl_184 vdd gnd cell_6t
Xbit_r185_c170 bl_170 br_170 wl_185 vdd gnd cell_6t
Xbit_r186_c170 bl_170 br_170 wl_186 vdd gnd cell_6t
Xbit_r187_c170 bl_170 br_170 wl_187 vdd gnd cell_6t
Xbit_r188_c170 bl_170 br_170 wl_188 vdd gnd cell_6t
Xbit_r189_c170 bl_170 br_170 wl_189 vdd gnd cell_6t
Xbit_r190_c170 bl_170 br_170 wl_190 vdd gnd cell_6t
Xbit_r191_c170 bl_170 br_170 wl_191 vdd gnd cell_6t
Xbit_r192_c170 bl_170 br_170 wl_192 vdd gnd cell_6t
Xbit_r193_c170 bl_170 br_170 wl_193 vdd gnd cell_6t
Xbit_r194_c170 bl_170 br_170 wl_194 vdd gnd cell_6t
Xbit_r195_c170 bl_170 br_170 wl_195 vdd gnd cell_6t
Xbit_r196_c170 bl_170 br_170 wl_196 vdd gnd cell_6t
Xbit_r197_c170 bl_170 br_170 wl_197 vdd gnd cell_6t
Xbit_r198_c170 bl_170 br_170 wl_198 vdd gnd cell_6t
Xbit_r199_c170 bl_170 br_170 wl_199 vdd gnd cell_6t
Xbit_r200_c170 bl_170 br_170 wl_200 vdd gnd cell_6t
Xbit_r201_c170 bl_170 br_170 wl_201 vdd gnd cell_6t
Xbit_r202_c170 bl_170 br_170 wl_202 vdd gnd cell_6t
Xbit_r203_c170 bl_170 br_170 wl_203 vdd gnd cell_6t
Xbit_r204_c170 bl_170 br_170 wl_204 vdd gnd cell_6t
Xbit_r205_c170 bl_170 br_170 wl_205 vdd gnd cell_6t
Xbit_r206_c170 bl_170 br_170 wl_206 vdd gnd cell_6t
Xbit_r207_c170 bl_170 br_170 wl_207 vdd gnd cell_6t
Xbit_r208_c170 bl_170 br_170 wl_208 vdd gnd cell_6t
Xbit_r209_c170 bl_170 br_170 wl_209 vdd gnd cell_6t
Xbit_r210_c170 bl_170 br_170 wl_210 vdd gnd cell_6t
Xbit_r211_c170 bl_170 br_170 wl_211 vdd gnd cell_6t
Xbit_r212_c170 bl_170 br_170 wl_212 vdd gnd cell_6t
Xbit_r213_c170 bl_170 br_170 wl_213 vdd gnd cell_6t
Xbit_r214_c170 bl_170 br_170 wl_214 vdd gnd cell_6t
Xbit_r215_c170 bl_170 br_170 wl_215 vdd gnd cell_6t
Xbit_r216_c170 bl_170 br_170 wl_216 vdd gnd cell_6t
Xbit_r217_c170 bl_170 br_170 wl_217 vdd gnd cell_6t
Xbit_r218_c170 bl_170 br_170 wl_218 vdd gnd cell_6t
Xbit_r219_c170 bl_170 br_170 wl_219 vdd gnd cell_6t
Xbit_r220_c170 bl_170 br_170 wl_220 vdd gnd cell_6t
Xbit_r221_c170 bl_170 br_170 wl_221 vdd gnd cell_6t
Xbit_r222_c170 bl_170 br_170 wl_222 vdd gnd cell_6t
Xbit_r223_c170 bl_170 br_170 wl_223 vdd gnd cell_6t
Xbit_r224_c170 bl_170 br_170 wl_224 vdd gnd cell_6t
Xbit_r225_c170 bl_170 br_170 wl_225 vdd gnd cell_6t
Xbit_r226_c170 bl_170 br_170 wl_226 vdd gnd cell_6t
Xbit_r227_c170 bl_170 br_170 wl_227 vdd gnd cell_6t
Xbit_r228_c170 bl_170 br_170 wl_228 vdd gnd cell_6t
Xbit_r229_c170 bl_170 br_170 wl_229 vdd gnd cell_6t
Xbit_r230_c170 bl_170 br_170 wl_230 vdd gnd cell_6t
Xbit_r231_c170 bl_170 br_170 wl_231 vdd gnd cell_6t
Xbit_r232_c170 bl_170 br_170 wl_232 vdd gnd cell_6t
Xbit_r233_c170 bl_170 br_170 wl_233 vdd gnd cell_6t
Xbit_r234_c170 bl_170 br_170 wl_234 vdd gnd cell_6t
Xbit_r235_c170 bl_170 br_170 wl_235 vdd gnd cell_6t
Xbit_r236_c170 bl_170 br_170 wl_236 vdd gnd cell_6t
Xbit_r237_c170 bl_170 br_170 wl_237 vdd gnd cell_6t
Xbit_r238_c170 bl_170 br_170 wl_238 vdd gnd cell_6t
Xbit_r239_c170 bl_170 br_170 wl_239 vdd gnd cell_6t
Xbit_r240_c170 bl_170 br_170 wl_240 vdd gnd cell_6t
Xbit_r241_c170 bl_170 br_170 wl_241 vdd gnd cell_6t
Xbit_r242_c170 bl_170 br_170 wl_242 vdd gnd cell_6t
Xbit_r243_c170 bl_170 br_170 wl_243 vdd gnd cell_6t
Xbit_r244_c170 bl_170 br_170 wl_244 vdd gnd cell_6t
Xbit_r245_c170 bl_170 br_170 wl_245 vdd gnd cell_6t
Xbit_r246_c170 bl_170 br_170 wl_246 vdd gnd cell_6t
Xbit_r247_c170 bl_170 br_170 wl_247 vdd gnd cell_6t
Xbit_r248_c170 bl_170 br_170 wl_248 vdd gnd cell_6t
Xbit_r249_c170 bl_170 br_170 wl_249 vdd gnd cell_6t
Xbit_r250_c170 bl_170 br_170 wl_250 vdd gnd cell_6t
Xbit_r251_c170 bl_170 br_170 wl_251 vdd gnd cell_6t
Xbit_r252_c170 bl_170 br_170 wl_252 vdd gnd cell_6t
Xbit_r253_c170 bl_170 br_170 wl_253 vdd gnd cell_6t
Xbit_r254_c170 bl_170 br_170 wl_254 vdd gnd cell_6t
Xbit_r255_c170 bl_170 br_170 wl_255 vdd gnd cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd cell_6t
Xbit_r1_c171 bl_171 br_171 wl_1 vdd gnd cell_6t
Xbit_r2_c171 bl_171 br_171 wl_2 vdd gnd cell_6t
Xbit_r3_c171 bl_171 br_171 wl_3 vdd gnd cell_6t
Xbit_r4_c171 bl_171 br_171 wl_4 vdd gnd cell_6t
Xbit_r5_c171 bl_171 br_171 wl_5 vdd gnd cell_6t
Xbit_r6_c171 bl_171 br_171 wl_6 vdd gnd cell_6t
Xbit_r7_c171 bl_171 br_171 wl_7 vdd gnd cell_6t
Xbit_r8_c171 bl_171 br_171 wl_8 vdd gnd cell_6t
Xbit_r9_c171 bl_171 br_171 wl_9 vdd gnd cell_6t
Xbit_r10_c171 bl_171 br_171 wl_10 vdd gnd cell_6t
Xbit_r11_c171 bl_171 br_171 wl_11 vdd gnd cell_6t
Xbit_r12_c171 bl_171 br_171 wl_12 vdd gnd cell_6t
Xbit_r13_c171 bl_171 br_171 wl_13 vdd gnd cell_6t
Xbit_r14_c171 bl_171 br_171 wl_14 vdd gnd cell_6t
Xbit_r15_c171 bl_171 br_171 wl_15 vdd gnd cell_6t
Xbit_r16_c171 bl_171 br_171 wl_16 vdd gnd cell_6t
Xbit_r17_c171 bl_171 br_171 wl_17 vdd gnd cell_6t
Xbit_r18_c171 bl_171 br_171 wl_18 vdd gnd cell_6t
Xbit_r19_c171 bl_171 br_171 wl_19 vdd gnd cell_6t
Xbit_r20_c171 bl_171 br_171 wl_20 vdd gnd cell_6t
Xbit_r21_c171 bl_171 br_171 wl_21 vdd gnd cell_6t
Xbit_r22_c171 bl_171 br_171 wl_22 vdd gnd cell_6t
Xbit_r23_c171 bl_171 br_171 wl_23 vdd gnd cell_6t
Xbit_r24_c171 bl_171 br_171 wl_24 vdd gnd cell_6t
Xbit_r25_c171 bl_171 br_171 wl_25 vdd gnd cell_6t
Xbit_r26_c171 bl_171 br_171 wl_26 vdd gnd cell_6t
Xbit_r27_c171 bl_171 br_171 wl_27 vdd gnd cell_6t
Xbit_r28_c171 bl_171 br_171 wl_28 vdd gnd cell_6t
Xbit_r29_c171 bl_171 br_171 wl_29 vdd gnd cell_6t
Xbit_r30_c171 bl_171 br_171 wl_30 vdd gnd cell_6t
Xbit_r31_c171 bl_171 br_171 wl_31 vdd gnd cell_6t
Xbit_r32_c171 bl_171 br_171 wl_32 vdd gnd cell_6t
Xbit_r33_c171 bl_171 br_171 wl_33 vdd gnd cell_6t
Xbit_r34_c171 bl_171 br_171 wl_34 vdd gnd cell_6t
Xbit_r35_c171 bl_171 br_171 wl_35 vdd gnd cell_6t
Xbit_r36_c171 bl_171 br_171 wl_36 vdd gnd cell_6t
Xbit_r37_c171 bl_171 br_171 wl_37 vdd gnd cell_6t
Xbit_r38_c171 bl_171 br_171 wl_38 vdd gnd cell_6t
Xbit_r39_c171 bl_171 br_171 wl_39 vdd gnd cell_6t
Xbit_r40_c171 bl_171 br_171 wl_40 vdd gnd cell_6t
Xbit_r41_c171 bl_171 br_171 wl_41 vdd gnd cell_6t
Xbit_r42_c171 bl_171 br_171 wl_42 vdd gnd cell_6t
Xbit_r43_c171 bl_171 br_171 wl_43 vdd gnd cell_6t
Xbit_r44_c171 bl_171 br_171 wl_44 vdd gnd cell_6t
Xbit_r45_c171 bl_171 br_171 wl_45 vdd gnd cell_6t
Xbit_r46_c171 bl_171 br_171 wl_46 vdd gnd cell_6t
Xbit_r47_c171 bl_171 br_171 wl_47 vdd gnd cell_6t
Xbit_r48_c171 bl_171 br_171 wl_48 vdd gnd cell_6t
Xbit_r49_c171 bl_171 br_171 wl_49 vdd gnd cell_6t
Xbit_r50_c171 bl_171 br_171 wl_50 vdd gnd cell_6t
Xbit_r51_c171 bl_171 br_171 wl_51 vdd gnd cell_6t
Xbit_r52_c171 bl_171 br_171 wl_52 vdd gnd cell_6t
Xbit_r53_c171 bl_171 br_171 wl_53 vdd gnd cell_6t
Xbit_r54_c171 bl_171 br_171 wl_54 vdd gnd cell_6t
Xbit_r55_c171 bl_171 br_171 wl_55 vdd gnd cell_6t
Xbit_r56_c171 bl_171 br_171 wl_56 vdd gnd cell_6t
Xbit_r57_c171 bl_171 br_171 wl_57 vdd gnd cell_6t
Xbit_r58_c171 bl_171 br_171 wl_58 vdd gnd cell_6t
Xbit_r59_c171 bl_171 br_171 wl_59 vdd gnd cell_6t
Xbit_r60_c171 bl_171 br_171 wl_60 vdd gnd cell_6t
Xbit_r61_c171 bl_171 br_171 wl_61 vdd gnd cell_6t
Xbit_r62_c171 bl_171 br_171 wl_62 vdd gnd cell_6t
Xbit_r63_c171 bl_171 br_171 wl_63 vdd gnd cell_6t
Xbit_r64_c171 bl_171 br_171 wl_64 vdd gnd cell_6t
Xbit_r65_c171 bl_171 br_171 wl_65 vdd gnd cell_6t
Xbit_r66_c171 bl_171 br_171 wl_66 vdd gnd cell_6t
Xbit_r67_c171 bl_171 br_171 wl_67 vdd gnd cell_6t
Xbit_r68_c171 bl_171 br_171 wl_68 vdd gnd cell_6t
Xbit_r69_c171 bl_171 br_171 wl_69 vdd gnd cell_6t
Xbit_r70_c171 bl_171 br_171 wl_70 vdd gnd cell_6t
Xbit_r71_c171 bl_171 br_171 wl_71 vdd gnd cell_6t
Xbit_r72_c171 bl_171 br_171 wl_72 vdd gnd cell_6t
Xbit_r73_c171 bl_171 br_171 wl_73 vdd gnd cell_6t
Xbit_r74_c171 bl_171 br_171 wl_74 vdd gnd cell_6t
Xbit_r75_c171 bl_171 br_171 wl_75 vdd gnd cell_6t
Xbit_r76_c171 bl_171 br_171 wl_76 vdd gnd cell_6t
Xbit_r77_c171 bl_171 br_171 wl_77 vdd gnd cell_6t
Xbit_r78_c171 bl_171 br_171 wl_78 vdd gnd cell_6t
Xbit_r79_c171 bl_171 br_171 wl_79 vdd gnd cell_6t
Xbit_r80_c171 bl_171 br_171 wl_80 vdd gnd cell_6t
Xbit_r81_c171 bl_171 br_171 wl_81 vdd gnd cell_6t
Xbit_r82_c171 bl_171 br_171 wl_82 vdd gnd cell_6t
Xbit_r83_c171 bl_171 br_171 wl_83 vdd gnd cell_6t
Xbit_r84_c171 bl_171 br_171 wl_84 vdd gnd cell_6t
Xbit_r85_c171 bl_171 br_171 wl_85 vdd gnd cell_6t
Xbit_r86_c171 bl_171 br_171 wl_86 vdd gnd cell_6t
Xbit_r87_c171 bl_171 br_171 wl_87 vdd gnd cell_6t
Xbit_r88_c171 bl_171 br_171 wl_88 vdd gnd cell_6t
Xbit_r89_c171 bl_171 br_171 wl_89 vdd gnd cell_6t
Xbit_r90_c171 bl_171 br_171 wl_90 vdd gnd cell_6t
Xbit_r91_c171 bl_171 br_171 wl_91 vdd gnd cell_6t
Xbit_r92_c171 bl_171 br_171 wl_92 vdd gnd cell_6t
Xbit_r93_c171 bl_171 br_171 wl_93 vdd gnd cell_6t
Xbit_r94_c171 bl_171 br_171 wl_94 vdd gnd cell_6t
Xbit_r95_c171 bl_171 br_171 wl_95 vdd gnd cell_6t
Xbit_r96_c171 bl_171 br_171 wl_96 vdd gnd cell_6t
Xbit_r97_c171 bl_171 br_171 wl_97 vdd gnd cell_6t
Xbit_r98_c171 bl_171 br_171 wl_98 vdd gnd cell_6t
Xbit_r99_c171 bl_171 br_171 wl_99 vdd gnd cell_6t
Xbit_r100_c171 bl_171 br_171 wl_100 vdd gnd cell_6t
Xbit_r101_c171 bl_171 br_171 wl_101 vdd gnd cell_6t
Xbit_r102_c171 bl_171 br_171 wl_102 vdd gnd cell_6t
Xbit_r103_c171 bl_171 br_171 wl_103 vdd gnd cell_6t
Xbit_r104_c171 bl_171 br_171 wl_104 vdd gnd cell_6t
Xbit_r105_c171 bl_171 br_171 wl_105 vdd gnd cell_6t
Xbit_r106_c171 bl_171 br_171 wl_106 vdd gnd cell_6t
Xbit_r107_c171 bl_171 br_171 wl_107 vdd gnd cell_6t
Xbit_r108_c171 bl_171 br_171 wl_108 vdd gnd cell_6t
Xbit_r109_c171 bl_171 br_171 wl_109 vdd gnd cell_6t
Xbit_r110_c171 bl_171 br_171 wl_110 vdd gnd cell_6t
Xbit_r111_c171 bl_171 br_171 wl_111 vdd gnd cell_6t
Xbit_r112_c171 bl_171 br_171 wl_112 vdd gnd cell_6t
Xbit_r113_c171 bl_171 br_171 wl_113 vdd gnd cell_6t
Xbit_r114_c171 bl_171 br_171 wl_114 vdd gnd cell_6t
Xbit_r115_c171 bl_171 br_171 wl_115 vdd gnd cell_6t
Xbit_r116_c171 bl_171 br_171 wl_116 vdd gnd cell_6t
Xbit_r117_c171 bl_171 br_171 wl_117 vdd gnd cell_6t
Xbit_r118_c171 bl_171 br_171 wl_118 vdd gnd cell_6t
Xbit_r119_c171 bl_171 br_171 wl_119 vdd gnd cell_6t
Xbit_r120_c171 bl_171 br_171 wl_120 vdd gnd cell_6t
Xbit_r121_c171 bl_171 br_171 wl_121 vdd gnd cell_6t
Xbit_r122_c171 bl_171 br_171 wl_122 vdd gnd cell_6t
Xbit_r123_c171 bl_171 br_171 wl_123 vdd gnd cell_6t
Xbit_r124_c171 bl_171 br_171 wl_124 vdd gnd cell_6t
Xbit_r125_c171 bl_171 br_171 wl_125 vdd gnd cell_6t
Xbit_r126_c171 bl_171 br_171 wl_126 vdd gnd cell_6t
Xbit_r127_c171 bl_171 br_171 wl_127 vdd gnd cell_6t
Xbit_r128_c171 bl_171 br_171 wl_128 vdd gnd cell_6t
Xbit_r129_c171 bl_171 br_171 wl_129 vdd gnd cell_6t
Xbit_r130_c171 bl_171 br_171 wl_130 vdd gnd cell_6t
Xbit_r131_c171 bl_171 br_171 wl_131 vdd gnd cell_6t
Xbit_r132_c171 bl_171 br_171 wl_132 vdd gnd cell_6t
Xbit_r133_c171 bl_171 br_171 wl_133 vdd gnd cell_6t
Xbit_r134_c171 bl_171 br_171 wl_134 vdd gnd cell_6t
Xbit_r135_c171 bl_171 br_171 wl_135 vdd gnd cell_6t
Xbit_r136_c171 bl_171 br_171 wl_136 vdd gnd cell_6t
Xbit_r137_c171 bl_171 br_171 wl_137 vdd gnd cell_6t
Xbit_r138_c171 bl_171 br_171 wl_138 vdd gnd cell_6t
Xbit_r139_c171 bl_171 br_171 wl_139 vdd gnd cell_6t
Xbit_r140_c171 bl_171 br_171 wl_140 vdd gnd cell_6t
Xbit_r141_c171 bl_171 br_171 wl_141 vdd gnd cell_6t
Xbit_r142_c171 bl_171 br_171 wl_142 vdd gnd cell_6t
Xbit_r143_c171 bl_171 br_171 wl_143 vdd gnd cell_6t
Xbit_r144_c171 bl_171 br_171 wl_144 vdd gnd cell_6t
Xbit_r145_c171 bl_171 br_171 wl_145 vdd gnd cell_6t
Xbit_r146_c171 bl_171 br_171 wl_146 vdd gnd cell_6t
Xbit_r147_c171 bl_171 br_171 wl_147 vdd gnd cell_6t
Xbit_r148_c171 bl_171 br_171 wl_148 vdd gnd cell_6t
Xbit_r149_c171 bl_171 br_171 wl_149 vdd gnd cell_6t
Xbit_r150_c171 bl_171 br_171 wl_150 vdd gnd cell_6t
Xbit_r151_c171 bl_171 br_171 wl_151 vdd gnd cell_6t
Xbit_r152_c171 bl_171 br_171 wl_152 vdd gnd cell_6t
Xbit_r153_c171 bl_171 br_171 wl_153 vdd gnd cell_6t
Xbit_r154_c171 bl_171 br_171 wl_154 vdd gnd cell_6t
Xbit_r155_c171 bl_171 br_171 wl_155 vdd gnd cell_6t
Xbit_r156_c171 bl_171 br_171 wl_156 vdd gnd cell_6t
Xbit_r157_c171 bl_171 br_171 wl_157 vdd gnd cell_6t
Xbit_r158_c171 bl_171 br_171 wl_158 vdd gnd cell_6t
Xbit_r159_c171 bl_171 br_171 wl_159 vdd gnd cell_6t
Xbit_r160_c171 bl_171 br_171 wl_160 vdd gnd cell_6t
Xbit_r161_c171 bl_171 br_171 wl_161 vdd gnd cell_6t
Xbit_r162_c171 bl_171 br_171 wl_162 vdd gnd cell_6t
Xbit_r163_c171 bl_171 br_171 wl_163 vdd gnd cell_6t
Xbit_r164_c171 bl_171 br_171 wl_164 vdd gnd cell_6t
Xbit_r165_c171 bl_171 br_171 wl_165 vdd gnd cell_6t
Xbit_r166_c171 bl_171 br_171 wl_166 vdd gnd cell_6t
Xbit_r167_c171 bl_171 br_171 wl_167 vdd gnd cell_6t
Xbit_r168_c171 bl_171 br_171 wl_168 vdd gnd cell_6t
Xbit_r169_c171 bl_171 br_171 wl_169 vdd gnd cell_6t
Xbit_r170_c171 bl_171 br_171 wl_170 vdd gnd cell_6t
Xbit_r171_c171 bl_171 br_171 wl_171 vdd gnd cell_6t
Xbit_r172_c171 bl_171 br_171 wl_172 vdd gnd cell_6t
Xbit_r173_c171 bl_171 br_171 wl_173 vdd gnd cell_6t
Xbit_r174_c171 bl_171 br_171 wl_174 vdd gnd cell_6t
Xbit_r175_c171 bl_171 br_171 wl_175 vdd gnd cell_6t
Xbit_r176_c171 bl_171 br_171 wl_176 vdd gnd cell_6t
Xbit_r177_c171 bl_171 br_171 wl_177 vdd gnd cell_6t
Xbit_r178_c171 bl_171 br_171 wl_178 vdd gnd cell_6t
Xbit_r179_c171 bl_171 br_171 wl_179 vdd gnd cell_6t
Xbit_r180_c171 bl_171 br_171 wl_180 vdd gnd cell_6t
Xbit_r181_c171 bl_171 br_171 wl_181 vdd gnd cell_6t
Xbit_r182_c171 bl_171 br_171 wl_182 vdd gnd cell_6t
Xbit_r183_c171 bl_171 br_171 wl_183 vdd gnd cell_6t
Xbit_r184_c171 bl_171 br_171 wl_184 vdd gnd cell_6t
Xbit_r185_c171 bl_171 br_171 wl_185 vdd gnd cell_6t
Xbit_r186_c171 bl_171 br_171 wl_186 vdd gnd cell_6t
Xbit_r187_c171 bl_171 br_171 wl_187 vdd gnd cell_6t
Xbit_r188_c171 bl_171 br_171 wl_188 vdd gnd cell_6t
Xbit_r189_c171 bl_171 br_171 wl_189 vdd gnd cell_6t
Xbit_r190_c171 bl_171 br_171 wl_190 vdd gnd cell_6t
Xbit_r191_c171 bl_171 br_171 wl_191 vdd gnd cell_6t
Xbit_r192_c171 bl_171 br_171 wl_192 vdd gnd cell_6t
Xbit_r193_c171 bl_171 br_171 wl_193 vdd gnd cell_6t
Xbit_r194_c171 bl_171 br_171 wl_194 vdd gnd cell_6t
Xbit_r195_c171 bl_171 br_171 wl_195 vdd gnd cell_6t
Xbit_r196_c171 bl_171 br_171 wl_196 vdd gnd cell_6t
Xbit_r197_c171 bl_171 br_171 wl_197 vdd gnd cell_6t
Xbit_r198_c171 bl_171 br_171 wl_198 vdd gnd cell_6t
Xbit_r199_c171 bl_171 br_171 wl_199 vdd gnd cell_6t
Xbit_r200_c171 bl_171 br_171 wl_200 vdd gnd cell_6t
Xbit_r201_c171 bl_171 br_171 wl_201 vdd gnd cell_6t
Xbit_r202_c171 bl_171 br_171 wl_202 vdd gnd cell_6t
Xbit_r203_c171 bl_171 br_171 wl_203 vdd gnd cell_6t
Xbit_r204_c171 bl_171 br_171 wl_204 vdd gnd cell_6t
Xbit_r205_c171 bl_171 br_171 wl_205 vdd gnd cell_6t
Xbit_r206_c171 bl_171 br_171 wl_206 vdd gnd cell_6t
Xbit_r207_c171 bl_171 br_171 wl_207 vdd gnd cell_6t
Xbit_r208_c171 bl_171 br_171 wl_208 vdd gnd cell_6t
Xbit_r209_c171 bl_171 br_171 wl_209 vdd gnd cell_6t
Xbit_r210_c171 bl_171 br_171 wl_210 vdd gnd cell_6t
Xbit_r211_c171 bl_171 br_171 wl_211 vdd gnd cell_6t
Xbit_r212_c171 bl_171 br_171 wl_212 vdd gnd cell_6t
Xbit_r213_c171 bl_171 br_171 wl_213 vdd gnd cell_6t
Xbit_r214_c171 bl_171 br_171 wl_214 vdd gnd cell_6t
Xbit_r215_c171 bl_171 br_171 wl_215 vdd gnd cell_6t
Xbit_r216_c171 bl_171 br_171 wl_216 vdd gnd cell_6t
Xbit_r217_c171 bl_171 br_171 wl_217 vdd gnd cell_6t
Xbit_r218_c171 bl_171 br_171 wl_218 vdd gnd cell_6t
Xbit_r219_c171 bl_171 br_171 wl_219 vdd gnd cell_6t
Xbit_r220_c171 bl_171 br_171 wl_220 vdd gnd cell_6t
Xbit_r221_c171 bl_171 br_171 wl_221 vdd gnd cell_6t
Xbit_r222_c171 bl_171 br_171 wl_222 vdd gnd cell_6t
Xbit_r223_c171 bl_171 br_171 wl_223 vdd gnd cell_6t
Xbit_r224_c171 bl_171 br_171 wl_224 vdd gnd cell_6t
Xbit_r225_c171 bl_171 br_171 wl_225 vdd gnd cell_6t
Xbit_r226_c171 bl_171 br_171 wl_226 vdd gnd cell_6t
Xbit_r227_c171 bl_171 br_171 wl_227 vdd gnd cell_6t
Xbit_r228_c171 bl_171 br_171 wl_228 vdd gnd cell_6t
Xbit_r229_c171 bl_171 br_171 wl_229 vdd gnd cell_6t
Xbit_r230_c171 bl_171 br_171 wl_230 vdd gnd cell_6t
Xbit_r231_c171 bl_171 br_171 wl_231 vdd gnd cell_6t
Xbit_r232_c171 bl_171 br_171 wl_232 vdd gnd cell_6t
Xbit_r233_c171 bl_171 br_171 wl_233 vdd gnd cell_6t
Xbit_r234_c171 bl_171 br_171 wl_234 vdd gnd cell_6t
Xbit_r235_c171 bl_171 br_171 wl_235 vdd gnd cell_6t
Xbit_r236_c171 bl_171 br_171 wl_236 vdd gnd cell_6t
Xbit_r237_c171 bl_171 br_171 wl_237 vdd gnd cell_6t
Xbit_r238_c171 bl_171 br_171 wl_238 vdd gnd cell_6t
Xbit_r239_c171 bl_171 br_171 wl_239 vdd gnd cell_6t
Xbit_r240_c171 bl_171 br_171 wl_240 vdd gnd cell_6t
Xbit_r241_c171 bl_171 br_171 wl_241 vdd gnd cell_6t
Xbit_r242_c171 bl_171 br_171 wl_242 vdd gnd cell_6t
Xbit_r243_c171 bl_171 br_171 wl_243 vdd gnd cell_6t
Xbit_r244_c171 bl_171 br_171 wl_244 vdd gnd cell_6t
Xbit_r245_c171 bl_171 br_171 wl_245 vdd gnd cell_6t
Xbit_r246_c171 bl_171 br_171 wl_246 vdd gnd cell_6t
Xbit_r247_c171 bl_171 br_171 wl_247 vdd gnd cell_6t
Xbit_r248_c171 bl_171 br_171 wl_248 vdd gnd cell_6t
Xbit_r249_c171 bl_171 br_171 wl_249 vdd gnd cell_6t
Xbit_r250_c171 bl_171 br_171 wl_250 vdd gnd cell_6t
Xbit_r251_c171 bl_171 br_171 wl_251 vdd gnd cell_6t
Xbit_r252_c171 bl_171 br_171 wl_252 vdd gnd cell_6t
Xbit_r253_c171 bl_171 br_171 wl_253 vdd gnd cell_6t
Xbit_r254_c171 bl_171 br_171 wl_254 vdd gnd cell_6t
Xbit_r255_c171 bl_171 br_171 wl_255 vdd gnd cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd cell_6t
Xbit_r1_c172 bl_172 br_172 wl_1 vdd gnd cell_6t
Xbit_r2_c172 bl_172 br_172 wl_2 vdd gnd cell_6t
Xbit_r3_c172 bl_172 br_172 wl_3 vdd gnd cell_6t
Xbit_r4_c172 bl_172 br_172 wl_4 vdd gnd cell_6t
Xbit_r5_c172 bl_172 br_172 wl_5 vdd gnd cell_6t
Xbit_r6_c172 bl_172 br_172 wl_6 vdd gnd cell_6t
Xbit_r7_c172 bl_172 br_172 wl_7 vdd gnd cell_6t
Xbit_r8_c172 bl_172 br_172 wl_8 vdd gnd cell_6t
Xbit_r9_c172 bl_172 br_172 wl_9 vdd gnd cell_6t
Xbit_r10_c172 bl_172 br_172 wl_10 vdd gnd cell_6t
Xbit_r11_c172 bl_172 br_172 wl_11 vdd gnd cell_6t
Xbit_r12_c172 bl_172 br_172 wl_12 vdd gnd cell_6t
Xbit_r13_c172 bl_172 br_172 wl_13 vdd gnd cell_6t
Xbit_r14_c172 bl_172 br_172 wl_14 vdd gnd cell_6t
Xbit_r15_c172 bl_172 br_172 wl_15 vdd gnd cell_6t
Xbit_r16_c172 bl_172 br_172 wl_16 vdd gnd cell_6t
Xbit_r17_c172 bl_172 br_172 wl_17 vdd gnd cell_6t
Xbit_r18_c172 bl_172 br_172 wl_18 vdd gnd cell_6t
Xbit_r19_c172 bl_172 br_172 wl_19 vdd gnd cell_6t
Xbit_r20_c172 bl_172 br_172 wl_20 vdd gnd cell_6t
Xbit_r21_c172 bl_172 br_172 wl_21 vdd gnd cell_6t
Xbit_r22_c172 bl_172 br_172 wl_22 vdd gnd cell_6t
Xbit_r23_c172 bl_172 br_172 wl_23 vdd gnd cell_6t
Xbit_r24_c172 bl_172 br_172 wl_24 vdd gnd cell_6t
Xbit_r25_c172 bl_172 br_172 wl_25 vdd gnd cell_6t
Xbit_r26_c172 bl_172 br_172 wl_26 vdd gnd cell_6t
Xbit_r27_c172 bl_172 br_172 wl_27 vdd gnd cell_6t
Xbit_r28_c172 bl_172 br_172 wl_28 vdd gnd cell_6t
Xbit_r29_c172 bl_172 br_172 wl_29 vdd gnd cell_6t
Xbit_r30_c172 bl_172 br_172 wl_30 vdd gnd cell_6t
Xbit_r31_c172 bl_172 br_172 wl_31 vdd gnd cell_6t
Xbit_r32_c172 bl_172 br_172 wl_32 vdd gnd cell_6t
Xbit_r33_c172 bl_172 br_172 wl_33 vdd gnd cell_6t
Xbit_r34_c172 bl_172 br_172 wl_34 vdd gnd cell_6t
Xbit_r35_c172 bl_172 br_172 wl_35 vdd gnd cell_6t
Xbit_r36_c172 bl_172 br_172 wl_36 vdd gnd cell_6t
Xbit_r37_c172 bl_172 br_172 wl_37 vdd gnd cell_6t
Xbit_r38_c172 bl_172 br_172 wl_38 vdd gnd cell_6t
Xbit_r39_c172 bl_172 br_172 wl_39 vdd gnd cell_6t
Xbit_r40_c172 bl_172 br_172 wl_40 vdd gnd cell_6t
Xbit_r41_c172 bl_172 br_172 wl_41 vdd gnd cell_6t
Xbit_r42_c172 bl_172 br_172 wl_42 vdd gnd cell_6t
Xbit_r43_c172 bl_172 br_172 wl_43 vdd gnd cell_6t
Xbit_r44_c172 bl_172 br_172 wl_44 vdd gnd cell_6t
Xbit_r45_c172 bl_172 br_172 wl_45 vdd gnd cell_6t
Xbit_r46_c172 bl_172 br_172 wl_46 vdd gnd cell_6t
Xbit_r47_c172 bl_172 br_172 wl_47 vdd gnd cell_6t
Xbit_r48_c172 bl_172 br_172 wl_48 vdd gnd cell_6t
Xbit_r49_c172 bl_172 br_172 wl_49 vdd gnd cell_6t
Xbit_r50_c172 bl_172 br_172 wl_50 vdd gnd cell_6t
Xbit_r51_c172 bl_172 br_172 wl_51 vdd gnd cell_6t
Xbit_r52_c172 bl_172 br_172 wl_52 vdd gnd cell_6t
Xbit_r53_c172 bl_172 br_172 wl_53 vdd gnd cell_6t
Xbit_r54_c172 bl_172 br_172 wl_54 vdd gnd cell_6t
Xbit_r55_c172 bl_172 br_172 wl_55 vdd gnd cell_6t
Xbit_r56_c172 bl_172 br_172 wl_56 vdd gnd cell_6t
Xbit_r57_c172 bl_172 br_172 wl_57 vdd gnd cell_6t
Xbit_r58_c172 bl_172 br_172 wl_58 vdd gnd cell_6t
Xbit_r59_c172 bl_172 br_172 wl_59 vdd gnd cell_6t
Xbit_r60_c172 bl_172 br_172 wl_60 vdd gnd cell_6t
Xbit_r61_c172 bl_172 br_172 wl_61 vdd gnd cell_6t
Xbit_r62_c172 bl_172 br_172 wl_62 vdd gnd cell_6t
Xbit_r63_c172 bl_172 br_172 wl_63 vdd gnd cell_6t
Xbit_r64_c172 bl_172 br_172 wl_64 vdd gnd cell_6t
Xbit_r65_c172 bl_172 br_172 wl_65 vdd gnd cell_6t
Xbit_r66_c172 bl_172 br_172 wl_66 vdd gnd cell_6t
Xbit_r67_c172 bl_172 br_172 wl_67 vdd gnd cell_6t
Xbit_r68_c172 bl_172 br_172 wl_68 vdd gnd cell_6t
Xbit_r69_c172 bl_172 br_172 wl_69 vdd gnd cell_6t
Xbit_r70_c172 bl_172 br_172 wl_70 vdd gnd cell_6t
Xbit_r71_c172 bl_172 br_172 wl_71 vdd gnd cell_6t
Xbit_r72_c172 bl_172 br_172 wl_72 vdd gnd cell_6t
Xbit_r73_c172 bl_172 br_172 wl_73 vdd gnd cell_6t
Xbit_r74_c172 bl_172 br_172 wl_74 vdd gnd cell_6t
Xbit_r75_c172 bl_172 br_172 wl_75 vdd gnd cell_6t
Xbit_r76_c172 bl_172 br_172 wl_76 vdd gnd cell_6t
Xbit_r77_c172 bl_172 br_172 wl_77 vdd gnd cell_6t
Xbit_r78_c172 bl_172 br_172 wl_78 vdd gnd cell_6t
Xbit_r79_c172 bl_172 br_172 wl_79 vdd gnd cell_6t
Xbit_r80_c172 bl_172 br_172 wl_80 vdd gnd cell_6t
Xbit_r81_c172 bl_172 br_172 wl_81 vdd gnd cell_6t
Xbit_r82_c172 bl_172 br_172 wl_82 vdd gnd cell_6t
Xbit_r83_c172 bl_172 br_172 wl_83 vdd gnd cell_6t
Xbit_r84_c172 bl_172 br_172 wl_84 vdd gnd cell_6t
Xbit_r85_c172 bl_172 br_172 wl_85 vdd gnd cell_6t
Xbit_r86_c172 bl_172 br_172 wl_86 vdd gnd cell_6t
Xbit_r87_c172 bl_172 br_172 wl_87 vdd gnd cell_6t
Xbit_r88_c172 bl_172 br_172 wl_88 vdd gnd cell_6t
Xbit_r89_c172 bl_172 br_172 wl_89 vdd gnd cell_6t
Xbit_r90_c172 bl_172 br_172 wl_90 vdd gnd cell_6t
Xbit_r91_c172 bl_172 br_172 wl_91 vdd gnd cell_6t
Xbit_r92_c172 bl_172 br_172 wl_92 vdd gnd cell_6t
Xbit_r93_c172 bl_172 br_172 wl_93 vdd gnd cell_6t
Xbit_r94_c172 bl_172 br_172 wl_94 vdd gnd cell_6t
Xbit_r95_c172 bl_172 br_172 wl_95 vdd gnd cell_6t
Xbit_r96_c172 bl_172 br_172 wl_96 vdd gnd cell_6t
Xbit_r97_c172 bl_172 br_172 wl_97 vdd gnd cell_6t
Xbit_r98_c172 bl_172 br_172 wl_98 vdd gnd cell_6t
Xbit_r99_c172 bl_172 br_172 wl_99 vdd gnd cell_6t
Xbit_r100_c172 bl_172 br_172 wl_100 vdd gnd cell_6t
Xbit_r101_c172 bl_172 br_172 wl_101 vdd gnd cell_6t
Xbit_r102_c172 bl_172 br_172 wl_102 vdd gnd cell_6t
Xbit_r103_c172 bl_172 br_172 wl_103 vdd gnd cell_6t
Xbit_r104_c172 bl_172 br_172 wl_104 vdd gnd cell_6t
Xbit_r105_c172 bl_172 br_172 wl_105 vdd gnd cell_6t
Xbit_r106_c172 bl_172 br_172 wl_106 vdd gnd cell_6t
Xbit_r107_c172 bl_172 br_172 wl_107 vdd gnd cell_6t
Xbit_r108_c172 bl_172 br_172 wl_108 vdd gnd cell_6t
Xbit_r109_c172 bl_172 br_172 wl_109 vdd gnd cell_6t
Xbit_r110_c172 bl_172 br_172 wl_110 vdd gnd cell_6t
Xbit_r111_c172 bl_172 br_172 wl_111 vdd gnd cell_6t
Xbit_r112_c172 bl_172 br_172 wl_112 vdd gnd cell_6t
Xbit_r113_c172 bl_172 br_172 wl_113 vdd gnd cell_6t
Xbit_r114_c172 bl_172 br_172 wl_114 vdd gnd cell_6t
Xbit_r115_c172 bl_172 br_172 wl_115 vdd gnd cell_6t
Xbit_r116_c172 bl_172 br_172 wl_116 vdd gnd cell_6t
Xbit_r117_c172 bl_172 br_172 wl_117 vdd gnd cell_6t
Xbit_r118_c172 bl_172 br_172 wl_118 vdd gnd cell_6t
Xbit_r119_c172 bl_172 br_172 wl_119 vdd gnd cell_6t
Xbit_r120_c172 bl_172 br_172 wl_120 vdd gnd cell_6t
Xbit_r121_c172 bl_172 br_172 wl_121 vdd gnd cell_6t
Xbit_r122_c172 bl_172 br_172 wl_122 vdd gnd cell_6t
Xbit_r123_c172 bl_172 br_172 wl_123 vdd gnd cell_6t
Xbit_r124_c172 bl_172 br_172 wl_124 vdd gnd cell_6t
Xbit_r125_c172 bl_172 br_172 wl_125 vdd gnd cell_6t
Xbit_r126_c172 bl_172 br_172 wl_126 vdd gnd cell_6t
Xbit_r127_c172 bl_172 br_172 wl_127 vdd gnd cell_6t
Xbit_r128_c172 bl_172 br_172 wl_128 vdd gnd cell_6t
Xbit_r129_c172 bl_172 br_172 wl_129 vdd gnd cell_6t
Xbit_r130_c172 bl_172 br_172 wl_130 vdd gnd cell_6t
Xbit_r131_c172 bl_172 br_172 wl_131 vdd gnd cell_6t
Xbit_r132_c172 bl_172 br_172 wl_132 vdd gnd cell_6t
Xbit_r133_c172 bl_172 br_172 wl_133 vdd gnd cell_6t
Xbit_r134_c172 bl_172 br_172 wl_134 vdd gnd cell_6t
Xbit_r135_c172 bl_172 br_172 wl_135 vdd gnd cell_6t
Xbit_r136_c172 bl_172 br_172 wl_136 vdd gnd cell_6t
Xbit_r137_c172 bl_172 br_172 wl_137 vdd gnd cell_6t
Xbit_r138_c172 bl_172 br_172 wl_138 vdd gnd cell_6t
Xbit_r139_c172 bl_172 br_172 wl_139 vdd gnd cell_6t
Xbit_r140_c172 bl_172 br_172 wl_140 vdd gnd cell_6t
Xbit_r141_c172 bl_172 br_172 wl_141 vdd gnd cell_6t
Xbit_r142_c172 bl_172 br_172 wl_142 vdd gnd cell_6t
Xbit_r143_c172 bl_172 br_172 wl_143 vdd gnd cell_6t
Xbit_r144_c172 bl_172 br_172 wl_144 vdd gnd cell_6t
Xbit_r145_c172 bl_172 br_172 wl_145 vdd gnd cell_6t
Xbit_r146_c172 bl_172 br_172 wl_146 vdd gnd cell_6t
Xbit_r147_c172 bl_172 br_172 wl_147 vdd gnd cell_6t
Xbit_r148_c172 bl_172 br_172 wl_148 vdd gnd cell_6t
Xbit_r149_c172 bl_172 br_172 wl_149 vdd gnd cell_6t
Xbit_r150_c172 bl_172 br_172 wl_150 vdd gnd cell_6t
Xbit_r151_c172 bl_172 br_172 wl_151 vdd gnd cell_6t
Xbit_r152_c172 bl_172 br_172 wl_152 vdd gnd cell_6t
Xbit_r153_c172 bl_172 br_172 wl_153 vdd gnd cell_6t
Xbit_r154_c172 bl_172 br_172 wl_154 vdd gnd cell_6t
Xbit_r155_c172 bl_172 br_172 wl_155 vdd gnd cell_6t
Xbit_r156_c172 bl_172 br_172 wl_156 vdd gnd cell_6t
Xbit_r157_c172 bl_172 br_172 wl_157 vdd gnd cell_6t
Xbit_r158_c172 bl_172 br_172 wl_158 vdd gnd cell_6t
Xbit_r159_c172 bl_172 br_172 wl_159 vdd gnd cell_6t
Xbit_r160_c172 bl_172 br_172 wl_160 vdd gnd cell_6t
Xbit_r161_c172 bl_172 br_172 wl_161 vdd gnd cell_6t
Xbit_r162_c172 bl_172 br_172 wl_162 vdd gnd cell_6t
Xbit_r163_c172 bl_172 br_172 wl_163 vdd gnd cell_6t
Xbit_r164_c172 bl_172 br_172 wl_164 vdd gnd cell_6t
Xbit_r165_c172 bl_172 br_172 wl_165 vdd gnd cell_6t
Xbit_r166_c172 bl_172 br_172 wl_166 vdd gnd cell_6t
Xbit_r167_c172 bl_172 br_172 wl_167 vdd gnd cell_6t
Xbit_r168_c172 bl_172 br_172 wl_168 vdd gnd cell_6t
Xbit_r169_c172 bl_172 br_172 wl_169 vdd gnd cell_6t
Xbit_r170_c172 bl_172 br_172 wl_170 vdd gnd cell_6t
Xbit_r171_c172 bl_172 br_172 wl_171 vdd gnd cell_6t
Xbit_r172_c172 bl_172 br_172 wl_172 vdd gnd cell_6t
Xbit_r173_c172 bl_172 br_172 wl_173 vdd gnd cell_6t
Xbit_r174_c172 bl_172 br_172 wl_174 vdd gnd cell_6t
Xbit_r175_c172 bl_172 br_172 wl_175 vdd gnd cell_6t
Xbit_r176_c172 bl_172 br_172 wl_176 vdd gnd cell_6t
Xbit_r177_c172 bl_172 br_172 wl_177 vdd gnd cell_6t
Xbit_r178_c172 bl_172 br_172 wl_178 vdd gnd cell_6t
Xbit_r179_c172 bl_172 br_172 wl_179 vdd gnd cell_6t
Xbit_r180_c172 bl_172 br_172 wl_180 vdd gnd cell_6t
Xbit_r181_c172 bl_172 br_172 wl_181 vdd gnd cell_6t
Xbit_r182_c172 bl_172 br_172 wl_182 vdd gnd cell_6t
Xbit_r183_c172 bl_172 br_172 wl_183 vdd gnd cell_6t
Xbit_r184_c172 bl_172 br_172 wl_184 vdd gnd cell_6t
Xbit_r185_c172 bl_172 br_172 wl_185 vdd gnd cell_6t
Xbit_r186_c172 bl_172 br_172 wl_186 vdd gnd cell_6t
Xbit_r187_c172 bl_172 br_172 wl_187 vdd gnd cell_6t
Xbit_r188_c172 bl_172 br_172 wl_188 vdd gnd cell_6t
Xbit_r189_c172 bl_172 br_172 wl_189 vdd gnd cell_6t
Xbit_r190_c172 bl_172 br_172 wl_190 vdd gnd cell_6t
Xbit_r191_c172 bl_172 br_172 wl_191 vdd gnd cell_6t
Xbit_r192_c172 bl_172 br_172 wl_192 vdd gnd cell_6t
Xbit_r193_c172 bl_172 br_172 wl_193 vdd gnd cell_6t
Xbit_r194_c172 bl_172 br_172 wl_194 vdd gnd cell_6t
Xbit_r195_c172 bl_172 br_172 wl_195 vdd gnd cell_6t
Xbit_r196_c172 bl_172 br_172 wl_196 vdd gnd cell_6t
Xbit_r197_c172 bl_172 br_172 wl_197 vdd gnd cell_6t
Xbit_r198_c172 bl_172 br_172 wl_198 vdd gnd cell_6t
Xbit_r199_c172 bl_172 br_172 wl_199 vdd gnd cell_6t
Xbit_r200_c172 bl_172 br_172 wl_200 vdd gnd cell_6t
Xbit_r201_c172 bl_172 br_172 wl_201 vdd gnd cell_6t
Xbit_r202_c172 bl_172 br_172 wl_202 vdd gnd cell_6t
Xbit_r203_c172 bl_172 br_172 wl_203 vdd gnd cell_6t
Xbit_r204_c172 bl_172 br_172 wl_204 vdd gnd cell_6t
Xbit_r205_c172 bl_172 br_172 wl_205 vdd gnd cell_6t
Xbit_r206_c172 bl_172 br_172 wl_206 vdd gnd cell_6t
Xbit_r207_c172 bl_172 br_172 wl_207 vdd gnd cell_6t
Xbit_r208_c172 bl_172 br_172 wl_208 vdd gnd cell_6t
Xbit_r209_c172 bl_172 br_172 wl_209 vdd gnd cell_6t
Xbit_r210_c172 bl_172 br_172 wl_210 vdd gnd cell_6t
Xbit_r211_c172 bl_172 br_172 wl_211 vdd gnd cell_6t
Xbit_r212_c172 bl_172 br_172 wl_212 vdd gnd cell_6t
Xbit_r213_c172 bl_172 br_172 wl_213 vdd gnd cell_6t
Xbit_r214_c172 bl_172 br_172 wl_214 vdd gnd cell_6t
Xbit_r215_c172 bl_172 br_172 wl_215 vdd gnd cell_6t
Xbit_r216_c172 bl_172 br_172 wl_216 vdd gnd cell_6t
Xbit_r217_c172 bl_172 br_172 wl_217 vdd gnd cell_6t
Xbit_r218_c172 bl_172 br_172 wl_218 vdd gnd cell_6t
Xbit_r219_c172 bl_172 br_172 wl_219 vdd gnd cell_6t
Xbit_r220_c172 bl_172 br_172 wl_220 vdd gnd cell_6t
Xbit_r221_c172 bl_172 br_172 wl_221 vdd gnd cell_6t
Xbit_r222_c172 bl_172 br_172 wl_222 vdd gnd cell_6t
Xbit_r223_c172 bl_172 br_172 wl_223 vdd gnd cell_6t
Xbit_r224_c172 bl_172 br_172 wl_224 vdd gnd cell_6t
Xbit_r225_c172 bl_172 br_172 wl_225 vdd gnd cell_6t
Xbit_r226_c172 bl_172 br_172 wl_226 vdd gnd cell_6t
Xbit_r227_c172 bl_172 br_172 wl_227 vdd gnd cell_6t
Xbit_r228_c172 bl_172 br_172 wl_228 vdd gnd cell_6t
Xbit_r229_c172 bl_172 br_172 wl_229 vdd gnd cell_6t
Xbit_r230_c172 bl_172 br_172 wl_230 vdd gnd cell_6t
Xbit_r231_c172 bl_172 br_172 wl_231 vdd gnd cell_6t
Xbit_r232_c172 bl_172 br_172 wl_232 vdd gnd cell_6t
Xbit_r233_c172 bl_172 br_172 wl_233 vdd gnd cell_6t
Xbit_r234_c172 bl_172 br_172 wl_234 vdd gnd cell_6t
Xbit_r235_c172 bl_172 br_172 wl_235 vdd gnd cell_6t
Xbit_r236_c172 bl_172 br_172 wl_236 vdd gnd cell_6t
Xbit_r237_c172 bl_172 br_172 wl_237 vdd gnd cell_6t
Xbit_r238_c172 bl_172 br_172 wl_238 vdd gnd cell_6t
Xbit_r239_c172 bl_172 br_172 wl_239 vdd gnd cell_6t
Xbit_r240_c172 bl_172 br_172 wl_240 vdd gnd cell_6t
Xbit_r241_c172 bl_172 br_172 wl_241 vdd gnd cell_6t
Xbit_r242_c172 bl_172 br_172 wl_242 vdd gnd cell_6t
Xbit_r243_c172 bl_172 br_172 wl_243 vdd gnd cell_6t
Xbit_r244_c172 bl_172 br_172 wl_244 vdd gnd cell_6t
Xbit_r245_c172 bl_172 br_172 wl_245 vdd gnd cell_6t
Xbit_r246_c172 bl_172 br_172 wl_246 vdd gnd cell_6t
Xbit_r247_c172 bl_172 br_172 wl_247 vdd gnd cell_6t
Xbit_r248_c172 bl_172 br_172 wl_248 vdd gnd cell_6t
Xbit_r249_c172 bl_172 br_172 wl_249 vdd gnd cell_6t
Xbit_r250_c172 bl_172 br_172 wl_250 vdd gnd cell_6t
Xbit_r251_c172 bl_172 br_172 wl_251 vdd gnd cell_6t
Xbit_r252_c172 bl_172 br_172 wl_252 vdd gnd cell_6t
Xbit_r253_c172 bl_172 br_172 wl_253 vdd gnd cell_6t
Xbit_r254_c172 bl_172 br_172 wl_254 vdd gnd cell_6t
Xbit_r255_c172 bl_172 br_172 wl_255 vdd gnd cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd cell_6t
Xbit_r1_c173 bl_173 br_173 wl_1 vdd gnd cell_6t
Xbit_r2_c173 bl_173 br_173 wl_2 vdd gnd cell_6t
Xbit_r3_c173 bl_173 br_173 wl_3 vdd gnd cell_6t
Xbit_r4_c173 bl_173 br_173 wl_4 vdd gnd cell_6t
Xbit_r5_c173 bl_173 br_173 wl_5 vdd gnd cell_6t
Xbit_r6_c173 bl_173 br_173 wl_6 vdd gnd cell_6t
Xbit_r7_c173 bl_173 br_173 wl_7 vdd gnd cell_6t
Xbit_r8_c173 bl_173 br_173 wl_8 vdd gnd cell_6t
Xbit_r9_c173 bl_173 br_173 wl_9 vdd gnd cell_6t
Xbit_r10_c173 bl_173 br_173 wl_10 vdd gnd cell_6t
Xbit_r11_c173 bl_173 br_173 wl_11 vdd gnd cell_6t
Xbit_r12_c173 bl_173 br_173 wl_12 vdd gnd cell_6t
Xbit_r13_c173 bl_173 br_173 wl_13 vdd gnd cell_6t
Xbit_r14_c173 bl_173 br_173 wl_14 vdd gnd cell_6t
Xbit_r15_c173 bl_173 br_173 wl_15 vdd gnd cell_6t
Xbit_r16_c173 bl_173 br_173 wl_16 vdd gnd cell_6t
Xbit_r17_c173 bl_173 br_173 wl_17 vdd gnd cell_6t
Xbit_r18_c173 bl_173 br_173 wl_18 vdd gnd cell_6t
Xbit_r19_c173 bl_173 br_173 wl_19 vdd gnd cell_6t
Xbit_r20_c173 bl_173 br_173 wl_20 vdd gnd cell_6t
Xbit_r21_c173 bl_173 br_173 wl_21 vdd gnd cell_6t
Xbit_r22_c173 bl_173 br_173 wl_22 vdd gnd cell_6t
Xbit_r23_c173 bl_173 br_173 wl_23 vdd gnd cell_6t
Xbit_r24_c173 bl_173 br_173 wl_24 vdd gnd cell_6t
Xbit_r25_c173 bl_173 br_173 wl_25 vdd gnd cell_6t
Xbit_r26_c173 bl_173 br_173 wl_26 vdd gnd cell_6t
Xbit_r27_c173 bl_173 br_173 wl_27 vdd gnd cell_6t
Xbit_r28_c173 bl_173 br_173 wl_28 vdd gnd cell_6t
Xbit_r29_c173 bl_173 br_173 wl_29 vdd gnd cell_6t
Xbit_r30_c173 bl_173 br_173 wl_30 vdd gnd cell_6t
Xbit_r31_c173 bl_173 br_173 wl_31 vdd gnd cell_6t
Xbit_r32_c173 bl_173 br_173 wl_32 vdd gnd cell_6t
Xbit_r33_c173 bl_173 br_173 wl_33 vdd gnd cell_6t
Xbit_r34_c173 bl_173 br_173 wl_34 vdd gnd cell_6t
Xbit_r35_c173 bl_173 br_173 wl_35 vdd gnd cell_6t
Xbit_r36_c173 bl_173 br_173 wl_36 vdd gnd cell_6t
Xbit_r37_c173 bl_173 br_173 wl_37 vdd gnd cell_6t
Xbit_r38_c173 bl_173 br_173 wl_38 vdd gnd cell_6t
Xbit_r39_c173 bl_173 br_173 wl_39 vdd gnd cell_6t
Xbit_r40_c173 bl_173 br_173 wl_40 vdd gnd cell_6t
Xbit_r41_c173 bl_173 br_173 wl_41 vdd gnd cell_6t
Xbit_r42_c173 bl_173 br_173 wl_42 vdd gnd cell_6t
Xbit_r43_c173 bl_173 br_173 wl_43 vdd gnd cell_6t
Xbit_r44_c173 bl_173 br_173 wl_44 vdd gnd cell_6t
Xbit_r45_c173 bl_173 br_173 wl_45 vdd gnd cell_6t
Xbit_r46_c173 bl_173 br_173 wl_46 vdd gnd cell_6t
Xbit_r47_c173 bl_173 br_173 wl_47 vdd gnd cell_6t
Xbit_r48_c173 bl_173 br_173 wl_48 vdd gnd cell_6t
Xbit_r49_c173 bl_173 br_173 wl_49 vdd gnd cell_6t
Xbit_r50_c173 bl_173 br_173 wl_50 vdd gnd cell_6t
Xbit_r51_c173 bl_173 br_173 wl_51 vdd gnd cell_6t
Xbit_r52_c173 bl_173 br_173 wl_52 vdd gnd cell_6t
Xbit_r53_c173 bl_173 br_173 wl_53 vdd gnd cell_6t
Xbit_r54_c173 bl_173 br_173 wl_54 vdd gnd cell_6t
Xbit_r55_c173 bl_173 br_173 wl_55 vdd gnd cell_6t
Xbit_r56_c173 bl_173 br_173 wl_56 vdd gnd cell_6t
Xbit_r57_c173 bl_173 br_173 wl_57 vdd gnd cell_6t
Xbit_r58_c173 bl_173 br_173 wl_58 vdd gnd cell_6t
Xbit_r59_c173 bl_173 br_173 wl_59 vdd gnd cell_6t
Xbit_r60_c173 bl_173 br_173 wl_60 vdd gnd cell_6t
Xbit_r61_c173 bl_173 br_173 wl_61 vdd gnd cell_6t
Xbit_r62_c173 bl_173 br_173 wl_62 vdd gnd cell_6t
Xbit_r63_c173 bl_173 br_173 wl_63 vdd gnd cell_6t
Xbit_r64_c173 bl_173 br_173 wl_64 vdd gnd cell_6t
Xbit_r65_c173 bl_173 br_173 wl_65 vdd gnd cell_6t
Xbit_r66_c173 bl_173 br_173 wl_66 vdd gnd cell_6t
Xbit_r67_c173 bl_173 br_173 wl_67 vdd gnd cell_6t
Xbit_r68_c173 bl_173 br_173 wl_68 vdd gnd cell_6t
Xbit_r69_c173 bl_173 br_173 wl_69 vdd gnd cell_6t
Xbit_r70_c173 bl_173 br_173 wl_70 vdd gnd cell_6t
Xbit_r71_c173 bl_173 br_173 wl_71 vdd gnd cell_6t
Xbit_r72_c173 bl_173 br_173 wl_72 vdd gnd cell_6t
Xbit_r73_c173 bl_173 br_173 wl_73 vdd gnd cell_6t
Xbit_r74_c173 bl_173 br_173 wl_74 vdd gnd cell_6t
Xbit_r75_c173 bl_173 br_173 wl_75 vdd gnd cell_6t
Xbit_r76_c173 bl_173 br_173 wl_76 vdd gnd cell_6t
Xbit_r77_c173 bl_173 br_173 wl_77 vdd gnd cell_6t
Xbit_r78_c173 bl_173 br_173 wl_78 vdd gnd cell_6t
Xbit_r79_c173 bl_173 br_173 wl_79 vdd gnd cell_6t
Xbit_r80_c173 bl_173 br_173 wl_80 vdd gnd cell_6t
Xbit_r81_c173 bl_173 br_173 wl_81 vdd gnd cell_6t
Xbit_r82_c173 bl_173 br_173 wl_82 vdd gnd cell_6t
Xbit_r83_c173 bl_173 br_173 wl_83 vdd gnd cell_6t
Xbit_r84_c173 bl_173 br_173 wl_84 vdd gnd cell_6t
Xbit_r85_c173 bl_173 br_173 wl_85 vdd gnd cell_6t
Xbit_r86_c173 bl_173 br_173 wl_86 vdd gnd cell_6t
Xbit_r87_c173 bl_173 br_173 wl_87 vdd gnd cell_6t
Xbit_r88_c173 bl_173 br_173 wl_88 vdd gnd cell_6t
Xbit_r89_c173 bl_173 br_173 wl_89 vdd gnd cell_6t
Xbit_r90_c173 bl_173 br_173 wl_90 vdd gnd cell_6t
Xbit_r91_c173 bl_173 br_173 wl_91 vdd gnd cell_6t
Xbit_r92_c173 bl_173 br_173 wl_92 vdd gnd cell_6t
Xbit_r93_c173 bl_173 br_173 wl_93 vdd gnd cell_6t
Xbit_r94_c173 bl_173 br_173 wl_94 vdd gnd cell_6t
Xbit_r95_c173 bl_173 br_173 wl_95 vdd gnd cell_6t
Xbit_r96_c173 bl_173 br_173 wl_96 vdd gnd cell_6t
Xbit_r97_c173 bl_173 br_173 wl_97 vdd gnd cell_6t
Xbit_r98_c173 bl_173 br_173 wl_98 vdd gnd cell_6t
Xbit_r99_c173 bl_173 br_173 wl_99 vdd gnd cell_6t
Xbit_r100_c173 bl_173 br_173 wl_100 vdd gnd cell_6t
Xbit_r101_c173 bl_173 br_173 wl_101 vdd gnd cell_6t
Xbit_r102_c173 bl_173 br_173 wl_102 vdd gnd cell_6t
Xbit_r103_c173 bl_173 br_173 wl_103 vdd gnd cell_6t
Xbit_r104_c173 bl_173 br_173 wl_104 vdd gnd cell_6t
Xbit_r105_c173 bl_173 br_173 wl_105 vdd gnd cell_6t
Xbit_r106_c173 bl_173 br_173 wl_106 vdd gnd cell_6t
Xbit_r107_c173 bl_173 br_173 wl_107 vdd gnd cell_6t
Xbit_r108_c173 bl_173 br_173 wl_108 vdd gnd cell_6t
Xbit_r109_c173 bl_173 br_173 wl_109 vdd gnd cell_6t
Xbit_r110_c173 bl_173 br_173 wl_110 vdd gnd cell_6t
Xbit_r111_c173 bl_173 br_173 wl_111 vdd gnd cell_6t
Xbit_r112_c173 bl_173 br_173 wl_112 vdd gnd cell_6t
Xbit_r113_c173 bl_173 br_173 wl_113 vdd gnd cell_6t
Xbit_r114_c173 bl_173 br_173 wl_114 vdd gnd cell_6t
Xbit_r115_c173 bl_173 br_173 wl_115 vdd gnd cell_6t
Xbit_r116_c173 bl_173 br_173 wl_116 vdd gnd cell_6t
Xbit_r117_c173 bl_173 br_173 wl_117 vdd gnd cell_6t
Xbit_r118_c173 bl_173 br_173 wl_118 vdd gnd cell_6t
Xbit_r119_c173 bl_173 br_173 wl_119 vdd gnd cell_6t
Xbit_r120_c173 bl_173 br_173 wl_120 vdd gnd cell_6t
Xbit_r121_c173 bl_173 br_173 wl_121 vdd gnd cell_6t
Xbit_r122_c173 bl_173 br_173 wl_122 vdd gnd cell_6t
Xbit_r123_c173 bl_173 br_173 wl_123 vdd gnd cell_6t
Xbit_r124_c173 bl_173 br_173 wl_124 vdd gnd cell_6t
Xbit_r125_c173 bl_173 br_173 wl_125 vdd gnd cell_6t
Xbit_r126_c173 bl_173 br_173 wl_126 vdd gnd cell_6t
Xbit_r127_c173 bl_173 br_173 wl_127 vdd gnd cell_6t
Xbit_r128_c173 bl_173 br_173 wl_128 vdd gnd cell_6t
Xbit_r129_c173 bl_173 br_173 wl_129 vdd gnd cell_6t
Xbit_r130_c173 bl_173 br_173 wl_130 vdd gnd cell_6t
Xbit_r131_c173 bl_173 br_173 wl_131 vdd gnd cell_6t
Xbit_r132_c173 bl_173 br_173 wl_132 vdd gnd cell_6t
Xbit_r133_c173 bl_173 br_173 wl_133 vdd gnd cell_6t
Xbit_r134_c173 bl_173 br_173 wl_134 vdd gnd cell_6t
Xbit_r135_c173 bl_173 br_173 wl_135 vdd gnd cell_6t
Xbit_r136_c173 bl_173 br_173 wl_136 vdd gnd cell_6t
Xbit_r137_c173 bl_173 br_173 wl_137 vdd gnd cell_6t
Xbit_r138_c173 bl_173 br_173 wl_138 vdd gnd cell_6t
Xbit_r139_c173 bl_173 br_173 wl_139 vdd gnd cell_6t
Xbit_r140_c173 bl_173 br_173 wl_140 vdd gnd cell_6t
Xbit_r141_c173 bl_173 br_173 wl_141 vdd gnd cell_6t
Xbit_r142_c173 bl_173 br_173 wl_142 vdd gnd cell_6t
Xbit_r143_c173 bl_173 br_173 wl_143 vdd gnd cell_6t
Xbit_r144_c173 bl_173 br_173 wl_144 vdd gnd cell_6t
Xbit_r145_c173 bl_173 br_173 wl_145 vdd gnd cell_6t
Xbit_r146_c173 bl_173 br_173 wl_146 vdd gnd cell_6t
Xbit_r147_c173 bl_173 br_173 wl_147 vdd gnd cell_6t
Xbit_r148_c173 bl_173 br_173 wl_148 vdd gnd cell_6t
Xbit_r149_c173 bl_173 br_173 wl_149 vdd gnd cell_6t
Xbit_r150_c173 bl_173 br_173 wl_150 vdd gnd cell_6t
Xbit_r151_c173 bl_173 br_173 wl_151 vdd gnd cell_6t
Xbit_r152_c173 bl_173 br_173 wl_152 vdd gnd cell_6t
Xbit_r153_c173 bl_173 br_173 wl_153 vdd gnd cell_6t
Xbit_r154_c173 bl_173 br_173 wl_154 vdd gnd cell_6t
Xbit_r155_c173 bl_173 br_173 wl_155 vdd gnd cell_6t
Xbit_r156_c173 bl_173 br_173 wl_156 vdd gnd cell_6t
Xbit_r157_c173 bl_173 br_173 wl_157 vdd gnd cell_6t
Xbit_r158_c173 bl_173 br_173 wl_158 vdd gnd cell_6t
Xbit_r159_c173 bl_173 br_173 wl_159 vdd gnd cell_6t
Xbit_r160_c173 bl_173 br_173 wl_160 vdd gnd cell_6t
Xbit_r161_c173 bl_173 br_173 wl_161 vdd gnd cell_6t
Xbit_r162_c173 bl_173 br_173 wl_162 vdd gnd cell_6t
Xbit_r163_c173 bl_173 br_173 wl_163 vdd gnd cell_6t
Xbit_r164_c173 bl_173 br_173 wl_164 vdd gnd cell_6t
Xbit_r165_c173 bl_173 br_173 wl_165 vdd gnd cell_6t
Xbit_r166_c173 bl_173 br_173 wl_166 vdd gnd cell_6t
Xbit_r167_c173 bl_173 br_173 wl_167 vdd gnd cell_6t
Xbit_r168_c173 bl_173 br_173 wl_168 vdd gnd cell_6t
Xbit_r169_c173 bl_173 br_173 wl_169 vdd gnd cell_6t
Xbit_r170_c173 bl_173 br_173 wl_170 vdd gnd cell_6t
Xbit_r171_c173 bl_173 br_173 wl_171 vdd gnd cell_6t
Xbit_r172_c173 bl_173 br_173 wl_172 vdd gnd cell_6t
Xbit_r173_c173 bl_173 br_173 wl_173 vdd gnd cell_6t
Xbit_r174_c173 bl_173 br_173 wl_174 vdd gnd cell_6t
Xbit_r175_c173 bl_173 br_173 wl_175 vdd gnd cell_6t
Xbit_r176_c173 bl_173 br_173 wl_176 vdd gnd cell_6t
Xbit_r177_c173 bl_173 br_173 wl_177 vdd gnd cell_6t
Xbit_r178_c173 bl_173 br_173 wl_178 vdd gnd cell_6t
Xbit_r179_c173 bl_173 br_173 wl_179 vdd gnd cell_6t
Xbit_r180_c173 bl_173 br_173 wl_180 vdd gnd cell_6t
Xbit_r181_c173 bl_173 br_173 wl_181 vdd gnd cell_6t
Xbit_r182_c173 bl_173 br_173 wl_182 vdd gnd cell_6t
Xbit_r183_c173 bl_173 br_173 wl_183 vdd gnd cell_6t
Xbit_r184_c173 bl_173 br_173 wl_184 vdd gnd cell_6t
Xbit_r185_c173 bl_173 br_173 wl_185 vdd gnd cell_6t
Xbit_r186_c173 bl_173 br_173 wl_186 vdd gnd cell_6t
Xbit_r187_c173 bl_173 br_173 wl_187 vdd gnd cell_6t
Xbit_r188_c173 bl_173 br_173 wl_188 vdd gnd cell_6t
Xbit_r189_c173 bl_173 br_173 wl_189 vdd gnd cell_6t
Xbit_r190_c173 bl_173 br_173 wl_190 vdd gnd cell_6t
Xbit_r191_c173 bl_173 br_173 wl_191 vdd gnd cell_6t
Xbit_r192_c173 bl_173 br_173 wl_192 vdd gnd cell_6t
Xbit_r193_c173 bl_173 br_173 wl_193 vdd gnd cell_6t
Xbit_r194_c173 bl_173 br_173 wl_194 vdd gnd cell_6t
Xbit_r195_c173 bl_173 br_173 wl_195 vdd gnd cell_6t
Xbit_r196_c173 bl_173 br_173 wl_196 vdd gnd cell_6t
Xbit_r197_c173 bl_173 br_173 wl_197 vdd gnd cell_6t
Xbit_r198_c173 bl_173 br_173 wl_198 vdd gnd cell_6t
Xbit_r199_c173 bl_173 br_173 wl_199 vdd gnd cell_6t
Xbit_r200_c173 bl_173 br_173 wl_200 vdd gnd cell_6t
Xbit_r201_c173 bl_173 br_173 wl_201 vdd gnd cell_6t
Xbit_r202_c173 bl_173 br_173 wl_202 vdd gnd cell_6t
Xbit_r203_c173 bl_173 br_173 wl_203 vdd gnd cell_6t
Xbit_r204_c173 bl_173 br_173 wl_204 vdd gnd cell_6t
Xbit_r205_c173 bl_173 br_173 wl_205 vdd gnd cell_6t
Xbit_r206_c173 bl_173 br_173 wl_206 vdd gnd cell_6t
Xbit_r207_c173 bl_173 br_173 wl_207 vdd gnd cell_6t
Xbit_r208_c173 bl_173 br_173 wl_208 vdd gnd cell_6t
Xbit_r209_c173 bl_173 br_173 wl_209 vdd gnd cell_6t
Xbit_r210_c173 bl_173 br_173 wl_210 vdd gnd cell_6t
Xbit_r211_c173 bl_173 br_173 wl_211 vdd gnd cell_6t
Xbit_r212_c173 bl_173 br_173 wl_212 vdd gnd cell_6t
Xbit_r213_c173 bl_173 br_173 wl_213 vdd gnd cell_6t
Xbit_r214_c173 bl_173 br_173 wl_214 vdd gnd cell_6t
Xbit_r215_c173 bl_173 br_173 wl_215 vdd gnd cell_6t
Xbit_r216_c173 bl_173 br_173 wl_216 vdd gnd cell_6t
Xbit_r217_c173 bl_173 br_173 wl_217 vdd gnd cell_6t
Xbit_r218_c173 bl_173 br_173 wl_218 vdd gnd cell_6t
Xbit_r219_c173 bl_173 br_173 wl_219 vdd gnd cell_6t
Xbit_r220_c173 bl_173 br_173 wl_220 vdd gnd cell_6t
Xbit_r221_c173 bl_173 br_173 wl_221 vdd gnd cell_6t
Xbit_r222_c173 bl_173 br_173 wl_222 vdd gnd cell_6t
Xbit_r223_c173 bl_173 br_173 wl_223 vdd gnd cell_6t
Xbit_r224_c173 bl_173 br_173 wl_224 vdd gnd cell_6t
Xbit_r225_c173 bl_173 br_173 wl_225 vdd gnd cell_6t
Xbit_r226_c173 bl_173 br_173 wl_226 vdd gnd cell_6t
Xbit_r227_c173 bl_173 br_173 wl_227 vdd gnd cell_6t
Xbit_r228_c173 bl_173 br_173 wl_228 vdd gnd cell_6t
Xbit_r229_c173 bl_173 br_173 wl_229 vdd gnd cell_6t
Xbit_r230_c173 bl_173 br_173 wl_230 vdd gnd cell_6t
Xbit_r231_c173 bl_173 br_173 wl_231 vdd gnd cell_6t
Xbit_r232_c173 bl_173 br_173 wl_232 vdd gnd cell_6t
Xbit_r233_c173 bl_173 br_173 wl_233 vdd gnd cell_6t
Xbit_r234_c173 bl_173 br_173 wl_234 vdd gnd cell_6t
Xbit_r235_c173 bl_173 br_173 wl_235 vdd gnd cell_6t
Xbit_r236_c173 bl_173 br_173 wl_236 vdd gnd cell_6t
Xbit_r237_c173 bl_173 br_173 wl_237 vdd gnd cell_6t
Xbit_r238_c173 bl_173 br_173 wl_238 vdd gnd cell_6t
Xbit_r239_c173 bl_173 br_173 wl_239 vdd gnd cell_6t
Xbit_r240_c173 bl_173 br_173 wl_240 vdd gnd cell_6t
Xbit_r241_c173 bl_173 br_173 wl_241 vdd gnd cell_6t
Xbit_r242_c173 bl_173 br_173 wl_242 vdd gnd cell_6t
Xbit_r243_c173 bl_173 br_173 wl_243 vdd gnd cell_6t
Xbit_r244_c173 bl_173 br_173 wl_244 vdd gnd cell_6t
Xbit_r245_c173 bl_173 br_173 wl_245 vdd gnd cell_6t
Xbit_r246_c173 bl_173 br_173 wl_246 vdd gnd cell_6t
Xbit_r247_c173 bl_173 br_173 wl_247 vdd gnd cell_6t
Xbit_r248_c173 bl_173 br_173 wl_248 vdd gnd cell_6t
Xbit_r249_c173 bl_173 br_173 wl_249 vdd gnd cell_6t
Xbit_r250_c173 bl_173 br_173 wl_250 vdd gnd cell_6t
Xbit_r251_c173 bl_173 br_173 wl_251 vdd gnd cell_6t
Xbit_r252_c173 bl_173 br_173 wl_252 vdd gnd cell_6t
Xbit_r253_c173 bl_173 br_173 wl_253 vdd gnd cell_6t
Xbit_r254_c173 bl_173 br_173 wl_254 vdd gnd cell_6t
Xbit_r255_c173 bl_173 br_173 wl_255 vdd gnd cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd cell_6t
Xbit_r1_c174 bl_174 br_174 wl_1 vdd gnd cell_6t
Xbit_r2_c174 bl_174 br_174 wl_2 vdd gnd cell_6t
Xbit_r3_c174 bl_174 br_174 wl_3 vdd gnd cell_6t
Xbit_r4_c174 bl_174 br_174 wl_4 vdd gnd cell_6t
Xbit_r5_c174 bl_174 br_174 wl_5 vdd gnd cell_6t
Xbit_r6_c174 bl_174 br_174 wl_6 vdd gnd cell_6t
Xbit_r7_c174 bl_174 br_174 wl_7 vdd gnd cell_6t
Xbit_r8_c174 bl_174 br_174 wl_8 vdd gnd cell_6t
Xbit_r9_c174 bl_174 br_174 wl_9 vdd gnd cell_6t
Xbit_r10_c174 bl_174 br_174 wl_10 vdd gnd cell_6t
Xbit_r11_c174 bl_174 br_174 wl_11 vdd gnd cell_6t
Xbit_r12_c174 bl_174 br_174 wl_12 vdd gnd cell_6t
Xbit_r13_c174 bl_174 br_174 wl_13 vdd gnd cell_6t
Xbit_r14_c174 bl_174 br_174 wl_14 vdd gnd cell_6t
Xbit_r15_c174 bl_174 br_174 wl_15 vdd gnd cell_6t
Xbit_r16_c174 bl_174 br_174 wl_16 vdd gnd cell_6t
Xbit_r17_c174 bl_174 br_174 wl_17 vdd gnd cell_6t
Xbit_r18_c174 bl_174 br_174 wl_18 vdd gnd cell_6t
Xbit_r19_c174 bl_174 br_174 wl_19 vdd gnd cell_6t
Xbit_r20_c174 bl_174 br_174 wl_20 vdd gnd cell_6t
Xbit_r21_c174 bl_174 br_174 wl_21 vdd gnd cell_6t
Xbit_r22_c174 bl_174 br_174 wl_22 vdd gnd cell_6t
Xbit_r23_c174 bl_174 br_174 wl_23 vdd gnd cell_6t
Xbit_r24_c174 bl_174 br_174 wl_24 vdd gnd cell_6t
Xbit_r25_c174 bl_174 br_174 wl_25 vdd gnd cell_6t
Xbit_r26_c174 bl_174 br_174 wl_26 vdd gnd cell_6t
Xbit_r27_c174 bl_174 br_174 wl_27 vdd gnd cell_6t
Xbit_r28_c174 bl_174 br_174 wl_28 vdd gnd cell_6t
Xbit_r29_c174 bl_174 br_174 wl_29 vdd gnd cell_6t
Xbit_r30_c174 bl_174 br_174 wl_30 vdd gnd cell_6t
Xbit_r31_c174 bl_174 br_174 wl_31 vdd gnd cell_6t
Xbit_r32_c174 bl_174 br_174 wl_32 vdd gnd cell_6t
Xbit_r33_c174 bl_174 br_174 wl_33 vdd gnd cell_6t
Xbit_r34_c174 bl_174 br_174 wl_34 vdd gnd cell_6t
Xbit_r35_c174 bl_174 br_174 wl_35 vdd gnd cell_6t
Xbit_r36_c174 bl_174 br_174 wl_36 vdd gnd cell_6t
Xbit_r37_c174 bl_174 br_174 wl_37 vdd gnd cell_6t
Xbit_r38_c174 bl_174 br_174 wl_38 vdd gnd cell_6t
Xbit_r39_c174 bl_174 br_174 wl_39 vdd gnd cell_6t
Xbit_r40_c174 bl_174 br_174 wl_40 vdd gnd cell_6t
Xbit_r41_c174 bl_174 br_174 wl_41 vdd gnd cell_6t
Xbit_r42_c174 bl_174 br_174 wl_42 vdd gnd cell_6t
Xbit_r43_c174 bl_174 br_174 wl_43 vdd gnd cell_6t
Xbit_r44_c174 bl_174 br_174 wl_44 vdd gnd cell_6t
Xbit_r45_c174 bl_174 br_174 wl_45 vdd gnd cell_6t
Xbit_r46_c174 bl_174 br_174 wl_46 vdd gnd cell_6t
Xbit_r47_c174 bl_174 br_174 wl_47 vdd gnd cell_6t
Xbit_r48_c174 bl_174 br_174 wl_48 vdd gnd cell_6t
Xbit_r49_c174 bl_174 br_174 wl_49 vdd gnd cell_6t
Xbit_r50_c174 bl_174 br_174 wl_50 vdd gnd cell_6t
Xbit_r51_c174 bl_174 br_174 wl_51 vdd gnd cell_6t
Xbit_r52_c174 bl_174 br_174 wl_52 vdd gnd cell_6t
Xbit_r53_c174 bl_174 br_174 wl_53 vdd gnd cell_6t
Xbit_r54_c174 bl_174 br_174 wl_54 vdd gnd cell_6t
Xbit_r55_c174 bl_174 br_174 wl_55 vdd gnd cell_6t
Xbit_r56_c174 bl_174 br_174 wl_56 vdd gnd cell_6t
Xbit_r57_c174 bl_174 br_174 wl_57 vdd gnd cell_6t
Xbit_r58_c174 bl_174 br_174 wl_58 vdd gnd cell_6t
Xbit_r59_c174 bl_174 br_174 wl_59 vdd gnd cell_6t
Xbit_r60_c174 bl_174 br_174 wl_60 vdd gnd cell_6t
Xbit_r61_c174 bl_174 br_174 wl_61 vdd gnd cell_6t
Xbit_r62_c174 bl_174 br_174 wl_62 vdd gnd cell_6t
Xbit_r63_c174 bl_174 br_174 wl_63 vdd gnd cell_6t
Xbit_r64_c174 bl_174 br_174 wl_64 vdd gnd cell_6t
Xbit_r65_c174 bl_174 br_174 wl_65 vdd gnd cell_6t
Xbit_r66_c174 bl_174 br_174 wl_66 vdd gnd cell_6t
Xbit_r67_c174 bl_174 br_174 wl_67 vdd gnd cell_6t
Xbit_r68_c174 bl_174 br_174 wl_68 vdd gnd cell_6t
Xbit_r69_c174 bl_174 br_174 wl_69 vdd gnd cell_6t
Xbit_r70_c174 bl_174 br_174 wl_70 vdd gnd cell_6t
Xbit_r71_c174 bl_174 br_174 wl_71 vdd gnd cell_6t
Xbit_r72_c174 bl_174 br_174 wl_72 vdd gnd cell_6t
Xbit_r73_c174 bl_174 br_174 wl_73 vdd gnd cell_6t
Xbit_r74_c174 bl_174 br_174 wl_74 vdd gnd cell_6t
Xbit_r75_c174 bl_174 br_174 wl_75 vdd gnd cell_6t
Xbit_r76_c174 bl_174 br_174 wl_76 vdd gnd cell_6t
Xbit_r77_c174 bl_174 br_174 wl_77 vdd gnd cell_6t
Xbit_r78_c174 bl_174 br_174 wl_78 vdd gnd cell_6t
Xbit_r79_c174 bl_174 br_174 wl_79 vdd gnd cell_6t
Xbit_r80_c174 bl_174 br_174 wl_80 vdd gnd cell_6t
Xbit_r81_c174 bl_174 br_174 wl_81 vdd gnd cell_6t
Xbit_r82_c174 bl_174 br_174 wl_82 vdd gnd cell_6t
Xbit_r83_c174 bl_174 br_174 wl_83 vdd gnd cell_6t
Xbit_r84_c174 bl_174 br_174 wl_84 vdd gnd cell_6t
Xbit_r85_c174 bl_174 br_174 wl_85 vdd gnd cell_6t
Xbit_r86_c174 bl_174 br_174 wl_86 vdd gnd cell_6t
Xbit_r87_c174 bl_174 br_174 wl_87 vdd gnd cell_6t
Xbit_r88_c174 bl_174 br_174 wl_88 vdd gnd cell_6t
Xbit_r89_c174 bl_174 br_174 wl_89 vdd gnd cell_6t
Xbit_r90_c174 bl_174 br_174 wl_90 vdd gnd cell_6t
Xbit_r91_c174 bl_174 br_174 wl_91 vdd gnd cell_6t
Xbit_r92_c174 bl_174 br_174 wl_92 vdd gnd cell_6t
Xbit_r93_c174 bl_174 br_174 wl_93 vdd gnd cell_6t
Xbit_r94_c174 bl_174 br_174 wl_94 vdd gnd cell_6t
Xbit_r95_c174 bl_174 br_174 wl_95 vdd gnd cell_6t
Xbit_r96_c174 bl_174 br_174 wl_96 vdd gnd cell_6t
Xbit_r97_c174 bl_174 br_174 wl_97 vdd gnd cell_6t
Xbit_r98_c174 bl_174 br_174 wl_98 vdd gnd cell_6t
Xbit_r99_c174 bl_174 br_174 wl_99 vdd gnd cell_6t
Xbit_r100_c174 bl_174 br_174 wl_100 vdd gnd cell_6t
Xbit_r101_c174 bl_174 br_174 wl_101 vdd gnd cell_6t
Xbit_r102_c174 bl_174 br_174 wl_102 vdd gnd cell_6t
Xbit_r103_c174 bl_174 br_174 wl_103 vdd gnd cell_6t
Xbit_r104_c174 bl_174 br_174 wl_104 vdd gnd cell_6t
Xbit_r105_c174 bl_174 br_174 wl_105 vdd gnd cell_6t
Xbit_r106_c174 bl_174 br_174 wl_106 vdd gnd cell_6t
Xbit_r107_c174 bl_174 br_174 wl_107 vdd gnd cell_6t
Xbit_r108_c174 bl_174 br_174 wl_108 vdd gnd cell_6t
Xbit_r109_c174 bl_174 br_174 wl_109 vdd gnd cell_6t
Xbit_r110_c174 bl_174 br_174 wl_110 vdd gnd cell_6t
Xbit_r111_c174 bl_174 br_174 wl_111 vdd gnd cell_6t
Xbit_r112_c174 bl_174 br_174 wl_112 vdd gnd cell_6t
Xbit_r113_c174 bl_174 br_174 wl_113 vdd gnd cell_6t
Xbit_r114_c174 bl_174 br_174 wl_114 vdd gnd cell_6t
Xbit_r115_c174 bl_174 br_174 wl_115 vdd gnd cell_6t
Xbit_r116_c174 bl_174 br_174 wl_116 vdd gnd cell_6t
Xbit_r117_c174 bl_174 br_174 wl_117 vdd gnd cell_6t
Xbit_r118_c174 bl_174 br_174 wl_118 vdd gnd cell_6t
Xbit_r119_c174 bl_174 br_174 wl_119 vdd gnd cell_6t
Xbit_r120_c174 bl_174 br_174 wl_120 vdd gnd cell_6t
Xbit_r121_c174 bl_174 br_174 wl_121 vdd gnd cell_6t
Xbit_r122_c174 bl_174 br_174 wl_122 vdd gnd cell_6t
Xbit_r123_c174 bl_174 br_174 wl_123 vdd gnd cell_6t
Xbit_r124_c174 bl_174 br_174 wl_124 vdd gnd cell_6t
Xbit_r125_c174 bl_174 br_174 wl_125 vdd gnd cell_6t
Xbit_r126_c174 bl_174 br_174 wl_126 vdd gnd cell_6t
Xbit_r127_c174 bl_174 br_174 wl_127 vdd gnd cell_6t
Xbit_r128_c174 bl_174 br_174 wl_128 vdd gnd cell_6t
Xbit_r129_c174 bl_174 br_174 wl_129 vdd gnd cell_6t
Xbit_r130_c174 bl_174 br_174 wl_130 vdd gnd cell_6t
Xbit_r131_c174 bl_174 br_174 wl_131 vdd gnd cell_6t
Xbit_r132_c174 bl_174 br_174 wl_132 vdd gnd cell_6t
Xbit_r133_c174 bl_174 br_174 wl_133 vdd gnd cell_6t
Xbit_r134_c174 bl_174 br_174 wl_134 vdd gnd cell_6t
Xbit_r135_c174 bl_174 br_174 wl_135 vdd gnd cell_6t
Xbit_r136_c174 bl_174 br_174 wl_136 vdd gnd cell_6t
Xbit_r137_c174 bl_174 br_174 wl_137 vdd gnd cell_6t
Xbit_r138_c174 bl_174 br_174 wl_138 vdd gnd cell_6t
Xbit_r139_c174 bl_174 br_174 wl_139 vdd gnd cell_6t
Xbit_r140_c174 bl_174 br_174 wl_140 vdd gnd cell_6t
Xbit_r141_c174 bl_174 br_174 wl_141 vdd gnd cell_6t
Xbit_r142_c174 bl_174 br_174 wl_142 vdd gnd cell_6t
Xbit_r143_c174 bl_174 br_174 wl_143 vdd gnd cell_6t
Xbit_r144_c174 bl_174 br_174 wl_144 vdd gnd cell_6t
Xbit_r145_c174 bl_174 br_174 wl_145 vdd gnd cell_6t
Xbit_r146_c174 bl_174 br_174 wl_146 vdd gnd cell_6t
Xbit_r147_c174 bl_174 br_174 wl_147 vdd gnd cell_6t
Xbit_r148_c174 bl_174 br_174 wl_148 vdd gnd cell_6t
Xbit_r149_c174 bl_174 br_174 wl_149 vdd gnd cell_6t
Xbit_r150_c174 bl_174 br_174 wl_150 vdd gnd cell_6t
Xbit_r151_c174 bl_174 br_174 wl_151 vdd gnd cell_6t
Xbit_r152_c174 bl_174 br_174 wl_152 vdd gnd cell_6t
Xbit_r153_c174 bl_174 br_174 wl_153 vdd gnd cell_6t
Xbit_r154_c174 bl_174 br_174 wl_154 vdd gnd cell_6t
Xbit_r155_c174 bl_174 br_174 wl_155 vdd gnd cell_6t
Xbit_r156_c174 bl_174 br_174 wl_156 vdd gnd cell_6t
Xbit_r157_c174 bl_174 br_174 wl_157 vdd gnd cell_6t
Xbit_r158_c174 bl_174 br_174 wl_158 vdd gnd cell_6t
Xbit_r159_c174 bl_174 br_174 wl_159 vdd gnd cell_6t
Xbit_r160_c174 bl_174 br_174 wl_160 vdd gnd cell_6t
Xbit_r161_c174 bl_174 br_174 wl_161 vdd gnd cell_6t
Xbit_r162_c174 bl_174 br_174 wl_162 vdd gnd cell_6t
Xbit_r163_c174 bl_174 br_174 wl_163 vdd gnd cell_6t
Xbit_r164_c174 bl_174 br_174 wl_164 vdd gnd cell_6t
Xbit_r165_c174 bl_174 br_174 wl_165 vdd gnd cell_6t
Xbit_r166_c174 bl_174 br_174 wl_166 vdd gnd cell_6t
Xbit_r167_c174 bl_174 br_174 wl_167 vdd gnd cell_6t
Xbit_r168_c174 bl_174 br_174 wl_168 vdd gnd cell_6t
Xbit_r169_c174 bl_174 br_174 wl_169 vdd gnd cell_6t
Xbit_r170_c174 bl_174 br_174 wl_170 vdd gnd cell_6t
Xbit_r171_c174 bl_174 br_174 wl_171 vdd gnd cell_6t
Xbit_r172_c174 bl_174 br_174 wl_172 vdd gnd cell_6t
Xbit_r173_c174 bl_174 br_174 wl_173 vdd gnd cell_6t
Xbit_r174_c174 bl_174 br_174 wl_174 vdd gnd cell_6t
Xbit_r175_c174 bl_174 br_174 wl_175 vdd gnd cell_6t
Xbit_r176_c174 bl_174 br_174 wl_176 vdd gnd cell_6t
Xbit_r177_c174 bl_174 br_174 wl_177 vdd gnd cell_6t
Xbit_r178_c174 bl_174 br_174 wl_178 vdd gnd cell_6t
Xbit_r179_c174 bl_174 br_174 wl_179 vdd gnd cell_6t
Xbit_r180_c174 bl_174 br_174 wl_180 vdd gnd cell_6t
Xbit_r181_c174 bl_174 br_174 wl_181 vdd gnd cell_6t
Xbit_r182_c174 bl_174 br_174 wl_182 vdd gnd cell_6t
Xbit_r183_c174 bl_174 br_174 wl_183 vdd gnd cell_6t
Xbit_r184_c174 bl_174 br_174 wl_184 vdd gnd cell_6t
Xbit_r185_c174 bl_174 br_174 wl_185 vdd gnd cell_6t
Xbit_r186_c174 bl_174 br_174 wl_186 vdd gnd cell_6t
Xbit_r187_c174 bl_174 br_174 wl_187 vdd gnd cell_6t
Xbit_r188_c174 bl_174 br_174 wl_188 vdd gnd cell_6t
Xbit_r189_c174 bl_174 br_174 wl_189 vdd gnd cell_6t
Xbit_r190_c174 bl_174 br_174 wl_190 vdd gnd cell_6t
Xbit_r191_c174 bl_174 br_174 wl_191 vdd gnd cell_6t
Xbit_r192_c174 bl_174 br_174 wl_192 vdd gnd cell_6t
Xbit_r193_c174 bl_174 br_174 wl_193 vdd gnd cell_6t
Xbit_r194_c174 bl_174 br_174 wl_194 vdd gnd cell_6t
Xbit_r195_c174 bl_174 br_174 wl_195 vdd gnd cell_6t
Xbit_r196_c174 bl_174 br_174 wl_196 vdd gnd cell_6t
Xbit_r197_c174 bl_174 br_174 wl_197 vdd gnd cell_6t
Xbit_r198_c174 bl_174 br_174 wl_198 vdd gnd cell_6t
Xbit_r199_c174 bl_174 br_174 wl_199 vdd gnd cell_6t
Xbit_r200_c174 bl_174 br_174 wl_200 vdd gnd cell_6t
Xbit_r201_c174 bl_174 br_174 wl_201 vdd gnd cell_6t
Xbit_r202_c174 bl_174 br_174 wl_202 vdd gnd cell_6t
Xbit_r203_c174 bl_174 br_174 wl_203 vdd gnd cell_6t
Xbit_r204_c174 bl_174 br_174 wl_204 vdd gnd cell_6t
Xbit_r205_c174 bl_174 br_174 wl_205 vdd gnd cell_6t
Xbit_r206_c174 bl_174 br_174 wl_206 vdd gnd cell_6t
Xbit_r207_c174 bl_174 br_174 wl_207 vdd gnd cell_6t
Xbit_r208_c174 bl_174 br_174 wl_208 vdd gnd cell_6t
Xbit_r209_c174 bl_174 br_174 wl_209 vdd gnd cell_6t
Xbit_r210_c174 bl_174 br_174 wl_210 vdd gnd cell_6t
Xbit_r211_c174 bl_174 br_174 wl_211 vdd gnd cell_6t
Xbit_r212_c174 bl_174 br_174 wl_212 vdd gnd cell_6t
Xbit_r213_c174 bl_174 br_174 wl_213 vdd gnd cell_6t
Xbit_r214_c174 bl_174 br_174 wl_214 vdd gnd cell_6t
Xbit_r215_c174 bl_174 br_174 wl_215 vdd gnd cell_6t
Xbit_r216_c174 bl_174 br_174 wl_216 vdd gnd cell_6t
Xbit_r217_c174 bl_174 br_174 wl_217 vdd gnd cell_6t
Xbit_r218_c174 bl_174 br_174 wl_218 vdd gnd cell_6t
Xbit_r219_c174 bl_174 br_174 wl_219 vdd gnd cell_6t
Xbit_r220_c174 bl_174 br_174 wl_220 vdd gnd cell_6t
Xbit_r221_c174 bl_174 br_174 wl_221 vdd gnd cell_6t
Xbit_r222_c174 bl_174 br_174 wl_222 vdd gnd cell_6t
Xbit_r223_c174 bl_174 br_174 wl_223 vdd gnd cell_6t
Xbit_r224_c174 bl_174 br_174 wl_224 vdd gnd cell_6t
Xbit_r225_c174 bl_174 br_174 wl_225 vdd gnd cell_6t
Xbit_r226_c174 bl_174 br_174 wl_226 vdd gnd cell_6t
Xbit_r227_c174 bl_174 br_174 wl_227 vdd gnd cell_6t
Xbit_r228_c174 bl_174 br_174 wl_228 vdd gnd cell_6t
Xbit_r229_c174 bl_174 br_174 wl_229 vdd gnd cell_6t
Xbit_r230_c174 bl_174 br_174 wl_230 vdd gnd cell_6t
Xbit_r231_c174 bl_174 br_174 wl_231 vdd gnd cell_6t
Xbit_r232_c174 bl_174 br_174 wl_232 vdd gnd cell_6t
Xbit_r233_c174 bl_174 br_174 wl_233 vdd gnd cell_6t
Xbit_r234_c174 bl_174 br_174 wl_234 vdd gnd cell_6t
Xbit_r235_c174 bl_174 br_174 wl_235 vdd gnd cell_6t
Xbit_r236_c174 bl_174 br_174 wl_236 vdd gnd cell_6t
Xbit_r237_c174 bl_174 br_174 wl_237 vdd gnd cell_6t
Xbit_r238_c174 bl_174 br_174 wl_238 vdd gnd cell_6t
Xbit_r239_c174 bl_174 br_174 wl_239 vdd gnd cell_6t
Xbit_r240_c174 bl_174 br_174 wl_240 vdd gnd cell_6t
Xbit_r241_c174 bl_174 br_174 wl_241 vdd gnd cell_6t
Xbit_r242_c174 bl_174 br_174 wl_242 vdd gnd cell_6t
Xbit_r243_c174 bl_174 br_174 wl_243 vdd gnd cell_6t
Xbit_r244_c174 bl_174 br_174 wl_244 vdd gnd cell_6t
Xbit_r245_c174 bl_174 br_174 wl_245 vdd gnd cell_6t
Xbit_r246_c174 bl_174 br_174 wl_246 vdd gnd cell_6t
Xbit_r247_c174 bl_174 br_174 wl_247 vdd gnd cell_6t
Xbit_r248_c174 bl_174 br_174 wl_248 vdd gnd cell_6t
Xbit_r249_c174 bl_174 br_174 wl_249 vdd gnd cell_6t
Xbit_r250_c174 bl_174 br_174 wl_250 vdd gnd cell_6t
Xbit_r251_c174 bl_174 br_174 wl_251 vdd gnd cell_6t
Xbit_r252_c174 bl_174 br_174 wl_252 vdd gnd cell_6t
Xbit_r253_c174 bl_174 br_174 wl_253 vdd gnd cell_6t
Xbit_r254_c174 bl_174 br_174 wl_254 vdd gnd cell_6t
Xbit_r255_c174 bl_174 br_174 wl_255 vdd gnd cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd cell_6t
Xbit_r1_c175 bl_175 br_175 wl_1 vdd gnd cell_6t
Xbit_r2_c175 bl_175 br_175 wl_2 vdd gnd cell_6t
Xbit_r3_c175 bl_175 br_175 wl_3 vdd gnd cell_6t
Xbit_r4_c175 bl_175 br_175 wl_4 vdd gnd cell_6t
Xbit_r5_c175 bl_175 br_175 wl_5 vdd gnd cell_6t
Xbit_r6_c175 bl_175 br_175 wl_6 vdd gnd cell_6t
Xbit_r7_c175 bl_175 br_175 wl_7 vdd gnd cell_6t
Xbit_r8_c175 bl_175 br_175 wl_8 vdd gnd cell_6t
Xbit_r9_c175 bl_175 br_175 wl_9 vdd gnd cell_6t
Xbit_r10_c175 bl_175 br_175 wl_10 vdd gnd cell_6t
Xbit_r11_c175 bl_175 br_175 wl_11 vdd gnd cell_6t
Xbit_r12_c175 bl_175 br_175 wl_12 vdd gnd cell_6t
Xbit_r13_c175 bl_175 br_175 wl_13 vdd gnd cell_6t
Xbit_r14_c175 bl_175 br_175 wl_14 vdd gnd cell_6t
Xbit_r15_c175 bl_175 br_175 wl_15 vdd gnd cell_6t
Xbit_r16_c175 bl_175 br_175 wl_16 vdd gnd cell_6t
Xbit_r17_c175 bl_175 br_175 wl_17 vdd gnd cell_6t
Xbit_r18_c175 bl_175 br_175 wl_18 vdd gnd cell_6t
Xbit_r19_c175 bl_175 br_175 wl_19 vdd gnd cell_6t
Xbit_r20_c175 bl_175 br_175 wl_20 vdd gnd cell_6t
Xbit_r21_c175 bl_175 br_175 wl_21 vdd gnd cell_6t
Xbit_r22_c175 bl_175 br_175 wl_22 vdd gnd cell_6t
Xbit_r23_c175 bl_175 br_175 wl_23 vdd gnd cell_6t
Xbit_r24_c175 bl_175 br_175 wl_24 vdd gnd cell_6t
Xbit_r25_c175 bl_175 br_175 wl_25 vdd gnd cell_6t
Xbit_r26_c175 bl_175 br_175 wl_26 vdd gnd cell_6t
Xbit_r27_c175 bl_175 br_175 wl_27 vdd gnd cell_6t
Xbit_r28_c175 bl_175 br_175 wl_28 vdd gnd cell_6t
Xbit_r29_c175 bl_175 br_175 wl_29 vdd gnd cell_6t
Xbit_r30_c175 bl_175 br_175 wl_30 vdd gnd cell_6t
Xbit_r31_c175 bl_175 br_175 wl_31 vdd gnd cell_6t
Xbit_r32_c175 bl_175 br_175 wl_32 vdd gnd cell_6t
Xbit_r33_c175 bl_175 br_175 wl_33 vdd gnd cell_6t
Xbit_r34_c175 bl_175 br_175 wl_34 vdd gnd cell_6t
Xbit_r35_c175 bl_175 br_175 wl_35 vdd gnd cell_6t
Xbit_r36_c175 bl_175 br_175 wl_36 vdd gnd cell_6t
Xbit_r37_c175 bl_175 br_175 wl_37 vdd gnd cell_6t
Xbit_r38_c175 bl_175 br_175 wl_38 vdd gnd cell_6t
Xbit_r39_c175 bl_175 br_175 wl_39 vdd gnd cell_6t
Xbit_r40_c175 bl_175 br_175 wl_40 vdd gnd cell_6t
Xbit_r41_c175 bl_175 br_175 wl_41 vdd gnd cell_6t
Xbit_r42_c175 bl_175 br_175 wl_42 vdd gnd cell_6t
Xbit_r43_c175 bl_175 br_175 wl_43 vdd gnd cell_6t
Xbit_r44_c175 bl_175 br_175 wl_44 vdd gnd cell_6t
Xbit_r45_c175 bl_175 br_175 wl_45 vdd gnd cell_6t
Xbit_r46_c175 bl_175 br_175 wl_46 vdd gnd cell_6t
Xbit_r47_c175 bl_175 br_175 wl_47 vdd gnd cell_6t
Xbit_r48_c175 bl_175 br_175 wl_48 vdd gnd cell_6t
Xbit_r49_c175 bl_175 br_175 wl_49 vdd gnd cell_6t
Xbit_r50_c175 bl_175 br_175 wl_50 vdd gnd cell_6t
Xbit_r51_c175 bl_175 br_175 wl_51 vdd gnd cell_6t
Xbit_r52_c175 bl_175 br_175 wl_52 vdd gnd cell_6t
Xbit_r53_c175 bl_175 br_175 wl_53 vdd gnd cell_6t
Xbit_r54_c175 bl_175 br_175 wl_54 vdd gnd cell_6t
Xbit_r55_c175 bl_175 br_175 wl_55 vdd gnd cell_6t
Xbit_r56_c175 bl_175 br_175 wl_56 vdd gnd cell_6t
Xbit_r57_c175 bl_175 br_175 wl_57 vdd gnd cell_6t
Xbit_r58_c175 bl_175 br_175 wl_58 vdd gnd cell_6t
Xbit_r59_c175 bl_175 br_175 wl_59 vdd gnd cell_6t
Xbit_r60_c175 bl_175 br_175 wl_60 vdd gnd cell_6t
Xbit_r61_c175 bl_175 br_175 wl_61 vdd gnd cell_6t
Xbit_r62_c175 bl_175 br_175 wl_62 vdd gnd cell_6t
Xbit_r63_c175 bl_175 br_175 wl_63 vdd gnd cell_6t
Xbit_r64_c175 bl_175 br_175 wl_64 vdd gnd cell_6t
Xbit_r65_c175 bl_175 br_175 wl_65 vdd gnd cell_6t
Xbit_r66_c175 bl_175 br_175 wl_66 vdd gnd cell_6t
Xbit_r67_c175 bl_175 br_175 wl_67 vdd gnd cell_6t
Xbit_r68_c175 bl_175 br_175 wl_68 vdd gnd cell_6t
Xbit_r69_c175 bl_175 br_175 wl_69 vdd gnd cell_6t
Xbit_r70_c175 bl_175 br_175 wl_70 vdd gnd cell_6t
Xbit_r71_c175 bl_175 br_175 wl_71 vdd gnd cell_6t
Xbit_r72_c175 bl_175 br_175 wl_72 vdd gnd cell_6t
Xbit_r73_c175 bl_175 br_175 wl_73 vdd gnd cell_6t
Xbit_r74_c175 bl_175 br_175 wl_74 vdd gnd cell_6t
Xbit_r75_c175 bl_175 br_175 wl_75 vdd gnd cell_6t
Xbit_r76_c175 bl_175 br_175 wl_76 vdd gnd cell_6t
Xbit_r77_c175 bl_175 br_175 wl_77 vdd gnd cell_6t
Xbit_r78_c175 bl_175 br_175 wl_78 vdd gnd cell_6t
Xbit_r79_c175 bl_175 br_175 wl_79 vdd gnd cell_6t
Xbit_r80_c175 bl_175 br_175 wl_80 vdd gnd cell_6t
Xbit_r81_c175 bl_175 br_175 wl_81 vdd gnd cell_6t
Xbit_r82_c175 bl_175 br_175 wl_82 vdd gnd cell_6t
Xbit_r83_c175 bl_175 br_175 wl_83 vdd gnd cell_6t
Xbit_r84_c175 bl_175 br_175 wl_84 vdd gnd cell_6t
Xbit_r85_c175 bl_175 br_175 wl_85 vdd gnd cell_6t
Xbit_r86_c175 bl_175 br_175 wl_86 vdd gnd cell_6t
Xbit_r87_c175 bl_175 br_175 wl_87 vdd gnd cell_6t
Xbit_r88_c175 bl_175 br_175 wl_88 vdd gnd cell_6t
Xbit_r89_c175 bl_175 br_175 wl_89 vdd gnd cell_6t
Xbit_r90_c175 bl_175 br_175 wl_90 vdd gnd cell_6t
Xbit_r91_c175 bl_175 br_175 wl_91 vdd gnd cell_6t
Xbit_r92_c175 bl_175 br_175 wl_92 vdd gnd cell_6t
Xbit_r93_c175 bl_175 br_175 wl_93 vdd gnd cell_6t
Xbit_r94_c175 bl_175 br_175 wl_94 vdd gnd cell_6t
Xbit_r95_c175 bl_175 br_175 wl_95 vdd gnd cell_6t
Xbit_r96_c175 bl_175 br_175 wl_96 vdd gnd cell_6t
Xbit_r97_c175 bl_175 br_175 wl_97 vdd gnd cell_6t
Xbit_r98_c175 bl_175 br_175 wl_98 vdd gnd cell_6t
Xbit_r99_c175 bl_175 br_175 wl_99 vdd gnd cell_6t
Xbit_r100_c175 bl_175 br_175 wl_100 vdd gnd cell_6t
Xbit_r101_c175 bl_175 br_175 wl_101 vdd gnd cell_6t
Xbit_r102_c175 bl_175 br_175 wl_102 vdd gnd cell_6t
Xbit_r103_c175 bl_175 br_175 wl_103 vdd gnd cell_6t
Xbit_r104_c175 bl_175 br_175 wl_104 vdd gnd cell_6t
Xbit_r105_c175 bl_175 br_175 wl_105 vdd gnd cell_6t
Xbit_r106_c175 bl_175 br_175 wl_106 vdd gnd cell_6t
Xbit_r107_c175 bl_175 br_175 wl_107 vdd gnd cell_6t
Xbit_r108_c175 bl_175 br_175 wl_108 vdd gnd cell_6t
Xbit_r109_c175 bl_175 br_175 wl_109 vdd gnd cell_6t
Xbit_r110_c175 bl_175 br_175 wl_110 vdd gnd cell_6t
Xbit_r111_c175 bl_175 br_175 wl_111 vdd gnd cell_6t
Xbit_r112_c175 bl_175 br_175 wl_112 vdd gnd cell_6t
Xbit_r113_c175 bl_175 br_175 wl_113 vdd gnd cell_6t
Xbit_r114_c175 bl_175 br_175 wl_114 vdd gnd cell_6t
Xbit_r115_c175 bl_175 br_175 wl_115 vdd gnd cell_6t
Xbit_r116_c175 bl_175 br_175 wl_116 vdd gnd cell_6t
Xbit_r117_c175 bl_175 br_175 wl_117 vdd gnd cell_6t
Xbit_r118_c175 bl_175 br_175 wl_118 vdd gnd cell_6t
Xbit_r119_c175 bl_175 br_175 wl_119 vdd gnd cell_6t
Xbit_r120_c175 bl_175 br_175 wl_120 vdd gnd cell_6t
Xbit_r121_c175 bl_175 br_175 wl_121 vdd gnd cell_6t
Xbit_r122_c175 bl_175 br_175 wl_122 vdd gnd cell_6t
Xbit_r123_c175 bl_175 br_175 wl_123 vdd gnd cell_6t
Xbit_r124_c175 bl_175 br_175 wl_124 vdd gnd cell_6t
Xbit_r125_c175 bl_175 br_175 wl_125 vdd gnd cell_6t
Xbit_r126_c175 bl_175 br_175 wl_126 vdd gnd cell_6t
Xbit_r127_c175 bl_175 br_175 wl_127 vdd gnd cell_6t
Xbit_r128_c175 bl_175 br_175 wl_128 vdd gnd cell_6t
Xbit_r129_c175 bl_175 br_175 wl_129 vdd gnd cell_6t
Xbit_r130_c175 bl_175 br_175 wl_130 vdd gnd cell_6t
Xbit_r131_c175 bl_175 br_175 wl_131 vdd gnd cell_6t
Xbit_r132_c175 bl_175 br_175 wl_132 vdd gnd cell_6t
Xbit_r133_c175 bl_175 br_175 wl_133 vdd gnd cell_6t
Xbit_r134_c175 bl_175 br_175 wl_134 vdd gnd cell_6t
Xbit_r135_c175 bl_175 br_175 wl_135 vdd gnd cell_6t
Xbit_r136_c175 bl_175 br_175 wl_136 vdd gnd cell_6t
Xbit_r137_c175 bl_175 br_175 wl_137 vdd gnd cell_6t
Xbit_r138_c175 bl_175 br_175 wl_138 vdd gnd cell_6t
Xbit_r139_c175 bl_175 br_175 wl_139 vdd gnd cell_6t
Xbit_r140_c175 bl_175 br_175 wl_140 vdd gnd cell_6t
Xbit_r141_c175 bl_175 br_175 wl_141 vdd gnd cell_6t
Xbit_r142_c175 bl_175 br_175 wl_142 vdd gnd cell_6t
Xbit_r143_c175 bl_175 br_175 wl_143 vdd gnd cell_6t
Xbit_r144_c175 bl_175 br_175 wl_144 vdd gnd cell_6t
Xbit_r145_c175 bl_175 br_175 wl_145 vdd gnd cell_6t
Xbit_r146_c175 bl_175 br_175 wl_146 vdd gnd cell_6t
Xbit_r147_c175 bl_175 br_175 wl_147 vdd gnd cell_6t
Xbit_r148_c175 bl_175 br_175 wl_148 vdd gnd cell_6t
Xbit_r149_c175 bl_175 br_175 wl_149 vdd gnd cell_6t
Xbit_r150_c175 bl_175 br_175 wl_150 vdd gnd cell_6t
Xbit_r151_c175 bl_175 br_175 wl_151 vdd gnd cell_6t
Xbit_r152_c175 bl_175 br_175 wl_152 vdd gnd cell_6t
Xbit_r153_c175 bl_175 br_175 wl_153 vdd gnd cell_6t
Xbit_r154_c175 bl_175 br_175 wl_154 vdd gnd cell_6t
Xbit_r155_c175 bl_175 br_175 wl_155 vdd gnd cell_6t
Xbit_r156_c175 bl_175 br_175 wl_156 vdd gnd cell_6t
Xbit_r157_c175 bl_175 br_175 wl_157 vdd gnd cell_6t
Xbit_r158_c175 bl_175 br_175 wl_158 vdd gnd cell_6t
Xbit_r159_c175 bl_175 br_175 wl_159 vdd gnd cell_6t
Xbit_r160_c175 bl_175 br_175 wl_160 vdd gnd cell_6t
Xbit_r161_c175 bl_175 br_175 wl_161 vdd gnd cell_6t
Xbit_r162_c175 bl_175 br_175 wl_162 vdd gnd cell_6t
Xbit_r163_c175 bl_175 br_175 wl_163 vdd gnd cell_6t
Xbit_r164_c175 bl_175 br_175 wl_164 vdd gnd cell_6t
Xbit_r165_c175 bl_175 br_175 wl_165 vdd gnd cell_6t
Xbit_r166_c175 bl_175 br_175 wl_166 vdd gnd cell_6t
Xbit_r167_c175 bl_175 br_175 wl_167 vdd gnd cell_6t
Xbit_r168_c175 bl_175 br_175 wl_168 vdd gnd cell_6t
Xbit_r169_c175 bl_175 br_175 wl_169 vdd gnd cell_6t
Xbit_r170_c175 bl_175 br_175 wl_170 vdd gnd cell_6t
Xbit_r171_c175 bl_175 br_175 wl_171 vdd gnd cell_6t
Xbit_r172_c175 bl_175 br_175 wl_172 vdd gnd cell_6t
Xbit_r173_c175 bl_175 br_175 wl_173 vdd gnd cell_6t
Xbit_r174_c175 bl_175 br_175 wl_174 vdd gnd cell_6t
Xbit_r175_c175 bl_175 br_175 wl_175 vdd gnd cell_6t
Xbit_r176_c175 bl_175 br_175 wl_176 vdd gnd cell_6t
Xbit_r177_c175 bl_175 br_175 wl_177 vdd gnd cell_6t
Xbit_r178_c175 bl_175 br_175 wl_178 vdd gnd cell_6t
Xbit_r179_c175 bl_175 br_175 wl_179 vdd gnd cell_6t
Xbit_r180_c175 bl_175 br_175 wl_180 vdd gnd cell_6t
Xbit_r181_c175 bl_175 br_175 wl_181 vdd gnd cell_6t
Xbit_r182_c175 bl_175 br_175 wl_182 vdd gnd cell_6t
Xbit_r183_c175 bl_175 br_175 wl_183 vdd gnd cell_6t
Xbit_r184_c175 bl_175 br_175 wl_184 vdd gnd cell_6t
Xbit_r185_c175 bl_175 br_175 wl_185 vdd gnd cell_6t
Xbit_r186_c175 bl_175 br_175 wl_186 vdd gnd cell_6t
Xbit_r187_c175 bl_175 br_175 wl_187 vdd gnd cell_6t
Xbit_r188_c175 bl_175 br_175 wl_188 vdd gnd cell_6t
Xbit_r189_c175 bl_175 br_175 wl_189 vdd gnd cell_6t
Xbit_r190_c175 bl_175 br_175 wl_190 vdd gnd cell_6t
Xbit_r191_c175 bl_175 br_175 wl_191 vdd gnd cell_6t
Xbit_r192_c175 bl_175 br_175 wl_192 vdd gnd cell_6t
Xbit_r193_c175 bl_175 br_175 wl_193 vdd gnd cell_6t
Xbit_r194_c175 bl_175 br_175 wl_194 vdd gnd cell_6t
Xbit_r195_c175 bl_175 br_175 wl_195 vdd gnd cell_6t
Xbit_r196_c175 bl_175 br_175 wl_196 vdd gnd cell_6t
Xbit_r197_c175 bl_175 br_175 wl_197 vdd gnd cell_6t
Xbit_r198_c175 bl_175 br_175 wl_198 vdd gnd cell_6t
Xbit_r199_c175 bl_175 br_175 wl_199 vdd gnd cell_6t
Xbit_r200_c175 bl_175 br_175 wl_200 vdd gnd cell_6t
Xbit_r201_c175 bl_175 br_175 wl_201 vdd gnd cell_6t
Xbit_r202_c175 bl_175 br_175 wl_202 vdd gnd cell_6t
Xbit_r203_c175 bl_175 br_175 wl_203 vdd gnd cell_6t
Xbit_r204_c175 bl_175 br_175 wl_204 vdd gnd cell_6t
Xbit_r205_c175 bl_175 br_175 wl_205 vdd gnd cell_6t
Xbit_r206_c175 bl_175 br_175 wl_206 vdd gnd cell_6t
Xbit_r207_c175 bl_175 br_175 wl_207 vdd gnd cell_6t
Xbit_r208_c175 bl_175 br_175 wl_208 vdd gnd cell_6t
Xbit_r209_c175 bl_175 br_175 wl_209 vdd gnd cell_6t
Xbit_r210_c175 bl_175 br_175 wl_210 vdd gnd cell_6t
Xbit_r211_c175 bl_175 br_175 wl_211 vdd gnd cell_6t
Xbit_r212_c175 bl_175 br_175 wl_212 vdd gnd cell_6t
Xbit_r213_c175 bl_175 br_175 wl_213 vdd gnd cell_6t
Xbit_r214_c175 bl_175 br_175 wl_214 vdd gnd cell_6t
Xbit_r215_c175 bl_175 br_175 wl_215 vdd gnd cell_6t
Xbit_r216_c175 bl_175 br_175 wl_216 vdd gnd cell_6t
Xbit_r217_c175 bl_175 br_175 wl_217 vdd gnd cell_6t
Xbit_r218_c175 bl_175 br_175 wl_218 vdd gnd cell_6t
Xbit_r219_c175 bl_175 br_175 wl_219 vdd gnd cell_6t
Xbit_r220_c175 bl_175 br_175 wl_220 vdd gnd cell_6t
Xbit_r221_c175 bl_175 br_175 wl_221 vdd gnd cell_6t
Xbit_r222_c175 bl_175 br_175 wl_222 vdd gnd cell_6t
Xbit_r223_c175 bl_175 br_175 wl_223 vdd gnd cell_6t
Xbit_r224_c175 bl_175 br_175 wl_224 vdd gnd cell_6t
Xbit_r225_c175 bl_175 br_175 wl_225 vdd gnd cell_6t
Xbit_r226_c175 bl_175 br_175 wl_226 vdd gnd cell_6t
Xbit_r227_c175 bl_175 br_175 wl_227 vdd gnd cell_6t
Xbit_r228_c175 bl_175 br_175 wl_228 vdd gnd cell_6t
Xbit_r229_c175 bl_175 br_175 wl_229 vdd gnd cell_6t
Xbit_r230_c175 bl_175 br_175 wl_230 vdd gnd cell_6t
Xbit_r231_c175 bl_175 br_175 wl_231 vdd gnd cell_6t
Xbit_r232_c175 bl_175 br_175 wl_232 vdd gnd cell_6t
Xbit_r233_c175 bl_175 br_175 wl_233 vdd gnd cell_6t
Xbit_r234_c175 bl_175 br_175 wl_234 vdd gnd cell_6t
Xbit_r235_c175 bl_175 br_175 wl_235 vdd gnd cell_6t
Xbit_r236_c175 bl_175 br_175 wl_236 vdd gnd cell_6t
Xbit_r237_c175 bl_175 br_175 wl_237 vdd gnd cell_6t
Xbit_r238_c175 bl_175 br_175 wl_238 vdd gnd cell_6t
Xbit_r239_c175 bl_175 br_175 wl_239 vdd gnd cell_6t
Xbit_r240_c175 bl_175 br_175 wl_240 vdd gnd cell_6t
Xbit_r241_c175 bl_175 br_175 wl_241 vdd gnd cell_6t
Xbit_r242_c175 bl_175 br_175 wl_242 vdd gnd cell_6t
Xbit_r243_c175 bl_175 br_175 wl_243 vdd gnd cell_6t
Xbit_r244_c175 bl_175 br_175 wl_244 vdd gnd cell_6t
Xbit_r245_c175 bl_175 br_175 wl_245 vdd gnd cell_6t
Xbit_r246_c175 bl_175 br_175 wl_246 vdd gnd cell_6t
Xbit_r247_c175 bl_175 br_175 wl_247 vdd gnd cell_6t
Xbit_r248_c175 bl_175 br_175 wl_248 vdd gnd cell_6t
Xbit_r249_c175 bl_175 br_175 wl_249 vdd gnd cell_6t
Xbit_r250_c175 bl_175 br_175 wl_250 vdd gnd cell_6t
Xbit_r251_c175 bl_175 br_175 wl_251 vdd gnd cell_6t
Xbit_r252_c175 bl_175 br_175 wl_252 vdd gnd cell_6t
Xbit_r253_c175 bl_175 br_175 wl_253 vdd gnd cell_6t
Xbit_r254_c175 bl_175 br_175 wl_254 vdd gnd cell_6t
Xbit_r255_c175 bl_175 br_175 wl_255 vdd gnd cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd cell_6t
Xbit_r1_c176 bl_176 br_176 wl_1 vdd gnd cell_6t
Xbit_r2_c176 bl_176 br_176 wl_2 vdd gnd cell_6t
Xbit_r3_c176 bl_176 br_176 wl_3 vdd gnd cell_6t
Xbit_r4_c176 bl_176 br_176 wl_4 vdd gnd cell_6t
Xbit_r5_c176 bl_176 br_176 wl_5 vdd gnd cell_6t
Xbit_r6_c176 bl_176 br_176 wl_6 vdd gnd cell_6t
Xbit_r7_c176 bl_176 br_176 wl_7 vdd gnd cell_6t
Xbit_r8_c176 bl_176 br_176 wl_8 vdd gnd cell_6t
Xbit_r9_c176 bl_176 br_176 wl_9 vdd gnd cell_6t
Xbit_r10_c176 bl_176 br_176 wl_10 vdd gnd cell_6t
Xbit_r11_c176 bl_176 br_176 wl_11 vdd gnd cell_6t
Xbit_r12_c176 bl_176 br_176 wl_12 vdd gnd cell_6t
Xbit_r13_c176 bl_176 br_176 wl_13 vdd gnd cell_6t
Xbit_r14_c176 bl_176 br_176 wl_14 vdd gnd cell_6t
Xbit_r15_c176 bl_176 br_176 wl_15 vdd gnd cell_6t
Xbit_r16_c176 bl_176 br_176 wl_16 vdd gnd cell_6t
Xbit_r17_c176 bl_176 br_176 wl_17 vdd gnd cell_6t
Xbit_r18_c176 bl_176 br_176 wl_18 vdd gnd cell_6t
Xbit_r19_c176 bl_176 br_176 wl_19 vdd gnd cell_6t
Xbit_r20_c176 bl_176 br_176 wl_20 vdd gnd cell_6t
Xbit_r21_c176 bl_176 br_176 wl_21 vdd gnd cell_6t
Xbit_r22_c176 bl_176 br_176 wl_22 vdd gnd cell_6t
Xbit_r23_c176 bl_176 br_176 wl_23 vdd gnd cell_6t
Xbit_r24_c176 bl_176 br_176 wl_24 vdd gnd cell_6t
Xbit_r25_c176 bl_176 br_176 wl_25 vdd gnd cell_6t
Xbit_r26_c176 bl_176 br_176 wl_26 vdd gnd cell_6t
Xbit_r27_c176 bl_176 br_176 wl_27 vdd gnd cell_6t
Xbit_r28_c176 bl_176 br_176 wl_28 vdd gnd cell_6t
Xbit_r29_c176 bl_176 br_176 wl_29 vdd gnd cell_6t
Xbit_r30_c176 bl_176 br_176 wl_30 vdd gnd cell_6t
Xbit_r31_c176 bl_176 br_176 wl_31 vdd gnd cell_6t
Xbit_r32_c176 bl_176 br_176 wl_32 vdd gnd cell_6t
Xbit_r33_c176 bl_176 br_176 wl_33 vdd gnd cell_6t
Xbit_r34_c176 bl_176 br_176 wl_34 vdd gnd cell_6t
Xbit_r35_c176 bl_176 br_176 wl_35 vdd gnd cell_6t
Xbit_r36_c176 bl_176 br_176 wl_36 vdd gnd cell_6t
Xbit_r37_c176 bl_176 br_176 wl_37 vdd gnd cell_6t
Xbit_r38_c176 bl_176 br_176 wl_38 vdd gnd cell_6t
Xbit_r39_c176 bl_176 br_176 wl_39 vdd gnd cell_6t
Xbit_r40_c176 bl_176 br_176 wl_40 vdd gnd cell_6t
Xbit_r41_c176 bl_176 br_176 wl_41 vdd gnd cell_6t
Xbit_r42_c176 bl_176 br_176 wl_42 vdd gnd cell_6t
Xbit_r43_c176 bl_176 br_176 wl_43 vdd gnd cell_6t
Xbit_r44_c176 bl_176 br_176 wl_44 vdd gnd cell_6t
Xbit_r45_c176 bl_176 br_176 wl_45 vdd gnd cell_6t
Xbit_r46_c176 bl_176 br_176 wl_46 vdd gnd cell_6t
Xbit_r47_c176 bl_176 br_176 wl_47 vdd gnd cell_6t
Xbit_r48_c176 bl_176 br_176 wl_48 vdd gnd cell_6t
Xbit_r49_c176 bl_176 br_176 wl_49 vdd gnd cell_6t
Xbit_r50_c176 bl_176 br_176 wl_50 vdd gnd cell_6t
Xbit_r51_c176 bl_176 br_176 wl_51 vdd gnd cell_6t
Xbit_r52_c176 bl_176 br_176 wl_52 vdd gnd cell_6t
Xbit_r53_c176 bl_176 br_176 wl_53 vdd gnd cell_6t
Xbit_r54_c176 bl_176 br_176 wl_54 vdd gnd cell_6t
Xbit_r55_c176 bl_176 br_176 wl_55 vdd gnd cell_6t
Xbit_r56_c176 bl_176 br_176 wl_56 vdd gnd cell_6t
Xbit_r57_c176 bl_176 br_176 wl_57 vdd gnd cell_6t
Xbit_r58_c176 bl_176 br_176 wl_58 vdd gnd cell_6t
Xbit_r59_c176 bl_176 br_176 wl_59 vdd gnd cell_6t
Xbit_r60_c176 bl_176 br_176 wl_60 vdd gnd cell_6t
Xbit_r61_c176 bl_176 br_176 wl_61 vdd gnd cell_6t
Xbit_r62_c176 bl_176 br_176 wl_62 vdd gnd cell_6t
Xbit_r63_c176 bl_176 br_176 wl_63 vdd gnd cell_6t
Xbit_r64_c176 bl_176 br_176 wl_64 vdd gnd cell_6t
Xbit_r65_c176 bl_176 br_176 wl_65 vdd gnd cell_6t
Xbit_r66_c176 bl_176 br_176 wl_66 vdd gnd cell_6t
Xbit_r67_c176 bl_176 br_176 wl_67 vdd gnd cell_6t
Xbit_r68_c176 bl_176 br_176 wl_68 vdd gnd cell_6t
Xbit_r69_c176 bl_176 br_176 wl_69 vdd gnd cell_6t
Xbit_r70_c176 bl_176 br_176 wl_70 vdd gnd cell_6t
Xbit_r71_c176 bl_176 br_176 wl_71 vdd gnd cell_6t
Xbit_r72_c176 bl_176 br_176 wl_72 vdd gnd cell_6t
Xbit_r73_c176 bl_176 br_176 wl_73 vdd gnd cell_6t
Xbit_r74_c176 bl_176 br_176 wl_74 vdd gnd cell_6t
Xbit_r75_c176 bl_176 br_176 wl_75 vdd gnd cell_6t
Xbit_r76_c176 bl_176 br_176 wl_76 vdd gnd cell_6t
Xbit_r77_c176 bl_176 br_176 wl_77 vdd gnd cell_6t
Xbit_r78_c176 bl_176 br_176 wl_78 vdd gnd cell_6t
Xbit_r79_c176 bl_176 br_176 wl_79 vdd gnd cell_6t
Xbit_r80_c176 bl_176 br_176 wl_80 vdd gnd cell_6t
Xbit_r81_c176 bl_176 br_176 wl_81 vdd gnd cell_6t
Xbit_r82_c176 bl_176 br_176 wl_82 vdd gnd cell_6t
Xbit_r83_c176 bl_176 br_176 wl_83 vdd gnd cell_6t
Xbit_r84_c176 bl_176 br_176 wl_84 vdd gnd cell_6t
Xbit_r85_c176 bl_176 br_176 wl_85 vdd gnd cell_6t
Xbit_r86_c176 bl_176 br_176 wl_86 vdd gnd cell_6t
Xbit_r87_c176 bl_176 br_176 wl_87 vdd gnd cell_6t
Xbit_r88_c176 bl_176 br_176 wl_88 vdd gnd cell_6t
Xbit_r89_c176 bl_176 br_176 wl_89 vdd gnd cell_6t
Xbit_r90_c176 bl_176 br_176 wl_90 vdd gnd cell_6t
Xbit_r91_c176 bl_176 br_176 wl_91 vdd gnd cell_6t
Xbit_r92_c176 bl_176 br_176 wl_92 vdd gnd cell_6t
Xbit_r93_c176 bl_176 br_176 wl_93 vdd gnd cell_6t
Xbit_r94_c176 bl_176 br_176 wl_94 vdd gnd cell_6t
Xbit_r95_c176 bl_176 br_176 wl_95 vdd gnd cell_6t
Xbit_r96_c176 bl_176 br_176 wl_96 vdd gnd cell_6t
Xbit_r97_c176 bl_176 br_176 wl_97 vdd gnd cell_6t
Xbit_r98_c176 bl_176 br_176 wl_98 vdd gnd cell_6t
Xbit_r99_c176 bl_176 br_176 wl_99 vdd gnd cell_6t
Xbit_r100_c176 bl_176 br_176 wl_100 vdd gnd cell_6t
Xbit_r101_c176 bl_176 br_176 wl_101 vdd gnd cell_6t
Xbit_r102_c176 bl_176 br_176 wl_102 vdd gnd cell_6t
Xbit_r103_c176 bl_176 br_176 wl_103 vdd gnd cell_6t
Xbit_r104_c176 bl_176 br_176 wl_104 vdd gnd cell_6t
Xbit_r105_c176 bl_176 br_176 wl_105 vdd gnd cell_6t
Xbit_r106_c176 bl_176 br_176 wl_106 vdd gnd cell_6t
Xbit_r107_c176 bl_176 br_176 wl_107 vdd gnd cell_6t
Xbit_r108_c176 bl_176 br_176 wl_108 vdd gnd cell_6t
Xbit_r109_c176 bl_176 br_176 wl_109 vdd gnd cell_6t
Xbit_r110_c176 bl_176 br_176 wl_110 vdd gnd cell_6t
Xbit_r111_c176 bl_176 br_176 wl_111 vdd gnd cell_6t
Xbit_r112_c176 bl_176 br_176 wl_112 vdd gnd cell_6t
Xbit_r113_c176 bl_176 br_176 wl_113 vdd gnd cell_6t
Xbit_r114_c176 bl_176 br_176 wl_114 vdd gnd cell_6t
Xbit_r115_c176 bl_176 br_176 wl_115 vdd gnd cell_6t
Xbit_r116_c176 bl_176 br_176 wl_116 vdd gnd cell_6t
Xbit_r117_c176 bl_176 br_176 wl_117 vdd gnd cell_6t
Xbit_r118_c176 bl_176 br_176 wl_118 vdd gnd cell_6t
Xbit_r119_c176 bl_176 br_176 wl_119 vdd gnd cell_6t
Xbit_r120_c176 bl_176 br_176 wl_120 vdd gnd cell_6t
Xbit_r121_c176 bl_176 br_176 wl_121 vdd gnd cell_6t
Xbit_r122_c176 bl_176 br_176 wl_122 vdd gnd cell_6t
Xbit_r123_c176 bl_176 br_176 wl_123 vdd gnd cell_6t
Xbit_r124_c176 bl_176 br_176 wl_124 vdd gnd cell_6t
Xbit_r125_c176 bl_176 br_176 wl_125 vdd gnd cell_6t
Xbit_r126_c176 bl_176 br_176 wl_126 vdd gnd cell_6t
Xbit_r127_c176 bl_176 br_176 wl_127 vdd gnd cell_6t
Xbit_r128_c176 bl_176 br_176 wl_128 vdd gnd cell_6t
Xbit_r129_c176 bl_176 br_176 wl_129 vdd gnd cell_6t
Xbit_r130_c176 bl_176 br_176 wl_130 vdd gnd cell_6t
Xbit_r131_c176 bl_176 br_176 wl_131 vdd gnd cell_6t
Xbit_r132_c176 bl_176 br_176 wl_132 vdd gnd cell_6t
Xbit_r133_c176 bl_176 br_176 wl_133 vdd gnd cell_6t
Xbit_r134_c176 bl_176 br_176 wl_134 vdd gnd cell_6t
Xbit_r135_c176 bl_176 br_176 wl_135 vdd gnd cell_6t
Xbit_r136_c176 bl_176 br_176 wl_136 vdd gnd cell_6t
Xbit_r137_c176 bl_176 br_176 wl_137 vdd gnd cell_6t
Xbit_r138_c176 bl_176 br_176 wl_138 vdd gnd cell_6t
Xbit_r139_c176 bl_176 br_176 wl_139 vdd gnd cell_6t
Xbit_r140_c176 bl_176 br_176 wl_140 vdd gnd cell_6t
Xbit_r141_c176 bl_176 br_176 wl_141 vdd gnd cell_6t
Xbit_r142_c176 bl_176 br_176 wl_142 vdd gnd cell_6t
Xbit_r143_c176 bl_176 br_176 wl_143 vdd gnd cell_6t
Xbit_r144_c176 bl_176 br_176 wl_144 vdd gnd cell_6t
Xbit_r145_c176 bl_176 br_176 wl_145 vdd gnd cell_6t
Xbit_r146_c176 bl_176 br_176 wl_146 vdd gnd cell_6t
Xbit_r147_c176 bl_176 br_176 wl_147 vdd gnd cell_6t
Xbit_r148_c176 bl_176 br_176 wl_148 vdd gnd cell_6t
Xbit_r149_c176 bl_176 br_176 wl_149 vdd gnd cell_6t
Xbit_r150_c176 bl_176 br_176 wl_150 vdd gnd cell_6t
Xbit_r151_c176 bl_176 br_176 wl_151 vdd gnd cell_6t
Xbit_r152_c176 bl_176 br_176 wl_152 vdd gnd cell_6t
Xbit_r153_c176 bl_176 br_176 wl_153 vdd gnd cell_6t
Xbit_r154_c176 bl_176 br_176 wl_154 vdd gnd cell_6t
Xbit_r155_c176 bl_176 br_176 wl_155 vdd gnd cell_6t
Xbit_r156_c176 bl_176 br_176 wl_156 vdd gnd cell_6t
Xbit_r157_c176 bl_176 br_176 wl_157 vdd gnd cell_6t
Xbit_r158_c176 bl_176 br_176 wl_158 vdd gnd cell_6t
Xbit_r159_c176 bl_176 br_176 wl_159 vdd gnd cell_6t
Xbit_r160_c176 bl_176 br_176 wl_160 vdd gnd cell_6t
Xbit_r161_c176 bl_176 br_176 wl_161 vdd gnd cell_6t
Xbit_r162_c176 bl_176 br_176 wl_162 vdd gnd cell_6t
Xbit_r163_c176 bl_176 br_176 wl_163 vdd gnd cell_6t
Xbit_r164_c176 bl_176 br_176 wl_164 vdd gnd cell_6t
Xbit_r165_c176 bl_176 br_176 wl_165 vdd gnd cell_6t
Xbit_r166_c176 bl_176 br_176 wl_166 vdd gnd cell_6t
Xbit_r167_c176 bl_176 br_176 wl_167 vdd gnd cell_6t
Xbit_r168_c176 bl_176 br_176 wl_168 vdd gnd cell_6t
Xbit_r169_c176 bl_176 br_176 wl_169 vdd gnd cell_6t
Xbit_r170_c176 bl_176 br_176 wl_170 vdd gnd cell_6t
Xbit_r171_c176 bl_176 br_176 wl_171 vdd gnd cell_6t
Xbit_r172_c176 bl_176 br_176 wl_172 vdd gnd cell_6t
Xbit_r173_c176 bl_176 br_176 wl_173 vdd gnd cell_6t
Xbit_r174_c176 bl_176 br_176 wl_174 vdd gnd cell_6t
Xbit_r175_c176 bl_176 br_176 wl_175 vdd gnd cell_6t
Xbit_r176_c176 bl_176 br_176 wl_176 vdd gnd cell_6t
Xbit_r177_c176 bl_176 br_176 wl_177 vdd gnd cell_6t
Xbit_r178_c176 bl_176 br_176 wl_178 vdd gnd cell_6t
Xbit_r179_c176 bl_176 br_176 wl_179 vdd gnd cell_6t
Xbit_r180_c176 bl_176 br_176 wl_180 vdd gnd cell_6t
Xbit_r181_c176 bl_176 br_176 wl_181 vdd gnd cell_6t
Xbit_r182_c176 bl_176 br_176 wl_182 vdd gnd cell_6t
Xbit_r183_c176 bl_176 br_176 wl_183 vdd gnd cell_6t
Xbit_r184_c176 bl_176 br_176 wl_184 vdd gnd cell_6t
Xbit_r185_c176 bl_176 br_176 wl_185 vdd gnd cell_6t
Xbit_r186_c176 bl_176 br_176 wl_186 vdd gnd cell_6t
Xbit_r187_c176 bl_176 br_176 wl_187 vdd gnd cell_6t
Xbit_r188_c176 bl_176 br_176 wl_188 vdd gnd cell_6t
Xbit_r189_c176 bl_176 br_176 wl_189 vdd gnd cell_6t
Xbit_r190_c176 bl_176 br_176 wl_190 vdd gnd cell_6t
Xbit_r191_c176 bl_176 br_176 wl_191 vdd gnd cell_6t
Xbit_r192_c176 bl_176 br_176 wl_192 vdd gnd cell_6t
Xbit_r193_c176 bl_176 br_176 wl_193 vdd gnd cell_6t
Xbit_r194_c176 bl_176 br_176 wl_194 vdd gnd cell_6t
Xbit_r195_c176 bl_176 br_176 wl_195 vdd gnd cell_6t
Xbit_r196_c176 bl_176 br_176 wl_196 vdd gnd cell_6t
Xbit_r197_c176 bl_176 br_176 wl_197 vdd gnd cell_6t
Xbit_r198_c176 bl_176 br_176 wl_198 vdd gnd cell_6t
Xbit_r199_c176 bl_176 br_176 wl_199 vdd gnd cell_6t
Xbit_r200_c176 bl_176 br_176 wl_200 vdd gnd cell_6t
Xbit_r201_c176 bl_176 br_176 wl_201 vdd gnd cell_6t
Xbit_r202_c176 bl_176 br_176 wl_202 vdd gnd cell_6t
Xbit_r203_c176 bl_176 br_176 wl_203 vdd gnd cell_6t
Xbit_r204_c176 bl_176 br_176 wl_204 vdd gnd cell_6t
Xbit_r205_c176 bl_176 br_176 wl_205 vdd gnd cell_6t
Xbit_r206_c176 bl_176 br_176 wl_206 vdd gnd cell_6t
Xbit_r207_c176 bl_176 br_176 wl_207 vdd gnd cell_6t
Xbit_r208_c176 bl_176 br_176 wl_208 vdd gnd cell_6t
Xbit_r209_c176 bl_176 br_176 wl_209 vdd gnd cell_6t
Xbit_r210_c176 bl_176 br_176 wl_210 vdd gnd cell_6t
Xbit_r211_c176 bl_176 br_176 wl_211 vdd gnd cell_6t
Xbit_r212_c176 bl_176 br_176 wl_212 vdd gnd cell_6t
Xbit_r213_c176 bl_176 br_176 wl_213 vdd gnd cell_6t
Xbit_r214_c176 bl_176 br_176 wl_214 vdd gnd cell_6t
Xbit_r215_c176 bl_176 br_176 wl_215 vdd gnd cell_6t
Xbit_r216_c176 bl_176 br_176 wl_216 vdd gnd cell_6t
Xbit_r217_c176 bl_176 br_176 wl_217 vdd gnd cell_6t
Xbit_r218_c176 bl_176 br_176 wl_218 vdd gnd cell_6t
Xbit_r219_c176 bl_176 br_176 wl_219 vdd gnd cell_6t
Xbit_r220_c176 bl_176 br_176 wl_220 vdd gnd cell_6t
Xbit_r221_c176 bl_176 br_176 wl_221 vdd gnd cell_6t
Xbit_r222_c176 bl_176 br_176 wl_222 vdd gnd cell_6t
Xbit_r223_c176 bl_176 br_176 wl_223 vdd gnd cell_6t
Xbit_r224_c176 bl_176 br_176 wl_224 vdd gnd cell_6t
Xbit_r225_c176 bl_176 br_176 wl_225 vdd gnd cell_6t
Xbit_r226_c176 bl_176 br_176 wl_226 vdd gnd cell_6t
Xbit_r227_c176 bl_176 br_176 wl_227 vdd gnd cell_6t
Xbit_r228_c176 bl_176 br_176 wl_228 vdd gnd cell_6t
Xbit_r229_c176 bl_176 br_176 wl_229 vdd gnd cell_6t
Xbit_r230_c176 bl_176 br_176 wl_230 vdd gnd cell_6t
Xbit_r231_c176 bl_176 br_176 wl_231 vdd gnd cell_6t
Xbit_r232_c176 bl_176 br_176 wl_232 vdd gnd cell_6t
Xbit_r233_c176 bl_176 br_176 wl_233 vdd gnd cell_6t
Xbit_r234_c176 bl_176 br_176 wl_234 vdd gnd cell_6t
Xbit_r235_c176 bl_176 br_176 wl_235 vdd gnd cell_6t
Xbit_r236_c176 bl_176 br_176 wl_236 vdd gnd cell_6t
Xbit_r237_c176 bl_176 br_176 wl_237 vdd gnd cell_6t
Xbit_r238_c176 bl_176 br_176 wl_238 vdd gnd cell_6t
Xbit_r239_c176 bl_176 br_176 wl_239 vdd gnd cell_6t
Xbit_r240_c176 bl_176 br_176 wl_240 vdd gnd cell_6t
Xbit_r241_c176 bl_176 br_176 wl_241 vdd gnd cell_6t
Xbit_r242_c176 bl_176 br_176 wl_242 vdd gnd cell_6t
Xbit_r243_c176 bl_176 br_176 wl_243 vdd gnd cell_6t
Xbit_r244_c176 bl_176 br_176 wl_244 vdd gnd cell_6t
Xbit_r245_c176 bl_176 br_176 wl_245 vdd gnd cell_6t
Xbit_r246_c176 bl_176 br_176 wl_246 vdd gnd cell_6t
Xbit_r247_c176 bl_176 br_176 wl_247 vdd gnd cell_6t
Xbit_r248_c176 bl_176 br_176 wl_248 vdd gnd cell_6t
Xbit_r249_c176 bl_176 br_176 wl_249 vdd gnd cell_6t
Xbit_r250_c176 bl_176 br_176 wl_250 vdd gnd cell_6t
Xbit_r251_c176 bl_176 br_176 wl_251 vdd gnd cell_6t
Xbit_r252_c176 bl_176 br_176 wl_252 vdd gnd cell_6t
Xbit_r253_c176 bl_176 br_176 wl_253 vdd gnd cell_6t
Xbit_r254_c176 bl_176 br_176 wl_254 vdd gnd cell_6t
Xbit_r255_c176 bl_176 br_176 wl_255 vdd gnd cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd cell_6t
Xbit_r1_c177 bl_177 br_177 wl_1 vdd gnd cell_6t
Xbit_r2_c177 bl_177 br_177 wl_2 vdd gnd cell_6t
Xbit_r3_c177 bl_177 br_177 wl_3 vdd gnd cell_6t
Xbit_r4_c177 bl_177 br_177 wl_4 vdd gnd cell_6t
Xbit_r5_c177 bl_177 br_177 wl_5 vdd gnd cell_6t
Xbit_r6_c177 bl_177 br_177 wl_6 vdd gnd cell_6t
Xbit_r7_c177 bl_177 br_177 wl_7 vdd gnd cell_6t
Xbit_r8_c177 bl_177 br_177 wl_8 vdd gnd cell_6t
Xbit_r9_c177 bl_177 br_177 wl_9 vdd gnd cell_6t
Xbit_r10_c177 bl_177 br_177 wl_10 vdd gnd cell_6t
Xbit_r11_c177 bl_177 br_177 wl_11 vdd gnd cell_6t
Xbit_r12_c177 bl_177 br_177 wl_12 vdd gnd cell_6t
Xbit_r13_c177 bl_177 br_177 wl_13 vdd gnd cell_6t
Xbit_r14_c177 bl_177 br_177 wl_14 vdd gnd cell_6t
Xbit_r15_c177 bl_177 br_177 wl_15 vdd gnd cell_6t
Xbit_r16_c177 bl_177 br_177 wl_16 vdd gnd cell_6t
Xbit_r17_c177 bl_177 br_177 wl_17 vdd gnd cell_6t
Xbit_r18_c177 bl_177 br_177 wl_18 vdd gnd cell_6t
Xbit_r19_c177 bl_177 br_177 wl_19 vdd gnd cell_6t
Xbit_r20_c177 bl_177 br_177 wl_20 vdd gnd cell_6t
Xbit_r21_c177 bl_177 br_177 wl_21 vdd gnd cell_6t
Xbit_r22_c177 bl_177 br_177 wl_22 vdd gnd cell_6t
Xbit_r23_c177 bl_177 br_177 wl_23 vdd gnd cell_6t
Xbit_r24_c177 bl_177 br_177 wl_24 vdd gnd cell_6t
Xbit_r25_c177 bl_177 br_177 wl_25 vdd gnd cell_6t
Xbit_r26_c177 bl_177 br_177 wl_26 vdd gnd cell_6t
Xbit_r27_c177 bl_177 br_177 wl_27 vdd gnd cell_6t
Xbit_r28_c177 bl_177 br_177 wl_28 vdd gnd cell_6t
Xbit_r29_c177 bl_177 br_177 wl_29 vdd gnd cell_6t
Xbit_r30_c177 bl_177 br_177 wl_30 vdd gnd cell_6t
Xbit_r31_c177 bl_177 br_177 wl_31 vdd gnd cell_6t
Xbit_r32_c177 bl_177 br_177 wl_32 vdd gnd cell_6t
Xbit_r33_c177 bl_177 br_177 wl_33 vdd gnd cell_6t
Xbit_r34_c177 bl_177 br_177 wl_34 vdd gnd cell_6t
Xbit_r35_c177 bl_177 br_177 wl_35 vdd gnd cell_6t
Xbit_r36_c177 bl_177 br_177 wl_36 vdd gnd cell_6t
Xbit_r37_c177 bl_177 br_177 wl_37 vdd gnd cell_6t
Xbit_r38_c177 bl_177 br_177 wl_38 vdd gnd cell_6t
Xbit_r39_c177 bl_177 br_177 wl_39 vdd gnd cell_6t
Xbit_r40_c177 bl_177 br_177 wl_40 vdd gnd cell_6t
Xbit_r41_c177 bl_177 br_177 wl_41 vdd gnd cell_6t
Xbit_r42_c177 bl_177 br_177 wl_42 vdd gnd cell_6t
Xbit_r43_c177 bl_177 br_177 wl_43 vdd gnd cell_6t
Xbit_r44_c177 bl_177 br_177 wl_44 vdd gnd cell_6t
Xbit_r45_c177 bl_177 br_177 wl_45 vdd gnd cell_6t
Xbit_r46_c177 bl_177 br_177 wl_46 vdd gnd cell_6t
Xbit_r47_c177 bl_177 br_177 wl_47 vdd gnd cell_6t
Xbit_r48_c177 bl_177 br_177 wl_48 vdd gnd cell_6t
Xbit_r49_c177 bl_177 br_177 wl_49 vdd gnd cell_6t
Xbit_r50_c177 bl_177 br_177 wl_50 vdd gnd cell_6t
Xbit_r51_c177 bl_177 br_177 wl_51 vdd gnd cell_6t
Xbit_r52_c177 bl_177 br_177 wl_52 vdd gnd cell_6t
Xbit_r53_c177 bl_177 br_177 wl_53 vdd gnd cell_6t
Xbit_r54_c177 bl_177 br_177 wl_54 vdd gnd cell_6t
Xbit_r55_c177 bl_177 br_177 wl_55 vdd gnd cell_6t
Xbit_r56_c177 bl_177 br_177 wl_56 vdd gnd cell_6t
Xbit_r57_c177 bl_177 br_177 wl_57 vdd gnd cell_6t
Xbit_r58_c177 bl_177 br_177 wl_58 vdd gnd cell_6t
Xbit_r59_c177 bl_177 br_177 wl_59 vdd gnd cell_6t
Xbit_r60_c177 bl_177 br_177 wl_60 vdd gnd cell_6t
Xbit_r61_c177 bl_177 br_177 wl_61 vdd gnd cell_6t
Xbit_r62_c177 bl_177 br_177 wl_62 vdd gnd cell_6t
Xbit_r63_c177 bl_177 br_177 wl_63 vdd gnd cell_6t
Xbit_r64_c177 bl_177 br_177 wl_64 vdd gnd cell_6t
Xbit_r65_c177 bl_177 br_177 wl_65 vdd gnd cell_6t
Xbit_r66_c177 bl_177 br_177 wl_66 vdd gnd cell_6t
Xbit_r67_c177 bl_177 br_177 wl_67 vdd gnd cell_6t
Xbit_r68_c177 bl_177 br_177 wl_68 vdd gnd cell_6t
Xbit_r69_c177 bl_177 br_177 wl_69 vdd gnd cell_6t
Xbit_r70_c177 bl_177 br_177 wl_70 vdd gnd cell_6t
Xbit_r71_c177 bl_177 br_177 wl_71 vdd gnd cell_6t
Xbit_r72_c177 bl_177 br_177 wl_72 vdd gnd cell_6t
Xbit_r73_c177 bl_177 br_177 wl_73 vdd gnd cell_6t
Xbit_r74_c177 bl_177 br_177 wl_74 vdd gnd cell_6t
Xbit_r75_c177 bl_177 br_177 wl_75 vdd gnd cell_6t
Xbit_r76_c177 bl_177 br_177 wl_76 vdd gnd cell_6t
Xbit_r77_c177 bl_177 br_177 wl_77 vdd gnd cell_6t
Xbit_r78_c177 bl_177 br_177 wl_78 vdd gnd cell_6t
Xbit_r79_c177 bl_177 br_177 wl_79 vdd gnd cell_6t
Xbit_r80_c177 bl_177 br_177 wl_80 vdd gnd cell_6t
Xbit_r81_c177 bl_177 br_177 wl_81 vdd gnd cell_6t
Xbit_r82_c177 bl_177 br_177 wl_82 vdd gnd cell_6t
Xbit_r83_c177 bl_177 br_177 wl_83 vdd gnd cell_6t
Xbit_r84_c177 bl_177 br_177 wl_84 vdd gnd cell_6t
Xbit_r85_c177 bl_177 br_177 wl_85 vdd gnd cell_6t
Xbit_r86_c177 bl_177 br_177 wl_86 vdd gnd cell_6t
Xbit_r87_c177 bl_177 br_177 wl_87 vdd gnd cell_6t
Xbit_r88_c177 bl_177 br_177 wl_88 vdd gnd cell_6t
Xbit_r89_c177 bl_177 br_177 wl_89 vdd gnd cell_6t
Xbit_r90_c177 bl_177 br_177 wl_90 vdd gnd cell_6t
Xbit_r91_c177 bl_177 br_177 wl_91 vdd gnd cell_6t
Xbit_r92_c177 bl_177 br_177 wl_92 vdd gnd cell_6t
Xbit_r93_c177 bl_177 br_177 wl_93 vdd gnd cell_6t
Xbit_r94_c177 bl_177 br_177 wl_94 vdd gnd cell_6t
Xbit_r95_c177 bl_177 br_177 wl_95 vdd gnd cell_6t
Xbit_r96_c177 bl_177 br_177 wl_96 vdd gnd cell_6t
Xbit_r97_c177 bl_177 br_177 wl_97 vdd gnd cell_6t
Xbit_r98_c177 bl_177 br_177 wl_98 vdd gnd cell_6t
Xbit_r99_c177 bl_177 br_177 wl_99 vdd gnd cell_6t
Xbit_r100_c177 bl_177 br_177 wl_100 vdd gnd cell_6t
Xbit_r101_c177 bl_177 br_177 wl_101 vdd gnd cell_6t
Xbit_r102_c177 bl_177 br_177 wl_102 vdd gnd cell_6t
Xbit_r103_c177 bl_177 br_177 wl_103 vdd gnd cell_6t
Xbit_r104_c177 bl_177 br_177 wl_104 vdd gnd cell_6t
Xbit_r105_c177 bl_177 br_177 wl_105 vdd gnd cell_6t
Xbit_r106_c177 bl_177 br_177 wl_106 vdd gnd cell_6t
Xbit_r107_c177 bl_177 br_177 wl_107 vdd gnd cell_6t
Xbit_r108_c177 bl_177 br_177 wl_108 vdd gnd cell_6t
Xbit_r109_c177 bl_177 br_177 wl_109 vdd gnd cell_6t
Xbit_r110_c177 bl_177 br_177 wl_110 vdd gnd cell_6t
Xbit_r111_c177 bl_177 br_177 wl_111 vdd gnd cell_6t
Xbit_r112_c177 bl_177 br_177 wl_112 vdd gnd cell_6t
Xbit_r113_c177 bl_177 br_177 wl_113 vdd gnd cell_6t
Xbit_r114_c177 bl_177 br_177 wl_114 vdd gnd cell_6t
Xbit_r115_c177 bl_177 br_177 wl_115 vdd gnd cell_6t
Xbit_r116_c177 bl_177 br_177 wl_116 vdd gnd cell_6t
Xbit_r117_c177 bl_177 br_177 wl_117 vdd gnd cell_6t
Xbit_r118_c177 bl_177 br_177 wl_118 vdd gnd cell_6t
Xbit_r119_c177 bl_177 br_177 wl_119 vdd gnd cell_6t
Xbit_r120_c177 bl_177 br_177 wl_120 vdd gnd cell_6t
Xbit_r121_c177 bl_177 br_177 wl_121 vdd gnd cell_6t
Xbit_r122_c177 bl_177 br_177 wl_122 vdd gnd cell_6t
Xbit_r123_c177 bl_177 br_177 wl_123 vdd gnd cell_6t
Xbit_r124_c177 bl_177 br_177 wl_124 vdd gnd cell_6t
Xbit_r125_c177 bl_177 br_177 wl_125 vdd gnd cell_6t
Xbit_r126_c177 bl_177 br_177 wl_126 vdd gnd cell_6t
Xbit_r127_c177 bl_177 br_177 wl_127 vdd gnd cell_6t
Xbit_r128_c177 bl_177 br_177 wl_128 vdd gnd cell_6t
Xbit_r129_c177 bl_177 br_177 wl_129 vdd gnd cell_6t
Xbit_r130_c177 bl_177 br_177 wl_130 vdd gnd cell_6t
Xbit_r131_c177 bl_177 br_177 wl_131 vdd gnd cell_6t
Xbit_r132_c177 bl_177 br_177 wl_132 vdd gnd cell_6t
Xbit_r133_c177 bl_177 br_177 wl_133 vdd gnd cell_6t
Xbit_r134_c177 bl_177 br_177 wl_134 vdd gnd cell_6t
Xbit_r135_c177 bl_177 br_177 wl_135 vdd gnd cell_6t
Xbit_r136_c177 bl_177 br_177 wl_136 vdd gnd cell_6t
Xbit_r137_c177 bl_177 br_177 wl_137 vdd gnd cell_6t
Xbit_r138_c177 bl_177 br_177 wl_138 vdd gnd cell_6t
Xbit_r139_c177 bl_177 br_177 wl_139 vdd gnd cell_6t
Xbit_r140_c177 bl_177 br_177 wl_140 vdd gnd cell_6t
Xbit_r141_c177 bl_177 br_177 wl_141 vdd gnd cell_6t
Xbit_r142_c177 bl_177 br_177 wl_142 vdd gnd cell_6t
Xbit_r143_c177 bl_177 br_177 wl_143 vdd gnd cell_6t
Xbit_r144_c177 bl_177 br_177 wl_144 vdd gnd cell_6t
Xbit_r145_c177 bl_177 br_177 wl_145 vdd gnd cell_6t
Xbit_r146_c177 bl_177 br_177 wl_146 vdd gnd cell_6t
Xbit_r147_c177 bl_177 br_177 wl_147 vdd gnd cell_6t
Xbit_r148_c177 bl_177 br_177 wl_148 vdd gnd cell_6t
Xbit_r149_c177 bl_177 br_177 wl_149 vdd gnd cell_6t
Xbit_r150_c177 bl_177 br_177 wl_150 vdd gnd cell_6t
Xbit_r151_c177 bl_177 br_177 wl_151 vdd gnd cell_6t
Xbit_r152_c177 bl_177 br_177 wl_152 vdd gnd cell_6t
Xbit_r153_c177 bl_177 br_177 wl_153 vdd gnd cell_6t
Xbit_r154_c177 bl_177 br_177 wl_154 vdd gnd cell_6t
Xbit_r155_c177 bl_177 br_177 wl_155 vdd gnd cell_6t
Xbit_r156_c177 bl_177 br_177 wl_156 vdd gnd cell_6t
Xbit_r157_c177 bl_177 br_177 wl_157 vdd gnd cell_6t
Xbit_r158_c177 bl_177 br_177 wl_158 vdd gnd cell_6t
Xbit_r159_c177 bl_177 br_177 wl_159 vdd gnd cell_6t
Xbit_r160_c177 bl_177 br_177 wl_160 vdd gnd cell_6t
Xbit_r161_c177 bl_177 br_177 wl_161 vdd gnd cell_6t
Xbit_r162_c177 bl_177 br_177 wl_162 vdd gnd cell_6t
Xbit_r163_c177 bl_177 br_177 wl_163 vdd gnd cell_6t
Xbit_r164_c177 bl_177 br_177 wl_164 vdd gnd cell_6t
Xbit_r165_c177 bl_177 br_177 wl_165 vdd gnd cell_6t
Xbit_r166_c177 bl_177 br_177 wl_166 vdd gnd cell_6t
Xbit_r167_c177 bl_177 br_177 wl_167 vdd gnd cell_6t
Xbit_r168_c177 bl_177 br_177 wl_168 vdd gnd cell_6t
Xbit_r169_c177 bl_177 br_177 wl_169 vdd gnd cell_6t
Xbit_r170_c177 bl_177 br_177 wl_170 vdd gnd cell_6t
Xbit_r171_c177 bl_177 br_177 wl_171 vdd gnd cell_6t
Xbit_r172_c177 bl_177 br_177 wl_172 vdd gnd cell_6t
Xbit_r173_c177 bl_177 br_177 wl_173 vdd gnd cell_6t
Xbit_r174_c177 bl_177 br_177 wl_174 vdd gnd cell_6t
Xbit_r175_c177 bl_177 br_177 wl_175 vdd gnd cell_6t
Xbit_r176_c177 bl_177 br_177 wl_176 vdd gnd cell_6t
Xbit_r177_c177 bl_177 br_177 wl_177 vdd gnd cell_6t
Xbit_r178_c177 bl_177 br_177 wl_178 vdd gnd cell_6t
Xbit_r179_c177 bl_177 br_177 wl_179 vdd gnd cell_6t
Xbit_r180_c177 bl_177 br_177 wl_180 vdd gnd cell_6t
Xbit_r181_c177 bl_177 br_177 wl_181 vdd gnd cell_6t
Xbit_r182_c177 bl_177 br_177 wl_182 vdd gnd cell_6t
Xbit_r183_c177 bl_177 br_177 wl_183 vdd gnd cell_6t
Xbit_r184_c177 bl_177 br_177 wl_184 vdd gnd cell_6t
Xbit_r185_c177 bl_177 br_177 wl_185 vdd gnd cell_6t
Xbit_r186_c177 bl_177 br_177 wl_186 vdd gnd cell_6t
Xbit_r187_c177 bl_177 br_177 wl_187 vdd gnd cell_6t
Xbit_r188_c177 bl_177 br_177 wl_188 vdd gnd cell_6t
Xbit_r189_c177 bl_177 br_177 wl_189 vdd gnd cell_6t
Xbit_r190_c177 bl_177 br_177 wl_190 vdd gnd cell_6t
Xbit_r191_c177 bl_177 br_177 wl_191 vdd gnd cell_6t
Xbit_r192_c177 bl_177 br_177 wl_192 vdd gnd cell_6t
Xbit_r193_c177 bl_177 br_177 wl_193 vdd gnd cell_6t
Xbit_r194_c177 bl_177 br_177 wl_194 vdd gnd cell_6t
Xbit_r195_c177 bl_177 br_177 wl_195 vdd gnd cell_6t
Xbit_r196_c177 bl_177 br_177 wl_196 vdd gnd cell_6t
Xbit_r197_c177 bl_177 br_177 wl_197 vdd gnd cell_6t
Xbit_r198_c177 bl_177 br_177 wl_198 vdd gnd cell_6t
Xbit_r199_c177 bl_177 br_177 wl_199 vdd gnd cell_6t
Xbit_r200_c177 bl_177 br_177 wl_200 vdd gnd cell_6t
Xbit_r201_c177 bl_177 br_177 wl_201 vdd gnd cell_6t
Xbit_r202_c177 bl_177 br_177 wl_202 vdd gnd cell_6t
Xbit_r203_c177 bl_177 br_177 wl_203 vdd gnd cell_6t
Xbit_r204_c177 bl_177 br_177 wl_204 vdd gnd cell_6t
Xbit_r205_c177 bl_177 br_177 wl_205 vdd gnd cell_6t
Xbit_r206_c177 bl_177 br_177 wl_206 vdd gnd cell_6t
Xbit_r207_c177 bl_177 br_177 wl_207 vdd gnd cell_6t
Xbit_r208_c177 bl_177 br_177 wl_208 vdd gnd cell_6t
Xbit_r209_c177 bl_177 br_177 wl_209 vdd gnd cell_6t
Xbit_r210_c177 bl_177 br_177 wl_210 vdd gnd cell_6t
Xbit_r211_c177 bl_177 br_177 wl_211 vdd gnd cell_6t
Xbit_r212_c177 bl_177 br_177 wl_212 vdd gnd cell_6t
Xbit_r213_c177 bl_177 br_177 wl_213 vdd gnd cell_6t
Xbit_r214_c177 bl_177 br_177 wl_214 vdd gnd cell_6t
Xbit_r215_c177 bl_177 br_177 wl_215 vdd gnd cell_6t
Xbit_r216_c177 bl_177 br_177 wl_216 vdd gnd cell_6t
Xbit_r217_c177 bl_177 br_177 wl_217 vdd gnd cell_6t
Xbit_r218_c177 bl_177 br_177 wl_218 vdd gnd cell_6t
Xbit_r219_c177 bl_177 br_177 wl_219 vdd gnd cell_6t
Xbit_r220_c177 bl_177 br_177 wl_220 vdd gnd cell_6t
Xbit_r221_c177 bl_177 br_177 wl_221 vdd gnd cell_6t
Xbit_r222_c177 bl_177 br_177 wl_222 vdd gnd cell_6t
Xbit_r223_c177 bl_177 br_177 wl_223 vdd gnd cell_6t
Xbit_r224_c177 bl_177 br_177 wl_224 vdd gnd cell_6t
Xbit_r225_c177 bl_177 br_177 wl_225 vdd gnd cell_6t
Xbit_r226_c177 bl_177 br_177 wl_226 vdd gnd cell_6t
Xbit_r227_c177 bl_177 br_177 wl_227 vdd gnd cell_6t
Xbit_r228_c177 bl_177 br_177 wl_228 vdd gnd cell_6t
Xbit_r229_c177 bl_177 br_177 wl_229 vdd gnd cell_6t
Xbit_r230_c177 bl_177 br_177 wl_230 vdd gnd cell_6t
Xbit_r231_c177 bl_177 br_177 wl_231 vdd gnd cell_6t
Xbit_r232_c177 bl_177 br_177 wl_232 vdd gnd cell_6t
Xbit_r233_c177 bl_177 br_177 wl_233 vdd gnd cell_6t
Xbit_r234_c177 bl_177 br_177 wl_234 vdd gnd cell_6t
Xbit_r235_c177 bl_177 br_177 wl_235 vdd gnd cell_6t
Xbit_r236_c177 bl_177 br_177 wl_236 vdd gnd cell_6t
Xbit_r237_c177 bl_177 br_177 wl_237 vdd gnd cell_6t
Xbit_r238_c177 bl_177 br_177 wl_238 vdd gnd cell_6t
Xbit_r239_c177 bl_177 br_177 wl_239 vdd gnd cell_6t
Xbit_r240_c177 bl_177 br_177 wl_240 vdd gnd cell_6t
Xbit_r241_c177 bl_177 br_177 wl_241 vdd gnd cell_6t
Xbit_r242_c177 bl_177 br_177 wl_242 vdd gnd cell_6t
Xbit_r243_c177 bl_177 br_177 wl_243 vdd gnd cell_6t
Xbit_r244_c177 bl_177 br_177 wl_244 vdd gnd cell_6t
Xbit_r245_c177 bl_177 br_177 wl_245 vdd gnd cell_6t
Xbit_r246_c177 bl_177 br_177 wl_246 vdd gnd cell_6t
Xbit_r247_c177 bl_177 br_177 wl_247 vdd gnd cell_6t
Xbit_r248_c177 bl_177 br_177 wl_248 vdd gnd cell_6t
Xbit_r249_c177 bl_177 br_177 wl_249 vdd gnd cell_6t
Xbit_r250_c177 bl_177 br_177 wl_250 vdd gnd cell_6t
Xbit_r251_c177 bl_177 br_177 wl_251 vdd gnd cell_6t
Xbit_r252_c177 bl_177 br_177 wl_252 vdd gnd cell_6t
Xbit_r253_c177 bl_177 br_177 wl_253 vdd gnd cell_6t
Xbit_r254_c177 bl_177 br_177 wl_254 vdd gnd cell_6t
Xbit_r255_c177 bl_177 br_177 wl_255 vdd gnd cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd cell_6t
Xbit_r1_c178 bl_178 br_178 wl_1 vdd gnd cell_6t
Xbit_r2_c178 bl_178 br_178 wl_2 vdd gnd cell_6t
Xbit_r3_c178 bl_178 br_178 wl_3 vdd gnd cell_6t
Xbit_r4_c178 bl_178 br_178 wl_4 vdd gnd cell_6t
Xbit_r5_c178 bl_178 br_178 wl_5 vdd gnd cell_6t
Xbit_r6_c178 bl_178 br_178 wl_6 vdd gnd cell_6t
Xbit_r7_c178 bl_178 br_178 wl_7 vdd gnd cell_6t
Xbit_r8_c178 bl_178 br_178 wl_8 vdd gnd cell_6t
Xbit_r9_c178 bl_178 br_178 wl_9 vdd gnd cell_6t
Xbit_r10_c178 bl_178 br_178 wl_10 vdd gnd cell_6t
Xbit_r11_c178 bl_178 br_178 wl_11 vdd gnd cell_6t
Xbit_r12_c178 bl_178 br_178 wl_12 vdd gnd cell_6t
Xbit_r13_c178 bl_178 br_178 wl_13 vdd gnd cell_6t
Xbit_r14_c178 bl_178 br_178 wl_14 vdd gnd cell_6t
Xbit_r15_c178 bl_178 br_178 wl_15 vdd gnd cell_6t
Xbit_r16_c178 bl_178 br_178 wl_16 vdd gnd cell_6t
Xbit_r17_c178 bl_178 br_178 wl_17 vdd gnd cell_6t
Xbit_r18_c178 bl_178 br_178 wl_18 vdd gnd cell_6t
Xbit_r19_c178 bl_178 br_178 wl_19 vdd gnd cell_6t
Xbit_r20_c178 bl_178 br_178 wl_20 vdd gnd cell_6t
Xbit_r21_c178 bl_178 br_178 wl_21 vdd gnd cell_6t
Xbit_r22_c178 bl_178 br_178 wl_22 vdd gnd cell_6t
Xbit_r23_c178 bl_178 br_178 wl_23 vdd gnd cell_6t
Xbit_r24_c178 bl_178 br_178 wl_24 vdd gnd cell_6t
Xbit_r25_c178 bl_178 br_178 wl_25 vdd gnd cell_6t
Xbit_r26_c178 bl_178 br_178 wl_26 vdd gnd cell_6t
Xbit_r27_c178 bl_178 br_178 wl_27 vdd gnd cell_6t
Xbit_r28_c178 bl_178 br_178 wl_28 vdd gnd cell_6t
Xbit_r29_c178 bl_178 br_178 wl_29 vdd gnd cell_6t
Xbit_r30_c178 bl_178 br_178 wl_30 vdd gnd cell_6t
Xbit_r31_c178 bl_178 br_178 wl_31 vdd gnd cell_6t
Xbit_r32_c178 bl_178 br_178 wl_32 vdd gnd cell_6t
Xbit_r33_c178 bl_178 br_178 wl_33 vdd gnd cell_6t
Xbit_r34_c178 bl_178 br_178 wl_34 vdd gnd cell_6t
Xbit_r35_c178 bl_178 br_178 wl_35 vdd gnd cell_6t
Xbit_r36_c178 bl_178 br_178 wl_36 vdd gnd cell_6t
Xbit_r37_c178 bl_178 br_178 wl_37 vdd gnd cell_6t
Xbit_r38_c178 bl_178 br_178 wl_38 vdd gnd cell_6t
Xbit_r39_c178 bl_178 br_178 wl_39 vdd gnd cell_6t
Xbit_r40_c178 bl_178 br_178 wl_40 vdd gnd cell_6t
Xbit_r41_c178 bl_178 br_178 wl_41 vdd gnd cell_6t
Xbit_r42_c178 bl_178 br_178 wl_42 vdd gnd cell_6t
Xbit_r43_c178 bl_178 br_178 wl_43 vdd gnd cell_6t
Xbit_r44_c178 bl_178 br_178 wl_44 vdd gnd cell_6t
Xbit_r45_c178 bl_178 br_178 wl_45 vdd gnd cell_6t
Xbit_r46_c178 bl_178 br_178 wl_46 vdd gnd cell_6t
Xbit_r47_c178 bl_178 br_178 wl_47 vdd gnd cell_6t
Xbit_r48_c178 bl_178 br_178 wl_48 vdd gnd cell_6t
Xbit_r49_c178 bl_178 br_178 wl_49 vdd gnd cell_6t
Xbit_r50_c178 bl_178 br_178 wl_50 vdd gnd cell_6t
Xbit_r51_c178 bl_178 br_178 wl_51 vdd gnd cell_6t
Xbit_r52_c178 bl_178 br_178 wl_52 vdd gnd cell_6t
Xbit_r53_c178 bl_178 br_178 wl_53 vdd gnd cell_6t
Xbit_r54_c178 bl_178 br_178 wl_54 vdd gnd cell_6t
Xbit_r55_c178 bl_178 br_178 wl_55 vdd gnd cell_6t
Xbit_r56_c178 bl_178 br_178 wl_56 vdd gnd cell_6t
Xbit_r57_c178 bl_178 br_178 wl_57 vdd gnd cell_6t
Xbit_r58_c178 bl_178 br_178 wl_58 vdd gnd cell_6t
Xbit_r59_c178 bl_178 br_178 wl_59 vdd gnd cell_6t
Xbit_r60_c178 bl_178 br_178 wl_60 vdd gnd cell_6t
Xbit_r61_c178 bl_178 br_178 wl_61 vdd gnd cell_6t
Xbit_r62_c178 bl_178 br_178 wl_62 vdd gnd cell_6t
Xbit_r63_c178 bl_178 br_178 wl_63 vdd gnd cell_6t
Xbit_r64_c178 bl_178 br_178 wl_64 vdd gnd cell_6t
Xbit_r65_c178 bl_178 br_178 wl_65 vdd gnd cell_6t
Xbit_r66_c178 bl_178 br_178 wl_66 vdd gnd cell_6t
Xbit_r67_c178 bl_178 br_178 wl_67 vdd gnd cell_6t
Xbit_r68_c178 bl_178 br_178 wl_68 vdd gnd cell_6t
Xbit_r69_c178 bl_178 br_178 wl_69 vdd gnd cell_6t
Xbit_r70_c178 bl_178 br_178 wl_70 vdd gnd cell_6t
Xbit_r71_c178 bl_178 br_178 wl_71 vdd gnd cell_6t
Xbit_r72_c178 bl_178 br_178 wl_72 vdd gnd cell_6t
Xbit_r73_c178 bl_178 br_178 wl_73 vdd gnd cell_6t
Xbit_r74_c178 bl_178 br_178 wl_74 vdd gnd cell_6t
Xbit_r75_c178 bl_178 br_178 wl_75 vdd gnd cell_6t
Xbit_r76_c178 bl_178 br_178 wl_76 vdd gnd cell_6t
Xbit_r77_c178 bl_178 br_178 wl_77 vdd gnd cell_6t
Xbit_r78_c178 bl_178 br_178 wl_78 vdd gnd cell_6t
Xbit_r79_c178 bl_178 br_178 wl_79 vdd gnd cell_6t
Xbit_r80_c178 bl_178 br_178 wl_80 vdd gnd cell_6t
Xbit_r81_c178 bl_178 br_178 wl_81 vdd gnd cell_6t
Xbit_r82_c178 bl_178 br_178 wl_82 vdd gnd cell_6t
Xbit_r83_c178 bl_178 br_178 wl_83 vdd gnd cell_6t
Xbit_r84_c178 bl_178 br_178 wl_84 vdd gnd cell_6t
Xbit_r85_c178 bl_178 br_178 wl_85 vdd gnd cell_6t
Xbit_r86_c178 bl_178 br_178 wl_86 vdd gnd cell_6t
Xbit_r87_c178 bl_178 br_178 wl_87 vdd gnd cell_6t
Xbit_r88_c178 bl_178 br_178 wl_88 vdd gnd cell_6t
Xbit_r89_c178 bl_178 br_178 wl_89 vdd gnd cell_6t
Xbit_r90_c178 bl_178 br_178 wl_90 vdd gnd cell_6t
Xbit_r91_c178 bl_178 br_178 wl_91 vdd gnd cell_6t
Xbit_r92_c178 bl_178 br_178 wl_92 vdd gnd cell_6t
Xbit_r93_c178 bl_178 br_178 wl_93 vdd gnd cell_6t
Xbit_r94_c178 bl_178 br_178 wl_94 vdd gnd cell_6t
Xbit_r95_c178 bl_178 br_178 wl_95 vdd gnd cell_6t
Xbit_r96_c178 bl_178 br_178 wl_96 vdd gnd cell_6t
Xbit_r97_c178 bl_178 br_178 wl_97 vdd gnd cell_6t
Xbit_r98_c178 bl_178 br_178 wl_98 vdd gnd cell_6t
Xbit_r99_c178 bl_178 br_178 wl_99 vdd gnd cell_6t
Xbit_r100_c178 bl_178 br_178 wl_100 vdd gnd cell_6t
Xbit_r101_c178 bl_178 br_178 wl_101 vdd gnd cell_6t
Xbit_r102_c178 bl_178 br_178 wl_102 vdd gnd cell_6t
Xbit_r103_c178 bl_178 br_178 wl_103 vdd gnd cell_6t
Xbit_r104_c178 bl_178 br_178 wl_104 vdd gnd cell_6t
Xbit_r105_c178 bl_178 br_178 wl_105 vdd gnd cell_6t
Xbit_r106_c178 bl_178 br_178 wl_106 vdd gnd cell_6t
Xbit_r107_c178 bl_178 br_178 wl_107 vdd gnd cell_6t
Xbit_r108_c178 bl_178 br_178 wl_108 vdd gnd cell_6t
Xbit_r109_c178 bl_178 br_178 wl_109 vdd gnd cell_6t
Xbit_r110_c178 bl_178 br_178 wl_110 vdd gnd cell_6t
Xbit_r111_c178 bl_178 br_178 wl_111 vdd gnd cell_6t
Xbit_r112_c178 bl_178 br_178 wl_112 vdd gnd cell_6t
Xbit_r113_c178 bl_178 br_178 wl_113 vdd gnd cell_6t
Xbit_r114_c178 bl_178 br_178 wl_114 vdd gnd cell_6t
Xbit_r115_c178 bl_178 br_178 wl_115 vdd gnd cell_6t
Xbit_r116_c178 bl_178 br_178 wl_116 vdd gnd cell_6t
Xbit_r117_c178 bl_178 br_178 wl_117 vdd gnd cell_6t
Xbit_r118_c178 bl_178 br_178 wl_118 vdd gnd cell_6t
Xbit_r119_c178 bl_178 br_178 wl_119 vdd gnd cell_6t
Xbit_r120_c178 bl_178 br_178 wl_120 vdd gnd cell_6t
Xbit_r121_c178 bl_178 br_178 wl_121 vdd gnd cell_6t
Xbit_r122_c178 bl_178 br_178 wl_122 vdd gnd cell_6t
Xbit_r123_c178 bl_178 br_178 wl_123 vdd gnd cell_6t
Xbit_r124_c178 bl_178 br_178 wl_124 vdd gnd cell_6t
Xbit_r125_c178 bl_178 br_178 wl_125 vdd gnd cell_6t
Xbit_r126_c178 bl_178 br_178 wl_126 vdd gnd cell_6t
Xbit_r127_c178 bl_178 br_178 wl_127 vdd gnd cell_6t
Xbit_r128_c178 bl_178 br_178 wl_128 vdd gnd cell_6t
Xbit_r129_c178 bl_178 br_178 wl_129 vdd gnd cell_6t
Xbit_r130_c178 bl_178 br_178 wl_130 vdd gnd cell_6t
Xbit_r131_c178 bl_178 br_178 wl_131 vdd gnd cell_6t
Xbit_r132_c178 bl_178 br_178 wl_132 vdd gnd cell_6t
Xbit_r133_c178 bl_178 br_178 wl_133 vdd gnd cell_6t
Xbit_r134_c178 bl_178 br_178 wl_134 vdd gnd cell_6t
Xbit_r135_c178 bl_178 br_178 wl_135 vdd gnd cell_6t
Xbit_r136_c178 bl_178 br_178 wl_136 vdd gnd cell_6t
Xbit_r137_c178 bl_178 br_178 wl_137 vdd gnd cell_6t
Xbit_r138_c178 bl_178 br_178 wl_138 vdd gnd cell_6t
Xbit_r139_c178 bl_178 br_178 wl_139 vdd gnd cell_6t
Xbit_r140_c178 bl_178 br_178 wl_140 vdd gnd cell_6t
Xbit_r141_c178 bl_178 br_178 wl_141 vdd gnd cell_6t
Xbit_r142_c178 bl_178 br_178 wl_142 vdd gnd cell_6t
Xbit_r143_c178 bl_178 br_178 wl_143 vdd gnd cell_6t
Xbit_r144_c178 bl_178 br_178 wl_144 vdd gnd cell_6t
Xbit_r145_c178 bl_178 br_178 wl_145 vdd gnd cell_6t
Xbit_r146_c178 bl_178 br_178 wl_146 vdd gnd cell_6t
Xbit_r147_c178 bl_178 br_178 wl_147 vdd gnd cell_6t
Xbit_r148_c178 bl_178 br_178 wl_148 vdd gnd cell_6t
Xbit_r149_c178 bl_178 br_178 wl_149 vdd gnd cell_6t
Xbit_r150_c178 bl_178 br_178 wl_150 vdd gnd cell_6t
Xbit_r151_c178 bl_178 br_178 wl_151 vdd gnd cell_6t
Xbit_r152_c178 bl_178 br_178 wl_152 vdd gnd cell_6t
Xbit_r153_c178 bl_178 br_178 wl_153 vdd gnd cell_6t
Xbit_r154_c178 bl_178 br_178 wl_154 vdd gnd cell_6t
Xbit_r155_c178 bl_178 br_178 wl_155 vdd gnd cell_6t
Xbit_r156_c178 bl_178 br_178 wl_156 vdd gnd cell_6t
Xbit_r157_c178 bl_178 br_178 wl_157 vdd gnd cell_6t
Xbit_r158_c178 bl_178 br_178 wl_158 vdd gnd cell_6t
Xbit_r159_c178 bl_178 br_178 wl_159 vdd gnd cell_6t
Xbit_r160_c178 bl_178 br_178 wl_160 vdd gnd cell_6t
Xbit_r161_c178 bl_178 br_178 wl_161 vdd gnd cell_6t
Xbit_r162_c178 bl_178 br_178 wl_162 vdd gnd cell_6t
Xbit_r163_c178 bl_178 br_178 wl_163 vdd gnd cell_6t
Xbit_r164_c178 bl_178 br_178 wl_164 vdd gnd cell_6t
Xbit_r165_c178 bl_178 br_178 wl_165 vdd gnd cell_6t
Xbit_r166_c178 bl_178 br_178 wl_166 vdd gnd cell_6t
Xbit_r167_c178 bl_178 br_178 wl_167 vdd gnd cell_6t
Xbit_r168_c178 bl_178 br_178 wl_168 vdd gnd cell_6t
Xbit_r169_c178 bl_178 br_178 wl_169 vdd gnd cell_6t
Xbit_r170_c178 bl_178 br_178 wl_170 vdd gnd cell_6t
Xbit_r171_c178 bl_178 br_178 wl_171 vdd gnd cell_6t
Xbit_r172_c178 bl_178 br_178 wl_172 vdd gnd cell_6t
Xbit_r173_c178 bl_178 br_178 wl_173 vdd gnd cell_6t
Xbit_r174_c178 bl_178 br_178 wl_174 vdd gnd cell_6t
Xbit_r175_c178 bl_178 br_178 wl_175 vdd gnd cell_6t
Xbit_r176_c178 bl_178 br_178 wl_176 vdd gnd cell_6t
Xbit_r177_c178 bl_178 br_178 wl_177 vdd gnd cell_6t
Xbit_r178_c178 bl_178 br_178 wl_178 vdd gnd cell_6t
Xbit_r179_c178 bl_178 br_178 wl_179 vdd gnd cell_6t
Xbit_r180_c178 bl_178 br_178 wl_180 vdd gnd cell_6t
Xbit_r181_c178 bl_178 br_178 wl_181 vdd gnd cell_6t
Xbit_r182_c178 bl_178 br_178 wl_182 vdd gnd cell_6t
Xbit_r183_c178 bl_178 br_178 wl_183 vdd gnd cell_6t
Xbit_r184_c178 bl_178 br_178 wl_184 vdd gnd cell_6t
Xbit_r185_c178 bl_178 br_178 wl_185 vdd gnd cell_6t
Xbit_r186_c178 bl_178 br_178 wl_186 vdd gnd cell_6t
Xbit_r187_c178 bl_178 br_178 wl_187 vdd gnd cell_6t
Xbit_r188_c178 bl_178 br_178 wl_188 vdd gnd cell_6t
Xbit_r189_c178 bl_178 br_178 wl_189 vdd gnd cell_6t
Xbit_r190_c178 bl_178 br_178 wl_190 vdd gnd cell_6t
Xbit_r191_c178 bl_178 br_178 wl_191 vdd gnd cell_6t
Xbit_r192_c178 bl_178 br_178 wl_192 vdd gnd cell_6t
Xbit_r193_c178 bl_178 br_178 wl_193 vdd gnd cell_6t
Xbit_r194_c178 bl_178 br_178 wl_194 vdd gnd cell_6t
Xbit_r195_c178 bl_178 br_178 wl_195 vdd gnd cell_6t
Xbit_r196_c178 bl_178 br_178 wl_196 vdd gnd cell_6t
Xbit_r197_c178 bl_178 br_178 wl_197 vdd gnd cell_6t
Xbit_r198_c178 bl_178 br_178 wl_198 vdd gnd cell_6t
Xbit_r199_c178 bl_178 br_178 wl_199 vdd gnd cell_6t
Xbit_r200_c178 bl_178 br_178 wl_200 vdd gnd cell_6t
Xbit_r201_c178 bl_178 br_178 wl_201 vdd gnd cell_6t
Xbit_r202_c178 bl_178 br_178 wl_202 vdd gnd cell_6t
Xbit_r203_c178 bl_178 br_178 wl_203 vdd gnd cell_6t
Xbit_r204_c178 bl_178 br_178 wl_204 vdd gnd cell_6t
Xbit_r205_c178 bl_178 br_178 wl_205 vdd gnd cell_6t
Xbit_r206_c178 bl_178 br_178 wl_206 vdd gnd cell_6t
Xbit_r207_c178 bl_178 br_178 wl_207 vdd gnd cell_6t
Xbit_r208_c178 bl_178 br_178 wl_208 vdd gnd cell_6t
Xbit_r209_c178 bl_178 br_178 wl_209 vdd gnd cell_6t
Xbit_r210_c178 bl_178 br_178 wl_210 vdd gnd cell_6t
Xbit_r211_c178 bl_178 br_178 wl_211 vdd gnd cell_6t
Xbit_r212_c178 bl_178 br_178 wl_212 vdd gnd cell_6t
Xbit_r213_c178 bl_178 br_178 wl_213 vdd gnd cell_6t
Xbit_r214_c178 bl_178 br_178 wl_214 vdd gnd cell_6t
Xbit_r215_c178 bl_178 br_178 wl_215 vdd gnd cell_6t
Xbit_r216_c178 bl_178 br_178 wl_216 vdd gnd cell_6t
Xbit_r217_c178 bl_178 br_178 wl_217 vdd gnd cell_6t
Xbit_r218_c178 bl_178 br_178 wl_218 vdd gnd cell_6t
Xbit_r219_c178 bl_178 br_178 wl_219 vdd gnd cell_6t
Xbit_r220_c178 bl_178 br_178 wl_220 vdd gnd cell_6t
Xbit_r221_c178 bl_178 br_178 wl_221 vdd gnd cell_6t
Xbit_r222_c178 bl_178 br_178 wl_222 vdd gnd cell_6t
Xbit_r223_c178 bl_178 br_178 wl_223 vdd gnd cell_6t
Xbit_r224_c178 bl_178 br_178 wl_224 vdd gnd cell_6t
Xbit_r225_c178 bl_178 br_178 wl_225 vdd gnd cell_6t
Xbit_r226_c178 bl_178 br_178 wl_226 vdd gnd cell_6t
Xbit_r227_c178 bl_178 br_178 wl_227 vdd gnd cell_6t
Xbit_r228_c178 bl_178 br_178 wl_228 vdd gnd cell_6t
Xbit_r229_c178 bl_178 br_178 wl_229 vdd gnd cell_6t
Xbit_r230_c178 bl_178 br_178 wl_230 vdd gnd cell_6t
Xbit_r231_c178 bl_178 br_178 wl_231 vdd gnd cell_6t
Xbit_r232_c178 bl_178 br_178 wl_232 vdd gnd cell_6t
Xbit_r233_c178 bl_178 br_178 wl_233 vdd gnd cell_6t
Xbit_r234_c178 bl_178 br_178 wl_234 vdd gnd cell_6t
Xbit_r235_c178 bl_178 br_178 wl_235 vdd gnd cell_6t
Xbit_r236_c178 bl_178 br_178 wl_236 vdd gnd cell_6t
Xbit_r237_c178 bl_178 br_178 wl_237 vdd gnd cell_6t
Xbit_r238_c178 bl_178 br_178 wl_238 vdd gnd cell_6t
Xbit_r239_c178 bl_178 br_178 wl_239 vdd gnd cell_6t
Xbit_r240_c178 bl_178 br_178 wl_240 vdd gnd cell_6t
Xbit_r241_c178 bl_178 br_178 wl_241 vdd gnd cell_6t
Xbit_r242_c178 bl_178 br_178 wl_242 vdd gnd cell_6t
Xbit_r243_c178 bl_178 br_178 wl_243 vdd gnd cell_6t
Xbit_r244_c178 bl_178 br_178 wl_244 vdd gnd cell_6t
Xbit_r245_c178 bl_178 br_178 wl_245 vdd gnd cell_6t
Xbit_r246_c178 bl_178 br_178 wl_246 vdd gnd cell_6t
Xbit_r247_c178 bl_178 br_178 wl_247 vdd gnd cell_6t
Xbit_r248_c178 bl_178 br_178 wl_248 vdd gnd cell_6t
Xbit_r249_c178 bl_178 br_178 wl_249 vdd gnd cell_6t
Xbit_r250_c178 bl_178 br_178 wl_250 vdd gnd cell_6t
Xbit_r251_c178 bl_178 br_178 wl_251 vdd gnd cell_6t
Xbit_r252_c178 bl_178 br_178 wl_252 vdd gnd cell_6t
Xbit_r253_c178 bl_178 br_178 wl_253 vdd gnd cell_6t
Xbit_r254_c178 bl_178 br_178 wl_254 vdd gnd cell_6t
Xbit_r255_c178 bl_178 br_178 wl_255 vdd gnd cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd cell_6t
Xbit_r1_c179 bl_179 br_179 wl_1 vdd gnd cell_6t
Xbit_r2_c179 bl_179 br_179 wl_2 vdd gnd cell_6t
Xbit_r3_c179 bl_179 br_179 wl_3 vdd gnd cell_6t
Xbit_r4_c179 bl_179 br_179 wl_4 vdd gnd cell_6t
Xbit_r5_c179 bl_179 br_179 wl_5 vdd gnd cell_6t
Xbit_r6_c179 bl_179 br_179 wl_6 vdd gnd cell_6t
Xbit_r7_c179 bl_179 br_179 wl_7 vdd gnd cell_6t
Xbit_r8_c179 bl_179 br_179 wl_8 vdd gnd cell_6t
Xbit_r9_c179 bl_179 br_179 wl_9 vdd gnd cell_6t
Xbit_r10_c179 bl_179 br_179 wl_10 vdd gnd cell_6t
Xbit_r11_c179 bl_179 br_179 wl_11 vdd gnd cell_6t
Xbit_r12_c179 bl_179 br_179 wl_12 vdd gnd cell_6t
Xbit_r13_c179 bl_179 br_179 wl_13 vdd gnd cell_6t
Xbit_r14_c179 bl_179 br_179 wl_14 vdd gnd cell_6t
Xbit_r15_c179 bl_179 br_179 wl_15 vdd gnd cell_6t
Xbit_r16_c179 bl_179 br_179 wl_16 vdd gnd cell_6t
Xbit_r17_c179 bl_179 br_179 wl_17 vdd gnd cell_6t
Xbit_r18_c179 bl_179 br_179 wl_18 vdd gnd cell_6t
Xbit_r19_c179 bl_179 br_179 wl_19 vdd gnd cell_6t
Xbit_r20_c179 bl_179 br_179 wl_20 vdd gnd cell_6t
Xbit_r21_c179 bl_179 br_179 wl_21 vdd gnd cell_6t
Xbit_r22_c179 bl_179 br_179 wl_22 vdd gnd cell_6t
Xbit_r23_c179 bl_179 br_179 wl_23 vdd gnd cell_6t
Xbit_r24_c179 bl_179 br_179 wl_24 vdd gnd cell_6t
Xbit_r25_c179 bl_179 br_179 wl_25 vdd gnd cell_6t
Xbit_r26_c179 bl_179 br_179 wl_26 vdd gnd cell_6t
Xbit_r27_c179 bl_179 br_179 wl_27 vdd gnd cell_6t
Xbit_r28_c179 bl_179 br_179 wl_28 vdd gnd cell_6t
Xbit_r29_c179 bl_179 br_179 wl_29 vdd gnd cell_6t
Xbit_r30_c179 bl_179 br_179 wl_30 vdd gnd cell_6t
Xbit_r31_c179 bl_179 br_179 wl_31 vdd gnd cell_6t
Xbit_r32_c179 bl_179 br_179 wl_32 vdd gnd cell_6t
Xbit_r33_c179 bl_179 br_179 wl_33 vdd gnd cell_6t
Xbit_r34_c179 bl_179 br_179 wl_34 vdd gnd cell_6t
Xbit_r35_c179 bl_179 br_179 wl_35 vdd gnd cell_6t
Xbit_r36_c179 bl_179 br_179 wl_36 vdd gnd cell_6t
Xbit_r37_c179 bl_179 br_179 wl_37 vdd gnd cell_6t
Xbit_r38_c179 bl_179 br_179 wl_38 vdd gnd cell_6t
Xbit_r39_c179 bl_179 br_179 wl_39 vdd gnd cell_6t
Xbit_r40_c179 bl_179 br_179 wl_40 vdd gnd cell_6t
Xbit_r41_c179 bl_179 br_179 wl_41 vdd gnd cell_6t
Xbit_r42_c179 bl_179 br_179 wl_42 vdd gnd cell_6t
Xbit_r43_c179 bl_179 br_179 wl_43 vdd gnd cell_6t
Xbit_r44_c179 bl_179 br_179 wl_44 vdd gnd cell_6t
Xbit_r45_c179 bl_179 br_179 wl_45 vdd gnd cell_6t
Xbit_r46_c179 bl_179 br_179 wl_46 vdd gnd cell_6t
Xbit_r47_c179 bl_179 br_179 wl_47 vdd gnd cell_6t
Xbit_r48_c179 bl_179 br_179 wl_48 vdd gnd cell_6t
Xbit_r49_c179 bl_179 br_179 wl_49 vdd gnd cell_6t
Xbit_r50_c179 bl_179 br_179 wl_50 vdd gnd cell_6t
Xbit_r51_c179 bl_179 br_179 wl_51 vdd gnd cell_6t
Xbit_r52_c179 bl_179 br_179 wl_52 vdd gnd cell_6t
Xbit_r53_c179 bl_179 br_179 wl_53 vdd gnd cell_6t
Xbit_r54_c179 bl_179 br_179 wl_54 vdd gnd cell_6t
Xbit_r55_c179 bl_179 br_179 wl_55 vdd gnd cell_6t
Xbit_r56_c179 bl_179 br_179 wl_56 vdd gnd cell_6t
Xbit_r57_c179 bl_179 br_179 wl_57 vdd gnd cell_6t
Xbit_r58_c179 bl_179 br_179 wl_58 vdd gnd cell_6t
Xbit_r59_c179 bl_179 br_179 wl_59 vdd gnd cell_6t
Xbit_r60_c179 bl_179 br_179 wl_60 vdd gnd cell_6t
Xbit_r61_c179 bl_179 br_179 wl_61 vdd gnd cell_6t
Xbit_r62_c179 bl_179 br_179 wl_62 vdd gnd cell_6t
Xbit_r63_c179 bl_179 br_179 wl_63 vdd gnd cell_6t
Xbit_r64_c179 bl_179 br_179 wl_64 vdd gnd cell_6t
Xbit_r65_c179 bl_179 br_179 wl_65 vdd gnd cell_6t
Xbit_r66_c179 bl_179 br_179 wl_66 vdd gnd cell_6t
Xbit_r67_c179 bl_179 br_179 wl_67 vdd gnd cell_6t
Xbit_r68_c179 bl_179 br_179 wl_68 vdd gnd cell_6t
Xbit_r69_c179 bl_179 br_179 wl_69 vdd gnd cell_6t
Xbit_r70_c179 bl_179 br_179 wl_70 vdd gnd cell_6t
Xbit_r71_c179 bl_179 br_179 wl_71 vdd gnd cell_6t
Xbit_r72_c179 bl_179 br_179 wl_72 vdd gnd cell_6t
Xbit_r73_c179 bl_179 br_179 wl_73 vdd gnd cell_6t
Xbit_r74_c179 bl_179 br_179 wl_74 vdd gnd cell_6t
Xbit_r75_c179 bl_179 br_179 wl_75 vdd gnd cell_6t
Xbit_r76_c179 bl_179 br_179 wl_76 vdd gnd cell_6t
Xbit_r77_c179 bl_179 br_179 wl_77 vdd gnd cell_6t
Xbit_r78_c179 bl_179 br_179 wl_78 vdd gnd cell_6t
Xbit_r79_c179 bl_179 br_179 wl_79 vdd gnd cell_6t
Xbit_r80_c179 bl_179 br_179 wl_80 vdd gnd cell_6t
Xbit_r81_c179 bl_179 br_179 wl_81 vdd gnd cell_6t
Xbit_r82_c179 bl_179 br_179 wl_82 vdd gnd cell_6t
Xbit_r83_c179 bl_179 br_179 wl_83 vdd gnd cell_6t
Xbit_r84_c179 bl_179 br_179 wl_84 vdd gnd cell_6t
Xbit_r85_c179 bl_179 br_179 wl_85 vdd gnd cell_6t
Xbit_r86_c179 bl_179 br_179 wl_86 vdd gnd cell_6t
Xbit_r87_c179 bl_179 br_179 wl_87 vdd gnd cell_6t
Xbit_r88_c179 bl_179 br_179 wl_88 vdd gnd cell_6t
Xbit_r89_c179 bl_179 br_179 wl_89 vdd gnd cell_6t
Xbit_r90_c179 bl_179 br_179 wl_90 vdd gnd cell_6t
Xbit_r91_c179 bl_179 br_179 wl_91 vdd gnd cell_6t
Xbit_r92_c179 bl_179 br_179 wl_92 vdd gnd cell_6t
Xbit_r93_c179 bl_179 br_179 wl_93 vdd gnd cell_6t
Xbit_r94_c179 bl_179 br_179 wl_94 vdd gnd cell_6t
Xbit_r95_c179 bl_179 br_179 wl_95 vdd gnd cell_6t
Xbit_r96_c179 bl_179 br_179 wl_96 vdd gnd cell_6t
Xbit_r97_c179 bl_179 br_179 wl_97 vdd gnd cell_6t
Xbit_r98_c179 bl_179 br_179 wl_98 vdd gnd cell_6t
Xbit_r99_c179 bl_179 br_179 wl_99 vdd gnd cell_6t
Xbit_r100_c179 bl_179 br_179 wl_100 vdd gnd cell_6t
Xbit_r101_c179 bl_179 br_179 wl_101 vdd gnd cell_6t
Xbit_r102_c179 bl_179 br_179 wl_102 vdd gnd cell_6t
Xbit_r103_c179 bl_179 br_179 wl_103 vdd gnd cell_6t
Xbit_r104_c179 bl_179 br_179 wl_104 vdd gnd cell_6t
Xbit_r105_c179 bl_179 br_179 wl_105 vdd gnd cell_6t
Xbit_r106_c179 bl_179 br_179 wl_106 vdd gnd cell_6t
Xbit_r107_c179 bl_179 br_179 wl_107 vdd gnd cell_6t
Xbit_r108_c179 bl_179 br_179 wl_108 vdd gnd cell_6t
Xbit_r109_c179 bl_179 br_179 wl_109 vdd gnd cell_6t
Xbit_r110_c179 bl_179 br_179 wl_110 vdd gnd cell_6t
Xbit_r111_c179 bl_179 br_179 wl_111 vdd gnd cell_6t
Xbit_r112_c179 bl_179 br_179 wl_112 vdd gnd cell_6t
Xbit_r113_c179 bl_179 br_179 wl_113 vdd gnd cell_6t
Xbit_r114_c179 bl_179 br_179 wl_114 vdd gnd cell_6t
Xbit_r115_c179 bl_179 br_179 wl_115 vdd gnd cell_6t
Xbit_r116_c179 bl_179 br_179 wl_116 vdd gnd cell_6t
Xbit_r117_c179 bl_179 br_179 wl_117 vdd gnd cell_6t
Xbit_r118_c179 bl_179 br_179 wl_118 vdd gnd cell_6t
Xbit_r119_c179 bl_179 br_179 wl_119 vdd gnd cell_6t
Xbit_r120_c179 bl_179 br_179 wl_120 vdd gnd cell_6t
Xbit_r121_c179 bl_179 br_179 wl_121 vdd gnd cell_6t
Xbit_r122_c179 bl_179 br_179 wl_122 vdd gnd cell_6t
Xbit_r123_c179 bl_179 br_179 wl_123 vdd gnd cell_6t
Xbit_r124_c179 bl_179 br_179 wl_124 vdd gnd cell_6t
Xbit_r125_c179 bl_179 br_179 wl_125 vdd gnd cell_6t
Xbit_r126_c179 bl_179 br_179 wl_126 vdd gnd cell_6t
Xbit_r127_c179 bl_179 br_179 wl_127 vdd gnd cell_6t
Xbit_r128_c179 bl_179 br_179 wl_128 vdd gnd cell_6t
Xbit_r129_c179 bl_179 br_179 wl_129 vdd gnd cell_6t
Xbit_r130_c179 bl_179 br_179 wl_130 vdd gnd cell_6t
Xbit_r131_c179 bl_179 br_179 wl_131 vdd gnd cell_6t
Xbit_r132_c179 bl_179 br_179 wl_132 vdd gnd cell_6t
Xbit_r133_c179 bl_179 br_179 wl_133 vdd gnd cell_6t
Xbit_r134_c179 bl_179 br_179 wl_134 vdd gnd cell_6t
Xbit_r135_c179 bl_179 br_179 wl_135 vdd gnd cell_6t
Xbit_r136_c179 bl_179 br_179 wl_136 vdd gnd cell_6t
Xbit_r137_c179 bl_179 br_179 wl_137 vdd gnd cell_6t
Xbit_r138_c179 bl_179 br_179 wl_138 vdd gnd cell_6t
Xbit_r139_c179 bl_179 br_179 wl_139 vdd gnd cell_6t
Xbit_r140_c179 bl_179 br_179 wl_140 vdd gnd cell_6t
Xbit_r141_c179 bl_179 br_179 wl_141 vdd gnd cell_6t
Xbit_r142_c179 bl_179 br_179 wl_142 vdd gnd cell_6t
Xbit_r143_c179 bl_179 br_179 wl_143 vdd gnd cell_6t
Xbit_r144_c179 bl_179 br_179 wl_144 vdd gnd cell_6t
Xbit_r145_c179 bl_179 br_179 wl_145 vdd gnd cell_6t
Xbit_r146_c179 bl_179 br_179 wl_146 vdd gnd cell_6t
Xbit_r147_c179 bl_179 br_179 wl_147 vdd gnd cell_6t
Xbit_r148_c179 bl_179 br_179 wl_148 vdd gnd cell_6t
Xbit_r149_c179 bl_179 br_179 wl_149 vdd gnd cell_6t
Xbit_r150_c179 bl_179 br_179 wl_150 vdd gnd cell_6t
Xbit_r151_c179 bl_179 br_179 wl_151 vdd gnd cell_6t
Xbit_r152_c179 bl_179 br_179 wl_152 vdd gnd cell_6t
Xbit_r153_c179 bl_179 br_179 wl_153 vdd gnd cell_6t
Xbit_r154_c179 bl_179 br_179 wl_154 vdd gnd cell_6t
Xbit_r155_c179 bl_179 br_179 wl_155 vdd gnd cell_6t
Xbit_r156_c179 bl_179 br_179 wl_156 vdd gnd cell_6t
Xbit_r157_c179 bl_179 br_179 wl_157 vdd gnd cell_6t
Xbit_r158_c179 bl_179 br_179 wl_158 vdd gnd cell_6t
Xbit_r159_c179 bl_179 br_179 wl_159 vdd gnd cell_6t
Xbit_r160_c179 bl_179 br_179 wl_160 vdd gnd cell_6t
Xbit_r161_c179 bl_179 br_179 wl_161 vdd gnd cell_6t
Xbit_r162_c179 bl_179 br_179 wl_162 vdd gnd cell_6t
Xbit_r163_c179 bl_179 br_179 wl_163 vdd gnd cell_6t
Xbit_r164_c179 bl_179 br_179 wl_164 vdd gnd cell_6t
Xbit_r165_c179 bl_179 br_179 wl_165 vdd gnd cell_6t
Xbit_r166_c179 bl_179 br_179 wl_166 vdd gnd cell_6t
Xbit_r167_c179 bl_179 br_179 wl_167 vdd gnd cell_6t
Xbit_r168_c179 bl_179 br_179 wl_168 vdd gnd cell_6t
Xbit_r169_c179 bl_179 br_179 wl_169 vdd gnd cell_6t
Xbit_r170_c179 bl_179 br_179 wl_170 vdd gnd cell_6t
Xbit_r171_c179 bl_179 br_179 wl_171 vdd gnd cell_6t
Xbit_r172_c179 bl_179 br_179 wl_172 vdd gnd cell_6t
Xbit_r173_c179 bl_179 br_179 wl_173 vdd gnd cell_6t
Xbit_r174_c179 bl_179 br_179 wl_174 vdd gnd cell_6t
Xbit_r175_c179 bl_179 br_179 wl_175 vdd gnd cell_6t
Xbit_r176_c179 bl_179 br_179 wl_176 vdd gnd cell_6t
Xbit_r177_c179 bl_179 br_179 wl_177 vdd gnd cell_6t
Xbit_r178_c179 bl_179 br_179 wl_178 vdd gnd cell_6t
Xbit_r179_c179 bl_179 br_179 wl_179 vdd gnd cell_6t
Xbit_r180_c179 bl_179 br_179 wl_180 vdd gnd cell_6t
Xbit_r181_c179 bl_179 br_179 wl_181 vdd gnd cell_6t
Xbit_r182_c179 bl_179 br_179 wl_182 vdd gnd cell_6t
Xbit_r183_c179 bl_179 br_179 wl_183 vdd gnd cell_6t
Xbit_r184_c179 bl_179 br_179 wl_184 vdd gnd cell_6t
Xbit_r185_c179 bl_179 br_179 wl_185 vdd gnd cell_6t
Xbit_r186_c179 bl_179 br_179 wl_186 vdd gnd cell_6t
Xbit_r187_c179 bl_179 br_179 wl_187 vdd gnd cell_6t
Xbit_r188_c179 bl_179 br_179 wl_188 vdd gnd cell_6t
Xbit_r189_c179 bl_179 br_179 wl_189 vdd gnd cell_6t
Xbit_r190_c179 bl_179 br_179 wl_190 vdd gnd cell_6t
Xbit_r191_c179 bl_179 br_179 wl_191 vdd gnd cell_6t
Xbit_r192_c179 bl_179 br_179 wl_192 vdd gnd cell_6t
Xbit_r193_c179 bl_179 br_179 wl_193 vdd gnd cell_6t
Xbit_r194_c179 bl_179 br_179 wl_194 vdd gnd cell_6t
Xbit_r195_c179 bl_179 br_179 wl_195 vdd gnd cell_6t
Xbit_r196_c179 bl_179 br_179 wl_196 vdd gnd cell_6t
Xbit_r197_c179 bl_179 br_179 wl_197 vdd gnd cell_6t
Xbit_r198_c179 bl_179 br_179 wl_198 vdd gnd cell_6t
Xbit_r199_c179 bl_179 br_179 wl_199 vdd gnd cell_6t
Xbit_r200_c179 bl_179 br_179 wl_200 vdd gnd cell_6t
Xbit_r201_c179 bl_179 br_179 wl_201 vdd gnd cell_6t
Xbit_r202_c179 bl_179 br_179 wl_202 vdd gnd cell_6t
Xbit_r203_c179 bl_179 br_179 wl_203 vdd gnd cell_6t
Xbit_r204_c179 bl_179 br_179 wl_204 vdd gnd cell_6t
Xbit_r205_c179 bl_179 br_179 wl_205 vdd gnd cell_6t
Xbit_r206_c179 bl_179 br_179 wl_206 vdd gnd cell_6t
Xbit_r207_c179 bl_179 br_179 wl_207 vdd gnd cell_6t
Xbit_r208_c179 bl_179 br_179 wl_208 vdd gnd cell_6t
Xbit_r209_c179 bl_179 br_179 wl_209 vdd gnd cell_6t
Xbit_r210_c179 bl_179 br_179 wl_210 vdd gnd cell_6t
Xbit_r211_c179 bl_179 br_179 wl_211 vdd gnd cell_6t
Xbit_r212_c179 bl_179 br_179 wl_212 vdd gnd cell_6t
Xbit_r213_c179 bl_179 br_179 wl_213 vdd gnd cell_6t
Xbit_r214_c179 bl_179 br_179 wl_214 vdd gnd cell_6t
Xbit_r215_c179 bl_179 br_179 wl_215 vdd gnd cell_6t
Xbit_r216_c179 bl_179 br_179 wl_216 vdd gnd cell_6t
Xbit_r217_c179 bl_179 br_179 wl_217 vdd gnd cell_6t
Xbit_r218_c179 bl_179 br_179 wl_218 vdd gnd cell_6t
Xbit_r219_c179 bl_179 br_179 wl_219 vdd gnd cell_6t
Xbit_r220_c179 bl_179 br_179 wl_220 vdd gnd cell_6t
Xbit_r221_c179 bl_179 br_179 wl_221 vdd gnd cell_6t
Xbit_r222_c179 bl_179 br_179 wl_222 vdd gnd cell_6t
Xbit_r223_c179 bl_179 br_179 wl_223 vdd gnd cell_6t
Xbit_r224_c179 bl_179 br_179 wl_224 vdd gnd cell_6t
Xbit_r225_c179 bl_179 br_179 wl_225 vdd gnd cell_6t
Xbit_r226_c179 bl_179 br_179 wl_226 vdd gnd cell_6t
Xbit_r227_c179 bl_179 br_179 wl_227 vdd gnd cell_6t
Xbit_r228_c179 bl_179 br_179 wl_228 vdd gnd cell_6t
Xbit_r229_c179 bl_179 br_179 wl_229 vdd gnd cell_6t
Xbit_r230_c179 bl_179 br_179 wl_230 vdd gnd cell_6t
Xbit_r231_c179 bl_179 br_179 wl_231 vdd gnd cell_6t
Xbit_r232_c179 bl_179 br_179 wl_232 vdd gnd cell_6t
Xbit_r233_c179 bl_179 br_179 wl_233 vdd gnd cell_6t
Xbit_r234_c179 bl_179 br_179 wl_234 vdd gnd cell_6t
Xbit_r235_c179 bl_179 br_179 wl_235 vdd gnd cell_6t
Xbit_r236_c179 bl_179 br_179 wl_236 vdd gnd cell_6t
Xbit_r237_c179 bl_179 br_179 wl_237 vdd gnd cell_6t
Xbit_r238_c179 bl_179 br_179 wl_238 vdd gnd cell_6t
Xbit_r239_c179 bl_179 br_179 wl_239 vdd gnd cell_6t
Xbit_r240_c179 bl_179 br_179 wl_240 vdd gnd cell_6t
Xbit_r241_c179 bl_179 br_179 wl_241 vdd gnd cell_6t
Xbit_r242_c179 bl_179 br_179 wl_242 vdd gnd cell_6t
Xbit_r243_c179 bl_179 br_179 wl_243 vdd gnd cell_6t
Xbit_r244_c179 bl_179 br_179 wl_244 vdd gnd cell_6t
Xbit_r245_c179 bl_179 br_179 wl_245 vdd gnd cell_6t
Xbit_r246_c179 bl_179 br_179 wl_246 vdd gnd cell_6t
Xbit_r247_c179 bl_179 br_179 wl_247 vdd gnd cell_6t
Xbit_r248_c179 bl_179 br_179 wl_248 vdd gnd cell_6t
Xbit_r249_c179 bl_179 br_179 wl_249 vdd gnd cell_6t
Xbit_r250_c179 bl_179 br_179 wl_250 vdd gnd cell_6t
Xbit_r251_c179 bl_179 br_179 wl_251 vdd gnd cell_6t
Xbit_r252_c179 bl_179 br_179 wl_252 vdd gnd cell_6t
Xbit_r253_c179 bl_179 br_179 wl_253 vdd gnd cell_6t
Xbit_r254_c179 bl_179 br_179 wl_254 vdd gnd cell_6t
Xbit_r255_c179 bl_179 br_179 wl_255 vdd gnd cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd cell_6t
Xbit_r1_c180 bl_180 br_180 wl_1 vdd gnd cell_6t
Xbit_r2_c180 bl_180 br_180 wl_2 vdd gnd cell_6t
Xbit_r3_c180 bl_180 br_180 wl_3 vdd gnd cell_6t
Xbit_r4_c180 bl_180 br_180 wl_4 vdd gnd cell_6t
Xbit_r5_c180 bl_180 br_180 wl_5 vdd gnd cell_6t
Xbit_r6_c180 bl_180 br_180 wl_6 vdd gnd cell_6t
Xbit_r7_c180 bl_180 br_180 wl_7 vdd gnd cell_6t
Xbit_r8_c180 bl_180 br_180 wl_8 vdd gnd cell_6t
Xbit_r9_c180 bl_180 br_180 wl_9 vdd gnd cell_6t
Xbit_r10_c180 bl_180 br_180 wl_10 vdd gnd cell_6t
Xbit_r11_c180 bl_180 br_180 wl_11 vdd gnd cell_6t
Xbit_r12_c180 bl_180 br_180 wl_12 vdd gnd cell_6t
Xbit_r13_c180 bl_180 br_180 wl_13 vdd gnd cell_6t
Xbit_r14_c180 bl_180 br_180 wl_14 vdd gnd cell_6t
Xbit_r15_c180 bl_180 br_180 wl_15 vdd gnd cell_6t
Xbit_r16_c180 bl_180 br_180 wl_16 vdd gnd cell_6t
Xbit_r17_c180 bl_180 br_180 wl_17 vdd gnd cell_6t
Xbit_r18_c180 bl_180 br_180 wl_18 vdd gnd cell_6t
Xbit_r19_c180 bl_180 br_180 wl_19 vdd gnd cell_6t
Xbit_r20_c180 bl_180 br_180 wl_20 vdd gnd cell_6t
Xbit_r21_c180 bl_180 br_180 wl_21 vdd gnd cell_6t
Xbit_r22_c180 bl_180 br_180 wl_22 vdd gnd cell_6t
Xbit_r23_c180 bl_180 br_180 wl_23 vdd gnd cell_6t
Xbit_r24_c180 bl_180 br_180 wl_24 vdd gnd cell_6t
Xbit_r25_c180 bl_180 br_180 wl_25 vdd gnd cell_6t
Xbit_r26_c180 bl_180 br_180 wl_26 vdd gnd cell_6t
Xbit_r27_c180 bl_180 br_180 wl_27 vdd gnd cell_6t
Xbit_r28_c180 bl_180 br_180 wl_28 vdd gnd cell_6t
Xbit_r29_c180 bl_180 br_180 wl_29 vdd gnd cell_6t
Xbit_r30_c180 bl_180 br_180 wl_30 vdd gnd cell_6t
Xbit_r31_c180 bl_180 br_180 wl_31 vdd gnd cell_6t
Xbit_r32_c180 bl_180 br_180 wl_32 vdd gnd cell_6t
Xbit_r33_c180 bl_180 br_180 wl_33 vdd gnd cell_6t
Xbit_r34_c180 bl_180 br_180 wl_34 vdd gnd cell_6t
Xbit_r35_c180 bl_180 br_180 wl_35 vdd gnd cell_6t
Xbit_r36_c180 bl_180 br_180 wl_36 vdd gnd cell_6t
Xbit_r37_c180 bl_180 br_180 wl_37 vdd gnd cell_6t
Xbit_r38_c180 bl_180 br_180 wl_38 vdd gnd cell_6t
Xbit_r39_c180 bl_180 br_180 wl_39 vdd gnd cell_6t
Xbit_r40_c180 bl_180 br_180 wl_40 vdd gnd cell_6t
Xbit_r41_c180 bl_180 br_180 wl_41 vdd gnd cell_6t
Xbit_r42_c180 bl_180 br_180 wl_42 vdd gnd cell_6t
Xbit_r43_c180 bl_180 br_180 wl_43 vdd gnd cell_6t
Xbit_r44_c180 bl_180 br_180 wl_44 vdd gnd cell_6t
Xbit_r45_c180 bl_180 br_180 wl_45 vdd gnd cell_6t
Xbit_r46_c180 bl_180 br_180 wl_46 vdd gnd cell_6t
Xbit_r47_c180 bl_180 br_180 wl_47 vdd gnd cell_6t
Xbit_r48_c180 bl_180 br_180 wl_48 vdd gnd cell_6t
Xbit_r49_c180 bl_180 br_180 wl_49 vdd gnd cell_6t
Xbit_r50_c180 bl_180 br_180 wl_50 vdd gnd cell_6t
Xbit_r51_c180 bl_180 br_180 wl_51 vdd gnd cell_6t
Xbit_r52_c180 bl_180 br_180 wl_52 vdd gnd cell_6t
Xbit_r53_c180 bl_180 br_180 wl_53 vdd gnd cell_6t
Xbit_r54_c180 bl_180 br_180 wl_54 vdd gnd cell_6t
Xbit_r55_c180 bl_180 br_180 wl_55 vdd gnd cell_6t
Xbit_r56_c180 bl_180 br_180 wl_56 vdd gnd cell_6t
Xbit_r57_c180 bl_180 br_180 wl_57 vdd gnd cell_6t
Xbit_r58_c180 bl_180 br_180 wl_58 vdd gnd cell_6t
Xbit_r59_c180 bl_180 br_180 wl_59 vdd gnd cell_6t
Xbit_r60_c180 bl_180 br_180 wl_60 vdd gnd cell_6t
Xbit_r61_c180 bl_180 br_180 wl_61 vdd gnd cell_6t
Xbit_r62_c180 bl_180 br_180 wl_62 vdd gnd cell_6t
Xbit_r63_c180 bl_180 br_180 wl_63 vdd gnd cell_6t
Xbit_r64_c180 bl_180 br_180 wl_64 vdd gnd cell_6t
Xbit_r65_c180 bl_180 br_180 wl_65 vdd gnd cell_6t
Xbit_r66_c180 bl_180 br_180 wl_66 vdd gnd cell_6t
Xbit_r67_c180 bl_180 br_180 wl_67 vdd gnd cell_6t
Xbit_r68_c180 bl_180 br_180 wl_68 vdd gnd cell_6t
Xbit_r69_c180 bl_180 br_180 wl_69 vdd gnd cell_6t
Xbit_r70_c180 bl_180 br_180 wl_70 vdd gnd cell_6t
Xbit_r71_c180 bl_180 br_180 wl_71 vdd gnd cell_6t
Xbit_r72_c180 bl_180 br_180 wl_72 vdd gnd cell_6t
Xbit_r73_c180 bl_180 br_180 wl_73 vdd gnd cell_6t
Xbit_r74_c180 bl_180 br_180 wl_74 vdd gnd cell_6t
Xbit_r75_c180 bl_180 br_180 wl_75 vdd gnd cell_6t
Xbit_r76_c180 bl_180 br_180 wl_76 vdd gnd cell_6t
Xbit_r77_c180 bl_180 br_180 wl_77 vdd gnd cell_6t
Xbit_r78_c180 bl_180 br_180 wl_78 vdd gnd cell_6t
Xbit_r79_c180 bl_180 br_180 wl_79 vdd gnd cell_6t
Xbit_r80_c180 bl_180 br_180 wl_80 vdd gnd cell_6t
Xbit_r81_c180 bl_180 br_180 wl_81 vdd gnd cell_6t
Xbit_r82_c180 bl_180 br_180 wl_82 vdd gnd cell_6t
Xbit_r83_c180 bl_180 br_180 wl_83 vdd gnd cell_6t
Xbit_r84_c180 bl_180 br_180 wl_84 vdd gnd cell_6t
Xbit_r85_c180 bl_180 br_180 wl_85 vdd gnd cell_6t
Xbit_r86_c180 bl_180 br_180 wl_86 vdd gnd cell_6t
Xbit_r87_c180 bl_180 br_180 wl_87 vdd gnd cell_6t
Xbit_r88_c180 bl_180 br_180 wl_88 vdd gnd cell_6t
Xbit_r89_c180 bl_180 br_180 wl_89 vdd gnd cell_6t
Xbit_r90_c180 bl_180 br_180 wl_90 vdd gnd cell_6t
Xbit_r91_c180 bl_180 br_180 wl_91 vdd gnd cell_6t
Xbit_r92_c180 bl_180 br_180 wl_92 vdd gnd cell_6t
Xbit_r93_c180 bl_180 br_180 wl_93 vdd gnd cell_6t
Xbit_r94_c180 bl_180 br_180 wl_94 vdd gnd cell_6t
Xbit_r95_c180 bl_180 br_180 wl_95 vdd gnd cell_6t
Xbit_r96_c180 bl_180 br_180 wl_96 vdd gnd cell_6t
Xbit_r97_c180 bl_180 br_180 wl_97 vdd gnd cell_6t
Xbit_r98_c180 bl_180 br_180 wl_98 vdd gnd cell_6t
Xbit_r99_c180 bl_180 br_180 wl_99 vdd gnd cell_6t
Xbit_r100_c180 bl_180 br_180 wl_100 vdd gnd cell_6t
Xbit_r101_c180 bl_180 br_180 wl_101 vdd gnd cell_6t
Xbit_r102_c180 bl_180 br_180 wl_102 vdd gnd cell_6t
Xbit_r103_c180 bl_180 br_180 wl_103 vdd gnd cell_6t
Xbit_r104_c180 bl_180 br_180 wl_104 vdd gnd cell_6t
Xbit_r105_c180 bl_180 br_180 wl_105 vdd gnd cell_6t
Xbit_r106_c180 bl_180 br_180 wl_106 vdd gnd cell_6t
Xbit_r107_c180 bl_180 br_180 wl_107 vdd gnd cell_6t
Xbit_r108_c180 bl_180 br_180 wl_108 vdd gnd cell_6t
Xbit_r109_c180 bl_180 br_180 wl_109 vdd gnd cell_6t
Xbit_r110_c180 bl_180 br_180 wl_110 vdd gnd cell_6t
Xbit_r111_c180 bl_180 br_180 wl_111 vdd gnd cell_6t
Xbit_r112_c180 bl_180 br_180 wl_112 vdd gnd cell_6t
Xbit_r113_c180 bl_180 br_180 wl_113 vdd gnd cell_6t
Xbit_r114_c180 bl_180 br_180 wl_114 vdd gnd cell_6t
Xbit_r115_c180 bl_180 br_180 wl_115 vdd gnd cell_6t
Xbit_r116_c180 bl_180 br_180 wl_116 vdd gnd cell_6t
Xbit_r117_c180 bl_180 br_180 wl_117 vdd gnd cell_6t
Xbit_r118_c180 bl_180 br_180 wl_118 vdd gnd cell_6t
Xbit_r119_c180 bl_180 br_180 wl_119 vdd gnd cell_6t
Xbit_r120_c180 bl_180 br_180 wl_120 vdd gnd cell_6t
Xbit_r121_c180 bl_180 br_180 wl_121 vdd gnd cell_6t
Xbit_r122_c180 bl_180 br_180 wl_122 vdd gnd cell_6t
Xbit_r123_c180 bl_180 br_180 wl_123 vdd gnd cell_6t
Xbit_r124_c180 bl_180 br_180 wl_124 vdd gnd cell_6t
Xbit_r125_c180 bl_180 br_180 wl_125 vdd gnd cell_6t
Xbit_r126_c180 bl_180 br_180 wl_126 vdd gnd cell_6t
Xbit_r127_c180 bl_180 br_180 wl_127 vdd gnd cell_6t
Xbit_r128_c180 bl_180 br_180 wl_128 vdd gnd cell_6t
Xbit_r129_c180 bl_180 br_180 wl_129 vdd gnd cell_6t
Xbit_r130_c180 bl_180 br_180 wl_130 vdd gnd cell_6t
Xbit_r131_c180 bl_180 br_180 wl_131 vdd gnd cell_6t
Xbit_r132_c180 bl_180 br_180 wl_132 vdd gnd cell_6t
Xbit_r133_c180 bl_180 br_180 wl_133 vdd gnd cell_6t
Xbit_r134_c180 bl_180 br_180 wl_134 vdd gnd cell_6t
Xbit_r135_c180 bl_180 br_180 wl_135 vdd gnd cell_6t
Xbit_r136_c180 bl_180 br_180 wl_136 vdd gnd cell_6t
Xbit_r137_c180 bl_180 br_180 wl_137 vdd gnd cell_6t
Xbit_r138_c180 bl_180 br_180 wl_138 vdd gnd cell_6t
Xbit_r139_c180 bl_180 br_180 wl_139 vdd gnd cell_6t
Xbit_r140_c180 bl_180 br_180 wl_140 vdd gnd cell_6t
Xbit_r141_c180 bl_180 br_180 wl_141 vdd gnd cell_6t
Xbit_r142_c180 bl_180 br_180 wl_142 vdd gnd cell_6t
Xbit_r143_c180 bl_180 br_180 wl_143 vdd gnd cell_6t
Xbit_r144_c180 bl_180 br_180 wl_144 vdd gnd cell_6t
Xbit_r145_c180 bl_180 br_180 wl_145 vdd gnd cell_6t
Xbit_r146_c180 bl_180 br_180 wl_146 vdd gnd cell_6t
Xbit_r147_c180 bl_180 br_180 wl_147 vdd gnd cell_6t
Xbit_r148_c180 bl_180 br_180 wl_148 vdd gnd cell_6t
Xbit_r149_c180 bl_180 br_180 wl_149 vdd gnd cell_6t
Xbit_r150_c180 bl_180 br_180 wl_150 vdd gnd cell_6t
Xbit_r151_c180 bl_180 br_180 wl_151 vdd gnd cell_6t
Xbit_r152_c180 bl_180 br_180 wl_152 vdd gnd cell_6t
Xbit_r153_c180 bl_180 br_180 wl_153 vdd gnd cell_6t
Xbit_r154_c180 bl_180 br_180 wl_154 vdd gnd cell_6t
Xbit_r155_c180 bl_180 br_180 wl_155 vdd gnd cell_6t
Xbit_r156_c180 bl_180 br_180 wl_156 vdd gnd cell_6t
Xbit_r157_c180 bl_180 br_180 wl_157 vdd gnd cell_6t
Xbit_r158_c180 bl_180 br_180 wl_158 vdd gnd cell_6t
Xbit_r159_c180 bl_180 br_180 wl_159 vdd gnd cell_6t
Xbit_r160_c180 bl_180 br_180 wl_160 vdd gnd cell_6t
Xbit_r161_c180 bl_180 br_180 wl_161 vdd gnd cell_6t
Xbit_r162_c180 bl_180 br_180 wl_162 vdd gnd cell_6t
Xbit_r163_c180 bl_180 br_180 wl_163 vdd gnd cell_6t
Xbit_r164_c180 bl_180 br_180 wl_164 vdd gnd cell_6t
Xbit_r165_c180 bl_180 br_180 wl_165 vdd gnd cell_6t
Xbit_r166_c180 bl_180 br_180 wl_166 vdd gnd cell_6t
Xbit_r167_c180 bl_180 br_180 wl_167 vdd gnd cell_6t
Xbit_r168_c180 bl_180 br_180 wl_168 vdd gnd cell_6t
Xbit_r169_c180 bl_180 br_180 wl_169 vdd gnd cell_6t
Xbit_r170_c180 bl_180 br_180 wl_170 vdd gnd cell_6t
Xbit_r171_c180 bl_180 br_180 wl_171 vdd gnd cell_6t
Xbit_r172_c180 bl_180 br_180 wl_172 vdd gnd cell_6t
Xbit_r173_c180 bl_180 br_180 wl_173 vdd gnd cell_6t
Xbit_r174_c180 bl_180 br_180 wl_174 vdd gnd cell_6t
Xbit_r175_c180 bl_180 br_180 wl_175 vdd gnd cell_6t
Xbit_r176_c180 bl_180 br_180 wl_176 vdd gnd cell_6t
Xbit_r177_c180 bl_180 br_180 wl_177 vdd gnd cell_6t
Xbit_r178_c180 bl_180 br_180 wl_178 vdd gnd cell_6t
Xbit_r179_c180 bl_180 br_180 wl_179 vdd gnd cell_6t
Xbit_r180_c180 bl_180 br_180 wl_180 vdd gnd cell_6t
Xbit_r181_c180 bl_180 br_180 wl_181 vdd gnd cell_6t
Xbit_r182_c180 bl_180 br_180 wl_182 vdd gnd cell_6t
Xbit_r183_c180 bl_180 br_180 wl_183 vdd gnd cell_6t
Xbit_r184_c180 bl_180 br_180 wl_184 vdd gnd cell_6t
Xbit_r185_c180 bl_180 br_180 wl_185 vdd gnd cell_6t
Xbit_r186_c180 bl_180 br_180 wl_186 vdd gnd cell_6t
Xbit_r187_c180 bl_180 br_180 wl_187 vdd gnd cell_6t
Xbit_r188_c180 bl_180 br_180 wl_188 vdd gnd cell_6t
Xbit_r189_c180 bl_180 br_180 wl_189 vdd gnd cell_6t
Xbit_r190_c180 bl_180 br_180 wl_190 vdd gnd cell_6t
Xbit_r191_c180 bl_180 br_180 wl_191 vdd gnd cell_6t
Xbit_r192_c180 bl_180 br_180 wl_192 vdd gnd cell_6t
Xbit_r193_c180 bl_180 br_180 wl_193 vdd gnd cell_6t
Xbit_r194_c180 bl_180 br_180 wl_194 vdd gnd cell_6t
Xbit_r195_c180 bl_180 br_180 wl_195 vdd gnd cell_6t
Xbit_r196_c180 bl_180 br_180 wl_196 vdd gnd cell_6t
Xbit_r197_c180 bl_180 br_180 wl_197 vdd gnd cell_6t
Xbit_r198_c180 bl_180 br_180 wl_198 vdd gnd cell_6t
Xbit_r199_c180 bl_180 br_180 wl_199 vdd gnd cell_6t
Xbit_r200_c180 bl_180 br_180 wl_200 vdd gnd cell_6t
Xbit_r201_c180 bl_180 br_180 wl_201 vdd gnd cell_6t
Xbit_r202_c180 bl_180 br_180 wl_202 vdd gnd cell_6t
Xbit_r203_c180 bl_180 br_180 wl_203 vdd gnd cell_6t
Xbit_r204_c180 bl_180 br_180 wl_204 vdd gnd cell_6t
Xbit_r205_c180 bl_180 br_180 wl_205 vdd gnd cell_6t
Xbit_r206_c180 bl_180 br_180 wl_206 vdd gnd cell_6t
Xbit_r207_c180 bl_180 br_180 wl_207 vdd gnd cell_6t
Xbit_r208_c180 bl_180 br_180 wl_208 vdd gnd cell_6t
Xbit_r209_c180 bl_180 br_180 wl_209 vdd gnd cell_6t
Xbit_r210_c180 bl_180 br_180 wl_210 vdd gnd cell_6t
Xbit_r211_c180 bl_180 br_180 wl_211 vdd gnd cell_6t
Xbit_r212_c180 bl_180 br_180 wl_212 vdd gnd cell_6t
Xbit_r213_c180 bl_180 br_180 wl_213 vdd gnd cell_6t
Xbit_r214_c180 bl_180 br_180 wl_214 vdd gnd cell_6t
Xbit_r215_c180 bl_180 br_180 wl_215 vdd gnd cell_6t
Xbit_r216_c180 bl_180 br_180 wl_216 vdd gnd cell_6t
Xbit_r217_c180 bl_180 br_180 wl_217 vdd gnd cell_6t
Xbit_r218_c180 bl_180 br_180 wl_218 vdd gnd cell_6t
Xbit_r219_c180 bl_180 br_180 wl_219 vdd gnd cell_6t
Xbit_r220_c180 bl_180 br_180 wl_220 vdd gnd cell_6t
Xbit_r221_c180 bl_180 br_180 wl_221 vdd gnd cell_6t
Xbit_r222_c180 bl_180 br_180 wl_222 vdd gnd cell_6t
Xbit_r223_c180 bl_180 br_180 wl_223 vdd gnd cell_6t
Xbit_r224_c180 bl_180 br_180 wl_224 vdd gnd cell_6t
Xbit_r225_c180 bl_180 br_180 wl_225 vdd gnd cell_6t
Xbit_r226_c180 bl_180 br_180 wl_226 vdd gnd cell_6t
Xbit_r227_c180 bl_180 br_180 wl_227 vdd gnd cell_6t
Xbit_r228_c180 bl_180 br_180 wl_228 vdd gnd cell_6t
Xbit_r229_c180 bl_180 br_180 wl_229 vdd gnd cell_6t
Xbit_r230_c180 bl_180 br_180 wl_230 vdd gnd cell_6t
Xbit_r231_c180 bl_180 br_180 wl_231 vdd gnd cell_6t
Xbit_r232_c180 bl_180 br_180 wl_232 vdd gnd cell_6t
Xbit_r233_c180 bl_180 br_180 wl_233 vdd gnd cell_6t
Xbit_r234_c180 bl_180 br_180 wl_234 vdd gnd cell_6t
Xbit_r235_c180 bl_180 br_180 wl_235 vdd gnd cell_6t
Xbit_r236_c180 bl_180 br_180 wl_236 vdd gnd cell_6t
Xbit_r237_c180 bl_180 br_180 wl_237 vdd gnd cell_6t
Xbit_r238_c180 bl_180 br_180 wl_238 vdd gnd cell_6t
Xbit_r239_c180 bl_180 br_180 wl_239 vdd gnd cell_6t
Xbit_r240_c180 bl_180 br_180 wl_240 vdd gnd cell_6t
Xbit_r241_c180 bl_180 br_180 wl_241 vdd gnd cell_6t
Xbit_r242_c180 bl_180 br_180 wl_242 vdd gnd cell_6t
Xbit_r243_c180 bl_180 br_180 wl_243 vdd gnd cell_6t
Xbit_r244_c180 bl_180 br_180 wl_244 vdd gnd cell_6t
Xbit_r245_c180 bl_180 br_180 wl_245 vdd gnd cell_6t
Xbit_r246_c180 bl_180 br_180 wl_246 vdd gnd cell_6t
Xbit_r247_c180 bl_180 br_180 wl_247 vdd gnd cell_6t
Xbit_r248_c180 bl_180 br_180 wl_248 vdd gnd cell_6t
Xbit_r249_c180 bl_180 br_180 wl_249 vdd gnd cell_6t
Xbit_r250_c180 bl_180 br_180 wl_250 vdd gnd cell_6t
Xbit_r251_c180 bl_180 br_180 wl_251 vdd gnd cell_6t
Xbit_r252_c180 bl_180 br_180 wl_252 vdd gnd cell_6t
Xbit_r253_c180 bl_180 br_180 wl_253 vdd gnd cell_6t
Xbit_r254_c180 bl_180 br_180 wl_254 vdd gnd cell_6t
Xbit_r255_c180 bl_180 br_180 wl_255 vdd gnd cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd cell_6t
Xbit_r1_c181 bl_181 br_181 wl_1 vdd gnd cell_6t
Xbit_r2_c181 bl_181 br_181 wl_2 vdd gnd cell_6t
Xbit_r3_c181 bl_181 br_181 wl_3 vdd gnd cell_6t
Xbit_r4_c181 bl_181 br_181 wl_4 vdd gnd cell_6t
Xbit_r5_c181 bl_181 br_181 wl_5 vdd gnd cell_6t
Xbit_r6_c181 bl_181 br_181 wl_6 vdd gnd cell_6t
Xbit_r7_c181 bl_181 br_181 wl_7 vdd gnd cell_6t
Xbit_r8_c181 bl_181 br_181 wl_8 vdd gnd cell_6t
Xbit_r9_c181 bl_181 br_181 wl_9 vdd gnd cell_6t
Xbit_r10_c181 bl_181 br_181 wl_10 vdd gnd cell_6t
Xbit_r11_c181 bl_181 br_181 wl_11 vdd gnd cell_6t
Xbit_r12_c181 bl_181 br_181 wl_12 vdd gnd cell_6t
Xbit_r13_c181 bl_181 br_181 wl_13 vdd gnd cell_6t
Xbit_r14_c181 bl_181 br_181 wl_14 vdd gnd cell_6t
Xbit_r15_c181 bl_181 br_181 wl_15 vdd gnd cell_6t
Xbit_r16_c181 bl_181 br_181 wl_16 vdd gnd cell_6t
Xbit_r17_c181 bl_181 br_181 wl_17 vdd gnd cell_6t
Xbit_r18_c181 bl_181 br_181 wl_18 vdd gnd cell_6t
Xbit_r19_c181 bl_181 br_181 wl_19 vdd gnd cell_6t
Xbit_r20_c181 bl_181 br_181 wl_20 vdd gnd cell_6t
Xbit_r21_c181 bl_181 br_181 wl_21 vdd gnd cell_6t
Xbit_r22_c181 bl_181 br_181 wl_22 vdd gnd cell_6t
Xbit_r23_c181 bl_181 br_181 wl_23 vdd gnd cell_6t
Xbit_r24_c181 bl_181 br_181 wl_24 vdd gnd cell_6t
Xbit_r25_c181 bl_181 br_181 wl_25 vdd gnd cell_6t
Xbit_r26_c181 bl_181 br_181 wl_26 vdd gnd cell_6t
Xbit_r27_c181 bl_181 br_181 wl_27 vdd gnd cell_6t
Xbit_r28_c181 bl_181 br_181 wl_28 vdd gnd cell_6t
Xbit_r29_c181 bl_181 br_181 wl_29 vdd gnd cell_6t
Xbit_r30_c181 bl_181 br_181 wl_30 vdd gnd cell_6t
Xbit_r31_c181 bl_181 br_181 wl_31 vdd gnd cell_6t
Xbit_r32_c181 bl_181 br_181 wl_32 vdd gnd cell_6t
Xbit_r33_c181 bl_181 br_181 wl_33 vdd gnd cell_6t
Xbit_r34_c181 bl_181 br_181 wl_34 vdd gnd cell_6t
Xbit_r35_c181 bl_181 br_181 wl_35 vdd gnd cell_6t
Xbit_r36_c181 bl_181 br_181 wl_36 vdd gnd cell_6t
Xbit_r37_c181 bl_181 br_181 wl_37 vdd gnd cell_6t
Xbit_r38_c181 bl_181 br_181 wl_38 vdd gnd cell_6t
Xbit_r39_c181 bl_181 br_181 wl_39 vdd gnd cell_6t
Xbit_r40_c181 bl_181 br_181 wl_40 vdd gnd cell_6t
Xbit_r41_c181 bl_181 br_181 wl_41 vdd gnd cell_6t
Xbit_r42_c181 bl_181 br_181 wl_42 vdd gnd cell_6t
Xbit_r43_c181 bl_181 br_181 wl_43 vdd gnd cell_6t
Xbit_r44_c181 bl_181 br_181 wl_44 vdd gnd cell_6t
Xbit_r45_c181 bl_181 br_181 wl_45 vdd gnd cell_6t
Xbit_r46_c181 bl_181 br_181 wl_46 vdd gnd cell_6t
Xbit_r47_c181 bl_181 br_181 wl_47 vdd gnd cell_6t
Xbit_r48_c181 bl_181 br_181 wl_48 vdd gnd cell_6t
Xbit_r49_c181 bl_181 br_181 wl_49 vdd gnd cell_6t
Xbit_r50_c181 bl_181 br_181 wl_50 vdd gnd cell_6t
Xbit_r51_c181 bl_181 br_181 wl_51 vdd gnd cell_6t
Xbit_r52_c181 bl_181 br_181 wl_52 vdd gnd cell_6t
Xbit_r53_c181 bl_181 br_181 wl_53 vdd gnd cell_6t
Xbit_r54_c181 bl_181 br_181 wl_54 vdd gnd cell_6t
Xbit_r55_c181 bl_181 br_181 wl_55 vdd gnd cell_6t
Xbit_r56_c181 bl_181 br_181 wl_56 vdd gnd cell_6t
Xbit_r57_c181 bl_181 br_181 wl_57 vdd gnd cell_6t
Xbit_r58_c181 bl_181 br_181 wl_58 vdd gnd cell_6t
Xbit_r59_c181 bl_181 br_181 wl_59 vdd gnd cell_6t
Xbit_r60_c181 bl_181 br_181 wl_60 vdd gnd cell_6t
Xbit_r61_c181 bl_181 br_181 wl_61 vdd gnd cell_6t
Xbit_r62_c181 bl_181 br_181 wl_62 vdd gnd cell_6t
Xbit_r63_c181 bl_181 br_181 wl_63 vdd gnd cell_6t
Xbit_r64_c181 bl_181 br_181 wl_64 vdd gnd cell_6t
Xbit_r65_c181 bl_181 br_181 wl_65 vdd gnd cell_6t
Xbit_r66_c181 bl_181 br_181 wl_66 vdd gnd cell_6t
Xbit_r67_c181 bl_181 br_181 wl_67 vdd gnd cell_6t
Xbit_r68_c181 bl_181 br_181 wl_68 vdd gnd cell_6t
Xbit_r69_c181 bl_181 br_181 wl_69 vdd gnd cell_6t
Xbit_r70_c181 bl_181 br_181 wl_70 vdd gnd cell_6t
Xbit_r71_c181 bl_181 br_181 wl_71 vdd gnd cell_6t
Xbit_r72_c181 bl_181 br_181 wl_72 vdd gnd cell_6t
Xbit_r73_c181 bl_181 br_181 wl_73 vdd gnd cell_6t
Xbit_r74_c181 bl_181 br_181 wl_74 vdd gnd cell_6t
Xbit_r75_c181 bl_181 br_181 wl_75 vdd gnd cell_6t
Xbit_r76_c181 bl_181 br_181 wl_76 vdd gnd cell_6t
Xbit_r77_c181 bl_181 br_181 wl_77 vdd gnd cell_6t
Xbit_r78_c181 bl_181 br_181 wl_78 vdd gnd cell_6t
Xbit_r79_c181 bl_181 br_181 wl_79 vdd gnd cell_6t
Xbit_r80_c181 bl_181 br_181 wl_80 vdd gnd cell_6t
Xbit_r81_c181 bl_181 br_181 wl_81 vdd gnd cell_6t
Xbit_r82_c181 bl_181 br_181 wl_82 vdd gnd cell_6t
Xbit_r83_c181 bl_181 br_181 wl_83 vdd gnd cell_6t
Xbit_r84_c181 bl_181 br_181 wl_84 vdd gnd cell_6t
Xbit_r85_c181 bl_181 br_181 wl_85 vdd gnd cell_6t
Xbit_r86_c181 bl_181 br_181 wl_86 vdd gnd cell_6t
Xbit_r87_c181 bl_181 br_181 wl_87 vdd gnd cell_6t
Xbit_r88_c181 bl_181 br_181 wl_88 vdd gnd cell_6t
Xbit_r89_c181 bl_181 br_181 wl_89 vdd gnd cell_6t
Xbit_r90_c181 bl_181 br_181 wl_90 vdd gnd cell_6t
Xbit_r91_c181 bl_181 br_181 wl_91 vdd gnd cell_6t
Xbit_r92_c181 bl_181 br_181 wl_92 vdd gnd cell_6t
Xbit_r93_c181 bl_181 br_181 wl_93 vdd gnd cell_6t
Xbit_r94_c181 bl_181 br_181 wl_94 vdd gnd cell_6t
Xbit_r95_c181 bl_181 br_181 wl_95 vdd gnd cell_6t
Xbit_r96_c181 bl_181 br_181 wl_96 vdd gnd cell_6t
Xbit_r97_c181 bl_181 br_181 wl_97 vdd gnd cell_6t
Xbit_r98_c181 bl_181 br_181 wl_98 vdd gnd cell_6t
Xbit_r99_c181 bl_181 br_181 wl_99 vdd gnd cell_6t
Xbit_r100_c181 bl_181 br_181 wl_100 vdd gnd cell_6t
Xbit_r101_c181 bl_181 br_181 wl_101 vdd gnd cell_6t
Xbit_r102_c181 bl_181 br_181 wl_102 vdd gnd cell_6t
Xbit_r103_c181 bl_181 br_181 wl_103 vdd gnd cell_6t
Xbit_r104_c181 bl_181 br_181 wl_104 vdd gnd cell_6t
Xbit_r105_c181 bl_181 br_181 wl_105 vdd gnd cell_6t
Xbit_r106_c181 bl_181 br_181 wl_106 vdd gnd cell_6t
Xbit_r107_c181 bl_181 br_181 wl_107 vdd gnd cell_6t
Xbit_r108_c181 bl_181 br_181 wl_108 vdd gnd cell_6t
Xbit_r109_c181 bl_181 br_181 wl_109 vdd gnd cell_6t
Xbit_r110_c181 bl_181 br_181 wl_110 vdd gnd cell_6t
Xbit_r111_c181 bl_181 br_181 wl_111 vdd gnd cell_6t
Xbit_r112_c181 bl_181 br_181 wl_112 vdd gnd cell_6t
Xbit_r113_c181 bl_181 br_181 wl_113 vdd gnd cell_6t
Xbit_r114_c181 bl_181 br_181 wl_114 vdd gnd cell_6t
Xbit_r115_c181 bl_181 br_181 wl_115 vdd gnd cell_6t
Xbit_r116_c181 bl_181 br_181 wl_116 vdd gnd cell_6t
Xbit_r117_c181 bl_181 br_181 wl_117 vdd gnd cell_6t
Xbit_r118_c181 bl_181 br_181 wl_118 vdd gnd cell_6t
Xbit_r119_c181 bl_181 br_181 wl_119 vdd gnd cell_6t
Xbit_r120_c181 bl_181 br_181 wl_120 vdd gnd cell_6t
Xbit_r121_c181 bl_181 br_181 wl_121 vdd gnd cell_6t
Xbit_r122_c181 bl_181 br_181 wl_122 vdd gnd cell_6t
Xbit_r123_c181 bl_181 br_181 wl_123 vdd gnd cell_6t
Xbit_r124_c181 bl_181 br_181 wl_124 vdd gnd cell_6t
Xbit_r125_c181 bl_181 br_181 wl_125 vdd gnd cell_6t
Xbit_r126_c181 bl_181 br_181 wl_126 vdd gnd cell_6t
Xbit_r127_c181 bl_181 br_181 wl_127 vdd gnd cell_6t
Xbit_r128_c181 bl_181 br_181 wl_128 vdd gnd cell_6t
Xbit_r129_c181 bl_181 br_181 wl_129 vdd gnd cell_6t
Xbit_r130_c181 bl_181 br_181 wl_130 vdd gnd cell_6t
Xbit_r131_c181 bl_181 br_181 wl_131 vdd gnd cell_6t
Xbit_r132_c181 bl_181 br_181 wl_132 vdd gnd cell_6t
Xbit_r133_c181 bl_181 br_181 wl_133 vdd gnd cell_6t
Xbit_r134_c181 bl_181 br_181 wl_134 vdd gnd cell_6t
Xbit_r135_c181 bl_181 br_181 wl_135 vdd gnd cell_6t
Xbit_r136_c181 bl_181 br_181 wl_136 vdd gnd cell_6t
Xbit_r137_c181 bl_181 br_181 wl_137 vdd gnd cell_6t
Xbit_r138_c181 bl_181 br_181 wl_138 vdd gnd cell_6t
Xbit_r139_c181 bl_181 br_181 wl_139 vdd gnd cell_6t
Xbit_r140_c181 bl_181 br_181 wl_140 vdd gnd cell_6t
Xbit_r141_c181 bl_181 br_181 wl_141 vdd gnd cell_6t
Xbit_r142_c181 bl_181 br_181 wl_142 vdd gnd cell_6t
Xbit_r143_c181 bl_181 br_181 wl_143 vdd gnd cell_6t
Xbit_r144_c181 bl_181 br_181 wl_144 vdd gnd cell_6t
Xbit_r145_c181 bl_181 br_181 wl_145 vdd gnd cell_6t
Xbit_r146_c181 bl_181 br_181 wl_146 vdd gnd cell_6t
Xbit_r147_c181 bl_181 br_181 wl_147 vdd gnd cell_6t
Xbit_r148_c181 bl_181 br_181 wl_148 vdd gnd cell_6t
Xbit_r149_c181 bl_181 br_181 wl_149 vdd gnd cell_6t
Xbit_r150_c181 bl_181 br_181 wl_150 vdd gnd cell_6t
Xbit_r151_c181 bl_181 br_181 wl_151 vdd gnd cell_6t
Xbit_r152_c181 bl_181 br_181 wl_152 vdd gnd cell_6t
Xbit_r153_c181 bl_181 br_181 wl_153 vdd gnd cell_6t
Xbit_r154_c181 bl_181 br_181 wl_154 vdd gnd cell_6t
Xbit_r155_c181 bl_181 br_181 wl_155 vdd gnd cell_6t
Xbit_r156_c181 bl_181 br_181 wl_156 vdd gnd cell_6t
Xbit_r157_c181 bl_181 br_181 wl_157 vdd gnd cell_6t
Xbit_r158_c181 bl_181 br_181 wl_158 vdd gnd cell_6t
Xbit_r159_c181 bl_181 br_181 wl_159 vdd gnd cell_6t
Xbit_r160_c181 bl_181 br_181 wl_160 vdd gnd cell_6t
Xbit_r161_c181 bl_181 br_181 wl_161 vdd gnd cell_6t
Xbit_r162_c181 bl_181 br_181 wl_162 vdd gnd cell_6t
Xbit_r163_c181 bl_181 br_181 wl_163 vdd gnd cell_6t
Xbit_r164_c181 bl_181 br_181 wl_164 vdd gnd cell_6t
Xbit_r165_c181 bl_181 br_181 wl_165 vdd gnd cell_6t
Xbit_r166_c181 bl_181 br_181 wl_166 vdd gnd cell_6t
Xbit_r167_c181 bl_181 br_181 wl_167 vdd gnd cell_6t
Xbit_r168_c181 bl_181 br_181 wl_168 vdd gnd cell_6t
Xbit_r169_c181 bl_181 br_181 wl_169 vdd gnd cell_6t
Xbit_r170_c181 bl_181 br_181 wl_170 vdd gnd cell_6t
Xbit_r171_c181 bl_181 br_181 wl_171 vdd gnd cell_6t
Xbit_r172_c181 bl_181 br_181 wl_172 vdd gnd cell_6t
Xbit_r173_c181 bl_181 br_181 wl_173 vdd gnd cell_6t
Xbit_r174_c181 bl_181 br_181 wl_174 vdd gnd cell_6t
Xbit_r175_c181 bl_181 br_181 wl_175 vdd gnd cell_6t
Xbit_r176_c181 bl_181 br_181 wl_176 vdd gnd cell_6t
Xbit_r177_c181 bl_181 br_181 wl_177 vdd gnd cell_6t
Xbit_r178_c181 bl_181 br_181 wl_178 vdd gnd cell_6t
Xbit_r179_c181 bl_181 br_181 wl_179 vdd gnd cell_6t
Xbit_r180_c181 bl_181 br_181 wl_180 vdd gnd cell_6t
Xbit_r181_c181 bl_181 br_181 wl_181 vdd gnd cell_6t
Xbit_r182_c181 bl_181 br_181 wl_182 vdd gnd cell_6t
Xbit_r183_c181 bl_181 br_181 wl_183 vdd gnd cell_6t
Xbit_r184_c181 bl_181 br_181 wl_184 vdd gnd cell_6t
Xbit_r185_c181 bl_181 br_181 wl_185 vdd gnd cell_6t
Xbit_r186_c181 bl_181 br_181 wl_186 vdd gnd cell_6t
Xbit_r187_c181 bl_181 br_181 wl_187 vdd gnd cell_6t
Xbit_r188_c181 bl_181 br_181 wl_188 vdd gnd cell_6t
Xbit_r189_c181 bl_181 br_181 wl_189 vdd gnd cell_6t
Xbit_r190_c181 bl_181 br_181 wl_190 vdd gnd cell_6t
Xbit_r191_c181 bl_181 br_181 wl_191 vdd gnd cell_6t
Xbit_r192_c181 bl_181 br_181 wl_192 vdd gnd cell_6t
Xbit_r193_c181 bl_181 br_181 wl_193 vdd gnd cell_6t
Xbit_r194_c181 bl_181 br_181 wl_194 vdd gnd cell_6t
Xbit_r195_c181 bl_181 br_181 wl_195 vdd gnd cell_6t
Xbit_r196_c181 bl_181 br_181 wl_196 vdd gnd cell_6t
Xbit_r197_c181 bl_181 br_181 wl_197 vdd gnd cell_6t
Xbit_r198_c181 bl_181 br_181 wl_198 vdd gnd cell_6t
Xbit_r199_c181 bl_181 br_181 wl_199 vdd gnd cell_6t
Xbit_r200_c181 bl_181 br_181 wl_200 vdd gnd cell_6t
Xbit_r201_c181 bl_181 br_181 wl_201 vdd gnd cell_6t
Xbit_r202_c181 bl_181 br_181 wl_202 vdd gnd cell_6t
Xbit_r203_c181 bl_181 br_181 wl_203 vdd gnd cell_6t
Xbit_r204_c181 bl_181 br_181 wl_204 vdd gnd cell_6t
Xbit_r205_c181 bl_181 br_181 wl_205 vdd gnd cell_6t
Xbit_r206_c181 bl_181 br_181 wl_206 vdd gnd cell_6t
Xbit_r207_c181 bl_181 br_181 wl_207 vdd gnd cell_6t
Xbit_r208_c181 bl_181 br_181 wl_208 vdd gnd cell_6t
Xbit_r209_c181 bl_181 br_181 wl_209 vdd gnd cell_6t
Xbit_r210_c181 bl_181 br_181 wl_210 vdd gnd cell_6t
Xbit_r211_c181 bl_181 br_181 wl_211 vdd gnd cell_6t
Xbit_r212_c181 bl_181 br_181 wl_212 vdd gnd cell_6t
Xbit_r213_c181 bl_181 br_181 wl_213 vdd gnd cell_6t
Xbit_r214_c181 bl_181 br_181 wl_214 vdd gnd cell_6t
Xbit_r215_c181 bl_181 br_181 wl_215 vdd gnd cell_6t
Xbit_r216_c181 bl_181 br_181 wl_216 vdd gnd cell_6t
Xbit_r217_c181 bl_181 br_181 wl_217 vdd gnd cell_6t
Xbit_r218_c181 bl_181 br_181 wl_218 vdd gnd cell_6t
Xbit_r219_c181 bl_181 br_181 wl_219 vdd gnd cell_6t
Xbit_r220_c181 bl_181 br_181 wl_220 vdd gnd cell_6t
Xbit_r221_c181 bl_181 br_181 wl_221 vdd gnd cell_6t
Xbit_r222_c181 bl_181 br_181 wl_222 vdd gnd cell_6t
Xbit_r223_c181 bl_181 br_181 wl_223 vdd gnd cell_6t
Xbit_r224_c181 bl_181 br_181 wl_224 vdd gnd cell_6t
Xbit_r225_c181 bl_181 br_181 wl_225 vdd gnd cell_6t
Xbit_r226_c181 bl_181 br_181 wl_226 vdd gnd cell_6t
Xbit_r227_c181 bl_181 br_181 wl_227 vdd gnd cell_6t
Xbit_r228_c181 bl_181 br_181 wl_228 vdd gnd cell_6t
Xbit_r229_c181 bl_181 br_181 wl_229 vdd gnd cell_6t
Xbit_r230_c181 bl_181 br_181 wl_230 vdd gnd cell_6t
Xbit_r231_c181 bl_181 br_181 wl_231 vdd gnd cell_6t
Xbit_r232_c181 bl_181 br_181 wl_232 vdd gnd cell_6t
Xbit_r233_c181 bl_181 br_181 wl_233 vdd gnd cell_6t
Xbit_r234_c181 bl_181 br_181 wl_234 vdd gnd cell_6t
Xbit_r235_c181 bl_181 br_181 wl_235 vdd gnd cell_6t
Xbit_r236_c181 bl_181 br_181 wl_236 vdd gnd cell_6t
Xbit_r237_c181 bl_181 br_181 wl_237 vdd gnd cell_6t
Xbit_r238_c181 bl_181 br_181 wl_238 vdd gnd cell_6t
Xbit_r239_c181 bl_181 br_181 wl_239 vdd gnd cell_6t
Xbit_r240_c181 bl_181 br_181 wl_240 vdd gnd cell_6t
Xbit_r241_c181 bl_181 br_181 wl_241 vdd gnd cell_6t
Xbit_r242_c181 bl_181 br_181 wl_242 vdd gnd cell_6t
Xbit_r243_c181 bl_181 br_181 wl_243 vdd gnd cell_6t
Xbit_r244_c181 bl_181 br_181 wl_244 vdd gnd cell_6t
Xbit_r245_c181 bl_181 br_181 wl_245 vdd gnd cell_6t
Xbit_r246_c181 bl_181 br_181 wl_246 vdd gnd cell_6t
Xbit_r247_c181 bl_181 br_181 wl_247 vdd gnd cell_6t
Xbit_r248_c181 bl_181 br_181 wl_248 vdd gnd cell_6t
Xbit_r249_c181 bl_181 br_181 wl_249 vdd gnd cell_6t
Xbit_r250_c181 bl_181 br_181 wl_250 vdd gnd cell_6t
Xbit_r251_c181 bl_181 br_181 wl_251 vdd gnd cell_6t
Xbit_r252_c181 bl_181 br_181 wl_252 vdd gnd cell_6t
Xbit_r253_c181 bl_181 br_181 wl_253 vdd gnd cell_6t
Xbit_r254_c181 bl_181 br_181 wl_254 vdd gnd cell_6t
Xbit_r255_c181 bl_181 br_181 wl_255 vdd gnd cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd cell_6t
Xbit_r1_c182 bl_182 br_182 wl_1 vdd gnd cell_6t
Xbit_r2_c182 bl_182 br_182 wl_2 vdd gnd cell_6t
Xbit_r3_c182 bl_182 br_182 wl_3 vdd gnd cell_6t
Xbit_r4_c182 bl_182 br_182 wl_4 vdd gnd cell_6t
Xbit_r5_c182 bl_182 br_182 wl_5 vdd gnd cell_6t
Xbit_r6_c182 bl_182 br_182 wl_6 vdd gnd cell_6t
Xbit_r7_c182 bl_182 br_182 wl_7 vdd gnd cell_6t
Xbit_r8_c182 bl_182 br_182 wl_8 vdd gnd cell_6t
Xbit_r9_c182 bl_182 br_182 wl_9 vdd gnd cell_6t
Xbit_r10_c182 bl_182 br_182 wl_10 vdd gnd cell_6t
Xbit_r11_c182 bl_182 br_182 wl_11 vdd gnd cell_6t
Xbit_r12_c182 bl_182 br_182 wl_12 vdd gnd cell_6t
Xbit_r13_c182 bl_182 br_182 wl_13 vdd gnd cell_6t
Xbit_r14_c182 bl_182 br_182 wl_14 vdd gnd cell_6t
Xbit_r15_c182 bl_182 br_182 wl_15 vdd gnd cell_6t
Xbit_r16_c182 bl_182 br_182 wl_16 vdd gnd cell_6t
Xbit_r17_c182 bl_182 br_182 wl_17 vdd gnd cell_6t
Xbit_r18_c182 bl_182 br_182 wl_18 vdd gnd cell_6t
Xbit_r19_c182 bl_182 br_182 wl_19 vdd gnd cell_6t
Xbit_r20_c182 bl_182 br_182 wl_20 vdd gnd cell_6t
Xbit_r21_c182 bl_182 br_182 wl_21 vdd gnd cell_6t
Xbit_r22_c182 bl_182 br_182 wl_22 vdd gnd cell_6t
Xbit_r23_c182 bl_182 br_182 wl_23 vdd gnd cell_6t
Xbit_r24_c182 bl_182 br_182 wl_24 vdd gnd cell_6t
Xbit_r25_c182 bl_182 br_182 wl_25 vdd gnd cell_6t
Xbit_r26_c182 bl_182 br_182 wl_26 vdd gnd cell_6t
Xbit_r27_c182 bl_182 br_182 wl_27 vdd gnd cell_6t
Xbit_r28_c182 bl_182 br_182 wl_28 vdd gnd cell_6t
Xbit_r29_c182 bl_182 br_182 wl_29 vdd gnd cell_6t
Xbit_r30_c182 bl_182 br_182 wl_30 vdd gnd cell_6t
Xbit_r31_c182 bl_182 br_182 wl_31 vdd gnd cell_6t
Xbit_r32_c182 bl_182 br_182 wl_32 vdd gnd cell_6t
Xbit_r33_c182 bl_182 br_182 wl_33 vdd gnd cell_6t
Xbit_r34_c182 bl_182 br_182 wl_34 vdd gnd cell_6t
Xbit_r35_c182 bl_182 br_182 wl_35 vdd gnd cell_6t
Xbit_r36_c182 bl_182 br_182 wl_36 vdd gnd cell_6t
Xbit_r37_c182 bl_182 br_182 wl_37 vdd gnd cell_6t
Xbit_r38_c182 bl_182 br_182 wl_38 vdd gnd cell_6t
Xbit_r39_c182 bl_182 br_182 wl_39 vdd gnd cell_6t
Xbit_r40_c182 bl_182 br_182 wl_40 vdd gnd cell_6t
Xbit_r41_c182 bl_182 br_182 wl_41 vdd gnd cell_6t
Xbit_r42_c182 bl_182 br_182 wl_42 vdd gnd cell_6t
Xbit_r43_c182 bl_182 br_182 wl_43 vdd gnd cell_6t
Xbit_r44_c182 bl_182 br_182 wl_44 vdd gnd cell_6t
Xbit_r45_c182 bl_182 br_182 wl_45 vdd gnd cell_6t
Xbit_r46_c182 bl_182 br_182 wl_46 vdd gnd cell_6t
Xbit_r47_c182 bl_182 br_182 wl_47 vdd gnd cell_6t
Xbit_r48_c182 bl_182 br_182 wl_48 vdd gnd cell_6t
Xbit_r49_c182 bl_182 br_182 wl_49 vdd gnd cell_6t
Xbit_r50_c182 bl_182 br_182 wl_50 vdd gnd cell_6t
Xbit_r51_c182 bl_182 br_182 wl_51 vdd gnd cell_6t
Xbit_r52_c182 bl_182 br_182 wl_52 vdd gnd cell_6t
Xbit_r53_c182 bl_182 br_182 wl_53 vdd gnd cell_6t
Xbit_r54_c182 bl_182 br_182 wl_54 vdd gnd cell_6t
Xbit_r55_c182 bl_182 br_182 wl_55 vdd gnd cell_6t
Xbit_r56_c182 bl_182 br_182 wl_56 vdd gnd cell_6t
Xbit_r57_c182 bl_182 br_182 wl_57 vdd gnd cell_6t
Xbit_r58_c182 bl_182 br_182 wl_58 vdd gnd cell_6t
Xbit_r59_c182 bl_182 br_182 wl_59 vdd gnd cell_6t
Xbit_r60_c182 bl_182 br_182 wl_60 vdd gnd cell_6t
Xbit_r61_c182 bl_182 br_182 wl_61 vdd gnd cell_6t
Xbit_r62_c182 bl_182 br_182 wl_62 vdd gnd cell_6t
Xbit_r63_c182 bl_182 br_182 wl_63 vdd gnd cell_6t
Xbit_r64_c182 bl_182 br_182 wl_64 vdd gnd cell_6t
Xbit_r65_c182 bl_182 br_182 wl_65 vdd gnd cell_6t
Xbit_r66_c182 bl_182 br_182 wl_66 vdd gnd cell_6t
Xbit_r67_c182 bl_182 br_182 wl_67 vdd gnd cell_6t
Xbit_r68_c182 bl_182 br_182 wl_68 vdd gnd cell_6t
Xbit_r69_c182 bl_182 br_182 wl_69 vdd gnd cell_6t
Xbit_r70_c182 bl_182 br_182 wl_70 vdd gnd cell_6t
Xbit_r71_c182 bl_182 br_182 wl_71 vdd gnd cell_6t
Xbit_r72_c182 bl_182 br_182 wl_72 vdd gnd cell_6t
Xbit_r73_c182 bl_182 br_182 wl_73 vdd gnd cell_6t
Xbit_r74_c182 bl_182 br_182 wl_74 vdd gnd cell_6t
Xbit_r75_c182 bl_182 br_182 wl_75 vdd gnd cell_6t
Xbit_r76_c182 bl_182 br_182 wl_76 vdd gnd cell_6t
Xbit_r77_c182 bl_182 br_182 wl_77 vdd gnd cell_6t
Xbit_r78_c182 bl_182 br_182 wl_78 vdd gnd cell_6t
Xbit_r79_c182 bl_182 br_182 wl_79 vdd gnd cell_6t
Xbit_r80_c182 bl_182 br_182 wl_80 vdd gnd cell_6t
Xbit_r81_c182 bl_182 br_182 wl_81 vdd gnd cell_6t
Xbit_r82_c182 bl_182 br_182 wl_82 vdd gnd cell_6t
Xbit_r83_c182 bl_182 br_182 wl_83 vdd gnd cell_6t
Xbit_r84_c182 bl_182 br_182 wl_84 vdd gnd cell_6t
Xbit_r85_c182 bl_182 br_182 wl_85 vdd gnd cell_6t
Xbit_r86_c182 bl_182 br_182 wl_86 vdd gnd cell_6t
Xbit_r87_c182 bl_182 br_182 wl_87 vdd gnd cell_6t
Xbit_r88_c182 bl_182 br_182 wl_88 vdd gnd cell_6t
Xbit_r89_c182 bl_182 br_182 wl_89 vdd gnd cell_6t
Xbit_r90_c182 bl_182 br_182 wl_90 vdd gnd cell_6t
Xbit_r91_c182 bl_182 br_182 wl_91 vdd gnd cell_6t
Xbit_r92_c182 bl_182 br_182 wl_92 vdd gnd cell_6t
Xbit_r93_c182 bl_182 br_182 wl_93 vdd gnd cell_6t
Xbit_r94_c182 bl_182 br_182 wl_94 vdd gnd cell_6t
Xbit_r95_c182 bl_182 br_182 wl_95 vdd gnd cell_6t
Xbit_r96_c182 bl_182 br_182 wl_96 vdd gnd cell_6t
Xbit_r97_c182 bl_182 br_182 wl_97 vdd gnd cell_6t
Xbit_r98_c182 bl_182 br_182 wl_98 vdd gnd cell_6t
Xbit_r99_c182 bl_182 br_182 wl_99 vdd gnd cell_6t
Xbit_r100_c182 bl_182 br_182 wl_100 vdd gnd cell_6t
Xbit_r101_c182 bl_182 br_182 wl_101 vdd gnd cell_6t
Xbit_r102_c182 bl_182 br_182 wl_102 vdd gnd cell_6t
Xbit_r103_c182 bl_182 br_182 wl_103 vdd gnd cell_6t
Xbit_r104_c182 bl_182 br_182 wl_104 vdd gnd cell_6t
Xbit_r105_c182 bl_182 br_182 wl_105 vdd gnd cell_6t
Xbit_r106_c182 bl_182 br_182 wl_106 vdd gnd cell_6t
Xbit_r107_c182 bl_182 br_182 wl_107 vdd gnd cell_6t
Xbit_r108_c182 bl_182 br_182 wl_108 vdd gnd cell_6t
Xbit_r109_c182 bl_182 br_182 wl_109 vdd gnd cell_6t
Xbit_r110_c182 bl_182 br_182 wl_110 vdd gnd cell_6t
Xbit_r111_c182 bl_182 br_182 wl_111 vdd gnd cell_6t
Xbit_r112_c182 bl_182 br_182 wl_112 vdd gnd cell_6t
Xbit_r113_c182 bl_182 br_182 wl_113 vdd gnd cell_6t
Xbit_r114_c182 bl_182 br_182 wl_114 vdd gnd cell_6t
Xbit_r115_c182 bl_182 br_182 wl_115 vdd gnd cell_6t
Xbit_r116_c182 bl_182 br_182 wl_116 vdd gnd cell_6t
Xbit_r117_c182 bl_182 br_182 wl_117 vdd gnd cell_6t
Xbit_r118_c182 bl_182 br_182 wl_118 vdd gnd cell_6t
Xbit_r119_c182 bl_182 br_182 wl_119 vdd gnd cell_6t
Xbit_r120_c182 bl_182 br_182 wl_120 vdd gnd cell_6t
Xbit_r121_c182 bl_182 br_182 wl_121 vdd gnd cell_6t
Xbit_r122_c182 bl_182 br_182 wl_122 vdd gnd cell_6t
Xbit_r123_c182 bl_182 br_182 wl_123 vdd gnd cell_6t
Xbit_r124_c182 bl_182 br_182 wl_124 vdd gnd cell_6t
Xbit_r125_c182 bl_182 br_182 wl_125 vdd gnd cell_6t
Xbit_r126_c182 bl_182 br_182 wl_126 vdd gnd cell_6t
Xbit_r127_c182 bl_182 br_182 wl_127 vdd gnd cell_6t
Xbit_r128_c182 bl_182 br_182 wl_128 vdd gnd cell_6t
Xbit_r129_c182 bl_182 br_182 wl_129 vdd gnd cell_6t
Xbit_r130_c182 bl_182 br_182 wl_130 vdd gnd cell_6t
Xbit_r131_c182 bl_182 br_182 wl_131 vdd gnd cell_6t
Xbit_r132_c182 bl_182 br_182 wl_132 vdd gnd cell_6t
Xbit_r133_c182 bl_182 br_182 wl_133 vdd gnd cell_6t
Xbit_r134_c182 bl_182 br_182 wl_134 vdd gnd cell_6t
Xbit_r135_c182 bl_182 br_182 wl_135 vdd gnd cell_6t
Xbit_r136_c182 bl_182 br_182 wl_136 vdd gnd cell_6t
Xbit_r137_c182 bl_182 br_182 wl_137 vdd gnd cell_6t
Xbit_r138_c182 bl_182 br_182 wl_138 vdd gnd cell_6t
Xbit_r139_c182 bl_182 br_182 wl_139 vdd gnd cell_6t
Xbit_r140_c182 bl_182 br_182 wl_140 vdd gnd cell_6t
Xbit_r141_c182 bl_182 br_182 wl_141 vdd gnd cell_6t
Xbit_r142_c182 bl_182 br_182 wl_142 vdd gnd cell_6t
Xbit_r143_c182 bl_182 br_182 wl_143 vdd gnd cell_6t
Xbit_r144_c182 bl_182 br_182 wl_144 vdd gnd cell_6t
Xbit_r145_c182 bl_182 br_182 wl_145 vdd gnd cell_6t
Xbit_r146_c182 bl_182 br_182 wl_146 vdd gnd cell_6t
Xbit_r147_c182 bl_182 br_182 wl_147 vdd gnd cell_6t
Xbit_r148_c182 bl_182 br_182 wl_148 vdd gnd cell_6t
Xbit_r149_c182 bl_182 br_182 wl_149 vdd gnd cell_6t
Xbit_r150_c182 bl_182 br_182 wl_150 vdd gnd cell_6t
Xbit_r151_c182 bl_182 br_182 wl_151 vdd gnd cell_6t
Xbit_r152_c182 bl_182 br_182 wl_152 vdd gnd cell_6t
Xbit_r153_c182 bl_182 br_182 wl_153 vdd gnd cell_6t
Xbit_r154_c182 bl_182 br_182 wl_154 vdd gnd cell_6t
Xbit_r155_c182 bl_182 br_182 wl_155 vdd gnd cell_6t
Xbit_r156_c182 bl_182 br_182 wl_156 vdd gnd cell_6t
Xbit_r157_c182 bl_182 br_182 wl_157 vdd gnd cell_6t
Xbit_r158_c182 bl_182 br_182 wl_158 vdd gnd cell_6t
Xbit_r159_c182 bl_182 br_182 wl_159 vdd gnd cell_6t
Xbit_r160_c182 bl_182 br_182 wl_160 vdd gnd cell_6t
Xbit_r161_c182 bl_182 br_182 wl_161 vdd gnd cell_6t
Xbit_r162_c182 bl_182 br_182 wl_162 vdd gnd cell_6t
Xbit_r163_c182 bl_182 br_182 wl_163 vdd gnd cell_6t
Xbit_r164_c182 bl_182 br_182 wl_164 vdd gnd cell_6t
Xbit_r165_c182 bl_182 br_182 wl_165 vdd gnd cell_6t
Xbit_r166_c182 bl_182 br_182 wl_166 vdd gnd cell_6t
Xbit_r167_c182 bl_182 br_182 wl_167 vdd gnd cell_6t
Xbit_r168_c182 bl_182 br_182 wl_168 vdd gnd cell_6t
Xbit_r169_c182 bl_182 br_182 wl_169 vdd gnd cell_6t
Xbit_r170_c182 bl_182 br_182 wl_170 vdd gnd cell_6t
Xbit_r171_c182 bl_182 br_182 wl_171 vdd gnd cell_6t
Xbit_r172_c182 bl_182 br_182 wl_172 vdd gnd cell_6t
Xbit_r173_c182 bl_182 br_182 wl_173 vdd gnd cell_6t
Xbit_r174_c182 bl_182 br_182 wl_174 vdd gnd cell_6t
Xbit_r175_c182 bl_182 br_182 wl_175 vdd gnd cell_6t
Xbit_r176_c182 bl_182 br_182 wl_176 vdd gnd cell_6t
Xbit_r177_c182 bl_182 br_182 wl_177 vdd gnd cell_6t
Xbit_r178_c182 bl_182 br_182 wl_178 vdd gnd cell_6t
Xbit_r179_c182 bl_182 br_182 wl_179 vdd gnd cell_6t
Xbit_r180_c182 bl_182 br_182 wl_180 vdd gnd cell_6t
Xbit_r181_c182 bl_182 br_182 wl_181 vdd gnd cell_6t
Xbit_r182_c182 bl_182 br_182 wl_182 vdd gnd cell_6t
Xbit_r183_c182 bl_182 br_182 wl_183 vdd gnd cell_6t
Xbit_r184_c182 bl_182 br_182 wl_184 vdd gnd cell_6t
Xbit_r185_c182 bl_182 br_182 wl_185 vdd gnd cell_6t
Xbit_r186_c182 bl_182 br_182 wl_186 vdd gnd cell_6t
Xbit_r187_c182 bl_182 br_182 wl_187 vdd gnd cell_6t
Xbit_r188_c182 bl_182 br_182 wl_188 vdd gnd cell_6t
Xbit_r189_c182 bl_182 br_182 wl_189 vdd gnd cell_6t
Xbit_r190_c182 bl_182 br_182 wl_190 vdd gnd cell_6t
Xbit_r191_c182 bl_182 br_182 wl_191 vdd gnd cell_6t
Xbit_r192_c182 bl_182 br_182 wl_192 vdd gnd cell_6t
Xbit_r193_c182 bl_182 br_182 wl_193 vdd gnd cell_6t
Xbit_r194_c182 bl_182 br_182 wl_194 vdd gnd cell_6t
Xbit_r195_c182 bl_182 br_182 wl_195 vdd gnd cell_6t
Xbit_r196_c182 bl_182 br_182 wl_196 vdd gnd cell_6t
Xbit_r197_c182 bl_182 br_182 wl_197 vdd gnd cell_6t
Xbit_r198_c182 bl_182 br_182 wl_198 vdd gnd cell_6t
Xbit_r199_c182 bl_182 br_182 wl_199 vdd gnd cell_6t
Xbit_r200_c182 bl_182 br_182 wl_200 vdd gnd cell_6t
Xbit_r201_c182 bl_182 br_182 wl_201 vdd gnd cell_6t
Xbit_r202_c182 bl_182 br_182 wl_202 vdd gnd cell_6t
Xbit_r203_c182 bl_182 br_182 wl_203 vdd gnd cell_6t
Xbit_r204_c182 bl_182 br_182 wl_204 vdd gnd cell_6t
Xbit_r205_c182 bl_182 br_182 wl_205 vdd gnd cell_6t
Xbit_r206_c182 bl_182 br_182 wl_206 vdd gnd cell_6t
Xbit_r207_c182 bl_182 br_182 wl_207 vdd gnd cell_6t
Xbit_r208_c182 bl_182 br_182 wl_208 vdd gnd cell_6t
Xbit_r209_c182 bl_182 br_182 wl_209 vdd gnd cell_6t
Xbit_r210_c182 bl_182 br_182 wl_210 vdd gnd cell_6t
Xbit_r211_c182 bl_182 br_182 wl_211 vdd gnd cell_6t
Xbit_r212_c182 bl_182 br_182 wl_212 vdd gnd cell_6t
Xbit_r213_c182 bl_182 br_182 wl_213 vdd gnd cell_6t
Xbit_r214_c182 bl_182 br_182 wl_214 vdd gnd cell_6t
Xbit_r215_c182 bl_182 br_182 wl_215 vdd gnd cell_6t
Xbit_r216_c182 bl_182 br_182 wl_216 vdd gnd cell_6t
Xbit_r217_c182 bl_182 br_182 wl_217 vdd gnd cell_6t
Xbit_r218_c182 bl_182 br_182 wl_218 vdd gnd cell_6t
Xbit_r219_c182 bl_182 br_182 wl_219 vdd gnd cell_6t
Xbit_r220_c182 bl_182 br_182 wl_220 vdd gnd cell_6t
Xbit_r221_c182 bl_182 br_182 wl_221 vdd gnd cell_6t
Xbit_r222_c182 bl_182 br_182 wl_222 vdd gnd cell_6t
Xbit_r223_c182 bl_182 br_182 wl_223 vdd gnd cell_6t
Xbit_r224_c182 bl_182 br_182 wl_224 vdd gnd cell_6t
Xbit_r225_c182 bl_182 br_182 wl_225 vdd gnd cell_6t
Xbit_r226_c182 bl_182 br_182 wl_226 vdd gnd cell_6t
Xbit_r227_c182 bl_182 br_182 wl_227 vdd gnd cell_6t
Xbit_r228_c182 bl_182 br_182 wl_228 vdd gnd cell_6t
Xbit_r229_c182 bl_182 br_182 wl_229 vdd gnd cell_6t
Xbit_r230_c182 bl_182 br_182 wl_230 vdd gnd cell_6t
Xbit_r231_c182 bl_182 br_182 wl_231 vdd gnd cell_6t
Xbit_r232_c182 bl_182 br_182 wl_232 vdd gnd cell_6t
Xbit_r233_c182 bl_182 br_182 wl_233 vdd gnd cell_6t
Xbit_r234_c182 bl_182 br_182 wl_234 vdd gnd cell_6t
Xbit_r235_c182 bl_182 br_182 wl_235 vdd gnd cell_6t
Xbit_r236_c182 bl_182 br_182 wl_236 vdd gnd cell_6t
Xbit_r237_c182 bl_182 br_182 wl_237 vdd gnd cell_6t
Xbit_r238_c182 bl_182 br_182 wl_238 vdd gnd cell_6t
Xbit_r239_c182 bl_182 br_182 wl_239 vdd gnd cell_6t
Xbit_r240_c182 bl_182 br_182 wl_240 vdd gnd cell_6t
Xbit_r241_c182 bl_182 br_182 wl_241 vdd gnd cell_6t
Xbit_r242_c182 bl_182 br_182 wl_242 vdd gnd cell_6t
Xbit_r243_c182 bl_182 br_182 wl_243 vdd gnd cell_6t
Xbit_r244_c182 bl_182 br_182 wl_244 vdd gnd cell_6t
Xbit_r245_c182 bl_182 br_182 wl_245 vdd gnd cell_6t
Xbit_r246_c182 bl_182 br_182 wl_246 vdd gnd cell_6t
Xbit_r247_c182 bl_182 br_182 wl_247 vdd gnd cell_6t
Xbit_r248_c182 bl_182 br_182 wl_248 vdd gnd cell_6t
Xbit_r249_c182 bl_182 br_182 wl_249 vdd gnd cell_6t
Xbit_r250_c182 bl_182 br_182 wl_250 vdd gnd cell_6t
Xbit_r251_c182 bl_182 br_182 wl_251 vdd gnd cell_6t
Xbit_r252_c182 bl_182 br_182 wl_252 vdd gnd cell_6t
Xbit_r253_c182 bl_182 br_182 wl_253 vdd gnd cell_6t
Xbit_r254_c182 bl_182 br_182 wl_254 vdd gnd cell_6t
Xbit_r255_c182 bl_182 br_182 wl_255 vdd gnd cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd cell_6t
Xbit_r1_c183 bl_183 br_183 wl_1 vdd gnd cell_6t
Xbit_r2_c183 bl_183 br_183 wl_2 vdd gnd cell_6t
Xbit_r3_c183 bl_183 br_183 wl_3 vdd gnd cell_6t
Xbit_r4_c183 bl_183 br_183 wl_4 vdd gnd cell_6t
Xbit_r5_c183 bl_183 br_183 wl_5 vdd gnd cell_6t
Xbit_r6_c183 bl_183 br_183 wl_6 vdd gnd cell_6t
Xbit_r7_c183 bl_183 br_183 wl_7 vdd gnd cell_6t
Xbit_r8_c183 bl_183 br_183 wl_8 vdd gnd cell_6t
Xbit_r9_c183 bl_183 br_183 wl_9 vdd gnd cell_6t
Xbit_r10_c183 bl_183 br_183 wl_10 vdd gnd cell_6t
Xbit_r11_c183 bl_183 br_183 wl_11 vdd gnd cell_6t
Xbit_r12_c183 bl_183 br_183 wl_12 vdd gnd cell_6t
Xbit_r13_c183 bl_183 br_183 wl_13 vdd gnd cell_6t
Xbit_r14_c183 bl_183 br_183 wl_14 vdd gnd cell_6t
Xbit_r15_c183 bl_183 br_183 wl_15 vdd gnd cell_6t
Xbit_r16_c183 bl_183 br_183 wl_16 vdd gnd cell_6t
Xbit_r17_c183 bl_183 br_183 wl_17 vdd gnd cell_6t
Xbit_r18_c183 bl_183 br_183 wl_18 vdd gnd cell_6t
Xbit_r19_c183 bl_183 br_183 wl_19 vdd gnd cell_6t
Xbit_r20_c183 bl_183 br_183 wl_20 vdd gnd cell_6t
Xbit_r21_c183 bl_183 br_183 wl_21 vdd gnd cell_6t
Xbit_r22_c183 bl_183 br_183 wl_22 vdd gnd cell_6t
Xbit_r23_c183 bl_183 br_183 wl_23 vdd gnd cell_6t
Xbit_r24_c183 bl_183 br_183 wl_24 vdd gnd cell_6t
Xbit_r25_c183 bl_183 br_183 wl_25 vdd gnd cell_6t
Xbit_r26_c183 bl_183 br_183 wl_26 vdd gnd cell_6t
Xbit_r27_c183 bl_183 br_183 wl_27 vdd gnd cell_6t
Xbit_r28_c183 bl_183 br_183 wl_28 vdd gnd cell_6t
Xbit_r29_c183 bl_183 br_183 wl_29 vdd gnd cell_6t
Xbit_r30_c183 bl_183 br_183 wl_30 vdd gnd cell_6t
Xbit_r31_c183 bl_183 br_183 wl_31 vdd gnd cell_6t
Xbit_r32_c183 bl_183 br_183 wl_32 vdd gnd cell_6t
Xbit_r33_c183 bl_183 br_183 wl_33 vdd gnd cell_6t
Xbit_r34_c183 bl_183 br_183 wl_34 vdd gnd cell_6t
Xbit_r35_c183 bl_183 br_183 wl_35 vdd gnd cell_6t
Xbit_r36_c183 bl_183 br_183 wl_36 vdd gnd cell_6t
Xbit_r37_c183 bl_183 br_183 wl_37 vdd gnd cell_6t
Xbit_r38_c183 bl_183 br_183 wl_38 vdd gnd cell_6t
Xbit_r39_c183 bl_183 br_183 wl_39 vdd gnd cell_6t
Xbit_r40_c183 bl_183 br_183 wl_40 vdd gnd cell_6t
Xbit_r41_c183 bl_183 br_183 wl_41 vdd gnd cell_6t
Xbit_r42_c183 bl_183 br_183 wl_42 vdd gnd cell_6t
Xbit_r43_c183 bl_183 br_183 wl_43 vdd gnd cell_6t
Xbit_r44_c183 bl_183 br_183 wl_44 vdd gnd cell_6t
Xbit_r45_c183 bl_183 br_183 wl_45 vdd gnd cell_6t
Xbit_r46_c183 bl_183 br_183 wl_46 vdd gnd cell_6t
Xbit_r47_c183 bl_183 br_183 wl_47 vdd gnd cell_6t
Xbit_r48_c183 bl_183 br_183 wl_48 vdd gnd cell_6t
Xbit_r49_c183 bl_183 br_183 wl_49 vdd gnd cell_6t
Xbit_r50_c183 bl_183 br_183 wl_50 vdd gnd cell_6t
Xbit_r51_c183 bl_183 br_183 wl_51 vdd gnd cell_6t
Xbit_r52_c183 bl_183 br_183 wl_52 vdd gnd cell_6t
Xbit_r53_c183 bl_183 br_183 wl_53 vdd gnd cell_6t
Xbit_r54_c183 bl_183 br_183 wl_54 vdd gnd cell_6t
Xbit_r55_c183 bl_183 br_183 wl_55 vdd gnd cell_6t
Xbit_r56_c183 bl_183 br_183 wl_56 vdd gnd cell_6t
Xbit_r57_c183 bl_183 br_183 wl_57 vdd gnd cell_6t
Xbit_r58_c183 bl_183 br_183 wl_58 vdd gnd cell_6t
Xbit_r59_c183 bl_183 br_183 wl_59 vdd gnd cell_6t
Xbit_r60_c183 bl_183 br_183 wl_60 vdd gnd cell_6t
Xbit_r61_c183 bl_183 br_183 wl_61 vdd gnd cell_6t
Xbit_r62_c183 bl_183 br_183 wl_62 vdd gnd cell_6t
Xbit_r63_c183 bl_183 br_183 wl_63 vdd gnd cell_6t
Xbit_r64_c183 bl_183 br_183 wl_64 vdd gnd cell_6t
Xbit_r65_c183 bl_183 br_183 wl_65 vdd gnd cell_6t
Xbit_r66_c183 bl_183 br_183 wl_66 vdd gnd cell_6t
Xbit_r67_c183 bl_183 br_183 wl_67 vdd gnd cell_6t
Xbit_r68_c183 bl_183 br_183 wl_68 vdd gnd cell_6t
Xbit_r69_c183 bl_183 br_183 wl_69 vdd gnd cell_6t
Xbit_r70_c183 bl_183 br_183 wl_70 vdd gnd cell_6t
Xbit_r71_c183 bl_183 br_183 wl_71 vdd gnd cell_6t
Xbit_r72_c183 bl_183 br_183 wl_72 vdd gnd cell_6t
Xbit_r73_c183 bl_183 br_183 wl_73 vdd gnd cell_6t
Xbit_r74_c183 bl_183 br_183 wl_74 vdd gnd cell_6t
Xbit_r75_c183 bl_183 br_183 wl_75 vdd gnd cell_6t
Xbit_r76_c183 bl_183 br_183 wl_76 vdd gnd cell_6t
Xbit_r77_c183 bl_183 br_183 wl_77 vdd gnd cell_6t
Xbit_r78_c183 bl_183 br_183 wl_78 vdd gnd cell_6t
Xbit_r79_c183 bl_183 br_183 wl_79 vdd gnd cell_6t
Xbit_r80_c183 bl_183 br_183 wl_80 vdd gnd cell_6t
Xbit_r81_c183 bl_183 br_183 wl_81 vdd gnd cell_6t
Xbit_r82_c183 bl_183 br_183 wl_82 vdd gnd cell_6t
Xbit_r83_c183 bl_183 br_183 wl_83 vdd gnd cell_6t
Xbit_r84_c183 bl_183 br_183 wl_84 vdd gnd cell_6t
Xbit_r85_c183 bl_183 br_183 wl_85 vdd gnd cell_6t
Xbit_r86_c183 bl_183 br_183 wl_86 vdd gnd cell_6t
Xbit_r87_c183 bl_183 br_183 wl_87 vdd gnd cell_6t
Xbit_r88_c183 bl_183 br_183 wl_88 vdd gnd cell_6t
Xbit_r89_c183 bl_183 br_183 wl_89 vdd gnd cell_6t
Xbit_r90_c183 bl_183 br_183 wl_90 vdd gnd cell_6t
Xbit_r91_c183 bl_183 br_183 wl_91 vdd gnd cell_6t
Xbit_r92_c183 bl_183 br_183 wl_92 vdd gnd cell_6t
Xbit_r93_c183 bl_183 br_183 wl_93 vdd gnd cell_6t
Xbit_r94_c183 bl_183 br_183 wl_94 vdd gnd cell_6t
Xbit_r95_c183 bl_183 br_183 wl_95 vdd gnd cell_6t
Xbit_r96_c183 bl_183 br_183 wl_96 vdd gnd cell_6t
Xbit_r97_c183 bl_183 br_183 wl_97 vdd gnd cell_6t
Xbit_r98_c183 bl_183 br_183 wl_98 vdd gnd cell_6t
Xbit_r99_c183 bl_183 br_183 wl_99 vdd gnd cell_6t
Xbit_r100_c183 bl_183 br_183 wl_100 vdd gnd cell_6t
Xbit_r101_c183 bl_183 br_183 wl_101 vdd gnd cell_6t
Xbit_r102_c183 bl_183 br_183 wl_102 vdd gnd cell_6t
Xbit_r103_c183 bl_183 br_183 wl_103 vdd gnd cell_6t
Xbit_r104_c183 bl_183 br_183 wl_104 vdd gnd cell_6t
Xbit_r105_c183 bl_183 br_183 wl_105 vdd gnd cell_6t
Xbit_r106_c183 bl_183 br_183 wl_106 vdd gnd cell_6t
Xbit_r107_c183 bl_183 br_183 wl_107 vdd gnd cell_6t
Xbit_r108_c183 bl_183 br_183 wl_108 vdd gnd cell_6t
Xbit_r109_c183 bl_183 br_183 wl_109 vdd gnd cell_6t
Xbit_r110_c183 bl_183 br_183 wl_110 vdd gnd cell_6t
Xbit_r111_c183 bl_183 br_183 wl_111 vdd gnd cell_6t
Xbit_r112_c183 bl_183 br_183 wl_112 vdd gnd cell_6t
Xbit_r113_c183 bl_183 br_183 wl_113 vdd gnd cell_6t
Xbit_r114_c183 bl_183 br_183 wl_114 vdd gnd cell_6t
Xbit_r115_c183 bl_183 br_183 wl_115 vdd gnd cell_6t
Xbit_r116_c183 bl_183 br_183 wl_116 vdd gnd cell_6t
Xbit_r117_c183 bl_183 br_183 wl_117 vdd gnd cell_6t
Xbit_r118_c183 bl_183 br_183 wl_118 vdd gnd cell_6t
Xbit_r119_c183 bl_183 br_183 wl_119 vdd gnd cell_6t
Xbit_r120_c183 bl_183 br_183 wl_120 vdd gnd cell_6t
Xbit_r121_c183 bl_183 br_183 wl_121 vdd gnd cell_6t
Xbit_r122_c183 bl_183 br_183 wl_122 vdd gnd cell_6t
Xbit_r123_c183 bl_183 br_183 wl_123 vdd gnd cell_6t
Xbit_r124_c183 bl_183 br_183 wl_124 vdd gnd cell_6t
Xbit_r125_c183 bl_183 br_183 wl_125 vdd gnd cell_6t
Xbit_r126_c183 bl_183 br_183 wl_126 vdd gnd cell_6t
Xbit_r127_c183 bl_183 br_183 wl_127 vdd gnd cell_6t
Xbit_r128_c183 bl_183 br_183 wl_128 vdd gnd cell_6t
Xbit_r129_c183 bl_183 br_183 wl_129 vdd gnd cell_6t
Xbit_r130_c183 bl_183 br_183 wl_130 vdd gnd cell_6t
Xbit_r131_c183 bl_183 br_183 wl_131 vdd gnd cell_6t
Xbit_r132_c183 bl_183 br_183 wl_132 vdd gnd cell_6t
Xbit_r133_c183 bl_183 br_183 wl_133 vdd gnd cell_6t
Xbit_r134_c183 bl_183 br_183 wl_134 vdd gnd cell_6t
Xbit_r135_c183 bl_183 br_183 wl_135 vdd gnd cell_6t
Xbit_r136_c183 bl_183 br_183 wl_136 vdd gnd cell_6t
Xbit_r137_c183 bl_183 br_183 wl_137 vdd gnd cell_6t
Xbit_r138_c183 bl_183 br_183 wl_138 vdd gnd cell_6t
Xbit_r139_c183 bl_183 br_183 wl_139 vdd gnd cell_6t
Xbit_r140_c183 bl_183 br_183 wl_140 vdd gnd cell_6t
Xbit_r141_c183 bl_183 br_183 wl_141 vdd gnd cell_6t
Xbit_r142_c183 bl_183 br_183 wl_142 vdd gnd cell_6t
Xbit_r143_c183 bl_183 br_183 wl_143 vdd gnd cell_6t
Xbit_r144_c183 bl_183 br_183 wl_144 vdd gnd cell_6t
Xbit_r145_c183 bl_183 br_183 wl_145 vdd gnd cell_6t
Xbit_r146_c183 bl_183 br_183 wl_146 vdd gnd cell_6t
Xbit_r147_c183 bl_183 br_183 wl_147 vdd gnd cell_6t
Xbit_r148_c183 bl_183 br_183 wl_148 vdd gnd cell_6t
Xbit_r149_c183 bl_183 br_183 wl_149 vdd gnd cell_6t
Xbit_r150_c183 bl_183 br_183 wl_150 vdd gnd cell_6t
Xbit_r151_c183 bl_183 br_183 wl_151 vdd gnd cell_6t
Xbit_r152_c183 bl_183 br_183 wl_152 vdd gnd cell_6t
Xbit_r153_c183 bl_183 br_183 wl_153 vdd gnd cell_6t
Xbit_r154_c183 bl_183 br_183 wl_154 vdd gnd cell_6t
Xbit_r155_c183 bl_183 br_183 wl_155 vdd gnd cell_6t
Xbit_r156_c183 bl_183 br_183 wl_156 vdd gnd cell_6t
Xbit_r157_c183 bl_183 br_183 wl_157 vdd gnd cell_6t
Xbit_r158_c183 bl_183 br_183 wl_158 vdd gnd cell_6t
Xbit_r159_c183 bl_183 br_183 wl_159 vdd gnd cell_6t
Xbit_r160_c183 bl_183 br_183 wl_160 vdd gnd cell_6t
Xbit_r161_c183 bl_183 br_183 wl_161 vdd gnd cell_6t
Xbit_r162_c183 bl_183 br_183 wl_162 vdd gnd cell_6t
Xbit_r163_c183 bl_183 br_183 wl_163 vdd gnd cell_6t
Xbit_r164_c183 bl_183 br_183 wl_164 vdd gnd cell_6t
Xbit_r165_c183 bl_183 br_183 wl_165 vdd gnd cell_6t
Xbit_r166_c183 bl_183 br_183 wl_166 vdd gnd cell_6t
Xbit_r167_c183 bl_183 br_183 wl_167 vdd gnd cell_6t
Xbit_r168_c183 bl_183 br_183 wl_168 vdd gnd cell_6t
Xbit_r169_c183 bl_183 br_183 wl_169 vdd gnd cell_6t
Xbit_r170_c183 bl_183 br_183 wl_170 vdd gnd cell_6t
Xbit_r171_c183 bl_183 br_183 wl_171 vdd gnd cell_6t
Xbit_r172_c183 bl_183 br_183 wl_172 vdd gnd cell_6t
Xbit_r173_c183 bl_183 br_183 wl_173 vdd gnd cell_6t
Xbit_r174_c183 bl_183 br_183 wl_174 vdd gnd cell_6t
Xbit_r175_c183 bl_183 br_183 wl_175 vdd gnd cell_6t
Xbit_r176_c183 bl_183 br_183 wl_176 vdd gnd cell_6t
Xbit_r177_c183 bl_183 br_183 wl_177 vdd gnd cell_6t
Xbit_r178_c183 bl_183 br_183 wl_178 vdd gnd cell_6t
Xbit_r179_c183 bl_183 br_183 wl_179 vdd gnd cell_6t
Xbit_r180_c183 bl_183 br_183 wl_180 vdd gnd cell_6t
Xbit_r181_c183 bl_183 br_183 wl_181 vdd gnd cell_6t
Xbit_r182_c183 bl_183 br_183 wl_182 vdd gnd cell_6t
Xbit_r183_c183 bl_183 br_183 wl_183 vdd gnd cell_6t
Xbit_r184_c183 bl_183 br_183 wl_184 vdd gnd cell_6t
Xbit_r185_c183 bl_183 br_183 wl_185 vdd gnd cell_6t
Xbit_r186_c183 bl_183 br_183 wl_186 vdd gnd cell_6t
Xbit_r187_c183 bl_183 br_183 wl_187 vdd gnd cell_6t
Xbit_r188_c183 bl_183 br_183 wl_188 vdd gnd cell_6t
Xbit_r189_c183 bl_183 br_183 wl_189 vdd gnd cell_6t
Xbit_r190_c183 bl_183 br_183 wl_190 vdd gnd cell_6t
Xbit_r191_c183 bl_183 br_183 wl_191 vdd gnd cell_6t
Xbit_r192_c183 bl_183 br_183 wl_192 vdd gnd cell_6t
Xbit_r193_c183 bl_183 br_183 wl_193 vdd gnd cell_6t
Xbit_r194_c183 bl_183 br_183 wl_194 vdd gnd cell_6t
Xbit_r195_c183 bl_183 br_183 wl_195 vdd gnd cell_6t
Xbit_r196_c183 bl_183 br_183 wl_196 vdd gnd cell_6t
Xbit_r197_c183 bl_183 br_183 wl_197 vdd gnd cell_6t
Xbit_r198_c183 bl_183 br_183 wl_198 vdd gnd cell_6t
Xbit_r199_c183 bl_183 br_183 wl_199 vdd gnd cell_6t
Xbit_r200_c183 bl_183 br_183 wl_200 vdd gnd cell_6t
Xbit_r201_c183 bl_183 br_183 wl_201 vdd gnd cell_6t
Xbit_r202_c183 bl_183 br_183 wl_202 vdd gnd cell_6t
Xbit_r203_c183 bl_183 br_183 wl_203 vdd gnd cell_6t
Xbit_r204_c183 bl_183 br_183 wl_204 vdd gnd cell_6t
Xbit_r205_c183 bl_183 br_183 wl_205 vdd gnd cell_6t
Xbit_r206_c183 bl_183 br_183 wl_206 vdd gnd cell_6t
Xbit_r207_c183 bl_183 br_183 wl_207 vdd gnd cell_6t
Xbit_r208_c183 bl_183 br_183 wl_208 vdd gnd cell_6t
Xbit_r209_c183 bl_183 br_183 wl_209 vdd gnd cell_6t
Xbit_r210_c183 bl_183 br_183 wl_210 vdd gnd cell_6t
Xbit_r211_c183 bl_183 br_183 wl_211 vdd gnd cell_6t
Xbit_r212_c183 bl_183 br_183 wl_212 vdd gnd cell_6t
Xbit_r213_c183 bl_183 br_183 wl_213 vdd gnd cell_6t
Xbit_r214_c183 bl_183 br_183 wl_214 vdd gnd cell_6t
Xbit_r215_c183 bl_183 br_183 wl_215 vdd gnd cell_6t
Xbit_r216_c183 bl_183 br_183 wl_216 vdd gnd cell_6t
Xbit_r217_c183 bl_183 br_183 wl_217 vdd gnd cell_6t
Xbit_r218_c183 bl_183 br_183 wl_218 vdd gnd cell_6t
Xbit_r219_c183 bl_183 br_183 wl_219 vdd gnd cell_6t
Xbit_r220_c183 bl_183 br_183 wl_220 vdd gnd cell_6t
Xbit_r221_c183 bl_183 br_183 wl_221 vdd gnd cell_6t
Xbit_r222_c183 bl_183 br_183 wl_222 vdd gnd cell_6t
Xbit_r223_c183 bl_183 br_183 wl_223 vdd gnd cell_6t
Xbit_r224_c183 bl_183 br_183 wl_224 vdd gnd cell_6t
Xbit_r225_c183 bl_183 br_183 wl_225 vdd gnd cell_6t
Xbit_r226_c183 bl_183 br_183 wl_226 vdd gnd cell_6t
Xbit_r227_c183 bl_183 br_183 wl_227 vdd gnd cell_6t
Xbit_r228_c183 bl_183 br_183 wl_228 vdd gnd cell_6t
Xbit_r229_c183 bl_183 br_183 wl_229 vdd gnd cell_6t
Xbit_r230_c183 bl_183 br_183 wl_230 vdd gnd cell_6t
Xbit_r231_c183 bl_183 br_183 wl_231 vdd gnd cell_6t
Xbit_r232_c183 bl_183 br_183 wl_232 vdd gnd cell_6t
Xbit_r233_c183 bl_183 br_183 wl_233 vdd gnd cell_6t
Xbit_r234_c183 bl_183 br_183 wl_234 vdd gnd cell_6t
Xbit_r235_c183 bl_183 br_183 wl_235 vdd gnd cell_6t
Xbit_r236_c183 bl_183 br_183 wl_236 vdd gnd cell_6t
Xbit_r237_c183 bl_183 br_183 wl_237 vdd gnd cell_6t
Xbit_r238_c183 bl_183 br_183 wl_238 vdd gnd cell_6t
Xbit_r239_c183 bl_183 br_183 wl_239 vdd gnd cell_6t
Xbit_r240_c183 bl_183 br_183 wl_240 vdd gnd cell_6t
Xbit_r241_c183 bl_183 br_183 wl_241 vdd gnd cell_6t
Xbit_r242_c183 bl_183 br_183 wl_242 vdd gnd cell_6t
Xbit_r243_c183 bl_183 br_183 wl_243 vdd gnd cell_6t
Xbit_r244_c183 bl_183 br_183 wl_244 vdd gnd cell_6t
Xbit_r245_c183 bl_183 br_183 wl_245 vdd gnd cell_6t
Xbit_r246_c183 bl_183 br_183 wl_246 vdd gnd cell_6t
Xbit_r247_c183 bl_183 br_183 wl_247 vdd gnd cell_6t
Xbit_r248_c183 bl_183 br_183 wl_248 vdd gnd cell_6t
Xbit_r249_c183 bl_183 br_183 wl_249 vdd gnd cell_6t
Xbit_r250_c183 bl_183 br_183 wl_250 vdd gnd cell_6t
Xbit_r251_c183 bl_183 br_183 wl_251 vdd gnd cell_6t
Xbit_r252_c183 bl_183 br_183 wl_252 vdd gnd cell_6t
Xbit_r253_c183 bl_183 br_183 wl_253 vdd gnd cell_6t
Xbit_r254_c183 bl_183 br_183 wl_254 vdd gnd cell_6t
Xbit_r255_c183 bl_183 br_183 wl_255 vdd gnd cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd cell_6t
Xbit_r1_c184 bl_184 br_184 wl_1 vdd gnd cell_6t
Xbit_r2_c184 bl_184 br_184 wl_2 vdd gnd cell_6t
Xbit_r3_c184 bl_184 br_184 wl_3 vdd gnd cell_6t
Xbit_r4_c184 bl_184 br_184 wl_4 vdd gnd cell_6t
Xbit_r5_c184 bl_184 br_184 wl_5 vdd gnd cell_6t
Xbit_r6_c184 bl_184 br_184 wl_6 vdd gnd cell_6t
Xbit_r7_c184 bl_184 br_184 wl_7 vdd gnd cell_6t
Xbit_r8_c184 bl_184 br_184 wl_8 vdd gnd cell_6t
Xbit_r9_c184 bl_184 br_184 wl_9 vdd gnd cell_6t
Xbit_r10_c184 bl_184 br_184 wl_10 vdd gnd cell_6t
Xbit_r11_c184 bl_184 br_184 wl_11 vdd gnd cell_6t
Xbit_r12_c184 bl_184 br_184 wl_12 vdd gnd cell_6t
Xbit_r13_c184 bl_184 br_184 wl_13 vdd gnd cell_6t
Xbit_r14_c184 bl_184 br_184 wl_14 vdd gnd cell_6t
Xbit_r15_c184 bl_184 br_184 wl_15 vdd gnd cell_6t
Xbit_r16_c184 bl_184 br_184 wl_16 vdd gnd cell_6t
Xbit_r17_c184 bl_184 br_184 wl_17 vdd gnd cell_6t
Xbit_r18_c184 bl_184 br_184 wl_18 vdd gnd cell_6t
Xbit_r19_c184 bl_184 br_184 wl_19 vdd gnd cell_6t
Xbit_r20_c184 bl_184 br_184 wl_20 vdd gnd cell_6t
Xbit_r21_c184 bl_184 br_184 wl_21 vdd gnd cell_6t
Xbit_r22_c184 bl_184 br_184 wl_22 vdd gnd cell_6t
Xbit_r23_c184 bl_184 br_184 wl_23 vdd gnd cell_6t
Xbit_r24_c184 bl_184 br_184 wl_24 vdd gnd cell_6t
Xbit_r25_c184 bl_184 br_184 wl_25 vdd gnd cell_6t
Xbit_r26_c184 bl_184 br_184 wl_26 vdd gnd cell_6t
Xbit_r27_c184 bl_184 br_184 wl_27 vdd gnd cell_6t
Xbit_r28_c184 bl_184 br_184 wl_28 vdd gnd cell_6t
Xbit_r29_c184 bl_184 br_184 wl_29 vdd gnd cell_6t
Xbit_r30_c184 bl_184 br_184 wl_30 vdd gnd cell_6t
Xbit_r31_c184 bl_184 br_184 wl_31 vdd gnd cell_6t
Xbit_r32_c184 bl_184 br_184 wl_32 vdd gnd cell_6t
Xbit_r33_c184 bl_184 br_184 wl_33 vdd gnd cell_6t
Xbit_r34_c184 bl_184 br_184 wl_34 vdd gnd cell_6t
Xbit_r35_c184 bl_184 br_184 wl_35 vdd gnd cell_6t
Xbit_r36_c184 bl_184 br_184 wl_36 vdd gnd cell_6t
Xbit_r37_c184 bl_184 br_184 wl_37 vdd gnd cell_6t
Xbit_r38_c184 bl_184 br_184 wl_38 vdd gnd cell_6t
Xbit_r39_c184 bl_184 br_184 wl_39 vdd gnd cell_6t
Xbit_r40_c184 bl_184 br_184 wl_40 vdd gnd cell_6t
Xbit_r41_c184 bl_184 br_184 wl_41 vdd gnd cell_6t
Xbit_r42_c184 bl_184 br_184 wl_42 vdd gnd cell_6t
Xbit_r43_c184 bl_184 br_184 wl_43 vdd gnd cell_6t
Xbit_r44_c184 bl_184 br_184 wl_44 vdd gnd cell_6t
Xbit_r45_c184 bl_184 br_184 wl_45 vdd gnd cell_6t
Xbit_r46_c184 bl_184 br_184 wl_46 vdd gnd cell_6t
Xbit_r47_c184 bl_184 br_184 wl_47 vdd gnd cell_6t
Xbit_r48_c184 bl_184 br_184 wl_48 vdd gnd cell_6t
Xbit_r49_c184 bl_184 br_184 wl_49 vdd gnd cell_6t
Xbit_r50_c184 bl_184 br_184 wl_50 vdd gnd cell_6t
Xbit_r51_c184 bl_184 br_184 wl_51 vdd gnd cell_6t
Xbit_r52_c184 bl_184 br_184 wl_52 vdd gnd cell_6t
Xbit_r53_c184 bl_184 br_184 wl_53 vdd gnd cell_6t
Xbit_r54_c184 bl_184 br_184 wl_54 vdd gnd cell_6t
Xbit_r55_c184 bl_184 br_184 wl_55 vdd gnd cell_6t
Xbit_r56_c184 bl_184 br_184 wl_56 vdd gnd cell_6t
Xbit_r57_c184 bl_184 br_184 wl_57 vdd gnd cell_6t
Xbit_r58_c184 bl_184 br_184 wl_58 vdd gnd cell_6t
Xbit_r59_c184 bl_184 br_184 wl_59 vdd gnd cell_6t
Xbit_r60_c184 bl_184 br_184 wl_60 vdd gnd cell_6t
Xbit_r61_c184 bl_184 br_184 wl_61 vdd gnd cell_6t
Xbit_r62_c184 bl_184 br_184 wl_62 vdd gnd cell_6t
Xbit_r63_c184 bl_184 br_184 wl_63 vdd gnd cell_6t
Xbit_r64_c184 bl_184 br_184 wl_64 vdd gnd cell_6t
Xbit_r65_c184 bl_184 br_184 wl_65 vdd gnd cell_6t
Xbit_r66_c184 bl_184 br_184 wl_66 vdd gnd cell_6t
Xbit_r67_c184 bl_184 br_184 wl_67 vdd gnd cell_6t
Xbit_r68_c184 bl_184 br_184 wl_68 vdd gnd cell_6t
Xbit_r69_c184 bl_184 br_184 wl_69 vdd gnd cell_6t
Xbit_r70_c184 bl_184 br_184 wl_70 vdd gnd cell_6t
Xbit_r71_c184 bl_184 br_184 wl_71 vdd gnd cell_6t
Xbit_r72_c184 bl_184 br_184 wl_72 vdd gnd cell_6t
Xbit_r73_c184 bl_184 br_184 wl_73 vdd gnd cell_6t
Xbit_r74_c184 bl_184 br_184 wl_74 vdd gnd cell_6t
Xbit_r75_c184 bl_184 br_184 wl_75 vdd gnd cell_6t
Xbit_r76_c184 bl_184 br_184 wl_76 vdd gnd cell_6t
Xbit_r77_c184 bl_184 br_184 wl_77 vdd gnd cell_6t
Xbit_r78_c184 bl_184 br_184 wl_78 vdd gnd cell_6t
Xbit_r79_c184 bl_184 br_184 wl_79 vdd gnd cell_6t
Xbit_r80_c184 bl_184 br_184 wl_80 vdd gnd cell_6t
Xbit_r81_c184 bl_184 br_184 wl_81 vdd gnd cell_6t
Xbit_r82_c184 bl_184 br_184 wl_82 vdd gnd cell_6t
Xbit_r83_c184 bl_184 br_184 wl_83 vdd gnd cell_6t
Xbit_r84_c184 bl_184 br_184 wl_84 vdd gnd cell_6t
Xbit_r85_c184 bl_184 br_184 wl_85 vdd gnd cell_6t
Xbit_r86_c184 bl_184 br_184 wl_86 vdd gnd cell_6t
Xbit_r87_c184 bl_184 br_184 wl_87 vdd gnd cell_6t
Xbit_r88_c184 bl_184 br_184 wl_88 vdd gnd cell_6t
Xbit_r89_c184 bl_184 br_184 wl_89 vdd gnd cell_6t
Xbit_r90_c184 bl_184 br_184 wl_90 vdd gnd cell_6t
Xbit_r91_c184 bl_184 br_184 wl_91 vdd gnd cell_6t
Xbit_r92_c184 bl_184 br_184 wl_92 vdd gnd cell_6t
Xbit_r93_c184 bl_184 br_184 wl_93 vdd gnd cell_6t
Xbit_r94_c184 bl_184 br_184 wl_94 vdd gnd cell_6t
Xbit_r95_c184 bl_184 br_184 wl_95 vdd gnd cell_6t
Xbit_r96_c184 bl_184 br_184 wl_96 vdd gnd cell_6t
Xbit_r97_c184 bl_184 br_184 wl_97 vdd gnd cell_6t
Xbit_r98_c184 bl_184 br_184 wl_98 vdd gnd cell_6t
Xbit_r99_c184 bl_184 br_184 wl_99 vdd gnd cell_6t
Xbit_r100_c184 bl_184 br_184 wl_100 vdd gnd cell_6t
Xbit_r101_c184 bl_184 br_184 wl_101 vdd gnd cell_6t
Xbit_r102_c184 bl_184 br_184 wl_102 vdd gnd cell_6t
Xbit_r103_c184 bl_184 br_184 wl_103 vdd gnd cell_6t
Xbit_r104_c184 bl_184 br_184 wl_104 vdd gnd cell_6t
Xbit_r105_c184 bl_184 br_184 wl_105 vdd gnd cell_6t
Xbit_r106_c184 bl_184 br_184 wl_106 vdd gnd cell_6t
Xbit_r107_c184 bl_184 br_184 wl_107 vdd gnd cell_6t
Xbit_r108_c184 bl_184 br_184 wl_108 vdd gnd cell_6t
Xbit_r109_c184 bl_184 br_184 wl_109 vdd gnd cell_6t
Xbit_r110_c184 bl_184 br_184 wl_110 vdd gnd cell_6t
Xbit_r111_c184 bl_184 br_184 wl_111 vdd gnd cell_6t
Xbit_r112_c184 bl_184 br_184 wl_112 vdd gnd cell_6t
Xbit_r113_c184 bl_184 br_184 wl_113 vdd gnd cell_6t
Xbit_r114_c184 bl_184 br_184 wl_114 vdd gnd cell_6t
Xbit_r115_c184 bl_184 br_184 wl_115 vdd gnd cell_6t
Xbit_r116_c184 bl_184 br_184 wl_116 vdd gnd cell_6t
Xbit_r117_c184 bl_184 br_184 wl_117 vdd gnd cell_6t
Xbit_r118_c184 bl_184 br_184 wl_118 vdd gnd cell_6t
Xbit_r119_c184 bl_184 br_184 wl_119 vdd gnd cell_6t
Xbit_r120_c184 bl_184 br_184 wl_120 vdd gnd cell_6t
Xbit_r121_c184 bl_184 br_184 wl_121 vdd gnd cell_6t
Xbit_r122_c184 bl_184 br_184 wl_122 vdd gnd cell_6t
Xbit_r123_c184 bl_184 br_184 wl_123 vdd gnd cell_6t
Xbit_r124_c184 bl_184 br_184 wl_124 vdd gnd cell_6t
Xbit_r125_c184 bl_184 br_184 wl_125 vdd gnd cell_6t
Xbit_r126_c184 bl_184 br_184 wl_126 vdd gnd cell_6t
Xbit_r127_c184 bl_184 br_184 wl_127 vdd gnd cell_6t
Xbit_r128_c184 bl_184 br_184 wl_128 vdd gnd cell_6t
Xbit_r129_c184 bl_184 br_184 wl_129 vdd gnd cell_6t
Xbit_r130_c184 bl_184 br_184 wl_130 vdd gnd cell_6t
Xbit_r131_c184 bl_184 br_184 wl_131 vdd gnd cell_6t
Xbit_r132_c184 bl_184 br_184 wl_132 vdd gnd cell_6t
Xbit_r133_c184 bl_184 br_184 wl_133 vdd gnd cell_6t
Xbit_r134_c184 bl_184 br_184 wl_134 vdd gnd cell_6t
Xbit_r135_c184 bl_184 br_184 wl_135 vdd gnd cell_6t
Xbit_r136_c184 bl_184 br_184 wl_136 vdd gnd cell_6t
Xbit_r137_c184 bl_184 br_184 wl_137 vdd gnd cell_6t
Xbit_r138_c184 bl_184 br_184 wl_138 vdd gnd cell_6t
Xbit_r139_c184 bl_184 br_184 wl_139 vdd gnd cell_6t
Xbit_r140_c184 bl_184 br_184 wl_140 vdd gnd cell_6t
Xbit_r141_c184 bl_184 br_184 wl_141 vdd gnd cell_6t
Xbit_r142_c184 bl_184 br_184 wl_142 vdd gnd cell_6t
Xbit_r143_c184 bl_184 br_184 wl_143 vdd gnd cell_6t
Xbit_r144_c184 bl_184 br_184 wl_144 vdd gnd cell_6t
Xbit_r145_c184 bl_184 br_184 wl_145 vdd gnd cell_6t
Xbit_r146_c184 bl_184 br_184 wl_146 vdd gnd cell_6t
Xbit_r147_c184 bl_184 br_184 wl_147 vdd gnd cell_6t
Xbit_r148_c184 bl_184 br_184 wl_148 vdd gnd cell_6t
Xbit_r149_c184 bl_184 br_184 wl_149 vdd gnd cell_6t
Xbit_r150_c184 bl_184 br_184 wl_150 vdd gnd cell_6t
Xbit_r151_c184 bl_184 br_184 wl_151 vdd gnd cell_6t
Xbit_r152_c184 bl_184 br_184 wl_152 vdd gnd cell_6t
Xbit_r153_c184 bl_184 br_184 wl_153 vdd gnd cell_6t
Xbit_r154_c184 bl_184 br_184 wl_154 vdd gnd cell_6t
Xbit_r155_c184 bl_184 br_184 wl_155 vdd gnd cell_6t
Xbit_r156_c184 bl_184 br_184 wl_156 vdd gnd cell_6t
Xbit_r157_c184 bl_184 br_184 wl_157 vdd gnd cell_6t
Xbit_r158_c184 bl_184 br_184 wl_158 vdd gnd cell_6t
Xbit_r159_c184 bl_184 br_184 wl_159 vdd gnd cell_6t
Xbit_r160_c184 bl_184 br_184 wl_160 vdd gnd cell_6t
Xbit_r161_c184 bl_184 br_184 wl_161 vdd gnd cell_6t
Xbit_r162_c184 bl_184 br_184 wl_162 vdd gnd cell_6t
Xbit_r163_c184 bl_184 br_184 wl_163 vdd gnd cell_6t
Xbit_r164_c184 bl_184 br_184 wl_164 vdd gnd cell_6t
Xbit_r165_c184 bl_184 br_184 wl_165 vdd gnd cell_6t
Xbit_r166_c184 bl_184 br_184 wl_166 vdd gnd cell_6t
Xbit_r167_c184 bl_184 br_184 wl_167 vdd gnd cell_6t
Xbit_r168_c184 bl_184 br_184 wl_168 vdd gnd cell_6t
Xbit_r169_c184 bl_184 br_184 wl_169 vdd gnd cell_6t
Xbit_r170_c184 bl_184 br_184 wl_170 vdd gnd cell_6t
Xbit_r171_c184 bl_184 br_184 wl_171 vdd gnd cell_6t
Xbit_r172_c184 bl_184 br_184 wl_172 vdd gnd cell_6t
Xbit_r173_c184 bl_184 br_184 wl_173 vdd gnd cell_6t
Xbit_r174_c184 bl_184 br_184 wl_174 vdd gnd cell_6t
Xbit_r175_c184 bl_184 br_184 wl_175 vdd gnd cell_6t
Xbit_r176_c184 bl_184 br_184 wl_176 vdd gnd cell_6t
Xbit_r177_c184 bl_184 br_184 wl_177 vdd gnd cell_6t
Xbit_r178_c184 bl_184 br_184 wl_178 vdd gnd cell_6t
Xbit_r179_c184 bl_184 br_184 wl_179 vdd gnd cell_6t
Xbit_r180_c184 bl_184 br_184 wl_180 vdd gnd cell_6t
Xbit_r181_c184 bl_184 br_184 wl_181 vdd gnd cell_6t
Xbit_r182_c184 bl_184 br_184 wl_182 vdd gnd cell_6t
Xbit_r183_c184 bl_184 br_184 wl_183 vdd gnd cell_6t
Xbit_r184_c184 bl_184 br_184 wl_184 vdd gnd cell_6t
Xbit_r185_c184 bl_184 br_184 wl_185 vdd gnd cell_6t
Xbit_r186_c184 bl_184 br_184 wl_186 vdd gnd cell_6t
Xbit_r187_c184 bl_184 br_184 wl_187 vdd gnd cell_6t
Xbit_r188_c184 bl_184 br_184 wl_188 vdd gnd cell_6t
Xbit_r189_c184 bl_184 br_184 wl_189 vdd gnd cell_6t
Xbit_r190_c184 bl_184 br_184 wl_190 vdd gnd cell_6t
Xbit_r191_c184 bl_184 br_184 wl_191 vdd gnd cell_6t
Xbit_r192_c184 bl_184 br_184 wl_192 vdd gnd cell_6t
Xbit_r193_c184 bl_184 br_184 wl_193 vdd gnd cell_6t
Xbit_r194_c184 bl_184 br_184 wl_194 vdd gnd cell_6t
Xbit_r195_c184 bl_184 br_184 wl_195 vdd gnd cell_6t
Xbit_r196_c184 bl_184 br_184 wl_196 vdd gnd cell_6t
Xbit_r197_c184 bl_184 br_184 wl_197 vdd gnd cell_6t
Xbit_r198_c184 bl_184 br_184 wl_198 vdd gnd cell_6t
Xbit_r199_c184 bl_184 br_184 wl_199 vdd gnd cell_6t
Xbit_r200_c184 bl_184 br_184 wl_200 vdd gnd cell_6t
Xbit_r201_c184 bl_184 br_184 wl_201 vdd gnd cell_6t
Xbit_r202_c184 bl_184 br_184 wl_202 vdd gnd cell_6t
Xbit_r203_c184 bl_184 br_184 wl_203 vdd gnd cell_6t
Xbit_r204_c184 bl_184 br_184 wl_204 vdd gnd cell_6t
Xbit_r205_c184 bl_184 br_184 wl_205 vdd gnd cell_6t
Xbit_r206_c184 bl_184 br_184 wl_206 vdd gnd cell_6t
Xbit_r207_c184 bl_184 br_184 wl_207 vdd gnd cell_6t
Xbit_r208_c184 bl_184 br_184 wl_208 vdd gnd cell_6t
Xbit_r209_c184 bl_184 br_184 wl_209 vdd gnd cell_6t
Xbit_r210_c184 bl_184 br_184 wl_210 vdd gnd cell_6t
Xbit_r211_c184 bl_184 br_184 wl_211 vdd gnd cell_6t
Xbit_r212_c184 bl_184 br_184 wl_212 vdd gnd cell_6t
Xbit_r213_c184 bl_184 br_184 wl_213 vdd gnd cell_6t
Xbit_r214_c184 bl_184 br_184 wl_214 vdd gnd cell_6t
Xbit_r215_c184 bl_184 br_184 wl_215 vdd gnd cell_6t
Xbit_r216_c184 bl_184 br_184 wl_216 vdd gnd cell_6t
Xbit_r217_c184 bl_184 br_184 wl_217 vdd gnd cell_6t
Xbit_r218_c184 bl_184 br_184 wl_218 vdd gnd cell_6t
Xbit_r219_c184 bl_184 br_184 wl_219 vdd gnd cell_6t
Xbit_r220_c184 bl_184 br_184 wl_220 vdd gnd cell_6t
Xbit_r221_c184 bl_184 br_184 wl_221 vdd gnd cell_6t
Xbit_r222_c184 bl_184 br_184 wl_222 vdd gnd cell_6t
Xbit_r223_c184 bl_184 br_184 wl_223 vdd gnd cell_6t
Xbit_r224_c184 bl_184 br_184 wl_224 vdd gnd cell_6t
Xbit_r225_c184 bl_184 br_184 wl_225 vdd gnd cell_6t
Xbit_r226_c184 bl_184 br_184 wl_226 vdd gnd cell_6t
Xbit_r227_c184 bl_184 br_184 wl_227 vdd gnd cell_6t
Xbit_r228_c184 bl_184 br_184 wl_228 vdd gnd cell_6t
Xbit_r229_c184 bl_184 br_184 wl_229 vdd gnd cell_6t
Xbit_r230_c184 bl_184 br_184 wl_230 vdd gnd cell_6t
Xbit_r231_c184 bl_184 br_184 wl_231 vdd gnd cell_6t
Xbit_r232_c184 bl_184 br_184 wl_232 vdd gnd cell_6t
Xbit_r233_c184 bl_184 br_184 wl_233 vdd gnd cell_6t
Xbit_r234_c184 bl_184 br_184 wl_234 vdd gnd cell_6t
Xbit_r235_c184 bl_184 br_184 wl_235 vdd gnd cell_6t
Xbit_r236_c184 bl_184 br_184 wl_236 vdd gnd cell_6t
Xbit_r237_c184 bl_184 br_184 wl_237 vdd gnd cell_6t
Xbit_r238_c184 bl_184 br_184 wl_238 vdd gnd cell_6t
Xbit_r239_c184 bl_184 br_184 wl_239 vdd gnd cell_6t
Xbit_r240_c184 bl_184 br_184 wl_240 vdd gnd cell_6t
Xbit_r241_c184 bl_184 br_184 wl_241 vdd gnd cell_6t
Xbit_r242_c184 bl_184 br_184 wl_242 vdd gnd cell_6t
Xbit_r243_c184 bl_184 br_184 wl_243 vdd gnd cell_6t
Xbit_r244_c184 bl_184 br_184 wl_244 vdd gnd cell_6t
Xbit_r245_c184 bl_184 br_184 wl_245 vdd gnd cell_6t
Xbit_r246_c184 bl_184 br_184 wl_246 vdd gnd cell_6t
Xbit_r247_c184 bl_184 br_184 wl_247 vdd gnd cell_6t
Xbit_r248_c184 bl_184 br_184 wl_248 vdd gnd cell_6t
Xbit_r249_c184 bl_184 br_184 wl_249 vdd gnd cell_6t
Xbit_r250_c184 bl_184 br_184 wl_250 vdd gnd cell_6t
Xbit_r251_c184 bl_184 br_184 wl_251 vdd gnd cell_6t
Xbit_r252_c184 bl_184 br_184 wl_252 vdd gnd cell_6t
Xbit_r253_c184 bl_184 br_184 wl_253 vdd gnd cell_6t
Xbit_r254_c184 bl_184 br_184 wl_254 vdd gnd cell_6t
Xbit_r255_c184 bl_184 br_184 wl_255 vdd gnd cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd cell_6t
Xbit_r1_c185 bl_185 br_185 wl_1 vdd gnd cell_6t
Xbit_r2_c185 bl_185 br_185 wl_2 vdd gnd cell_6t
Xbit_r3_c185 bl_185 br_185 wl_3 vdd gnd cell_6t
Xbit_r4_c185 bl_185 br_185 wl_4 vdd gnd cell_6t
Xbit_r5_c185 bl_185 br_185 wl_5 vdd gnd cell_6t
Xbit_r6_c185 bl_185 br_185 wl_6 vdd gnd cell_6t
Xbit_r7_c185 bl_185 br_185 wl_7 vdd gnd cell_6t
Xbit_r8_c185 bl_185 br_185 wl_8 vdd gnd cell_6t
Xbit_r9_c185 bl_185 br_185 wl_9 vdd gnd cell_6t
Xbit_r10_c185 bl_185 br_185 wl_10 vdd gnd cell_6t
Xbit_r11_c185 bl_185 br_185 wl_11 vdd gnd cell_6t
Xbit_r12_c185 bl_185 br_185 wl_12 vdd gnd cell_6t
Xbit_r13_c185 bl_185 br_185 wl_13 vdd gnd cell_6t
Xbit_r14_c185 bl_185 br_185 wl_14 vdd gnd cell_6t
Xbit_r15_c185 bl_185 br_185 wl_15 vdd gnd cell_6t
Xbit_r16_c185 bl_185 br_185 wl_16 vdd gnd cell_6t
Xbit_r17_c185 bl_185 br_185 wl_17 vdd gnd cell_6t
Xbit_r18_c185 bl_185 br_185 wl_18 vdd gnd cell_6t
Xbit_r19_c185 bl_185 br_185 wl_19 vdd gnd cell_6t
Xbit_r20_c185 bl_185 br_185 wl_20 vdd gnd cell_6t
Xbit_r21_c185 bl_185 br_185 wl_21 vdd gnd cell_6t
Xbit_r22_c185 bl_185 br_185 wl_22 vdd gnd cell_6t
Xbit_r23_c185 bl_185 br_185 wl_23 vdd gnd cell_6t
Xbit_r24_c185 bl_185 br_185 wl_24 vdd gnd cell_6t
Xbit_r25_c185 bl_185 br_185 wl_25 vdd gnd cell_6t
Xbit_r26_c185 bl_185 br_185 wl_26 vdd gnd cell_6t
Xbit_r27_c185 bl_185 br_185 wl_27 vdd gnd cell_6t
Xbit_r28_c185 bl_185 br_185 wl_28 vdd gnd cell_6t
Xbit_r29_c185 bl_185 br_185 wl_29 vdd gnd cell_6t
Xbit_r30_c185 bl_185 br_185 wl_30 vdd gnd cell_6t
Xbit_r31_c185 bl_185 br_185 wl_31 vdd gnd cell_6t
Xbit_r32_c185 bl_185 br_185 wl_32 vdd gnd cell_6t
Xbit_r33_c185 bl_185 br_185 wl_33 vdd gnd cell_6t
Xbit_r34_c185 bl_185 br_185 wl_34 vdd gnd cell_6t
Xbit_r35_c185 bl_185 br_185 wl_35 vdd gnd cell_6t
Xbit_r36_c185 bl_185 br_185 wl_36 vdd gnd cell_6t
Xbit_r37_c185 bl_185 br_185 wl_37 vdd gnd cell_6t
Xbit_r38_c185 bl_185 br_185 wl_38 vdd gnd cell_6t
Xbit_r39_c185 bl_185 br_185 wl_39 vdd gnd cell_6t
Xbit_r40_c185 bl_185 br_185 wl_40 vdd gnd cell_6t
Xbit_r41_c185 bl_185 br_185 wl_41 vdd gnd cell_6t
Xbit_r42_c185 bl_185 br_185 wl_42 vdd gnd cell_6t
Xbit_r43_c185 bl_185 br_185 wl_43 vdd gnd cell_6t
Xbit_r44_c185 bl_185 br_185 wl_44 vdd gnd cell_6t
Xbit_r45_c185 bl_185 br_185 wl_45 vdd gnd cell_6t
Xbit_r46_c185 bl_185 br_185 wl_46 vdd gnd cell_6t
Xbit_r47_c185 bl_185 br_185 wl_47 vdd gnd cell_6t
Xbit_r48_c185 bl_185 br_185 wl_48 vdd gnd cell_6t
Xbit_r49_c185 bl_185 br_185 wl_49 vdd gnd cell_6t
Xbit_r50_c185 bl_185 br_185 wl_50 vdd gnd cell_6t
Xbit_r51_c185 bl_185 br_185 wl_51 vdd gnd cell_6t
Xbit_r52_c185 bl_185 br_185 wl_52 vdd gnd cell_6t
Xbit_r53_c185 bl_185 br_185 wl_53 vdd gnd cell_6t
Xbit_r54_c185 bl_185 br_185 wl_54 vdd gnd cell_6t
Xbit_r55_c185 bl_185 br_185 wl_55 vdd gnd cell_6t
Xbit_r56_c185 bl_185 br_185 wl_56 vdd gnd cell_6t
Xbit_r57_c185 bl_185 br_185 wl_57 vdd gnd cell_6t
Xbit_r58_c185 bl_185 br_185 wl_58 vdd gnd cell_6t
Xbit_r59_c185 bl_185 br_185 wl_59 vdd gnd cell_6t
Xbit_r60_c185 bl_185 br_185 wl_60 vdd gnd cell_6t
Xbit_r61_c185 bl_185 br_185 wl_61 vdd gnd cell_6t
Xbit_r62_c185 bl_185 br_185 wl_62 vdd gnd cell_6t
Xbit_r63_c185 bl_185 br_185 wl_63 vdd gnd cell_6t
Xbit_r64_c185 bl_185 br_185 wl_64 vdd gnd cell_6t
Xbit_r65_c185 bl_185 br_185 wl_65 vdd gnd cell_6t
Xbit_r66_c185 bl_185 br_185 wl_66 vdd gnd cell_6t
Xbit_r67_c185 bl_185 br_185 wl_67 vdd gnd cell_6t
Xbit_r68_c185 bl_185 br_185 wl_68 vdd gnd cell_6t
Xbit_r69_c185 bl_185 br_185 wl_69 vdd gnd cell_6t
Xbit_r70_c185 bl_185 br_185 wl_70 vdd gnd cell_6t
Xbit_r71_c185 bl_185 br_185 wl_71 vdd gnd cell_6t
Xbit_r72_c185 bl_185 br_185 wl_72 vdd gnd cell_6t
Xbit_r73_c185 bl_185 br_185 wl_73 vdd gnd cell_6t
Xbit_r74_c185 bl_185 br_185 wl_74 vdd gnd cell_6t
Xbit_r75_c185 bl_185 br_185 wl_75 vdd gnd cell_6t
Xbit_r76_c185 bl_185 br_185 wl_76 vdd gnd cell_6t
Xbit_r77_c185 bl_185 br_185 wl_77 vdd gnd cell_6t
Xbit_r78_c185 bl_185 br_185 wl_78 vdd gnd cell_6t
Xbit_r79_c185 bl_185 br_185 wl_79 vdd gnd cell_6t
Xbit_r80_c185 bl_185 br_185 wl_80 vdd gnd cell_6t
Xbit_r81_c185 bl_185 br_185 wl_81 vdd gnd cell_6t
Xbit_r82_c185 bl_185 br_185 wl_82 vdd gnd cell_6t
Xbit_r83_c185 bl_185 br_185 wl_83 vdd gnd cell_6t
Xbit_r84_c185 bl_185 br_185 wl_84 vdd gnd cell_6t
Xbit_r85_c185 bl_185 br_185 wl_85 vdd gnd cell_6t
Xbit_r86_c185 bl_185 br_185 wl_86 vdd gnd cell_6t
Xbit_r87_c185 bl_185 br_185 wl_87 vdd gnd cell_6t
Xbit_r88_c185 bl_185 br_185 wl_88 vdd gnd cell_6t
Xbit_r89_c185 bl_185 br_185 wl_89 vdd gnd cell_6t
Xbit_r90_c185 bl_185 br_185 wl_90 vdd gnd cell_6t
Xbit_r91_c185 bl_185 br_185 wl_91 vdd gnd cell_6t
Xbit_r92_c185 bl_185 br_185 wl_92 vdd gnd cell_6t
Xbit_r93_c185 bl_185 br_185 wl_93 vdd gnd cell_6t
Xbit_r94_c185 bl_185 br_185 wl_94 vdd gnd cell_6t
Xbit_r95_c185 bl_185 br_185 wl_95 vdd gnd cell_6t
Xbit_r96_c185 bl_185 br_185 wl_96 vdd gnd cell_6t
Xbit_r97_c185 bl_185 br_185 wl_97 vdd gnd cell_6t
Xbit_r98_c185 bl_185 br_185 wl_98 vdd gnd cell_6t
Xbit_r99_c185 bl_185 br_185 wl_99 vdd gnd cell_6t
Xbit_r100_c185 bl_185 br_185 wl_100 vdd gnd cell_6t
Xbit_r101_c185 bl_185 br_185 wl_101 vdd gnd cell_6t
Xbit_r102_c185 bl_185 br_185 wl_102 vdd gnd cell_6t
Xbit_r103_c185 bl_185 br_185 wl_103 vdd gnd cell_6t
Xbit_r104_c185 bl_185 br_185 wl_104 vdd gnd cell_6t
Xbit_r105_c185 bl_185 br_185 wl_105 vdd gnd cell_6t
Xbit_r106_c185 bl_185 br_185 wl_106 vdd gnd cell_6t
Xbit_r107_c185 bl_185 br_185 wl_107 vdd gnd cell_6t
Xbit_r108_c185 bl_185 br_185 wl_108 vdd gnd cell_6t
Xbit_r109_c185 bl_185 br_185 wl_109 vdd gnd cell_6t
Xbit_r110_c185 bl_185 br_185 wl_110 vdd gnd cell_6t
Xbit_r111_c185 bl_185 br_185 wl_111 vdd gnd cell_6t
Xbit_r112_c185 bl_185 br_185 wl_112 vdd gnd cell_6t
Xbit_r113_c185 bl_185 br_185 wl_113 vdd gnd cell_6t
Xbit_r114_c185 bl_185 br_185 wl_114 vdd gnd cell_6t
Xbit_r115_c185 bl_185 br_185 wl_115 vdd gnd cell_6t
Xbit_r116_c185 bl_185 br_185 wl_116 vdd gnd cell_6t
Xbit_r117_c185 bl_185 br_185 wl_117 vdd gnd cell_6t
Xbit_r118_c185 bl_185 br_185 wl_118 vdd gnd cell_6t
Xbit_r119_c185 bl_185 br_185 wl_119 vdd gnd cell_6t
Xbit_r120_c185 bl_185 br_185 wl_120 vdd gnd cell_6t
Xbit_r121_c185 bl_185 br_185 wl_121 vdd gnd cell_6t
Xbit_r122_c185 bl_185 br_185 wl_122 vdd gnd cell_6t
Xbit_r123_c185 bl_185 br_185 wl_123 vdd gnd cell_6t
Xbit_r124_c185 bl_185 br_185 wl_124 vdd gnd cell_6t
Xbit_r125_c185 bl_185 br_185 wl_125 vdd gnd cell_6t
Xbit_r126_c185 bl_185 br_185 wl_126 vdd gnd cell_6t
Xbit_r127_c185 bl_185 br_185 wl_127 vdd gnd cell_6t
Xbit_r128_c185 bl_185 br_185 wl_128 vdd gnd cell_6t
Xbit_r129_c185 bl_185 br_185 wl_129 vdd gnd cell_6t
Xbit_r130_c185 bl_185 br_185 wl_130 vdd gnd cell_6t
Xbit_r131_c185 bl_185 br_185 wl_131 vdd gnd cell_6t
Xbit_r132_c185 bl_185 br_185 wl_132 vdd gnd cell_6t
Xbit_r133_c185 bl_185 br_185 wl_133 vdd gnd cell_6t
Xbit_r134_c185 bl_185 br_185 wl_134 vdd gnd cell_6t
Xbit_r135_c185 bl_185 br_185 wl_135 vdd gnd cell_6t
Xbit_r136_c185 bl_185 br_185 wl_136 vdd gnd cell_6t
Xbit_r137_c185 bl_185 br_185 wl_137 vdd gnd cell_6t
Xbit_r138_c185 bl_185 br_185 wl_138 vdd gnd cell_6t
Xbit_r139_c185 bl_185 br_185 wl_139 vdd gnd cell_6t
Xbit_r140_c185 bl_185 br_185 wl_140 vdd gnd cell_6t
Xbit_r141_c185 bl_185 br_185 wl_141 vdd gnd cell_6t
Xbit_r142_c185 bl_185 br_185 wl_142 vdd gnd cell_6t
Xbit_r143_c185 bl_185 br_185 wl_143 vdd gnd cell_6t
Xbit_r144_c185 bl_185 br_185 wl_144 vdd gnd cell_6t
Xbit_r145_c185 bl_185 br_185 wl_145 vdd gnd cell_6t
Xbit_r146_c185 bl_185 br_185 wl_146 vdd gnd cell_6t
Xbit_r147_c185 bl_185 br_185 wl_147 vdd gnd cell_6t
Xbit_r148_c185 bl_185 br_185 wl_148 vdd gnd cell_6t
Xbit_r149_c185 bl_185 br_185 wl_149 vdd gnd cell_6t
Xbit_r150_c185 bl_185 br_185 wl_150 vdd gnd cell_6t
Xbit_r151_c185 bl_185 br_185 wl_151 vdd gnd cell_6t
Xbit_r152_c185 bl_185 br_185 wl_152 vdd gnd cell_6t
Xbit_r153_c185 bl_185 br_185 wl_153 vdd gnd cell_6t
Xbit_r154_c185 bl_185 br_185 wl_154 vdd gnd cell_6t
Xbit_r155_c185 bl_185 br_185 wl_155 vdd gnd cell_6t
Xbit_r156_c185 bl_185 br_185 wl_156 vdd gnd cell_6t
Xbit_r157_c185 bl_185 br_185 wl_157 vdd gnd cell_6t
Xbit_r158_c185 bl_185 br_185 wl_158 vdd gnd cell_6t
Xbit_r159_c185 bl_185 br_185 wl_159 vdd gnd cell_6t
Xbit_r160_c185 bl_185 br_185 wl_160 vdd gnd cell_6t
Xbit_r161_c185 bl_185 br_185 wl_161 vdd gnd cell_6t
Xbit_r162_c185 bl_185 br_185 wl_162 vdd gnd cell_6t
Xbit_r163_c185 bl_185 br_185 wl_163 vdd gnd cell_6t
Xbit_r164_c185 bl_185 br_185 wl_164 vdd gnd cell_6t
Xbit_r165_c185 bl_185 br_185 wl_165 vdd gnd cell_6t
Xbit_r166_c185 bl_185 br_185 wl_166 vdd gnd cell_6t
Xbit_r167_c185 bl_185 br_185 wl_167 vdd gnd cell_6t
Xbit_r168_c185 bl_185 br_185 wl_168 vdd gnd cell_6t
Xbit_r169_c185 bl_185 br_185 wl_169 vdd gnd cell_6t
Xbit_r170_c185 bl_185 br_185 wl_170 vdd gnd cell_6t
Xbit_r171_c185 bl_185 br_185 wl_171 vdd gnd cell_6t
Xbit_r172_c185 bl_185 br_185 wl_172 vdd gnd cell_6t
Xbit_r173_c185 bl_185 br_185 wl_173 vdd gnd cell_6t
Xbit_r174_c185 bl_185 br_185 wl_174 vdd gnd cell_6t
Xbit_r175_c185 bl_185 br_185 wl_175 vdd gnd cell_6t
Xbit_r176_c185 bl_185 br_185 wl_176 vdd gnd cell_6t
Xbit_r177_c185 bl_185 br_185 wl_177 vdd gnd cell_6t
Xbit_r178_c185 bl_185 br_185 wl_178 vdd gnd cell_6t
Xbit_r179_c185 bl_185 br_185 wl_179 vdd gnd cell_6t
Xbit_r180_c185 bl_185 br_185 wl_180 vdd gnd cell_6t
Xbit_r181_c185 bl_185 br_185 wl_181 vdd gnd cell_6t
Xbit_r182_c185 bl_185 br_185 wl_182 vdd gnd cell_6t
Xbit_r183_c185 bl_185 br_185 wl_183 vdd gnd cell_6t
Xbit_r184_c185 bl_185 br_185 wl_184 vdd gnd cell_6t
Xbit_r185_c185 bl_185 br_185 wl_185 vdd gnd cell_6t
Xbit_r186_c185 bl_185 br_185 wl_186 vdd gnd cell_6t
Xbit_r187_c185 bl_185 br_185 wl_187 vdd gnd cell_6t
Xbit_r188_c185 bl_185 br_185 wl_188 vdd gnd cell_6t
Xbit_r189_c185 bl_185 br_185 wl_189 vdd gnd cell_6t
Xbit_r190_c185 bl_185 br_185 wl_190 vdd gnd cell_6t
Xbit_r191_c185 bl_185 br_185 wl_191 vdd gnd cell_6t
Xbit_r192_c185 bl_185 br_185 wl_192 vdd gnd cell_6t
Xbit_r193_c185 bl_185 br_185 wl_193 vdd gnd cell_6t
Xbit_r194_c185 bl_185 br_185 wl_194 vdd gnd cell_6t
Xbit_r195_c185 bl_185 br_185 wl_195 vdd gnd cell_6t
Xbit_r196_c185 bl_185 br_185 wl_196 vdd gnd cell_6t
Xbit_r197_c185 bl_185 br_185 wl_197 vdd gnd cell_6t
Xbit_r198_c185 bl_185 br_185 wl_198 vdd gnd cell_6t
Xbit_r199_c185 bl_185 br_185 wl_199 vdd gnd cell_6t
Xbit_r200_c185 bl_185 br_185 wl_200 vdd gnd cell_6t
Xbit_r201_c185 bl_185 br_185 wl_201 vdd gnd cell_6t
Xbit_r202_c185 bl_185 br_185 wl_202 vdd gnd cell_6t
Xbit_r203_c185 bl_185 br_185 wl_203 vdd gnd cell_6t
Xbit_r204_c185 bl_185 br_185 wl_204 vdd gnd cell_6t
Xbit_r205_c185 bl_185 br_185 wl_205 vdd gnd cell_6t
Xbit_r206_c185 bl_185 br_185 wl_206 vdd gnd cell_6t
Xbit_r207_c185 bl_185 br_185 wl_207 vdd gnd cell_6t
Xbit_r208_c185 bl_185 br_185 wl_208 vdd gnd cell_6t
Xbit_r209_c185 bl_185 br_185 wl_209 vdd gnd cell_6t
Xbit_r210_c185 bl_185 br_185 wl_210 vdd gnd cell_6t
Xbit_r211_c185 bl_185 br_185 wl_211 vdd gnd cell_6t
Xbit_r212_c185 bl_185 br_185 wl_212 vdd gnd cell_6t
Xbit_r213_c185 bl_185 br_185 wl_213 vdd gnd cell_6t
Xbit_r214_c185 bl_185 br_185 wl_214 vdd gnd cell_6t
Xbit_r215_c185 bl_185 br_185 wl_215 vdd gnd cell_6t
Xbit_r216_c185 bl_185 br_185 wl_216 vdd gnd cell_6t
Xbit_r217_c185 bl_185 br_185 wl_217 vdd gnd cell_6t
Xbit_r218_c185 bl_185 br_185 wl_218 vdd gnd cell_6t
Xbit_r219_c185 bl_185 br_185 wl_219 vdd gnd cell_6t
Xbit_r220_c185 bl_185 br_185 wl_220 vdd gnd cell_6t
Xbit_r221_c185 bl_185 br_185 wl_221 vdd gnd cell_6t
Xbit_r222_c185 bl_185 br_185 wl_222 vdd gnd cell_6t
Xbit_r223_c185 bl_185 br_185 wl_223 vdd gnd cell_6t
Xbit_r224_c185 bl_185 br_185 wl_224 vdd gnd cell_6t
Xbit_r225_c185 bl_185 br_185 wl_225 vdd gnd cell_6t
Xbit_r226_c185 bl_185 br_185 wl_226 vdd gnd cell_6t
Xbit_r227_c185 bl_185 br_185 wl_227 vdd gnd cell_6t
Xbit_r228_c185 bl_185 br_185 wl_228 vdd gnd cell_6t
Xbit_r229_c185 bl_185 br_185 wl_229 vdd gnd cell_6t
Xbit_r230_c185 bl_185 br_185 wl_230 vdd gnd cell_6t
Xbit_r231_c185 bl_185 br_185 wl_231 vdd gnd cell_6t
Xbit_r232_c185 bl_185 br_185 wl_232 vdd gnd cell_6t
Xbit_r233_c185 bl_185 br_185 wl_233 vdd gnd cell_6t
Xbit_r234_c185 bl_185 br_185 wl_234 vdd gnd cell_6t
Xbit_r235_c185 bl_185 br_185 wl_235 vdd gnd cell_6t
Xbit_r236_c185 bl_185 br_185 wl_236 vdd gnd cell_6t
Xbit_r237_c185 bl_185 br_185 wl_237 vdd gnd cell_6t
Xbit_r238_c185 bl_185 br_185 wl_238 vdd gnd cell_6t
Xbit_r239_c185 bl_185 br_185 wl_239 vdd gnd cell_6t
Xbit_r240_c185 bl_185 br_185 wl_240 vdd gnd cell_6t
Xbit_r241_c185 bl_185 br_185 wl_241 vdd gnd cell_6t
Xbit_r242_c185 bl_185 br_185 wl_242 vdd gnd cell_6t
Xbit_r243_c185 bl_185 br_185 wl_243 vdd gnd cell_6t
Xbit_r244_c185 bl_185 br_185 wl_244 vdd gnd cell_6t
Xbit_r245_c185 bl_185 br_185 wl_245 vdd gnd cell_6t
Xbit_r246_c185 bl_185 br_185 wl_246 vdd gnd cell_6t
Xbit_r247_c185 bl_185 br_185 wl_247 vdd gnd cell_6t
Xbit_r248_c185 bl_185 br_185 wl_248 vdd gnd cell_6t
Xbit_r249_c185 bl_185 br_185 wl_249 vdd gnd cell_6t
Xbit_r250_c185 bl_185 br_185 wl_250 vdd gnd cell_6t
Xbit_r251_c185 bl_185 br_185 wl_251 vdd gnd cell_6t
Xbit_r252_c185 bl_185 br_185 wl_252 vdd gnd cell_6t
Xbit_r253_c185 bl_185 br_185 wl_253 vdd gnd cell_6t
Xbit_r254_c185 bl_185 br_185 wl_254 vdd gnd cell_6t
Xbit_r255_c185 bl_185 br_185 wl_255 vdd gnd cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd cell_6t
Xbit_r1_c186 bl_186 br_186 wl_1 vdd gnd cell_6t
Xbit_r2_c186 bl_186 br_186 wl_2 vdd gnd cell_6t
Xbit_r3_c186 bl_186 br_186 wl_3 vdd gnd cell_6t
Xbit_r4_c186 bl_186 br_186 wl_4 vdd gnd cell_6t
Xbit_r5_c186 bl_186 br_186 wl_5 vdd gnd cell_6t
Xbit_r6_c186 bl_186 br_186 wl_6 vdd gnd cell_6t
Xbit_r7_c186 bl_186 br_186 wl_7 vdd gnd cell_6t
Xbit_r8_c186 bl_186 br_186 wl_8 vdd gnd cell_6t
Xbit_r9_c186 bl_186 br_186 wl_9 vdd gnd cell_6t
Xbit_r10_c186 bl_186 br_186 wl_10 vdd gnd cell_6t
Xbit_r11_c186 bl_186 br_186 wl_11 vdd gnd cell_6t
Xbit_r12_c186 bl_186 br_186 wl_12 vdd gnd cell_6t
Xbit_r13_c186 bl_186 br_186 wl_13 vdd gnd cell_6t
Xbit_r14_c186 bl_186 br_186 wl_14 vdd gnd cell_6t
Xbit_r15_c186 bl_186 br_186 wl_15 vdd gnd cell_6t
Xbit_r16_c186 bl_186 br_186 wl_16 vdd gnd cell_6t
Xbit_r17_c186 bl_186 br_186 wl_17 vdd gnd cell_6t
Xbit_r18_c186 bl_186 br_186 wl_18 vdd gnd cell_6t
Xbit_r19_c186 bl_186 br_186 wl_19 vdd gnd cell_6t
Xbit_r20_c186 bl_186 br_186 wl_20 vdd gnd cell_6t
Xbit_r21_c186 bl_186 br_186 wl_21 vdd gnd cell_6t
Xbit_r22_c186 bl_186 br_186 wl_22 vdd gnd cell_6t
Xbit_r23_c186 bl_186 br_186 wl_23 vdd gnd cell_6t
Xbit_r24_c186 bl_186 br_186 wl_24 vdd gnd cell_6t
Xbit_r25_c186 bl_186 br_186 wl_25 vdd gnd cell_6t
Xbit_r26_c186 bl_186 br_186 wl_26 vdd gnd cell_6t
Xbit_r27_c186 bl_186 br_186 wl_27 vdd gnd cell_6t
Xbit_r28_c186 bl_186 br_186 wl_28 vdd gnd cell_6t
Xbit_r29_c186 bl_186 br_186 wl_29 vdd gnd cell_6t
Xbit_r30_c186 bl_186 br_186 wl_30 vdd gnd cell_6t
Xbit_r31_c186 bl_186 br_186 wl_31 vdd gnd cell_6t
Xbit_r32_c186 bl_186 br_186 wl_32 vdd gnd cell_6t
Xbit_r33_c186 bl_186 br_186 wl_33 vdd gnd cell_6t
Xbit_r34_c186 bl_186 br_186 wl_34 vdd gnd cell_6t
Xbit_r35_c186 bl_186 br_186 wl_35 vdd gnd cell_6t
Xbit_r36_c186 bl_186 br_186 wl_36 vdd gnd cell_6t
Xbit_r37_c186 bl_186 br_186 wl_37 vdd gnd cell_6t
Xbit_r38_c186 bl_186 br_186 wl_38 vdd gnd cell_6t
Xbit_r39_c186 bl_186 br_186 wl_39 vdd gnd cell_6t
Xbit_r40_c186 bl_186 br_186 wl_40 vdd gnd cell_6t
Xbit_r41_c186 bl_186 br_186 wl_41 vdd gnd cell_6t
Xbit_r42_c186 bl_186 br_186 wl_42 vdd gnd cell_6t
Xbit_r43_c186 bl_186 br_186 wl_43 vdd gnd cell_6t
Xbit_r44_c186 bl_186 br_186 wl_44 vdd gnd cell_6t
Xbit_r45_c186 bl_186 br_186 wl_45 vdd gnd cell_6t
Xbit_r46_c186 bl_186 br_186 wl_46 vdd gnd cell_6t
Xbit_r47_c186 bl_186 br_186 wl_47 vdd gnd cell_6t
Xbit_r48_c186 bl_186 br_186 wl_48 vdd gnd cell_6t
Xbit_r49_c186 bl_186 br_186 wl_49 vdd gnd cell_6t
Xbit_r50_c186 bl_186 br_186 wl_50 vdd gnd cell_6t
Xbit_r51_c186 bl_186 br_186 wl_51 vdd gnd cell_6t
Xbit_r52_c186 bl_186 br_186 wl_52 vdd gnd cell_6t
Xbit_r53_c186 bl_186 br_186 wl_53 vdd gnd cell_6t
Xbit_r54_c186 bl_186 br_186 wl_54 vdd gnd cell_6t
Xbit_r55_c186 bl_186 br_186 wl_55 vdd gnd cell_6t
Xbit_r56_c186 bl_186 br_186 wl_56 vdd gnd cell_6t
Xbit_r57_c186 bl_186 br_186 wl_57 vdd gnd cell_6t
Xbit_r58_c186 bl_186 br_186 wl_58 vdd gnd cell_6t
Xbit_r59_c186 bl_186 br_186 wl_59 vdd gnd cell_6t
Xbit_r60_c186 bl_186 br_186 wl_60 vdd gnd cell_6t
Xbit_r61_c186 bl_186 br_186 wl_61 vdd gnd cell_6t
Xbit_r62_c186 bl_186 br_186 wl_62 vdd gnd cell_6t
Xbit_r63_c186 bl_186 br_186 wl_63 vdd gnd cell_6t
Xbit_r64_c186 bl_186 br_186 wl_64 vdd gnd cell_6t
Xbit_r65_c186 bl_186 br_186 wl_65 vdd gnd cell_6t
Xbit_r66_c186 bl_186 br_186 wl_66 vdd gnd cell_6t
Xbit_r67_c186 bl_186 br_186 wl_67 vdd gnd cell_6t
Xbit_r68_c186 bl_186 br_186 wl_68 vdd gnd cell_6t
Xbit_r69_c186 bl_186 br_186 wl_69 vdd gnd cell_6t
Xbit_r70_c186 bl_186 br_186 wl_70 vdd gnd cell_6t
Xbit_r71_c186 bl_186 br_186 wl_71 vdd gnd cell_6t
Xbit_r72_c186 bl_186 br_186 wl_72 vdd gnd cell_6t
Xbit_r73_c186 bl_186 br_186 wl_73 vdd gnd cell_6t
Xbit_r74_c186 bl_186 br_186 wl_74 vdd gnd cell_6t
Xbit_r75_c186 bl_186 br_186 wl_75 vdd gnd cell_6t
Xbit_r76_c186 bl_186 br_186 wl_76 vdd gnd cell_6t
Xbit_r77_c186 bl_186 br_186 wl_77 vdd gnd cell_6t
Xbit_r78_c186 bl_186 br_186 wl_78 vdd gnd cell_6t
Xbit_r79_c186 bl_186 br_186 wl_79 vdd gnd cell_6t
Xbit_r80_c186 bl_186 br_186 wl_80 vdd gnd cell_6t
Xbit_r81_c186 bl_186 br_186 wl_81 vdd gnd cell_6t
Xbit_r82_c186 bl_186 br_186 wl_82 vdd gnd cell_6t
Xbit_r83_c186 bl_186 br_186 wl_83 vdd gnd cell_6t
Xbit_r84_c186 bl_186 br_186 wl_84 vdd gnd cell_6t
Xbit_r85_c186 bl_186 br_186 wl_85 vdd gnd cell_6t
Xbit_r86_c186 bl_186 br_186 wl_86 vdd gnd cell_6t
Xbit_r87_c186 bl_186 br_186 wl_87 vdd gnd cell_6t
Xbit_r88_c186 bl_186 br_186 wl_88 vdd gnd cell_6t
Xbit_r89_c186 bl_186 br_186 wl_89 vdd gnd cell_6t
Xbit_r90_c186 bl_186 br_186 wl_90 vdd gnd cell_6t
Xbit_r91_c186 bl_186 br_186 wl_91 vdd gnd cell_6t
Xbit_r92_c186 bl_186 br_186 wl_92 vdd gnd cell_6t
Xbit_r93_c186 bl_186 br_186 wl_93 vdd gnd cell_6t
Xbit_r94_c186 bl_186 br_186 wl_94 vdd gnd cell_6t
Xbit_r95_c186 bl_186 br_186 wl_95 vdd gnd cell_6t
Xbit_r96_c186 bl_186 br_186 wl_96 vdd gnd cell_6t
Xbit_r97_c186 bl_186 br_186 wl_97 vdd gnd cell_6t
Xbit_r98_c186 bl_186 br_186 wl_98 vdd gnd cell_6t
Xbit_r99_c186 bl_186 br_186 wl_99 vdd gnd cell_6t
Xbit_r100_c186 bl_186 br_186 wl_100 vdd gnd cell_6t
Xbit_r101_c186 bl_186 br_186 wl_101 vdd gnd cell_6t
Xbit_r102_c186 bl_186 br_186 wl_102 vdd gnd cell_6t
Xbit_r103_c186 bl_186 br_186 wl_103 vdd gnd cell_6t
Xbit_r104_c186 bl_186 br_186 wl_104 vdd gnd cell_6t
Xbit_r105_c186 bl_186 br_186 wl_105 vdd gnd cell_6t
Xbit_r106_c186 bl_186 br_186 wl_106 vdd gnd cell_6t
Xbit_r107_c186 bl_186 br_186 wl_107 vdd gnd cell_6t
Xbit_r108_c186 bl_186 br_186 wl_108 vdd gnd cell_6t
Xbit_r109_c186 bl_186 br_186 wl_109 vdd gnd cell_6t
Xbit_r110_c186 bl_186 br_186 wl_110 vdd gnd cell_6t
Xbit_r111_c186 bl_186 br_186 wl_111 vdd gnd cell_6t
Xbit_r112_c186 bl_186 br_186 wl_112 vdd gnd cell_6t
Xbit_r113_c186 bl_186 br_186 wl_113 vdd gnd cell_6t
Xbit_r114_c186 bl_186 br_186 wl_114 vdd gnd cell_6t
Xbit_r115_c186 bl_186 br_186 wl_115 vdd gnd cell_6t
Xbit_r116_c186 bl_186 br_186 wl_116 vdd gnd cell_6t
Xbit_r117_c186 bl_186 br_186 wl_117 vdd gnd cell_6t
Xbit_r118_c186 bl_186 br_186 wl_118 vdd gnd cell_6t
Xbit_r119_c186 bl_186 br_186 wl_119 vdd gnd cell_6t
Xbit_r120_c186 bl_186 br_186 wl_120 vdd gnd cell_6t
Xbit_r121_c186 bl_186 br_186 wl_121 vdd gnd cell_6t
Xbit_r122_c186 bl_186 br_186 wl_122 vdd gnd cell_6t
Xbit_r123_c186 bl_186 br_186 wl_123 vdd gnd cell_6t
Xbit_r124_c186 bl_186 br_186 wl_124 vdd gnd cell_6t
Xbit_r125_c186 bl_186 br_186 wl_125 vdd gnd cell_6t
Xbit_r126_c186 bl_186 br_186 wl_126 vdd gnd cell_6t
Xbit_r127_c186 bl_186 br_186 wl_127 vdd gnd cell_6t
Xbit_r128_c186 bl_186 br_186 wl_128 vdd gnd cell_6t
Xbit_r129_c186 bl_186 br_186 wl_129 vdd gnd cell_6t
Xbit_r130_c186 bl_186 br_186 wl_130 vdd gnd cell_6t
Xbit_r131_c186 bl_186 br_186 wl_131 vdd gnd cell_6t
Xbit_r132_c186 bl_186 br_186 wl_132 vdd gnd cell_6t
Xbit_r133_c186 bl_186 br_186 wl_133 vdd gnd cell_6t
Xbit_r134_c186 bl_186 br_186 wl_134 vdd gnd cell_6t
Xbit_r135_c186 bl_186 br_186 wl_135 vdd gnd cell_6t
Xbit_r136_c186 bl_186 br_186 wl_136 vdd gnd cell_6t
Xbit_r137_c186 bl_186 br_186 wl_137 vdd gnd cell_6t
Xbit_r138_c186 bl_186 br_186 wl_138 vdd gnd cell_6t
Xbit_r139_c186 bl_186 br_186 wl_139 vdd gnd cell_6t
Xbit_r140_c186 bl_186 br_186 wl_140 vdd gnd cell_6t
Xbit_r141_c186 bl_186 br_186 wl_141 vdd gnd cell_6t
Xbit_r142_c186 bl_186 br_186 wl_142 vdd gnd cell_6t
Xbit_r143_c186 bl_186 br_186 wl_143 vdd gnd cell_6t
Xbit_r144_c186 bl_186 br_186 wl_144 vdd gnd cell_6t
Xbit_r145_c186 bl_186 br_186 wl_145 vdd gnd cell_6t
Xbit_r146_c186 bl_186 br_186 wl_146 vdd gnd cell_6t
Xbit_r147_c186 bl_186 br_186 wl_147 vdd gnd cell_6t
Xbit_r148_c186 bl_186 br_186 wl_148 vdd gnd cell_6t
Xbit_r149_c186 bl_186 br_186 wl_149 vdd gnd cell_6t
Xbit_r150_c186 bl_186 br_186 wl_150 vdd gnd cell_6t
Xbit_r151_c186 bl_186 br_186 wl_151 vdd gnd cell_6t
Xbit_r152_c186 bl_186 br_186 wl_152 vdd gnd cell_6t
Xbit_r153_c186 bl_186 br_186 wl_153 vdd gnd cell_6t
Xbit_r154_c186 bl_186 br_186 wl_154 vdd gnd cell_6t
Xbit_r155_c186 bl_186 br_186 wl_155 vdd gnd cell_6t
Xbit_r156_c186 bl_186 br_186 wl_156 vdd gnd cell_6t
Xbit_r157_c186 bl_186 br_186 wl_157 vdd gnd cell_6t
Xbit_r158_c186 bl_186 br_186 wl_158 vdd gnd cell_6t
Xbit_r159_c186 bl_186 br_186 wl_159 vdd gnd cell_6t
Xbit_r160_c186 bl_186 br_186 wl_160 vdd gnd cell_6t
Xbit_r161_c186 bl_186 br_186 wl_161 vdd gnd cell_6t
Xbit_r162_c186 bl_186 br_186 wl_162 vdd gnd cell_6t
Xbit_r163_c186 bl_186 br_186 wl_163 vdd gnd cell_6t
Xbit_r164_c186 bl_186 br_186 wl_164 vdd gnd cell_6t
Xbit_r165_c186 bl_186 br_186 wl_165 vdd gnd cell_6t
Xbit_r166_c186 bl_186 br_186 wl_166 vdd gnd cell_6t
Xbit_r167_c186 bl_186 br_186 wl_167 vdd gnd cell_6t
Xbit_r168_c186 bl_186 br_186 wl_168 vdd gnd cell_6t
Xbit_r169_c186 bl_186 br_186 wl_169 vdd gnd cell_6t
Xbit_r170_c186 bl_186 br_186 wl_170 vdd gnd cell_6t
Xbit_r171_c186 bl_186 br_186 wl_171 vdd gnd cell_6t
Xbit_r172_c186 bl_186 br_186 wl_172 vdd gnd cell_6t
Xbit_r173_c186 bl_186 br_186 wl_173 vdd gnd cell_6t
Xbit_r174_c186 bl_186 br_186 wl_174 vdd gnd cell_6t
Xbit_r175_c186 bl_186 br_186 wl_175 vdd gnd cell_6t
Xbit_r176_c186 bl_186 br_186 wl_176 vdd gnd cell_6t
Xbit_r177_c186 bl_186 br_186 wl_177 vdd gnd cell_6t
Xbit_r178_c186 bl_186 br_186 wl_178 vdd gnd cell_6t
Xbit_r179_c186 bl_186 br_186 wl_179 vdd gnd cell_6t
Xbit_r180_c186 bl_186 br_186 wl_180 vdd gnd cell_6t
Xbit_r181_c186 bl_186 br_186 wl_181 vdd gnd cell_6t
Xbit_r182_c186 bl_186 br_186 wl_182 vdd gnd cell_6t
Xbit_r183_c186 bl_186 br_186 wl_183 vdd gnd cell_6t
Xbit_r184_c186 bl_186 br_186 wl_184 vdd gnd cell_6t
Xbit_r185_c186 bl_186 br_186 wl_185 vdd gnd cell_6t
Xbit_r186_c186 bl_186 br_186 wl_186 vdd gnd cell_6t
Xbit_r187_c186 bl_186 br_186 wl_187 vdd gnd cell_6t
Xbit_r188_c186 bl_186 br_186 wl_188 vdd gnd cell_6t
Xbit_r189_c186 bl_186 br_186 wl_189 vdd gnd cell_6t
Xbit_r190_c186 bl_186 br_186 wl_190 vdd gnd cell_6t
Xbit_r191_c186 bl_186 br_186 wl_191 vdd gnd cell_6t
Xbit_r192_c186 bl_186 br_186 wl_192 vdd gnd cell_6t
Xbit_r193_c186 bl_186 br_186 wl_193 vdd gnd cell_6t
Xbit_r194_c186 bl_186 br_186 wl_194 vdd gnd cell_6t
Xbit_r195_c186 bl_186 br_186 wl_195 vdd gnd cell_6t
Xbit_r196_c186 bl_186 br_186 wl_196 vdd gnd cell_6t
Xbit_r197_c186 bl_186 br_186 wl_197 vdd gnd cell_6t
Xbit_r198_c186 bl_186 br_186 wl_198 vdd gnd cell_6t
Xbit_r199_c186 bl_186 br_186 wl_199 vdd gnd cell_6t
Xbit_r200_c186 bl_186 br_186 wl_200 vdd gnd cell_6t
Xbit_r201_c186 bl_186 br_186 wl_201 vdd gnd cell_6t
Xbit_r202_c186 bl_186 br_186 wl_202 vdd gnd cell_6t
Xbit_r203_c186 bl_186 br_186 wl_203 vdd gnd cell_6t
Xbit_r204_c186 bl_186 br_186 wl_204 vdd gnd cell_6t
Xbit_r205_c186 bl_186 br_186 wl_205 vdd gnd cell_6t
Xbit_r206_c186 bl_186 br_186 wl_206 vdd gnd cell_6t
Xbit_r207_c186 bl_186 br_186 wl_207 vdd gnd cell_6t
Xbit_r208_c186 bl_186 br_186 wl_208 vdd gnd cell_6t
Xbit_r209_c186 bl_186 br_186 wl_209 vdd gnd cell_6t
Xbit_r210_c186 bl_186 br_186 wl_210 vdd gnd cell_6t
Xbit_r211_c186 bl_186 br_186 wl_211 vdd gnd cell_6t
Xbit_r212_c186 bl_186 br_186 wl_212 vdd gnd cell_6t
Xbit_r213_c186 bl_186 br_186 wl_213 vdd gnd cell_6t
Xbit_r214_c186 bl_186 br_186 wl_214 vdd gnd cell_6t
Xbit_r215_c186 bl_186 br_186 wl_215 vdd gnd cell_6t
Xbit_r216_c186 bl_186 br_186 wl_216 vdd gnd cell_6t
Xbit_r217_c186 bl_186 br_186 wl_217 vdd gnd cell_6t
Xbit_r218_c186 bl_186 br_186 wl_218 vdd gnd cell_6t
Xbit_r219_c186 bl_186 br_186 wl_219 vdd gnd cell_6t
Xbit_r220_c186 bl_186 br_186 wl_220 vdd gnd cell_6t
Xbit_r221_c186 bl_186 br_186 wl_221 vdd gnd cell_6t
Xbit_r222_c186 bl_186 br_186 wl_222 vdd gnd cell_6t
Xbit_r223_c186 bl_186 br_186 wl_223 vdd gnd cell_6t
Xbit_r224_c186 bl_186 br_186 wl_224 vdd gnd cell_6t
Xbit_r225_c186 bl_186 br_186 wl_225 vdd gnd cell_6t
Xbit_r226_c186 bl_186 br_186 wl_226 vdd gnd cell_6t
Xbit_r227_c186 bl_186 br_186 wl_227 vdd gnd cell_6t
Xbit_r228_c186 bl_186 br_186 wl_228 vdd gnd cell_6t
Xbit_r229_c186 bl_186 br_186 wl_229 vdd gnd cell_6t
Xbit_r230_c186 bl_186 br_186 wl_230 vdd gnd cell_6t
Xbit_r231_c186 bl_186 br_186 wl_231 vdd gnd cell_6t
Xbit_r232_c186 bl_186 br_186 wl_232 vdd gnd cell_6t
Xbit_r233_c186 bl_186 br_186 wl_233 vdd gnd cell_6t
Xbit_r234_c186 bl_186 br_186 wl_234 vdd gnd cell_6t
Xbit_r235_c186 bl_186 br_186 wl_235 vdd gnd cell_6t
Xbit_r236_c186 bl_186 br_186 wl_236 vdd gnd cell_6t
Xbit_r237_c186 bl_186 br_186 wl_237 vdd gnd cell_6t
Xbit_r238_c186 bl_186 br_186 wl_238 vdd gnd cell_6t
Xbit_r239_c186 bl_186 br_186 wl_239 vdd gnd cell_6t
Xbit_r240_c186 bl_186 br_186 wl_240 vdd gnd cell_6t
Xbit_r241_c186 bl_186 br_186 wl_241 vdd gnd cell_6t
Xbit_r242_c186 bl_186 br_186 wl_242 vdd gnd cell_6t
Xbit_r243_c186 bl_186 br_186 wl_243 vdd gnd cell_6t
Xbit_r244_c186 bl_186 br_186 wl_244 vdd gnd cell_6t
Xbit_r245_c186 bl_186 br_186 wl_245 vdd gnd cell_6t
Xbit_r246_c186 bl_186 br_186 wl_246 vdd gnd cell_6t
Xbit_r247_c186 bl_186 br_186 wl_247 vdd gnd cell_6t
Xbit_r248_c186 bl_186 br_186 wl_248 vdd gnd cell_6t
Xbit_r249_c186 bl_186 br_186 wl_249 vdd gnd cell_6t
Xbit_r250_c186 bl_186 br_186 wl_250 vdd gnd cell_6t
Xbit_r251_c186 bl_186 br_186 wl_251 vdd gnd cell_6t
Xbit_r252_c186 bl_186 br_186 wl_252 vdd gnd cell_6t
Xbit_r253_c186 bl_186 br_186 wl_253 vdd gnd cell_6t
Xbit_r254_c186 bl_186 br_186 wl_254 vdd gnd cell_6t
Xbit_r255_c186 bl_186 br_186 wl_255 vdd gnd cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd cell_6t
Xbit_r1_c187 bl_187 br_187 wl_1 vdd gnd cell_6t
Xbit_r2_c187 bl_187 br_187 wl_2 vdd gnd cell_6t
Xbit_r3_c187 bl_187 br_187 wl_3 vdd gnd cell_6t
Xbit_r4_c187 bl_187 br_187 wl_4 vdd gnd cell_6t
Xbit_r5_c187 bl_187 br_187 wl_5 vdd gnd cell_6t
Xbit_r6_c187 bl_187 br_187 wl_6 vdd gnd cell_6t
Xbit_r7_c187 bl_187 br_187 wl_7 vdd gnd cell_6t
Xbit_r8_c187 bl_187 br_187 wl_8 vdd gnd cell_6t
Xbit_r9_c187 bl_187 br_187 wl_9 vdd gnd cell_6t
Xbit_r10_c187 bl_187 br_187 wl_10 vdd gnd cell_6t
Xbit_r11_c187 bl_187 br_187 wl_11 vdd gnd cell_6t
Xbit_r12_c187 bl_187 br_187 wl_12 vdd gnd cell_6t
Xbit_r13_c187 bl_187 br_187 wl_13 vdd gnd cell_6t
Xbit_r14_c187 bl_187 br_187 wl_14 vdd gnd cell_6t
Xbit_r15_c187 bl_187 br_187 wl_15 vdd gnd cell_6t
Xbit_r16_c187 bl_187 br_187 wl_16 vdd gnd cell_6t
Xbit_r17_c187 bl_187 br_187 wl_17 vdd gnd cell_6t
Xbit_r18_c187 bl_187 br_187 wl_18 vdd gnd cell_6t
Xbit_r19_c187 bl_187 br_187 wl_19 vdd gnd cell_6t
Xbit_r20_c187 bl_187 br_187 wl_20 vdd gnd cell_6t
Xbit_r21_c187 bl_187 br_187 wl_21 vdd gnd cell_6t
Xbit_r22_c187 bl_187 br_187 wl_22 vdd gnd cell_6t
Xbit_r23_c187 bl_187 br_187 wl_23 vdd gnd cell_6t
Xbit_r24_c187 bl_187 br_187 wl_24 vdd gnd cell_6t
Xbit_r25_c187 bl_187 br_187 wl_25 vdd gnd cell_6t
Xbit_r26_c187 bl_187 br_187 wl_26 vdd gnd cell_6t
Xbit_r27_c187 bl_187 br_187 wl_27 vdd gnd cell_6t
Xbit_r28_c187 bl_187 br_187 wl_28 vdd gnd cell_6t
Xbit_r29_c187 bl_187 br_187 wl_29 vdd gnd cell_6t
Xbit_r30_c187 bl_187 br_187 wl_30 vdd gnd cell_6t
Xbit_r31_c187 bl_187 br_187 wl_31 vdd gnd cell_6t
Xbit_r32_c187 bl_187 br_187 wl_32 vdd gnd cell_6t
Xbit_r33_c187 bl_187 br_187 wl_33 vdd gnd cell_6t
Xbit_r34_c187 bl_187 br_187 wl_34 vdd gnd cell_6t
Xbit_r35_c187 bl_187 br_187 wl_35 vdd gnd cell_6t
Xbit_r36_c187 bl_187 br_187 wl_36 vdd gnd cell_6t
Xbit_r37_c187 bl_187 br_187 wl_37 vdd gnd cell_6t
Xbit_r38_c187 bl_187 br_187 wl_38 vdd gnd cell_6t
Xbit_r39_c187 bl_187 br_187 wl_39 vdd gnd cell_6t
Xbit_r40_c187 bl_187 br_187 wl_40 vdd gnd cell_6t
Xbit_r41_c187 bl_187 br_187 wl_41 vdd gnd cell_6t
Xbit_r42_c187 bl_187 br_187 wl_42 vdd gnd cell_6t
Xbit_r43_c187 bl_187 br_187 wl_43 vdd gnd cell_6t
Xbit_r44_c187 bl_187 br_187 wl_44 vdd gnd cell_6t
Xbit_r45_c187 bl_187 br_187 wl_45 vdd gnd cell_6t
Xbit_r46_c187 bl_187 br_187 wl_46 vdd gnd cell_6t
Xbit_r47_c187 bl_187 br_187 wl_47 vdd gnd cell_6t
Xbit_r48_c187 bl_187 br_187 wl_48 vdd gnd cell_6t
Xbit_r49_c187 bl_187 br_187 wl_49 vdd gnd cell_6t
Xbit_r50_c187 bl_187 br_187 wl_50 vdd gnd cell_6t
Xbit_r51_c187 bl_187 br_187 wl_51 vdd gnd cell_6t
Xbit_r52_c187 bl_187 br_187 wl_52 vdd gnd cell_6t
Xbit_r53_c187 bl_187 br_187 wl_53 vdd gnd cell_6t
Xbit_r54_c187 bl_187 br_187 wl_54 vdd gnd cell_6t
Xbit_r55_c187 bl_187 br_187 wl_55 vdd gnd cell_6t
Xbit_r56_c187 bl_187 br_187 wl_56 vdd gnd cell_6t
Xbit_r57_c187 bl_187 br_187 wl_57 vdd gnd cell_6t
Xbit_r58_c187 bl_187 br_187 wl_58 vdd gnd cell_6t
Xbit_r59_c187 bl_187 br_187 wl_59 vdd gnd cell_6t
Xbit_r60_c187 bl_187 br_187 wl_60 vdd gnd cell_6t
Xbit_r61_c187 bl_187 br_187 wl_61 vdd gnd cell_6t
Xbit_r62_c187 bl_187 br_187 wl_62 vdd gnd cell_6t
Xbit_r63_c187 bl_187 br_187 wl_63 vdd gnd cell_6t
Xbit_r64_c187 bl_187 br_187 wl_64 vdd gnd cell_6t
Xbit_r65_c187 bl_187 br_187 wl_65 vdd gnd cell_6t
Xbit_r66_c187 bl_187 br_187 wl_66 vdd gnd cell_6t
Xbit_r67_c187 bl_187 br_187 wl_67 vdd gnd cell_6t
Xbit_r68_c187 bl_187 br_187 wl_68 vdd gnd cell_6t
Xbit_r69_c187 bl_187 br_187 wl_69 vdd gnd cell_6t
Xbit_r70_c187 bl_187 br_187 wl_70 vdd gnd cell_6t
Xbit_r71_c187 bl_187 br_187 wl_71 vdd gnd cell_6t
Xbit_r72_c187 bl_187 br_187 wl_72 vdd gnd cell_6t
Xbit_r73_c187 bl_187 br_187 wl_73 vdd gnd cell_6t
Xbit_r74_c187 bl_187 br_187 wl_74 vdd gnd cell_6t
Xbit_r75_c187 bl_187 br_187 wl_75 vdd gnd cell_6t
Xbit_r76_c187 bl_187 br_187 wl_76 vdd gnd cell_6t
Xbit_r77_c187 bl_187 br_187 wl_77 vdd gnd cell_6t
Xbit_r78_c187 bl_187 br_187 wl_78 vdd gnd cell_6t
Xbit_r79_c187 bl_187 br_187 wl_79 vdd gnd cell_6t
Xbit_r80_c187 bl_187 br_187 wl_80 vdd gnd cell_6t
Xbit_r81_c187 bl_187 br_187 wl_81 vdd gnd cell_6t
Xbit_r82_c187 bl_187 br_187 wl_82 vdd gnd cell_6t
Xbit_r83_c187 bl_187 br_187 wl_83 vdd gnd cell_6t
Xbit_r84_c187 bl_187 br_187 wl_84 vdd gnd cell_6t
Xbit_r85_c187 bl_187 br_187 wl_85 vdd gnd cell_6t
Xbit_r86_c187 bl_187 br_187 wl_86 vdd gnd cell_6t
Xbit_r87_c187 bl_187 br_187 wl_87 vdd gnd cell_6t
Xbit_r88_c187 bl_187 br_187 wl_88 vdd gnd cell_6t
Xbit_r89_c187 bl_187 br_187 wl_89 vdd gnd cell_6t
Xbit_r90_c187 bl_187 br_187 wl_90 vdd gnd cell_6t
Xbit_r91_c187 bl_187 br_187 wl_91 vdd gnd cell_6t
Xbit_r92_c187 bl_187 br_187 wl_92 vdd gnd cell_6t
Xbit_r93_c187 bl_187 br_187 wl_93 vdd gnd cell_6t
Xbit_r94_c187 bl_187 br_187 wl_94 vdd gnd cell_6t
Xbit_r95_c187 bl_187 br_187 wl_95 vdd gnd cell_6t
Xbit_r96_c187 bl_187 br_187 wl_96 vdd gnd cell_6t
Xbit_r97_c187 bl_187 br_187 wl_97 vdd gnd cell_6t
Xbit_r98_c187 bl_187 br_187 wl_98 vdd gnd cell_6t
Xbit_r99_c187 bl_187 br_187 wl_99 vdd gnd cell_6t
Xbit_r100_c187 bl_187 br_187 wl_100 vdd gnd cell_6t
Xbit_r101_c187 bl_187 br_187 wl_101 vdd gnd cell_6t
Xbit_r102_c187 bl_187 br_187 wl_102 vdd gnd cell_6t
Xbit_r103_c187 bl_187 br_187 wl_103 vdd gnd cell_6t
Xbit_r104_c187 bl_187 br_187 wl_104 vdd gnd cell_6t
Xbit_r105_c187 bl_187 br_187 wl_105 vdd gnd cell_6t
Xbit_r106_c187 bl_187 br_187 wl_106 vdd gnd cell_6t
Xbit_r107_c187 bl_187 br_187 wl_107 vdd gnd cell_6t
Xbit_r108_c187 bl_187 br_187 wl_108 vdd gnd cell_6t
Xbit_r109_c187 bl_187 br_187 wl_109 vdd gnd cell_6t
Xbit_r110_c187 bl_187 br_187 wl_110 vdd gnd cell_6t
Xbit_r111_c187 bl_187 br_187 wl_111 vdd gnd cell_6t
Xbit_r112_c187 bl_187 br_187 wl_112 vdd gnd cell_6t
Xbit_r113_c187 bl_187 br_187 wl_113 vdd gnd cell_6t
Xbit_r114_c187 bl_187 br_187 wl_114 vdd gnd cell_6t
Xbit_r115_c187 bl_187 br_187 wl_115 vdd gnd cell_6t
Xbit_r116_c187 bl_187 br_187 wl_116 vdd gnd cell_6t
Xbit_r117_c187 bl_187 br_187 wl_117 vdd gnd cell_6t
Xbit_r118_c187 bl_187 br_187 wl_118 vdd gnd cell_6t
Xbit_r119_c187 bl_187 br_187 wl_119 vdd gnd cell_6t
Xbit_r120_c187 bl_187 br_187 wl_120 vdd gnd cell_6t
Xbit_r121_c187 bl_187 br_187 wl_121 vdd gnd cell_6t
Xbit_r122_c187 bl_187 br_187 wl_122 vdd gnd cell_6t
Xbit_r123_c187 bl_187 br_187 wl_123 vdd gnd cell_6t
Xbit_r124_c187 bl_187 br_187 wl_124 vdd gnd cell_6t
Xbit_r125_c187 bl_187 br_187 wl_125 vdd gnd cell_6t
Xbit_r126_c187 bl_187 br_187 wl_126 vdd gnd cell_6t
Xbit_r127_c187 bl_187 br_187 wl_127 vdd gnd cell_6t
Xbit_r128_c187 bl_187 br_187 wl_128 vdd gnd cell_6t
Xbit_r129_c187 bl_187 br_187 wl_129 vdd gnd cell_6t
Xbit_r130_c187 bl_187 br_187 wl_130 vdd gnd cell_6t
Xbit_r131_c187 bl_187 br_187 wl_131 vdd gnd cell_6t
Xbit_r132_c187 bl_187 br_187 wl_132 vdd gnd cell_6t
Xbit_r133_c187 bl_187 br_187 wl_133 vdd gnd cell_6t
Xbit_r134_c187 bl_187 br_187 wl_134 vdd gnd cell_6t
Xbit_r135_c187 bl_187 br_187 wl_135 vdd gnd cell_6t
Xbit_r136_c187 bl_187 br_187 wl_136 vdd gnd cell_6t
Xbit_r137_c187 bl_187 br_187 wl_137 vdd gnd cell_6t
Xbit_r138_c187 bl_187 br_187 wl_138 vdd gnd cell_6t
Xbit_r139_c187 bl_187 br_187 wl_139 vdd gnd cell_6t
Xbit_r140_c187 bl_187 br_187 wl_140 vdd gnd cell_6t
Xbit_r141_c187 bl_187 br_187 wl_141 vdd gnd cell_6t
Xbit_r142_c187 bl_187 br_187 wl_142 vdd gnd cell_6t
Xbit_r143_c187 bl_187 br_187 wl_143 vdd gnd cell_6t
Xbit_r144_c187 bl_187 br_187 wl_144 vdd gnd cell_6t
Xbit_r145_c187 bl_187 br_187 wl_145 vdd gnd cell_6t
Xbit_r146_c187 bl_187 br_187 wl_146 vdd gnd cell_6t
Xbit_r147_c187 bl_187 br_187 wl_147 vdd gnd cell_6t
Xbit_r148_c187 bl_187 br_187 wl_148 vdd gnd cell_6t
Xbit_r149_c187 bl_187 br_187 wl_149 vdd gnd cell_6t
Xbit_r150_c187 bl_187 br_187 wl_150 vdd gnd cell_6t
Xbit_r151_c187 bl_187 br_187 wl_151 vdd gnd cell_6t
Xbit_r152_c187 bl_187 br_187 wl_152 vdd gnd cell_6t
Xbit_r153_c187 bl_187 br_187 wl_153 vdd gnd cell_6t
Xbit_r154_c187 bl_187 br_187 wl_154 vdd gnd cell_6t
Xbit_r155_c187 bl_187 br_187 wl_155 vdd gnd cell_6t
Xbit_r156_c187 bl_187 br_187 wl_156 vdd gnd cell_6t
Xbit_r157_c187 bl_187 br_187 wl_157 vdd gnd cell_6t
Xbit_r158_c187 bl_187 br_187 wl_158 vdd gnd cell_6t
Xbit_r159_c187 bl_187 br_187 wl_159 vdd gnd cell_6t
Xbit_r160_c187 bl_187 br_187 wl_160 vdd gnd cell_6t
Xbit_r161_c187 bl_187 br_187 wl_161 vdd gnd cell_6t
Xbit_r162_c187 bl_187 br_187 wl_162 vdd gnd cell_6t
Xbit_r163_c187 bl_187 br_187 wl_163 vdd gnd cell_6t
Xbit_r164_c187 bl_187 br_187 wl_164 vdd gnd cell_6t
Xbit_r165_c187 bl_187 br_187 wl_165 vdd gnd cell_6t
Xbit_r166_c187 bl_187 br_187 wl_166 vdd gnd cell_6t
Xbit_r167_c187 bl_187 br_187 wl_167 vdd gnd cell_6t
Xbit_r168_c187 bl_187 br_187 wl_168 vdd gnd cell_6t
Xbit_r169_c187 bl_187 br_187 wl_169 vdd gnd cell_6t
Xbit_r170_c187 bl_187 br_187 wl_170 vdd gnd cell_6t
Xbit_r171_c187 bl_187 br_187 wl_171 vdd gnd cell_6t
Xbit_r172_c187 bl_187 br_187 wl_172 vdd gnd cell_6t
Xbit_r173_c187 bl_187 br_187 wl_173 vdd gnd cell_6t
Xbit_r174_c187 bl_187 br_187 wl_174 vdd gnd cell_6t
Xbit_r175_c187 bl_187 br_187 wl_175 vdd gnd cell_6t
Xbit_r176_c187 bl_187 br_187 wl_176 vdd gnd cell_6t
Xbit_r177_c187 bl_187 br_187 wl_177 vdd gnd cell_6t
Xbit_r178_c187 bl_187 br_187 wl_178 vdd gnd cell_6t
Xbit_r179_c187 bl_187 br_187 wl_179 vdd gnd cell_6t
Xbit_r180_c187 bl_187 br_187 wl_180 vdd gnd cell_6t
Xbit_r181_c187 bl_187 br_187 wl_181 vdd gnd cell_6t
Xbit_r182_c187 bl_187 br_187 wl_182 vdd gnd cell_6t
Xbit_r183_c187 bl_187 br_187 wl_183 vdd gnd cell_6t
Xbit_r184_c187 bl_187 br_187 wl_184 vdd gnd cell_6t
Xbit_r185_c187 bl_187 br_187 wl_185 vdd gnd cell_6t
Xbit_r186_c187 bl_187 br_187 wl_186 vdd gnd cell_6t
Xbit_r187_c187 bl_187 br_187 wl_187 vdd gnd cell_6t
Xbit_r188_c187 bl_187 br_187 wl_188 vdd gnd cell_6t
Xbit_r189_c187 bl_187 br_187 wl_189 vdd gnd cell_6t
Xbit_r190_c187 bl_187 br_187 wl_190 vdd gnd cell_6t
Xbit_r191_c187 bl_187 br_187 wl_191 vdd gnd cell_6t
Xbit_r192_c187 bl_187 br_187 wl_192 vdd gnd cell_6t
Xbit_r193_c187 bl_187 br_187 wl_193 vdd gnd cell_6t
Xbit_r194_c187 bl_187 br_187 wl_194 vdd gnd cell_6t
Xbit_r195_c187 bl_187 br_187 wl_195 vdd gnd cell_6t
Xbit_r196_c187 bl_187 br_187 wl_196 vdd gnd cell_6t
Xbit_r197_c187 bl_187 br_187 wl_197 vdd gnd cell_6t
Xbit_r198_c187 bl_187 br_187 wl_198 vdd gnd cell_6t
Xbit_r199_c187 bl_187 br_187 wl_199 vdd gnd cell_6t
Xbit_r200_c187 bl_187 br_187 wl_200 vdd gnd cell_6t
Xbit_r201_c187 bl_187 br_187 wl_201 vdd gnd cell_6t
Xbit_r202_c187 bl_187 br_187 wl_202 vdd gnd cell_6t
Xbit_r203_c187 bl_187 br_187 wl_203 vdd gnd cell_6t
Xbit_r204_c187 bl_187 br_187 wl_204 vdd gnd cell_6t
Xbit_r205_c187 bl_187 br_187 wl_205 vdd gnd cell_6t
Xbit_r206_c187 bl_187 br_187 wl_206 vdd gnd cell_6t
Xbit_r207_c187 bl_187 br_187 wl_207 vdd gnd cell_6t
Xbit_r208_c187 bl_187 br_187 wl_208 vdd gnd cell_6t
Xbit_r209_c187 bl_187 br_187 wl_209 vdd gnd cell_6t
Xbit_r210_c187 bl_187 br_187 wl_210 vdd gnd cell_6t
Xbit_r211_c187 bl_187 br_187 wl_211 vdd gnd cell_6t
Xbit_r212_c187 bl_187 br_187 wl_212 vdd gnd cell_6t
Xbit_r213_c187 bl_187 br_187 wl_213 vdd gnd cell_6t
Xbit_r214_c187 bl_187 br_187 wl_214 vdd gnd cell_6t
Xbit_r215_c187 bl_187 br_187 wl_215 vdd gnd cell_6t
Xbit_r216_c187 bl_187 br_187 wl_216 vdd gnd cell_6t
Xbit_r217_c187 bl_187 br_187 wl_217 vdd gnd cell_6t
Xbit_r218_c187 bl_187 br_187 wl_218 vdd gnd cell_6t
Xbit_r219_c187 bl_187 br_187 wl_219 vdd gnd cell_6t
Xbit_r220_c187 bl_187 br_187 wl_220 vdd gnd cell_6t
Xbit_r221_c187 bl_187 br_187 wl_221 vdd gnd cell_6t
Xbit_r222_c187 bl_187 br_187 wl_222 vdd gnd cell_6t
Xbit_r223_c187 bl_187 br_187 wl_223 vdd gnd cell_6t
Xbit_r224_c187 bl_187 br_187 wl_224 vdd gnd cell_6t
Xbit_r225_c187 bl_187 br_187 wl_225 vdd gnd cell_6t
Xbit_r226_c187 bl_187 br_187 wl_226 vdd gnd cell_6t
Xbit_r227_c187 bl_187 br_187 wl_227 vdd gnd cell_6t
Xbit_r228_c187 bl_187 br_187 wl_228 vdd gnd cell_6t
Xbit_r229_c187 bl_187 br_187 wl_229 vdd gnd cell_6t
Xbit_r230_c187 bl_187 br_187 wl_230 vdd gnd cell_6t
Xbit_r231_c187 bl_187 br_187 wl_231 vdd gnd cell_6t
Xbit_r232_c187 bl_187 br_187 wl_232 vdd gnd cell_6t
Xbit_r233_c187 bl_187 br_187 wl_233 vdd gnd cell_6t
Xbit_r234_c187 bl_187 br_187 wl_234 vdd gnd cell_6t
Xbit_r235_c187 bl_187 br_187 wl_235 vdd gnd cell_6t
Xbit_r236_c187 bl_187 br_187 wl_236 vdd gnd cell_6t
Xbit_r237_c187 bl_187 br_187 wl_237 vdd gnd cell_6t
Xbit_r238_c187 bl_187 br_187 wl_238 vdd gnd cell_6t
Xbit_r239_c187 bl_187 br_187 wl_239 vdd gnd cell_6t
Xbit_r240_c187 bl_187 br_187 wl_240 vdd gnd cell_6t
Xbit_r241_c187 bl_187 br_187 wl_241 vdd gnd cell_6t
Xbit_r242_c187 bl_187 br_187 wl_242 vdd gnd cell_6t
Xbit_r243_c187 bl_187 br_187 wl_243 vdd gnd cell_6t
Xbit_r244_c187 bl_187 br_187 wl_244 vdd gnd cell_6t
Xbit_r245_c187 bl_187 br_187 wl_245 vdd gnd cell_6t
Xbit_r246_c187 bl_187 br_187 wl_246 vdd gnd cell_6t
Xbit_r247_c187 bl_187 br_187 wl_247 vdd gnd cell_6t
Xbit_r248_c187 bl_187 br_187 wl_248 vdd gnd cell_6t
Xbit_r249_c187 bl_187 br_187 wl_249 vdd gnd cell_6t
Xbit_r250_c187 bl_187 br_187 wl_250 vdd gnd cell_6t
Xbit_r251_c187 bl_187 br_187 wl_251 vdd gnd cell_6t
Xbit_r252_c187 bl_187 br_187 wl_252 vdd gnd cell_6t
Xbit_r253_c187 bl_187 br_187 wl_253 vdd gnd cell_6t
Xbit_r254_c187 bl_187 br_187 wl_254 vdd gnd cell_6t
Xbit_r255_c187 bl_187 br_187 wl_255 vdd gnd cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd cell_6t
Xbit_r1_c188 bl_188 br_188 wl_1 vdd gnd cell_6t
Xbit_r2_c188 bl_188 br_188 wl_2 vdd gnd cell_6t
Xbit_r3_c188 bl_188 br_188 wl_3 vdd gnd cell_6t
Xbit_r4_c188 bl_188 br_188 wl_4 vdd gnd cell_6t
Xbit_r5_c188 bl_188 br_188 wl_5 vdd gnd cell_6t
Xbit_r6_c188 bl_188 br_188 wl_6 vdd gnd cell_6t
Xbit_r7_c188 bl_188 br_188 wl_7 vdd gnd cell_6t
Xbit_r8_c188 bl_188 br_188 wl_8 vdd gnd cell_6t
Xbit_r9_c188 bl_188 br_188 wl_9 vdd gnd cell_6t
Xbit_r10_c188 bl_188 br_188 wl_10 vdd gnd cell_6t
Xbit_r11_c188 bl_188 br_188 wl_11 vdd gnd cell_6t
Xbit_r12_c188 bl_188 br_188 wl_12 vdd gnd cell_6t
Xbit_r13_c188 bl_188 br_188 wl_13 vdd gnd cell_6t
Xbit_r14_c188 bl_188 br_188 wl_14 vdd gnd cell_6t
Xbit_r15_c188 bl_188 br_188 wl_15 vdd gnd cell_6t
Xbit_r16_c188 bl_188 br_188 wl_16 vdd gnd cell_6t
Xbit_r17_c188 bl_188 br_188 wl_17 vdd gnd cell_6t
Xbit_r18_c188 bl_188 br_188 wl_18 vdd gnd cell_6t
Xbit_r19_c188 bl_188 br_188 wl_19 vdd gnd cell_6t
Xbit_r20_c188 bl_188 br_188 wl_20 vdd gnd cell_6t
Xbit_r21_c188 bl_188 br_188 wl_21 vdd gnd cell_6t
Xbit_r22_c188 bl_188 br_188 wl_22 vdd gnd cell_6t
Xbit_r23_c188 bl_188 br_188 wl_23 vdd gnd cell_6t
Xbit_r24_c188 bl_188 br_188 wl_24 vdd gnd cell_6t
Xbit_r25_c188 bl_188 br_188 wl_25 vdd gnd cell_6t
Xbit_r26_c188 bl_188 br_188 wl_26 vdd gnd cell_6t
Xbit_r27_c188 bl_188 br_188 wl_27 vdd gnd cell_6t
Xbit_r28_c188 bl_188 br_188 wl_28 vdd gnd cell_6t
Xbit_r29_c188 bl_188 br_188 wl_29 vdd gnd cell_6t
Xbit_r30_c188 bl_188 br_188 wl_30 vdd gnd cell_6t
Xbit_r31_c188 bl_188 br_188 wl_31 vdd gnd cell_6t
Xbit_r32_c188 bl_188 br_188 wl_32 vdd gnd cell_6t
Xbit_r33_c188 bl_188 br_188 wl_33 vdd gnd cell_6t
Xbit_r34_c188 bl_188 br_188 wl_34 vdd gnd cell_6t
Xbit_r35_c188 bl_188 br_188 wl_35 vdd gnd cell_6t
Xbit_r36_c188 bl_188 br_188 wl_36 vdd gnd cell_6t
Xbit_r37_c188 bl_188 br_188 wl_37 vdd gnd cell_6t
Xbit_r38_c188 bl_188 br_188 wl_38 vdd gnd cell_6t
Xbit_r39_c188 bl_188 br_188 wl_39 vdd gnd cell_6t
Xbit_r40_c188 bl_188 br_188 wl_40 vdd gnd cell_6t
Xbit_r41_c188 bl_188 br_188 wl_41 vdd gnd cell_6t
Xbit_r42_c188 bl_188 br_188 wl_42 vdd gnd cell_6t
Xbit_r43_c188 bl_188 br_188 wl_43 vdd gnd cell_6t
Xbit_r44_c188 bl_188 br_188 wl_44 vdd gnd cell_6t
Xbit_r45_c188 bl_188 br_188 wl_45 vdd gnd cell_6t
Xbit_r46_c188 bl_188 br_188 wl_46 vdd gnd cell_6t
Xbit_r47_c188 bl_188 br_188 wl_47 vdd gnd cell_6t
Xbit_r48_c188 bl_188 br_188 wl_48 vdd gnd cell_6t
Xbit_r49_c188 bl_188 br_188 wl_49 vdd gnd cell_6t
Xbit_r50_c188 bl_188 br_188 wl_50 vdd gnd cell_6t
Xbit_r51_c188 bl_188 br_188 wl_51 vdd gnd cell_6t
Xbit_r52_c188 bl_188 br_188 wl_52 vdd gnd cell_6t
Xbit_r53_c188 bl_188 br_188 wl_53 vdd gnd cell_6t
Xbit_r54_c188 bl_188 br_188 wl_54 vdd gnd cell_6t
Xbit_r55_c188 bl_188 br_188 wl_55 vdd gnd cell_6t
Xbit_r56_c188 bl_188 br_188 wl_56 vdd gnd cell_6t
Xbit_r57_c188 bl_188 br_188 wl_57 vdd gnd cell_6t
Xbit_r58_c188 bl_188 br_188 wl_58 vdd gnd cell_6t
Xbit_r59_c188 bl_188 br_188 wl_59 vdd gnd cell_6t
Xbit_r60_c188 bl_188 br_188 wl_60 vdd gnd cell_6t
Xbit_r61_c188 bl_188 br_188 wl_61 vdd gnd cell_6t
Xbit_r62_c188 bl_188 br_188 wl_62 vdd gnd cell_6t
Xbit_r63_c188 bl_188 br_188 wl_63 vdd gnd cell_6t
Xbit_r64_c188 bl_188 br_188 wl_64 vdd gnd cell_6t
Xbit_r65_c188 bl_188 br_188 wl_65 vdd gnd cell_6t
Xbit_r66_c188 bl_188 br_188 wl_66 vdd gnd cell_6t
Xbit_r67_c188 bl_188 br_188 wl_67 vdd gnd cell_6t
Xbit_r68_c188 bl_188 br_188 wl_68 vdd gnd cell_6t
Xbit_r69_c188 bl_188 br_188 wl_69 vdd gnd cell_6t
Xbit_r70_c188 bl_188 br_188 wl_70 vdd gnd cell_6t
Xbit_r71_c188 bl_188 br_188 wl_71 vdd gnd cell_6t
Xbit_r72_c188 bl_188 br_188 wl_72 vdd gnd cell_6t
Xbit_r73_c188 bl_188 br_188 wl_73 vdd gnd cell_6t
Xbit_r74_c188 bl_188 br_188 wl_74 vdd gnd cell_6t
Xbit_r75_c188 bl_188 br_188 wl_75 vdd gnd cell_6t
Xbit_r76_c188 bl_188 br_188 wl_76 vdd gnd cell_6t
Xbit_r77_c188 bl_188 br_188 wl_77 vdd gnd cell_6t
Xbit_r78_c188 bl_188 br_188 wl_78 vdd gnd cell_6t
Xbit_r79_c188 bl_188 br_188 wl_79 vdd gnd cell_6t
Xbit_r80_c188 bl_188 br_188 wl_80 vdd gnd cell_6t
Xbit_r81_c188 bl_188 br_188 wl_81 vdd gnd cell_6t
Xbit_r82_c188 bl_188 br_188 wl_82 vdd gnd cell_6t
Xbit_r83_c188 bl_188 br_188 wl_83 vdd gnd cell_6t
Xbit_r84_c188 bl_188 br_188 wl_84 vdd gnd cell_6t
Xbit_r85_c188 bl_188 br_188 wl_85 vdd gnd cell_6t
Xbit_r86_c188 bl_188 br_188 wl_86 vdd gnd cell_6t
Xbit_r87_c188 bl_188 br_188 wl_87 vdd gnd cell_6t
Xbit_r88_c188 bl_188 br_188 wl_88 vdd gnd cell_6t
Xbit_r89_c188 bl_188 br_188 wl_89 vdd gnd cell_6t
Xbit_r90_c188 bl_188 br_188 wl_90 vdd gnd cell_6t
Xbit_r91_c188 bl_188 br_188 wl_91 vdd gnd cell_6t
Xbit_r92_c188 bl_188 br_188 wl_92 vdd gnd cell_6t
Xbit_r93_c188 bl_188 br_188 wl_93 vdd gnd cell_6t
Xbit_r94_c188 bl_188 br_188 wl_94 vdd gnd cell_6t
Xbit_r95_c188 bl_188 br_188 wl_95 vdd gnd cell_6t
Xbit_r96_c188 bl_188 br_188 wl_96 vdd gnd cell_6t
Xbit_r97_c188 bl_188 br_188 wl_97 vdd gnd cell_6t
Xbit_r98_c188 bl_188 br_188 wl_98 vdd gnd cell_6t
Xbit_r99_c188 bl_188 br_188 wl_99 vdd gnd cell_6t
Xbit_r100_c188 bl_188 br_188 wl_100 vdd gnd cell_6t
Xbit_r101_c188 bl_188 br_188 wl_101 vdd gnd cell_6t
Xbit_r102_c188 bl_188 br_188 wl_102 vdd gnd cell_6t
Xbit_r103_c188 bl_188 br_188 wl_103 vdd gnd cell_6t
Xbit_r104_c188 bl_188 br_188 wl_104 vdd gnd cell_6t
Xbit_r105_c188 bl_188 br_188 wl_105 vdd gnd cell_6t
Xbit_r106_c188 bl_188 br_188 wl_106 vdd gnd cell_6t
Xbit_r107_c188 bl_188 br_188 wl_107 vdd gnd cell_6t
Xbit_r108_c188 bl_188 br_188 wl_108 vdd gnd cell_6t
Xbit_r109_c188 bl_188 br_188 wl_109 vdd gnd cell_6t
Xbit_r110_c188 bl_188 br_188 wl_110 vdd gnd cell_6t
Xbit_r111_c188 bl_188 br_188 wl_111 vdd gnd cell_6t
Xbit_r112_c188 bl_188 br_188 wl_112 vdd gnd cell_6t
Xbit_r113_c188 bl_188 br_188 wl_113 vdd gnd cell_6t
Xbit_r114_c188 bl_188 br_188 wl_114 vdd gnd cell_6t
Xbit_r115_c188 bl_188 br_188 wl_115 vdd gnd cell_6t
Xbit_r116_c188 bl_188 br_188 wl_116 vdd gnd cell_6t
Xbit_r117_c188 bl_188 br_188 wl_117 vdd gnd cell_6t
Xbit_r118_c188 bl_188 br_188 wl_118 vdd gnd cell_6t
Xbit_r119_c188 bl_188 br_188 wl_119 vdd gnd cell_6t
Xbit_r120_c188 bl_188 br_188 wl_120 vdd gnd cell_6t
Xbit_r121_c188 bl_188 br_188 wl_121 vdd gnd cell_6t
Xbit_r122_c188 bl_188 br_188 wl_122 vdd gnd cell_6t
Xbit_r123_c188 bl_188 br_188 wl_123 vdd gnd cell_6t
Xbit_r124_c188 bl_188 br_188 wl_124 vdd gnd cell_6t
Xbit_r125_c188 bl_188 br_188 wl_125 vdd gnd cell_6t
Xbit_r126_c188 bl_188 br_188 wl_126 vdd gnd cell_6t
Xbit_r127_c188 bl_188 br_188 wl_127 vdd gnd cell_6t
Xbit_r128_c188 bl_188 br_188 wl_128 vdd gnd cell_6t
Xbit_r129_c188 bl_188 br_188 wl_129 vdd gnd cell_6t
Xbit_r130_c188 bl_188 br_188 wl_130 vdd gnd cell_6t
Xbit_r131_c188 bl_188 br_188 wl_131 vdd gnd cell_6t
Xbit_r132_c188 bl_188 br_188 wl_132 vdd gnd cell_6t
Xbit_r133_c188 bl_188 br_188 wl_133 vdd gnd cell_6t
Xbit_r134_c188 bl_188 br_188 wl_134 vdd gnd cell_6t
Xbit_r135_c188 bl_188 br_188 wl_135 vdd gnd cell_6t
Xbit_r136_c188 bl_188 br_188 wl_136 vdd gnd cell_6t
Xbit_r137_c188 bl_188 br_188 wl_137 vdd gnd cell_6t
Xbit_r138_c188 bl_188 br_188 wl_138 vdd gnd cell_6t
Xbit_r139_c188 bl_188 br_188 wl_139 vdd gnd cell_6t
Xbit_r140_c188 bl_188 br_188 wl_140 vdd gnd cell_6t
Xbit_r141_c188 bl_188 br_188 wl_141 vdd gnd cell_6t
Xbit_r142_c188 bl_188 br_188 wl_142 vdd gnd cell_6t
Xbit_r143_c188 bl_188 br_188 wl_143 vdd gnd cell_6t
Xbit_r144_c188 bl_188 br_188 wl_144 vdd gnd cell_6t
Xbit_r145_c188 bl_188 br_188 wl_145 vdd gnd cell_6t
Xbit_r146_c188 bl_188 br_188 wl_146 vdd gnd cell_6t
Xbit_r147_c188 bl_188 br_188 wl_147 vdd gnd cell_6t
Xbit_r148_c188 bl_188 br_188 wl_148 vdd gnd cell_6t
Xbit_r149_c188 bl_188 br_188 wl_149 vdd gnd cell_6t
Xbit_r150_c188 bl_188 br_188 wl_150 vdd gnd cell_6t
Xbit_r151_c188 bl_188 br_188 wl_151 vdd gnd cell_6t
Xbit_r152_c188 bl_188 br_188 wl_152 vdd gnd cell_6t
Xbit_r153_c188 bl_188 br_188 wl_153 vdd gnd cell_6t
Xbit_r154_c188 bl_188 br_188 wl_154 vdd gnd cell_6t
Xbit_r155_c188 bl_188 br_188 wl_155 vdd gnd cell_6t
Xbit_r156_c188 bl_188 br_188 wl_156 vdd gnd cell_6t
Xbit_r157_c188 bl_188 br_188 wl_157 vdd gnd cell_6t
Xbit_r158_c188 bl_188 br_188 wl_158 vdd gnd cell_6t
Xbit_r159_c188 bl_188 br_188 wl_159 vdd gnd cell_6t
Xbit_r160_c188 bl_188 br_188 wl_160 vdd gnd cell_6t
Xbit_r161_c188 bl_188 br_188 wl_161 vdd gnd cell_6t
Xbit_r162_c188 bl_188 br_188 wl_162 vdd gnd cell_6t
Xbit_r163_c188 bl_188 br_188 wl_163 vdd gnd cell_6t
Xbit_r164_c188 bl_188 br_188 wl_164 vdd gnd cell_6t
Xbit_r165_c188 bl_188 br_188 wl_165 vdd gnd cell_6t
Xbit_r166_c188 bl_188 br_188 wl_166 vdd gnd cell_6t
Xbit_r167_c188 bl_188 br_188 wl_167 vdd gnd cell_6t
Xbit_r168_c188 bl_188 br_188 wl_168 vdd gnd cell_6t
Xbit_r169_c188 bl_188 br_188 wl_169 vdd gnd cell_6t
Xbit_r170_c188 bl_188 br_188 wl_170 vdd gnd cell_6t
Xbit_r171_c188 bl_188 br_188 wl_171 vdd gnd cell_6t
Xbit_r172_c188 bl_188 br_188 wl_172 vdd gnd cell_6t
Xbit_r173_c188 bl_188 br_188 wl_173 vdd gnd cell_6t
Xbit_r174_c188 bl_188 br_188 wl_174 vdd gnd cell_6t
Xbit_r175_c188 bl_188 br_188 wl_175 vdd gnd cell_6t
Xbit_r176_c188 bl_188 br_188 wl_176 vdd gnd cell_6t
Xbit_r177_c188 bl_188 br_188 wl_177 vdd gnd cell_6t
Xbit_r178_c188 bl_188 br_188 wl_178 vdd gnd cell_6t
Xbit_r179_c188 bl_188 br_188 wl_179 vdd gnd cell_6t
Xbit_r180_c188 bl_188 br_188 wl_180 vdd gnd cell_6t
Xbit_r181_c188 bl_188 br_188 wl_181 vdd gnd cell_6t
Xbit_r182_c188 bl_188 br_188 wl_182 vdd gnd cell_6t
Xbit_r183_c188 bl_188 br_188 wl_183 vdd gnd cell_6t
Xbit_r184_c188 bl_188 br_188 wl_184 vdd gnd cell_6t
Xbit_r185_c188 bl_188 br_188 wl_185 vdd gnd cell_6t
Xbit_r186_c188 bl_188 br_188 wl_186 vdd gnd cell_6t
Xbit_r187_c188 bl_188 br_188 wl_187 vdd gnd cell_6t
Xbit_r188_c188 bl_188 br_188 wl_188 vdd gnd cell_6t
Xbit_r189_c188 bl_188 br_188 wl_189 vdd gnd cell_6t
Xbit_r190_c188 bl_188 br_188 wl_190 vdd gnd cell_6t
Xbit_r191_c188 bl_188 br_188 wl_191 vdd gnd cell_6t
Xbit_r192_c188 bl_188 br_188 wl_192 vdd gnd cell_6t
Xbit_r193_c188 bl_188 br_188 wl_193 vdd gnd cell_6t
Xbit_r194_c188 bl_188 br_188 wl_194 vdd gnd cell_6t
Xbit_r195_c188 bl_188 br_188 wl_195 vdd gnd cell_6t
Xbit_r196_c188 bl_188 br_188 wl_196 vdd gnd cell_6t
Xbit_r197_c188 bl_188 br_188 wl_197 vdd gnd cell_6t
Xbit_r198_c188 bl_188 br_188 wl_198 vdd gnd cell_6t
Xbit_r199_c188 bl_188 br_188 wl_199 vdd gnd cell_6t
Xbit_r200_c188 bl_188 br_188 wl_200 vdd gnd cell_6t
Xbit_r201_c188 bl_188 br_188 wl_201 vdd gnd cell_6t
Xbit_r202_c188 bl_188 br_188 wl_202 vdd gnd cell_6t
Xbit_r203_c188 bl_188 br_188 wl_203 vdd gnd cell_6t
Xbit_r204_c188 bl_188 br_188 wl_204 vdd gnd cell_6t
Xbit_r205_c188 bl_188 br_188 wl_205 vdd gnd cell_6t
Xbit_r206_c188 bl_188 br_188 wl_206 vdd gnd cell_6t
Xbit_r207_c188 bl_188 br_188 wl_207 vdd gnd cell_6t
Xbit_r208_c188 bl_188 br_188 wl_208 vdd gnd cell_6t
Xbit_r209_c188 bl_188 br_188 wl_209 vdd gnd cell_6t
Xbit_r210_c188 bl_188 br_188 wl_210 vdd gnd cell_6t
Xbit_r211_c188 bl_188 br_188 wl_211 vdd gnd cell_6t
Xbit_r212_c188 bl_188 br_188 wl_212 vdd gnd cell_6t
Xbit_r213_c188 bl_188 br_188 wl_213 vdd gnd cell_6t
Xbit_r214_c188 bl_188 br_188 wl_214 vdd gnd cell_6t
Xbit_r215_c188 bl_188 br_188 wl_215 vdd gnd cell_6t
Xbit_r216_c188 bl_188 br_188 wl_216 vdd gnd cell_6t
Xbit_r217_c188 bl_188 br_188 wl_217 vdd gnd cell_6t
Xbit_r218_c188 bl_188 br_188 wl_218 vdd gnd cell_6t
Xbit_r219_c188 bl_188 br_188 wl_219 vdd gnd cell_6t
Xbit_r220_c188 bl_188 br_188 wl_220 vdd gnd cell_6t
Xbit_r221_c188 bl_188 br_188 wl_221 vdd gnd cell_6t
Xbit_r222_c188 bl_188 br_188 wl_222 vdd gnd cell_6t
Xbit_r223_c188 bl_188 br_188 wl_223 vdd gnd cell_6t
Xbit_r224_c188 bl_188 br_188 wl_224 vdd gnd cell_6t
Xbit_r225_c188 bl_188 br_188 wl_225 vdd gnd cell_6t
Xbit_r226_c188 bl_188 br_188 wl_226 vdd gnd cell_6t
Xbit_r227_c188 bl_188 br_188 wl_227 vdd gnd cell_6t
Xbit_r228_c188 bl_188 br_188 wl_228 vdd gnd cell_6t
Xbit_r229_c188 bl_188 br_188 wl_229 vdd gnd cell_6t
Xbit_r230_c188 bl_188 br_188 wl_230 vdd gnd cell_6t
Xbit_r231_c188 bl_188 br_188 wl_231 vdd gnd cell_6t
Xbit_r232_c188 bl_188 br_188 wl_232 vdd gnd cell_6t
Xbit_r233_c188 bl_188 br_188 wl_233 vdd gnd cell_6t
Xbit_r234_c188 bl_188 br_188 wl_234 vdd gnd cell_6t
Xbit_r235_c188 bl_188 br_188 wl_235 vdd gnd cell_6t
Xbit_r236_c188 bl_188 br_188 wl_236 vdd gnd cell_6t
Xbit_r237_c188 bl_188 br_188 wl_237 vdd gnd cell_6t
Xbit_r238_c188 bl_188 br_188 wl_238 vdd gnd cell_6t
Xbit_r239_c188 bl_188 br_188 wl_239 vdd gnd cell_6t
Xbit_r240_c188 bl_188 br_188 wl_240 vdd gnd cell_6t
Xbit_r241_c188 bl_188 br_188 wl_241 vdd gnd cell_6t
Xbit_r242_c188 bl_188 br_188 wl_242 vdd gnd cell_6t
Xbit_r243_c188 bl_188 br_188 wl_243 vdd gnd cell_6t
Xbit_r244_c188 bl_188 br_188 wl_244 vdd gnd cell_6t
Xbit_r245_c188 bl_188 br_188 wl_245 vdd gnd cell_6t
Xbit_r246_c188 bl_188 br_188 wl_246 vdd gnd cell_6t
Xbit_r247_c188 bl_188 br_188 wl_247 vdd gnd cell_6t
Xbit_r248_c188 bl_188 br_188 wl_248 vdd gnd cell_6t
Xbit_r249_c188 bl_188 br_188 wl_249 vdd gnd cell_6t
Xbit_r250_c188 bl_188 br_188 wl_250 vdd gnd cell_6t
Xbit_r251_c188 bl_188 br_188 wl_251 vdd gnd cell_6t
Xbit_r252_c188 bl_188 br_188 wl_252 vdd gnd cell_6t
Xbit_r253_c188 bl_188 br_188 wl_253 vdd gnd cell_6t
Xbit_r254_c188 bl_188 br_188 wl_254 vdd gnd cell_6t
Xbit_r255_c188 bl_188 br_188 wl_255 vdd gnd cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd cell_6t
Xbit_r1_c189 bl_189 br_189 wl_1 vdd gnd cell_6t
Xbit_r2_c189 bl_189 br_189 wl_2 vdd gnd cell_6t
Xbit_r3_c189 bl_189 br_189 wl_3 vdd gnd cell_6t
Xbit_r4_c189 bl_189 br_189 wl_4 vdd gnd cell_6t
Xbit_r5_c189 bl_189 br_189 wl_5 vdd gnd cell_6t
Xbit_r6_c189 bl_189 br_189 wl_6 vdd gnd cell_6t
Xbit_r7_c189 bl_189 br_189 wl_7 vdd gnd cell_6t
Xbit_r8_c189 bl_189 br_189 wl_8 vdd gnd cell_6t
Xbit_r9_c189 bl_189 br_189 wl_9 vdd gnd cell_6t
Xbit_r10_c189 bl_189 br_189 wl_10 vdd gnd cell_6t
Xbit_r11_c189 bl_189 br_189 wl_11 vdd gnd cell_6t
Xbit_r12_c189 bl_189 br_189 wl_12 vdd gnd cell_6t
Xbit_r13_c189 bl_189 br_189 wl_13 vdd gnd cell_6t
Xbit_r14_c189 bl_189 br_189 wl_14 vdd gnd cell_6t
Xbit_r15_c189 bl_189 br_189 wl_15 vdd gnd cell_6t
Xbit_r16_c189 bl_189 br_189 wl_16 vdd gnd cell_6t
Xbit_r17_c189 bl_189 br_189 wl_17 vdd gnd cell_6t
Xbit_r18_c189 bl_189 br_189 wl_18 vdd gnd cell_6t
Xbit_r19_c189 bl_189 br_189 wl_19 vdd gnd cell_6t
Xbit_r20_c189 bl_189 br_189 wl_20 vdd gnd cell_6t
Xbit_r21_c189 bl_189 br_189 wl_21 vdd gnd cell_6t
Xbit_r22_c189 bl_189 br_189 wl_22 vdd gnd cell_6t
Xbit_r23_c189 bl_189 br_189 wl_23 vdd gnd cell_6t
Xbit_r24_c189 bl_189 br_189 wl_24 vdd gnd cell_6t
Xbit_r25_c189 bl_189 br_189 wl_25 vdd gnd cell_6t
Xbit_r26_c189 bl_189 br_189 wl_26 vdd gnd cell_6t
Xbit_r27_c189 bl_189 br_189 wl_27 vdd gnd cell_6t
Xbit_r28_c189 bl_189 br_189 wl_28 vdd gnd cell_6t
Xbit_r29_c189 bl_189 br_189 wl_29 vdd gnd cell_6t
Xbit_r30_c189 bl_189 br_189 wl_30 vdd gnd cell_6t
Xbit_r31_c189 bl_189 br_189 wl_31 vdd gnd cell_6t
Xbit_r32_c189 bl_189 br_189 wl_32 vdd gnd cell_6t
Xbit_r33_c189 bl_189 br_189 wl_33 vdd gnd cell_6t
Xbit_r34_c189 bl_189 br_189 wl_34 vdd gnd cell_6t
Xbit_r35_c189 bl_189 br_189 wl_35 vdd gnd cell_6t
Xbit_r36_c189 bl_189 br_189 wl_36 vdd gnd cell_6t
Xbit_r37_c189 bl_189 br_189 wl_37 vdd gnd cell_6t
Xbit_r38_c189 bl_189 br_189 wl_38 vdd gnd cell_6t
Xbit_r39_c189 bl_189 br_189 wl_39 vdd gnd cell_6t
Xbit_r40_c189 bl_189 br_189 wl_40 vdd gnd cell_6t
Xbit_r41_c189 bl_189 br_189 wl_41 vdd gnd cell_6t
Xbit_r42_c189 bl_189 br_189 wl_42 vdd gnd cell_6t
Xbit_r43_c189 bl_189 br_189 wl_43 vdd gnd cell_6t
Xbit_r44_c189 bl_189 br_189 wl_44 vdd gnd cell_6t
Xbit_r45_c189 bl_189 br_189 wl_45 vdd gnd cell_6t
Xbit_r46_c189 bl_189 br_189 wl_46 vdd gnd cell_6t
Xbit_r47_c189 bl_189 br_189 wl_47 vdd gnd cell_6t
Xbit_r48_c189 bl_189 br_189 wl_48 vdd gnd cell_6t
Xbit_r49_c189 bl_189 br_189 wl_49 vdd gnd cell_6t
Xbit_r50_c189 bl_189 br_189 wl_50 vdd gnd cell_6t
Xbit_r51_c189 bl_189 br_189 wl_51 vdd gnd cell_6t
Xbit_r52_c189 bl_189 br_189 wl_52 vdd gnd cell_6t
Xbit_r53_c189 bl_189 br_189 wl_53 vdd gnd cell_6t
Xbit_r54_c189 bl_189 br_189 wl_54 vdd gnd cell_6t
Xbit_r55_c189 bl_189 br_189 wl_55 vdd gnd cell_6t
Xbit_r56_c189 bl_189 br_189 wl_56 vdd gnd cell_6t
Xbit_r57_c189 bl_189 br_189 wl_57 vdd gnd cell_6t
Xbit_r58_c189 bl_189 br_189 wl_58 vdd gnd cell_6t
Xbit_r59_c189 bl_189 br_189 wl_59 vdd gnd cell_6t
Xbit_r60_c189 bl_189 br_189 wl_60 vdd gnd cell_6t
Xbit_r61_c189 bl_189 br_189 wl_61 vdd gnd cell_6t
Xbit_r62_c189 bl_189 br_189 wl_62 vdd gnd cell_6t
Xbit_r63_c189 bl_189 br_189 wl_63 vdd gnd cell_6t
Xbit_r64_c189 bl_189 br_189 wl_64 vdd gnd cell_6t
Xbit_r65_c189 bl_189 br_189 wl_65 vdd gnd cell_6t
Xbit_r66_c189 bl_189 br_189 wl_66 vdd gnd cell_6t
Xbit_r67_c189 bl_189 br_189 wl_67 vdd gnd cell_6t
Xbit_r68_c189 bl_189 br_189 wl_68 vdd gnd cell_6t
Xbit_r69_c189 bl_189 br_189 wl_69 vdd gnd cell_6t
Xbit_r70_c189 bl_189 br_189 wl_70 vdd gnd cell_6t
Xbit_r71_c189 bl_189 br_189 wl_71 vdd gnd cell_6t
Xbit_r72_c189 bl_189 br_189 wl_72 vdd gnd cell_6t
Xbit_r73_c189 bl_189 br_189 wl_73 vdd gnd cell_6t
Xbit_r74_c189 bl_189 br_189 wl_74 vdd gnd cell_6t
Xbit_r75_c189 bl_189 br_189 wl_75 vdd gnd cell_6t
Xbit_r76_c189 bl_189 br_189 wl_76 vdd gnd cell_6t
Xbit_r77_c189 bl_189 br_189 wl_77 vdd gnd cell_6t
Xbit_r78_c189 bl_189 br_189 wl_78 vdd gnd cell_6t
Xbit_r79_c189 bl_189 br_189 wl_79 vdd gnd cell_6t
Xbit_r80_c189 bl_189 br_189 wl_80 vdd gnd cell_6t
Xbit_r81_c189 bl_189 br_189 wl_81 vdd gnd cell_6t
Xbit_r82_c189 bl_189 br_189 wl_82 vdd gnd cell_6t
Xbit_r83_c189 bl_189 br_189 wl_83 vdd gnd cell_6t
Xbit_r84_c189 bl_189 br_189 wl_84 vdd gnd cell_6t
Xbit_r85_c189 bl_189 br_189 wl_85 vdd gnd cell_6t
Xbit_r86_c189 bl_189 br_189 wl_86 vdd gnd cell_6t
Xbit_r87_c189 bl_189 br_189 wl_87 vdd gnd cell_6t
Xbit_r88_c189 bl_189 br_189 wl_88 vdd gnd cell_6t
Xbit_r89_c189 bl_189 br_189 wl_89 vdd gnd cell_6t
Xbit_r90_c189 bl_189 br_189 wl_90 vdd gnd cell_6t
Xbit_r91_c189 bl_189 br_189 wl_91 vdd gnd cell_6t
Xbit_r92_c189 bl_189 br_189 wl_92 vdd gnd cell_6t
Xbit_r93_c189 bl_189 br_189 wl_93 vdd gnd cell_6t
Xbit_r94_c189 bl_189 br_189 wl_94 vdd gnd cell_6t
Xbit_r95_c189 bl_189 br_189 wl_95 vdd gnd cell_6t
Xbit_r96_c189 bl_189 br_189 wl_96 vdd gnd cell_6t
Xbit_r97_c189 bl_189 br_189 wl_97 vdd gnd cell_6t
Xbit_r98_c189 bl_189 br_189 wl_98 vdd gnd cell_6t
Xbit_r99_c189 bl_189 br_189 wl_99 vdd gnd cell_6t
Xbit_r100_c189 bl_189 br_189 wl_100 vdd gnd cell_6t
Xbit_r101_c189 bl_189 br_189 wl_101 vdd gnd cell_6t
Xbit_r102_c189 bl_189 br_189 wl_102 vdd gnd cell_6t
Xbit_r103_c189 bl_189 br_189 wl_103 vdd gnd cell_6t
Xbit_r104_c189 bl_189 br_189 wl_104 vdd gnd cell_6t
Xbit_r105_c189 bl_189 br_189 wl_105 vdd gnd cell_6t
Xbit_r106_c189 bl_189 br_189 wl_106 vdd gnd cell_6t
Xbit_r107_c189 bl_189 br_189 wl_107 vdd gnd cell_6t
Xbit_r108_c189 bl_189 br_189 wl_108 vdd gnd cell_6t
Xbit_r109_c189 bl_189 br_189 wl_109 vdd gnd cell_6t
Xbit_r110_c189 bl_189 br_189 wl_110 vdd gnd cell_6t
Xbit_r111_c189 bl_189 br_189 wl_111 vdd gnd cell_6t
Xbit_r112_c189 bl_189 br_189 wl_112 vdd gnd cell_6t
Xbit_r113_c189 bl_189 br_189 wl_113 vdd gnd cell_6t
Xbit_r114_c189 bl_189 br_189 wl_114 vdd gnd cell_6t
Xbit_r115_c189 bl_189 br_189 wl_115 vdd gnd cell_6t
Xbit_r116_c189 bl_189 br_189 wl_116 vdd gnd cell_6t
Xbit_r117_c189 bl_189 br_189 wl_117 vdd gnd cell_6t
Xbit_r118_c189 bl_189 br_189 wl_118 vdd gnd cell_6t
Xbit_r119_c189 bl_189 br_189 wl_119 vdd gnd cell_6t
Xbit_r120_c189 bl_189 br_189 wl_120 vdd gnd cell_6t
Xbit_r121_c189 bl_189 br_189 wl_121 vdd gnd cell_6t
Xbit_r122_c189 bl_189 br_189 wl_122 vdd gnd cell_6t
Xbit_r123_c189 bl_189 br_189 wl_123 vdd gnd cell_6t
Xbit_r124_c189 bl_189 br_189 wl_124 vdd gnd cell_6t
Xbit_r125_c189 bl_189 br_189 wl_125 vdd gnd cell_6t
Xbit_r126_c189 bl_189 br_189 wl_126 vdd gnd cell_6t
Xbit_r127_c189 bl_189 br_189 wl_127 vdd gnd cell_6t
Xbit_r128_c189 bl_189 br_189 wl_128 vdd gnd cell_6t
Xbit_r129_c189 bl_189 br_189 wl_129 vdd gnd cell_6t
Xbit_r130_c189 bl_189 br_189 wl_130 vdd gnd cell_6t
Xbit_r131_c189 bl_189 br_189 wl_131 vdd gnd cell_6t
Xbit_r132_c189 bl_189 br_189 wl_132 vdd gnd cell_6t
Xbit_r133_c189 bl_189 br_189 wl_133 vdd gnd cell_6t
Xbit_r134_c189 bl_189 br_189 wl_134 vdd gnd cell_6t
Xbit_r135_c189 bl_189 br_189 wl_135 vdd gnd cell_6t
Xbit_r136_c189 bl_189 br_189 wl_136 vdd gnd cell_6t
Xbit_r137_c189 bl_189 br_189 wl_137 vdd gnd cell_6t
Xbit_r138_c189 bl_189 br_189 wl_138 vdd gnd cell_6t
Xbit_r139_c189 bl_189 br_189 wl_139 vdd gnd cell_6t
Xbit_r140_c189 bl_189 br_189 wl_140 vdd gnd cell_6t
Xbit_r141_c189 bl_189 br_189 wl_141 vdd gnd cell_6t
Xbit_r142_c189 bl_189 br_189 wl_142 vdd gnd cell_6t
Xbit_r143_c189 bl_189 br_189 wl_143 vdd gnd cell_6t
Xbit_r144_c189 bl_189 br_189 wl_144 vdd gnd cell_6t
Xbit_r145_c189 bl_189 br_189 wl_145 vdd gnd cell_6t
Xbit_r146_c189 bl_189 br_189 wl_146 vdd gnd cell_6t
Xbit_r147_c189 bl_189 br_189 wl_147 vdd gnd cell_6t
Xbit_r148_c189 bl_189 br_189 wl_148 vdd gnd cell_6t
Xbit_r149_c189 bl_189 br_189 wl_149 vdd gnd cell_6t
Xbit_r150_c189 bl_189 br_189 wl_150 vdd gnd cell_6t
Xbit_r151_c189 bl_189 br_189 wl_151 vdd gnd cell_6t
Xbit_r152_c189 bl_189 br_189 wl_152 vdd gnd cell_6t
Xbit_r153_c189 bl_189 br_189 wl_153 vdd gnd cell_6t
Xbit_r154_c189 bl_189 br_189 wl_154 vdd gnd cell_6t
Xbit_r155_c189 bl_189 br_189 wl_155 vdd gnd cell_6t
Xbit_r156_c189 bl_189 br_189 wl_156 vdd gnd cell_6t
Xbit_r157_c189 bl_189 br_189 wl_157 vdd gnd cell_6t
Xbit_r158_c189 bl_189 br_189 wl_158 vdd gnd cell_6t
Xbit_r159_c189 bl_189 br_189 wl_159 vdd gnd cell_6t
Xbit_r160_c189 bl_189 br_189 wl_160 vdd gnd cell_6t
Xbit_r161_c189 bl_189 br_189 wl_161 vdd gnd cell_6t
Xbit_r162_c189 bl_189 br_189 wl_162 vdd gnd cell_6t
Xbit_r163_c189 bl_189 br_189 wl_163 vdd gnd cell_6t
Xbit_r164_c189 bl_189 br_189 wl_164 vdd gnd cell_6t
Xbit_r165_c189 bl_189 br_189 wl_165 vdd gnd cell_6t
Xbit_r166_c189 bl_189 br_189 wl_166 vdd gnd cell_6t
Xbit_r167_c189 bl_189 br_189 wl_167 vdd gnd cell_6t
Xbit_r168_c189 bl_189 br_189 wl_168 vdd gnd cell_6t
Xbit_r169_c189 bl_189 br_189 wl_169 vdd gnd cell_6t
Xbit_r170_c189 bl_189 br_189 wl_170 vdd gnd cell_6t
Xbit_r171_c189 bl_189 br_189 wl_171 vdd gnd cell_6t
Xbit_r172_c189 bl_189 br_189 wl_172 vdd gnd cell_6t
Xbit_r173_c189 bl_189 br_189 wl_173 vdd gnd cell_6t
Xbit_r174_c189 bl_189 br_189 wl_174 vdd gnd cell_6t
Xbit_r175_c189 bl_189 br_189 wl_175 vdd gnd cell_6t
Xbit_r176_c189 bl_189 br_189 wl_176 vdd gnd cell_6t
Xbit_r177_c189 bl_189 br_189 wl_177 vdd gnd cell_6t
Xbit_r178_c189 bl_189 br_189 wl_178 vdd gnd cell_6t
Xbit_r179_c189 bl_189 br_189 wl_179 vdd gnd cell_6t
Xbit_r180_c189 bl_189 br_189 wl_180 vdd gnd cell_6t
Xbit_r181_c189 bl_189 br_189 wl_181 vdd gnd cell_6t
Xbit_r182_c189 bl_189 br_189 wl_182 vdd gnd cell_6t
Xbit_r183_c189 bl_189 br_189 wl_183 vdd gnd cell_6t
Xbit_r184_c189 bl_189 br_189 wl_184 vdd gnd cell_6t
Xbit_r185_c189 bl_189 br_189 wl_185 vdd gnd cell_6t
Xbit_r186_c189 bl_189 br_189 wl_186 vdd gnd cell_6t
Xbit_r187_c189 bl_189 br_189 wl_187 vdd gnd cell_6t
Xbit_r188_c189 bl_189 br_189 wl_188 vdd gnd cell_6t
Xbit_r189_c189 bl_189 br_189 wl_189 vdd gnd cell_6t
Xbit_r190_c189 bl_189 br_189 wl_190 vdd gnd cell_6t
Xbit_r191_c189 bl_189 br_189 wl_191 vdd gnd cell_6t
Xbit_r192_c189 bl_189 br_189 wl_192 vdd gnd cell_6t
Xbit_r193_c189 bl_189 br_189 wl_193 vdd gnd cell_6t
Xbit_r194_c189 bl_189 br_189 wl_194 vdd gnd cell_6t
Xbit_r195_c189 bl_189 br_189 wl_195 vdd gnd cell_6t
Xbit_r196_c189 bl_189 br_189 wl_196 vdd gnd cell_6t
Xbit_r197_c189 bl_189 br_189 wl_197 vdd gnd cell_6t
Xbit_r198_c189 bl_189 br_189 wl_198 vdd gnd cell_6t
Xbit_r199_c189 bl_189 br_189 wl_199 vdd gnd cell_6t
Xbit_r200_c189 bl_189 br_189 wl_200 vdd gnd cell_6t
Xbit_r201_c189 bl_189 br_189 wl_201 vdd gnd cell_6t
Xbit_r202_c189 bl_189 br_189 wl_202 vdd gnd cell_6t
Xbit_r203_c189 bl_189 br_189 wl_203 vdd gnd cell_6t
Xbit_r204_c189 bl_189 br_189 wl_204 vdd gnd cell_6t
Xbit_r205_c189 bl_189 br_189 wl_205 vdd gnd cell_6t
Xbit_r206_c189 bl_189 br_189 wl_206 vdd gnd cell_6t
Xbit_r207_c189 bl_189 br_189 wl_207 vdd gnd cell_6t
Xbit_r208_c189 bl_189 br_189 wl_208 vdd gnd cell_6t
Xbit_r209_c189 bl_189 br_189 wl_209 vdd gnd cell_6t
Xbit_r210_c189 bl_189 br_189 wl_210 vdd gnd cell_6t
Xbit_r211_c189 bl_189 br_189 wl_211 vdd gnd cell_6t
Xbit_r212_c189 bl_189 br_189 wl_212 vdd gnd cell_6t
Xbit_r213_c189 bl_189 br_189 wl_213 vdd gnd cell_6t
Xbit_r214_c189 bl_189 br_189 wl_214 vdd gnd cell_6t
Xbit_r215_c189 bl_189 br_189 wl_215 vdd gnd cell_6t
Xbit_r216_c189 bl_189 br_189 wl_216 vdd gnd cell_6t
Xbit_r217_c189 bl_189 br_189 wl_217 vdd gnd cell_6t
Xbit_r218_c189 bl_189 br_189 wl_218 vdd gnd cell_6t
Xbit_r219_c189 bl_189 br_189 wl_219 vdd gnd cell_6t
Xbit_r220_c189 bl_189 br_189 wl_220 vdd gnd cell_6t
Xbit_r221_c189 bl_189 br_189 wl_221 vdd gnd cell_6t
Xbit_r222_c189 bl_189 br_189 wl_222 vdd gnd cell_6t
Xbit_r223_c189 bl_189 br_189 wl_223 vdd gnd cell_6t
Xbit_r224_c189 bl_189 br_189 wl_224 vdd gnd cell_6t
Xbit_r225_c189 bl_189 br_189 wl_225 vdd gnd cell_6t
Xbit_r226_c189 bl_189 br_189 wl_226 vdd gnd cell_6t
Xbit_r227_c189 bl_189 br_189 wl_227 vdd gnd cell_6t
Xbit_r228_c189 bl_189 br_189 wl_228 vdd gnd cell_6t
Xbit_r229_c189 bl_189 br_189 wl_229 vdd gnd cell_6t
Xbit_r230_c189 bl_189 br_189 wl_230 vdd gnd cell_6t
Xbit_r231_c189 bl_189 br_189 wl_231 vdd gnd cell_6t
Xbit_r232_c189 bl_189 br_189 wl_232 vdd gnd cell_6t
Xbit_r233_c189 bl_189 br_189 wl_233 vdd gnd cell_6t
Xbit_r234_c189 bl_189 br_189 wl_234 vdd gnd cell_6t
Xbit_r235_c189 bl_189 br_189 wl_235 vdd gnd cell_6t
Xbit_r236_c189 bl_189 br_189 wl_236 vdd gnd cell_6t
Xbit_r237_c189 bl_189 br_189 wl_237 vdd gnd cell_6t
Xbit_r238_c189 bl_189 br_189 wl_238 vdd gnd cell_6t
Xbit_r239_c189 bl_189 br_189 wl_239 vdd gnd cell_6t
Xbit_r240_c189 bl_189 br_189 wl_240 vdd gnd cell_6t
Xbit_r241_c189 bl_189 br_189 wl_241 vdd gnd cell_6t
Xbit_r242_c189 bl_189 br_189 wl_242 vdd gnd cell_6t
Xbit_r243_c189 bl_189 br_189 wl_243 vdd gnd cell_6t
Xbit_r244_c189 bl_189 br_189 wl_244 vdd gnd cell_6t
Xbit_r245_c189 bl_189 br_189 wl_245 vdd gnd cell_6t
Xbit_r246_c189 bl_189 br_189 wl_246 vdd gnd cell_6t
Xbit_r247_c189 bl_189 br_189 wl_247 vdd gnd cell_6t
Xbit_r248_c189 bl_189 br_189 wl_248 vdd gnd cell_6t
Xbit_r249_c189 bl_189 br_189 wl_249 vdd gnd cell_6t
Xbit_r250_c189 bl_189 br_189 wl_250 vdd gnd cell_6t
Xbit_r251_c189 bl_189 br_189 wl_251 vdd gnd cell_6t
Xbit_r252_c189 bl_189 br_189 wl_252 vdd gnd cell_6t
Xbit_r253_c189 bl_189 br_189 wl_253 vdd gnd cell_6t
Xbit_r254_c189 bl_189 br_189 wl_254 vdd gnd cell_6t
Xbit_r255_c189 bl_189 br_189 wl_255 vdd gnd cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd cell_6t
Xbit_r1_c190 bl_190 br_190 wl_1 vdd gnd cell_6t
Xbit_r2_c190 bl_190 br_190 wl_2 vdd gnd cell_6t
Xbit_r3_c190 bl_190 br_190 wl_3 vdd gnd cell_6t
Xbit_r4_c190 bl_190 br_190 wl_4 vdd gnd cell_6t
Xbit_r5_c190 bl_190 br_190 wl_5 vdd gnd cell_6t
Xbit_r6_c190 bl_190 br_190 wl_6 vdd gnd cell_6t
Xbit_r7_c190 bl_190 br_190 wl_7 vdd gnd cell_6t
Xbit_r8_c190 bl_190 br_190 wl_8 vdd gnd cell_6t
Xbit_r9_c190 bl_190 br_190 wl_9 vdd gnd cell_6t
Xbit_r10_c190 bl_190 br_190 wl_10 vdd gnd cell_6t
Xbit_r11_c190 bl_190 br_190 wl_11 vdd gnd cell_6t
Xbit_r12_c190 bl_190 br_190 wl_12 vdd gnd cell_6t
Xbit_r13_c190 bl_190 br_190 wl_13 vdd gnd cell_6t
Xbit_r14_c190 bl_190 br_190 wl_14 vdd gnd cell_6t
Xbit_r15_c190 bl_190 br_190 wl_15 vdd gnd cell_6t
Xbit_r16_c190 bl_190 br_190 wl_16 vdd gnd cell_6t
Xbit_r17_c190 bl_190 br_190 wl_17 vdd gnd cell_6t
Xbit_r18_c190 bl_190 br_190 wl_18 vdd gnd cell_6t
Xbit_r19_c190 bl_190 br_190 wl_19 vdd gnd cell_6t
Xbit_r20_c190 bl_190 br_190 wl_20 vdd gnd cell_6t
Xbit_r21_c190 bl_190 br_190 wl_21 vdd gnd cell_6t
Xbit_r22_c190 bl_190 br_190 wl_22 vdd gnd cell_6t
Xbit_r23_c190 bl_190 br_190 wl_23 vdd gnd cell_6t
Xbit_r24_c190 bl_190 br_190 wl_24 vdd gnd cell_6t
Xbit_r25_c190 bl_190 br_190 wl_25 vdd gnd cell_6t
Xbit_r26_c190 bl_190 br_190 wl_26 vdd gnd cell_6t
Xbit_r27_c190 bl_190 br_190 wl_27 vdd gnd cell_6t
Xbit_r28_c190 bl_190 br_190 wl_28 vdd gnd cell_6t
Xbit_r29_c190 bl_190 br_190 wl_29 vdd gnd cell_6t
Xbit_r30_c190 bl_190 br_190 wl_30 vdd gnd cell_6t
Xbit_r31_c190 bl_190 br_190 wl_31 vdd gnd cell_6t
Xbit_r32_c190 bl_190 br_190 wl_32 vdd gnd cell_6t
Xbit_r33_c190 bl_190 br_190 wl_33 vdd gnd cell_6t
Xbit_r34_c190 bl_190 br_190 wl_34 vdd gnd cell_6t
Xbit_r35_c190 bl_190 br_190 wl_35 vdd gnd cell_6t
Xbit_r36_c190 bl_190 br_190 wl_36 vdd gnd cell_6t
Xbit_r37_c190 bl_190 br_190 wl_37 vdd gnd cell_6t
Xbit_r38_c190 bl_190 br_190 wl_38 vdd gnd cell_6t
Xbit_r39_c190 bl_190 br_190 wl_39 vdd gnd cell_6t
Xbit_r40_c190 bl_190 br_190 wl_40 vdd gnd cell_6t
Xbit_r41_c190 bl_190 br_190 wl_41 vdd gnd cell_6t
Xbit_r42_c190 bl_190 br_190 wl_42 vdd gnd cell_6t
Xbit_r43_c190 bl_190 br_190 wl_43 vdd gnd cell_6t
Xbit_r44_c190 bl_190 br_190 wl_44 vdd gnd cell_6t
Xbit_r45_c190 bl_190 br_190 wl_45 vdd gnd cell_6t
Xbit_r46_c190 bl_190 br_190 wl_46 vdd gnd cell_6t
Xbit_r47_c190 bl_190 br_190 wl_47 vdd gnd cell_6t
Xbit_r48_c190 bl_190 br_190 wl_48 vdd gnd cell_6t
Xbit_r49_c190 bl_190 br_190 wl_49 vdd gnd cell_6t
Xbit_r50_c190 bl_190 br_190 wl_50 vdd gnd cell_6t
Xbit_r51_c190 bl_190 br_190 wl_51 vdd gnd cell_6t
Xbit_r52_c190 bl_190 br_190 wl_52 vdd gnd cell_6t
Xbit_r53_c190 bl_190 br_190 wl_53 vdd gnd cell_6t
Xbit_r54_c190 bl_190 br_190 wl_54 vdd gnd cell_6t
Xbit_r55_c190 bl_190 br_190 wl_55 vdd gnd cell_6t
Xbit_r56_c190 bl_190 br_190 wl_56 vdd gnd cell_6t
Xbit_r57_c190 bl_190 br_190 wl_57 vdd gnd cell_6t
Xbit_r58_c190 bl_190 br_190 wl_58 vdd gnd cell_6t
Xbit_r59_c190 bl_190 br_190 wl_59 vdd gnd cell_6t
Xbit_r60_c190 bl_190 br_190 wl_60 vdd gnd cell_6t
Xbit_r61_c190 bl_190 br_190 wl_61 vdd gnd cell_6t
Xbit_r62_c190 bl_190 br_190 wl_62 vdd gnd cell_6t
Xbit_r63_c190 bl_190 br_190 wl_63 vdd gnd cell_6t
Xbit_r64_c190 bl_190 br_190 wl_64 vdd gnd cell_6t
Xbit_r65_c190 bl_190 br_190 wl_65 vdd gnd cell_6t
Xbit_r66_c190 bl_190 br_190 wl_66 vdd gnd cell_6t
Xbit_r67_c190 bl_190 br_190 wl_67 vdd gnd cell_6t
Xbit_r68_c190 bl_190 br_190 wl_68 vdd gnd cell_6t
Xbit_r69_c190 bl_190 br_190 wl_69 vdd gnd cell_6t
Xbit_r70_c190 bl_190 br_190 wl_70 vdd gnd cell_6t
Xbit_r71_c190 bl_190 br_190 wl_71 vdd gnd cell_6t
Xbit_r72_c190 bl_190 br_190 wl_72 vdd gnd cell_6t
Xbit_r73_c190 bl_190 br_190 wl_73 vdd gnd cell_6t
Xbit_r74_c190 bl_190 br_190 wl_74 vdd gnd cell_6t
Xbit_r75_c190 bl_190 br_190 wl_75 vdd gnd cell_6t
Xbit_r76_c190 bl_190 br_190 wl_76 vdd gnd cell_6t
Xbit_r77_c190 bl_190 br_190 wl_77 vdd gnd cell_6t
Xbit_r78_c190 bl_190 br_190 wl_78 vdd gnd cell_6t
Xbit_r79_c190 bl_190 br_190 wl_79 vdd gnd cell_6t
Xbit_r80_c190 bl_190 br_190 wl_80 vdd gnd cell_6t
Xbit_r81_c190 bl_190 br_190 wl_81 vdd gnd cell_6t
Xbit_r82_c190 bl_190 br_190 wl_82 vdd gnd cell_6t
Xbit_r83_c190 bl_190 br_190 wl_83 vdd gnd cell_6t
Xbit_r84_c190 bl_190 br_190 wl_84 vdd gnd cell_6t
Xbit_r85_c190 bl_190 br_190 wl_85 vdd gnd cell_6t
Xbit_r86_c190 bl_190 br_190 wl_86 vdd gnd cell_6t
Xbit_r87_c190 bl_190 br_190 wl_87 vdd gnd cell_6t
Xbit_r88_c190 bl_190 br_190 wl_88 vdd gnd cell_6t
Xbit_r89_c190 bl_190 br_190 wl_89 vdd gnd cell_6t
Xbit_r90_c190 bl_190 br_190 wl_90 vdd gnd cell_6t
Xbit_r91_c190 bl_190 br_190 wl_91 vdd gnd cell_6t
Xbit_r92_c190 bl_190 br_190 wl_92 vdd gnd cell_6t
Xbit_r93_c190 bl_190 br_190 wl_93 vdd gnd cell_6t
Xbit_r94_c190 bl_190 br_190 wl_94 vdd gnd cell_6t
Xbit_r95_c190 bl_190 br_190 wl_95 vdd gnd cell_6t
Xbit_r96_c190 bl_190 br_190 wl_96 vdd gnd cell_6t
Xbit_r97_c190 bl_190 br_190 wl_97 vdd gnd cell_6t
Xbit_r98_c190 bl_190 br_190 wl_98 vdd gnd cell_6t
Xbit_r99_c190 bl_190 br_190 wl_99 vdd gnd cell_6t
Xbit_r100_c190 bl_190 br_190 wl_100 vdd gnd cell_6t
Xbit_r101_c190 bl_190 br_190 wl_101 vdd gnd cell_6t
Xbit_r102_c190 bl_190 br_190 wl_102 vdd gnd cell_6t
Xbit_r103_c190 bl_190 br_190 wl_103 vdd gnd cell_6t
Xbit_r104_c190 bl_190 br_190 wl_104 vdd gnd cell_6t
Xbit_r105_c190 bl_190 br_190 wl_105 vdd gnd cell_6t
Xbit_r106_c190 bl_190 br_190 wl_106 vdd gnd cell_6t
Xbit_r107_c190 bl_190 br_190 wl_107 vdd gnd cell_6t
Xbit_r108_c190 bl_190 br_190 wl_108 vdd gnd cell_6t
Xbit_r109_c190 bl_190 br_190 wl_109 vdd gnd cell_6t
Xbit_r110_c190 bl_190 br_190 wl_110 vdd gnd cell_6t
Xbit_r111_c190 bl_190 br_190 wl_111 vdd gnd cell_6t
Xbit_r112_c190 bl_190 br_190 wl_112 vdd gnd cell_6t
Xbit_r113_c190 bl_190 br_190 wl_113 vdd gnd cell_6t
Xbit_r114_c190 bl_190 br_190 wl_114 vdd gnd cell_6t
Xbit_r115_c190 bl_190 br_190 wl_115 vdd gnd cell_6t
Xbit_r116_c190 bl_190 br_190 wl_116 vdd gnd cell_6t
Xbit_r117_c190 bl_190 br_190 wl_117 vdd gnd cell_6t
Xbit_r118_c190 bl_190 br_190 wl_118 vdd gnd cell_6t
Xbit_r119_c190 bl_190 br_190 wl_119 vdd gnd cell_6t
Xbit_r120_c190 bl_190 br_190 wl_120 vdd gnd cell_6t
Xbit_r121_c190 bl_190 br_190 wl_121 vdd gnd cell_6t
Xbit_r122_c190 bl_190 br_190 wl_122 vdd gnd cell_6t
Xbit_r123_c190 bl_190 br_190 wl_123 vdd gnd cell_6t
Xbit_r124_c190 bl_190 br_190 wl_124 vdd gnd cell_6t
Xbit_r125_c190 bl_190 br_190 wl_125 vdd gnd cell_6t
Xbit_r126_c190 bl_190 br_190 wl_126 vdd gnd cell_6t
Xbit_r127_c190 bl_190 br_190 wl_127 vdd gnd cell_6t
Xbit_r128_c190 bl_190 br_190 wl_128 vdd gnd cell_6t
Xbit_r129_c190 bl_190 br_190 wl_129 vdd gnd cell_6t
Xbit_r130_c190 bl_190 br_190 wl_130 vdd gnd cell_6t
Xbit_r131_c190 bl_190 br_190 wl_131 vdd gnd cell_6t
Xbit_r132_c190 bl_190 br_190 wl_132 vdd gnd cell_6t
Xbit_r133_c190 bl_190 br_190 wl_133 vdd gnd cell_6t
Xbit_r134_c190 bl_190 br_190 wl_134 vdd gnd cell_6t
Xbit_r135_c190 bl_190 br_190 wl_135 vdd gnd cell_6t
Xbit_r136_c190 bl_190 br_190 wl_136 vdd gnd cell_6t
Xbit_r137_c190 bl_190 br_190 wl_137 vdd gnd cell_6t
Xbit_r138_c190 bl_190 br_190 wl_138 vdd gnd cell_6t
Xbit_r139_c190 bl_190 br_190 wl_139 vdd gnd cell_6t
Xbit_r140_c190 bl_190 br_190 wl_140 vdd gnd cell_6t
Xbit_r141_c190 bl_190 br_190 wl_141 vdd gnd cell_6t
Xbit_r142_c190 bl_190 br_190 wl_142 vdd gnd cell_6t
Xbit_r143_c190 bl_190 br_190 wl_143 vdd gnd cell_6t
Xbit_r144_c190 bl_190 br_190 wl_144 vdd gnd cell_6t
Xbit_r145_c190 bl_190 br_190 wl_145 vdd gnd cell_6t
Xbit_r146_c190 bl_190 br_190 wl_146 vdd gnd cell_6t
Xbit_r147_c190 bl_190 br_190 wl_147 vdd gnd cell_6t
Xbit_r148_c190 bl_190 br_190 wl_148 vdd gnd cell_6t
Xbit_r149_c190 bl_190 br_190 wl_149 vdd gnd cell_6t
Xbit_r150_c190 bl_190 br_190 wl_150 vdd gnd cell_6t
Xbit_r151_c190 bl_190 br_190 wl_151 vdd gnd cell_6t
Xbit_r152_c190 bl_190 br_190 wl_152 vdd gnd cell_6t
Xbit_r153_c190 bl_190 br_190 wl_153 vdd gnd cell_6t
Xbit_r154_c190 bl_190 br_190 wl_154 vdd gnd cell_6t
Xbit_r155_c190 bl_190 br_190 wl_155 vdd gnd cell_6t
Xbit_r156_c190 bl_190 br_190 wl_156 vdd gnd cell_6t
Xbit_r157_c190 bl_190 br_190 wl_157 vdd gnd cell_6t
Xbit_r158_c190 bl_190 br_190 wl_158 vdd gnd cell_6t
Xbit_r159_c190 bl_190 br_190 wl_159 vdd gnd cell_6t
Xbit_r160_c190 bl_190 br_190 wl_160 vdd gnd cell_6t
Xbit_r161_c190 bl_190 br_190 wl_161 vdd gnd cell_6t
Xbit_r162_c190 bl_190 br_190 wl_162 vdd gnd cell_6t
Xbit_r163_c190 bl_190 br_190 wl_163 vdd gnd cell_6t
Xbit_r164_c190 bl_190 br_190 wl_164 vdd gnd cell_6t
Xbit_r165_c190 bl_190 br_190 wl_165 vdd gnd cell_6t
Xbit_r166_c190 bl_190 br_190 wl_166 vdd gnd cell_6t
Xbit_r167_c190 bl_190 br_190 wl_167 vdd gnd cell_6t
Xbit_r168_c190 bl_190 br_190 wl_168 vdd gnd cell_6t
Xbit_r169_c190 bl_190 br_190 wl_169 vdd gnd cell_6t
Xbit_r170_c190 bl_190 br_190 wl_170 vdd gnd cell_6t
Xbit_r171_c190 bl_190 br_190 wl_171 vdd gnd cell_6t
Xbit_r172_c190 bl_190 br_190 wl_172 vdd gnd cell_6t
Xbit_r173_c190 bl_190 br_190 wl_173 vdd gnd cell_6t
Xbit_r174_c190 bl_190 br_190 wl_174 vdd gnd cell_6t
Xbit_r175_c190 bl_190 br_190 wl_175 vdd gnd cell_6t
Xbit_r176_c190 bl_190 br_190 wl_176 vdd gnd cell_6t
Xbit_r177_c190 bl_190 br_190 wl_177 vdd gnd cell_6t
Xbit_r178_c190 bl_190 br_190 wl_178 vdd gnd cell_6t
Xbit_r179_c190 bl_190 br_190 wl_179 vdd gnd cell_6t
Xbit_r180_c190 bl_190 br_190 wl_180 vdd gnd cell_6t
Xbit_r181_c190 bl_190 br_190 wl_181 vdd gnd cell_6t
Xbit_r182_c190 bl_190 br_190 wl_182 vdd gnd cell_6t
Xbit_r183_c190 bl_190 br_190 wl_183 vdd gnd cell_6t
Xbit_r184_c190 bl_190 br_190 wl_184 vdd gnd cell_6t
Xbit_r185_c190 bl_190 br_190 wl_185 vdd gnd cell_6t
Xbit_r186_c190 bl_190 br_190 wl_186 vdd gnd cell_6t
Xbit_r187_c190 bl_190 br_190 wl_187 vdd gnd cell_6t
Xbit_r188_c190 bl_190 br_190 wl_188 vdd gnd cell_6t
Xbit_r189_c190 bl_190 br_190 wl_189 vdd gnd cell_6t
Xbit_r190_c190 bl_190 br_190 wl_190 vdd gnd cell_6t
Xbit_r191_c190 bl_190 br_190 wl_191 vdd gnd cell_6t
Xbit_r192_c190 bl_190 br_190 wl_192 vdd gnd cell_6t
Xbit_r193_c190 bl_190 br_190 wl_193 vdd gnd cell_6t
Xbit_r194_c190 bl_190 br_190 wl_194 vdd gnd cell_6t
Xbit_r195_c190 bl_190 br_190 wl_195 vdd gnd cell_6t
Xbit_r196_c190 bl_190 br_190 wl_196 vdd gnd cell_6t
Xbit_r197_c190 bl_190 br_190 wl_197 vdd gnd cell_6t
Xbit_r198_c190 bl_190 br_190 wl_198 vdd gnd cell_6t
Xbit_r199_c190 bl_190 br_190 wl_199 vdd gnd cell_6t
Xbit_r200_c190 bl_190 br_190 wl_200 vdd gnd cell_6t
Xbit_r201_c190 bl_190 br_190 wl_201 vdd gnd cell_6t
Xbit_r202_c190 bl_190 br_190 wl_202 vdd gnd cell_6t
Xbit_r203_c190 bl_190 br_190 wl_203 vdd gnd cell_6t
Xbit_r204_c190 bl_190 br_190 wl_204 vdd gnd cell_6t
Xbit_r205_c190 bl_190 br_190 wl_205 vdd gnd cell_6t
Xbit_r206_c190 bl_190 br_190 wl_206 vdd gnd cell_6t
Xbit_r207_c190 bl_190 br_190 wl_207 vdd gnd cell_6t
Xbit_r208_c190 bl_190 br_190 wl_208 vdd gnd cell_6t
Xbit_r209_c190 bl_190 br_190 wl_209 vdd gnd cell_6t
Xbit_r210_c190 bl_190 br_190 wl_210 vdd gnd cell_6t
Xbit_r211_c190 bl_190 br_190 wl_211 vdd gnd cell_6t
Xbit_r212_c190 bl_190 br_190 wl_212 vdd gnd cell_6t
Xbit_r213_c190 bl_190 br_190 wl_213 vdd gnd cell_6t
Xbit_r214_c190 bl_190 br_190 wl_214 vdd gnd cell_6t
Xbit_r215_c190 bl_190 br_190 wl_215 vdd gnd cell_6t
Xbit_r216_c190 bl_190 br_190 wl_216 vdd gnd cell_6t
Xbit_r217_c190 bl_190 br_190 wl_217 vdd gnd cell_6t
Xbit_r218_c190 bl_190 br_190 wl_218 vdd gnd cell_6t
Xbit_r219_c190 bl_190 br_190 wl_219 vdd gnd cell_6t
Xbit_r220_c190 bl_190 br_190 wl_220 vdd gnd cell_6t
Xbit_r221_c190 bl_190 br_190 wl_221 vdd gnd cell_6t
Xbit_r222_c190 bl_190 br_190 wl_222 vdd gnd cell_6t
Xbit_r223_c190 bl_190 br_190 wl_223 vdd gnd cell_6t
Xbit_r224_c190 bl_190 br_190 wl_224 vdd gnd cell_6t
Xbit_r225_c190 bl_190 br_190 wl_225 vdd gnd cell_6t
Xbit_r226_c190 bl_190 br_190 wl_226 vdd gnd cell_6t
Xbit_r227_c190 bl_190 br_190 wl_227 vdd gnd cell_6t
Xbit_r228_c190 bl_190 br_190 wl_228 vdd gnd cell_6t
Xbit_r229_c190 bl_190 br_190 wl_229 vdd gnd cell_6t
Xbit_r230_c190 bl_190 br_190 wl_230 vdd gnd cell_6t
Xbit_r231_c190 bl_190 br_190 wl_231 vdd gnd cell_6t
Xbit_r232_c190 bl_190 br_190 wl_232 vdd gnd cell_6t
Xbit_r233_c190 bl_190 br_190 wl_233 vdd gnd cell_6t
Xbit_r234_c190 bl_190 br_190 wl_234 vdd gnd cell_6t
Xbit_r235_c190 bl_190 br_190 wl_235 vdd gnd cell_6t
Xbit_r236_c190 bl_190 br_190 wl_236 vdd gnd cell_6t
Xbit_r237_c190 bl_190 br_190 wl_237 vdd gnd cell_6t
Xbit_r238_c190 bl_190 br_190 wl_238 vdd gnd cell_6t
Xbit_r239_c190 bl_190 br_190 wl_239 vdd gnd cell_6t
Xbit_r240_c190 bl_190 br_190 wl_240 vdd gnd cell_6t
Xbit_r241_c190 bl_190 br_190 wl_241 vdd gnd cell_6t
Xbit_r242_c190 bl_190 br_190 wl_242 vdd gnd cell_6t
Xbit_r243_c190 bl_190 br_190 wl_243 vdd gnd cell_6t
Xbit_r244_c190 bl_190 br_190 wl_244 vdd gnd cell_6t
Xbit_r245_c190 bl_190 br_190 wl_245 vdd gnd cell_6t
Xbit_r246_c190 bl_190 br_190 wl_246 vdd gnd cell_6t
Xbit_r247_c190 bl_190 br_190 wl_247 vdd gnd cell_6t
Xbit_r248_c190 bl_190 br_190 wl_248 vdd gnd cell_6t
Xbit_r249_c190 bl_190 br_190 wl_249 vdd gnd cell_6t
Xbit_r250_c190 bl_190 br_190 wl_250 vdd gnd cell_6t
Xbit_r251_c190 bl_190 br_190 wl_251 vdd gnd cell_6t
Xbit_r252_c190 bl_190 br_190 wl_252 vdd gnd cell_6t
Xbit_r253_c190 bl_190 br_190 wl_253 vdd gnd cell_6t
Xbit_r254_c190 bl_190 br_190 wl_254 vdd gnd cell_6t
Xbit_r255_c190 bl_190 br_190 wl_255 vdd gnd cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd cell_6t
Xbit_r1_c191 bl_191 br_191 wl_1 vdd gnd cell_6t
Xbit_r2_c191 bl_191 br_191 wl_2 vdd gnd cell_6t
Xbit_r3_c191 bl_191 br_191 wl_3 vdd gnd cell_6t
Xbit_r4_c191 bl_191 br_191 wl_4 vdd gnd cell_6t
Xbit_r5_c191 bl_191 br_191 wl_5 vdd gnd cell_6t
Xbit_r6_c191 bl_191 br_191 wl_6 vdd gnd cell_6t
Xbit_r7_c191 bl_191 br_191 wl_7 vdd gnd cell_6t
Xbit_r8_c191 bl_191 br_191 wl_8 vdd gnd cell_6t
Xbit_r9_c191 bl_191 br_191 wl_9 vdd gnd cell_6t
Xbit_r10_c191 bl_191 br_191 wl_10 vdd gnd cell_6t
Xbit_r11_c191 bl_191 br_191 wl_11 vdd gnd cell_6t
Xbit_r12_c191 bl_191 br_191 wl_12 vdd gnd cell_6t
Xbit_r13_c191 bl_191 br_191 wl_13 vdd gnd cell_6t
Xbit_r14_c191 bl_191 br_191 wl_14 vdd gnd cell_6t
Xbit_r15_c191 bl_191 br_191 wl_15 vdd gnd cell_6t
Xbit_r16_c191 bl_191 br_191 wl_16 vdd gnd cell_6t
Xbit_r17_c191 bl_191 br_191 wl_17 vdd gnd cell_6t
Xbit_r18_c191 bl_191 br_191 wl_18 vdd gnd cell_6t
Xbit_r19_c191 bl_191 br_191 wl_19 vdd gnd cell_6t
Xbit_r20_c191 bl_191 br_191 wl_20 vdd gnd cell_6t
Xbit_r21_c191 bl_191 br_191 wl_21 vdd gnd cell_6t
Xbit_r22_c191 bl_191 br_191 wl_22 vdd gnd cell_6t
Xbit_r23_c191 bl_191 br_191 wl_23 vdd gnd cell_6t
Xbit_r24_c191 bl_191 br_191 wl_24 vdd gnd cell_6t
Xbit_r25_c191 bl_191 br_191 wl_25 vdd gnd cell_6t
Xbit_r26_c191 bl_191 br_191 wl_26 vdd gnd cell_6t
Xbit_r27_c191 bl_191 br_191 wl_27 vdd gnd cell_6t
Xbit_r28_c191 bl_191 br_191 wl_28 vdd gnd cell_6t
Xbit_r29_c191 bl_191 br_191 wl_29 vdd gnd cell_6t
Xbit_r30_c191 bl_191 br_191 wl_30 vdd gnd cell_6t
Xbit_r31_c191 bl_191 br_191 wl_31 vdd gnd cell_6t
Xbit_r32_c191 bl_191 br_191 wl_32 vdd gnd cell_6t
Xbit_r33_c191 bl_191 br_191 wl_33 vdd gnd cell_6t
Xbit_r34_c191 bl_191 br_191 wl_34 vdd gnd cell_6t
Xbit_r35_c191 bl_191 br_191 wl_35 vdd gnd cell_6t
Xbit_r36_c191 bl_191 br_191 wl_36 vdd gnd cell_6t
Xbit_r37_c191 bl_191 br_191 wl_37 vdd gnd cell_6t
Xbit_r38_c191 bl_191 br_191 wl_38 vdd gnd cell_6t
Xbit_r39_c191 bl_191 br_191 wl_39 vdd gnd cell_6t
Xbit_r40_c191 bl_191 br_191 wl_40 vdd gnd cell_6t
Xbit_r41_c191 bl_191 br_191 wl_41 vdd gnd cell_6t
Xbit_r42_c191 bl_191 br_191 wl_42 vdd gnd cell_6t
Xbit_r43_c191 bl_191 br_191 wl_43 vdd gnd cell_6t
Xbit_r44_c191 bl_191 br_191 wl_44 vdd gnd cell_6t
Xbit_r45_c191 bl_191 br_191 wl_45 vdd gnd cell_6t
Xbit_r46_c191 bl_191 br_191 wl_46 vdd gnd cell_6t
Xbit_r47_c191 bl_191 br_191 wl_47 vdd gnd cell_6t
Xbit_r48_c191 bl_191 br_191 wl_48 vdd gnd cell_6t
Xbit_r49_c191 bl_191 br_191 wl_49 vdd gnd cell_6t
Xbit_r50_c191 bl_191 br_191 wl_50 vdd gnd cell_6t
Xbit_r51_c191 bl_191 br_191 wl_51 vdd gnd cell_6t
Xbit_r52_c191 bl_191 br_191 wl_52 vdd gnd cell_6t
Xbit_r53_c191 bl_191 br_191 wl_53 vdd gnd cell_6t
Xbit_r54_c191 bl_191 br_191 wl_54 vdd gnd cell_6t
Xbit_r55_c191 bl_191 br_191 wl_55 vdd gnd cell_6t
Xbit_r56_c191 bl_191 br_191 wl_56 vdd gnd cell_6t
Xbit_r57_c191 bl_191 br_191 wl_57 vdd gnd cell_6t
Xbit_r58_c191 bl_191 br_191 wl_58 vdd gnd cell_6t
Xbit_r59_c191 bl_191 br_191 wl_59 vdd gnd cell_6t
Xbit_r60_c191 bl_191 br_191 wl_60 vdd gnd cell_6t
Xbit_r61_c191 bl_191 br_191 wl_61 vdd gnd cell_6t
Xbit_r62_c191 bl_191 br_191 wl_62 vdd gnd cell_6t
Xbit_r63_c191 bl_191 br_191 wl_63 vdd gnd cell_6t
Xbit_r64_c191 bl_191 br_191 wl_64 vdd gnd cell_6t
Xbit_r65_c191 bl_191 br_191 wl_65 vdd gnd cell_6t
Xbit_r66_c191 bl_191 br_191 wl_66 vdd gnd cell_6t
Xbit_r67_c191 bl_191 br_191 wl_67 vdd gnd cell_6t
Xbit_r68_c191 bl_191 br_191 wl_68 vdd gnd cell_6t
Xbit_r69_c191 bl_191 br_191 wl_69 vdd gnd cell_6t
Xbit_r70_c191 bl_191 br_191 wl_70 vdd gnd cell_6t
Xbit_r71_c191 bl_191 br_191 wl_71 vdd gnd cell_6t
Xbit_r72_c191 bl_191 br_191 wl_72 vdd gnd cell_6t
Xbit_r73_c191 bl_191 br_191 wl_73 vdd gnd cell_6t
Xbit_r74_c191 bl_191 br_191 wl_74 vdd gnd cell_6t
Xbit_r75_c191 bl_191 br_191 wl_75 vdd gnd cell_6t
Xbit_r76_c191 bl_191 br_191 wl_76 vdd gnd cell_6t
Xbit_r77_c191 bl_191 br_191 wl_77 vdd gnd cell_6t
Xbit_r78_c191 bl_191 br_191 wl_78 vdd gnd cell_6t
Xbit_r79_c191 bl_191 br_191 wl_79 vdd gnd cell_6t
Xbit_r80_c191 bl_191 br_191 wl_80 vdd gnd cell_6t
Xbit_r81_c191 bl_191 br_191 wl_81 vdd gnd cell_6t
Xbit_r82_c191 bl_191 br_191 wl_82 vdd gnd cell_6t
Xbit_r83_c191 bl_191 br_191 wl_83 vdd gnd cell_6t
Xbit_r84_c191 bl_191 br_191 wl_84 vdd gnd cell_6t
Xbit_r85_c191 bl_191 br_191 wl_85 vdd gnd cell_6t
Xbit_r86_c191 bl_191 br_191 wl_86 vdd gnd cell_6t
Xbit_r87_c191 bl_191 br_191 wl_87 vdd gnd cell_6t
Xbit_r88_c191 bl_191 br_191 wl_88 vdd gnd cell_6t
Xbit_r89_c191 bl_191 br_191 wl_89 vdd gnd cell_6t
Xbit_r90_c191 bl_191 br_191 wl_90 vdd gnd cell_6t
Xbit_r91_c191 bl_191 br_191 wl_91 vdd gnd cell_6t
Xbit_r92_c191 bl_191 br_191 wl_92 vdd gnd cell_6t
Xbit_r93_c191 bl_191 br_191 wl_93 vdd gnd cell_6t
Xbit_r94_c191 bl_191 br_191 wl_94 vdd gnd cell_6t
Xbit_r95_c191 bl_191 br_191 wl_95 vdd gnd cell_6t
Xbit_r96_c191 bl_191 br_191 wl_96 vdd gnd cell_6t
Xbit_r97_c191 bl_191 br_191 wl_97 vdd gnd cell_6t
Xbit_r98_c191 bl_191 br_191 wl_98 vdd gnd cell_6t
Xbit_r99_c191 bl_191 br_191 wl_99 vdd gnd cell_6t
Xbit_r100_c191 bl_191 br_191 wl_100 vdd gnd cell_6t
Xbit_r101_c191 bl_191 br_191 wl_101 vdd gnd cell_6t
Xbit_r102_c191 bl_191 br_191 wl_102 vdd gnd cell_6t
Xbit_r103_c191 bl_191 br_191 wl_103 vdd gnd cell_6t
Xbit_r104_c191 bl_191 br_191 wl_104 vdd gnd cell_6t
Xbit_r105_c191 bl_191 br_191 wl_105 vdd gnd cell_6t
Xbit_r106_c191 bl_191 br_191 wl_106 vdd gnd cell_6t
Xbit_r107_c191 bl_191 br_191 wl_107 vdd gnd cell_6t
Xbit_r108_c191 bl_191 br_191 wl_108 vdd gnd cell_6t
Xbit_r109_c191 bl_191 br_191 wl_109 vdd gnd cell_6t
Xbit_r110_c191 bl_191 br_191 wl_110 vdd gnd cell_6t
Xbit_r111_c191 bl_191 br_191 wl_111 vdd gnd cell_6t
Xbit_r112_c191 bl_191 br_191 wl_112 vdd gnd cell_6t
Xbit_r113_c191 bl_191 br_191 wl_113 vdd gnd cell_6t
Xbit_r114_c191 bl_191 br_191 wl_114 vdd gnd cell_6t
Xbit_r115_c191 bl_191 br_191 wl_115 vdd gnd cell_6t
Xbit_r116_c191 bl_191 br_191 wl_116 vdd gnd cell_6t
Xbit_r117_c191 bl_191 br_191 wl_117 vdd gnd cell_6t
Xbit_r118_c191 bl_191 br_191 wl_118 vdd gnd cell_6t
Xbit_r119_c191 bl_191 br_191 wl_119 vdd gnd cell_6t
Xbit_r120_c191 bl_191 br_191 wl_120 vdd gnd cell_6t
Xbit_r121_c191 bl_191 br_191 wl_121 vdd gnd cell_6t
Xbit_r122_c191 bl_191 br_191 wl_122 vdd gnd cell_6t
Xbit_r123_c191 bl_191 br_191 wl_123 vdd gnd cell_6t
Xbit_r124_c191 bl_191 br_191 wl_124 vdd gnd cell_6t
Xbit_r125_c191 bl_191 br_191 wl_125 vdd gnd cell_6t
Xbit_r126_c191 bl_191 br_191 wl_126 vdd gnd cell_6t
Xbit_r127_c191 bl_191 br_191 wl_127 vdd gnd cell_6t
Xbit_r128_c191 bl_191 br_191 wl_128 vdd gnd cell_6t
Xbit_r129_c191 bl_191 br_191 wl_129 vdd gnd cell_6t
Xbit_r130_c191 bl_191 br_191 wl_130 vdd gnd cell_6t
Xbit_r131_c191 bl_191 br_191 wl_131 vdd gnd cell_6t
Xbit_r132_c191 bl_191 br_191 wl_132 vdd gnd cell_6t
Xbit_r133_c191 bl_191 br_191 wl_133 vdd gnd cell_6t
Xbit_r134_c191 bl_191 br_191 wl_134 vdd gnd cell_6t
Xbit_r135_c191 bl_191 br_191 wl_135 vdd gnd cell_6t
Xbit_r136_c191 bl_191 br_191 wl_136 vdd gnd cell_6t
Xbit_r137_c191 bl_191 br_191 wl_137 vdd gnd cell_6t
Xbit_r138_c191 bl_191 br_191 wl_138 vdd gnd cell_6t
Xbit_r139_c191 bl_191 br_191 wl_139 vdd gnd cell_6t
Xbit_r140_c191 bl_191 br_191 wl_140 vdd gnd cell_6t
Xbit_r141_c191 bl_191 br_191 wl_141 vdd gnd cell_6t
Xbit_r142_c191 bl_191 br_191 wl_142 vdd gnd cell_6t
Xbit_r143_c191 bl_191 br_191 wl_143 vdd gnd cell_6t
Xbit_r144_c191 bl_191 br_191 wl_144 vdd gnd cell_6t
Xbit_r145_c191 bl_191 br_191 wl_145 vdd gnd cell_6t
Xbit_r146_c191 bl_191 br_191 wl_146 vdd gnd cell_6t
Xbit_r147_c191 bl_191 br_191 wl_147 vdd gnd cell_6t
Xbit_r148_c191 bl_191 br_191 wl_148 vdd gnd cell_6t
Xbit_r149_c191 bl_191 br_191 wl_149 vdd gnd cell_6t
Xbit_r150_c191 bl_191 br_191 wl_150 vdd gnd cell_6t
Xbit_r151_c191 bl_191 br_191 wl_151 vdd gnd cell_6t
Xbit_r152_c191 bl_191 br_191 wl_152 vdd gnd cell_6t
Xbit_r153_c191 bl_191 br_191 wl_153 vdd gnd cell_6t
Xbit_r154_c191 bl_191 br_191 wl_154 vdd gnd cell_6t
Xbit_r155_c191 bl_191 br_191 wl_155 vdd gnd cell_6t
Xbit_r156_c191 bl_191 br_191 wl_156 vdd gnd cell_6t
Xbit_r157_c191 bl_191 br_191 wl_157 vdd gnd cell_6t
Xbit_r158_c191 bl_191 br_191 wl_158 vdd gnd cell_6t
Xbit_r159_c191 bl_191 br_191 wl_159 vdd gnd cell_6t
Xbit_r160_c191 bl_191 br_191 wl_160 vdd gnd cell_6t
Xbit_r161_c191 bl_191 br_191 wl_161 vdd gnd cell_6t
Xbit_r162_c191 bl_191 br_191 wl_162 vdd gnd cell_6t
Xbit_r163_c191 bl_191 br_191 wl_163 vdd gnd cell_6t
Xbit_r164_c191 bl_191 br_191 wl_164 vdd gnd cell_6t
Xbit_r165_c191 bl_191 br_191 wl_165 vdd gnd cell_6t
Xbit_r166_c191 bl_191 br_191 wl_166 vdd gnd cell_6t
Xbit_r167_c191 bl_191 br_191 wl_167 vdd gnd cell_6t
Xbit_r168_c191 bl_191 br_191 wl_168 vdd gnd cell_6t
Xbit_r169_c191 bl_191 br_191 wl_169 vdd gnd cell_6t
Xbit_r170_c191 bl_191 br_191 wl_170 vdd gnd cell_6t
Xbit_r171_c191 bl_191 br_191 wl_171 vdd gnd cell_6t
Xbit_r172_c191 bl_191 br_191 wl_172 vdd gnd cell_6t
Xbit_r173_c191 bl_191 br_191 wl_173 vdd gnd cell_6t
Xbit_r174_c191 bl_191 br_191 wl_174 vdd gnd cell_6t
Xbit_r175_c191 bl_191 br_191 wl_175 vdd gnd cell_6t
Xbit_r176_c191 bl_191 br_191 wl_176 vdd gnd cell_6t
Xbit_r177_c191 bl_191 br_191 wl_177 vdd gnd cell_6t
Xbit_r178_c191 bl_191 br_191 wl_178 vdd gnd cell_6t
Xbit_r179_c191 bl_191 br_191 wl_179 vdd gnd cell_6t
Xbit_r180_c191 bl_191 br_191 wl_180 vdd gnd cell_6t
Xbit_r181_c191 bl_191 br_191 wl_181 vdd gnd cell_6t
Xbit_r182_c191 bl_191 br_191 wl_182 vdd gnd cell_6t
Xbit_r183_c191 bl_191 br_191 wl_183 vdd gnd cell_6t
Xbit_r184_c191 bl_191 br_191 wl_184 vdd gnd cell_6t
Xbit_r185_c191 bl_191 br_191 wl_185 vdd gnd cell_6t
Xbit_r186_c191 bl_191 br_191 wl_186 vdd gnd cell_6t
Xbit_r187_c191 bl_191 br_191 wl_187 vdd gnd cell_6t
Xbit_r188_c191 bl_191 br_191 wl_188 vdd gnd cell_6t
Xbit_r189_c191 bl_191 br_191 wl_189 vdd gnd cell_6t
Xbit_r190_c191 bl_191 br_191 wl_190 vdd gnd cell_6t
Xbit_r191_c191 bl_191 br_191 wl_191 vdd gnd cell_6t
Xbit_r192_c191 bl_191 br_191 wl_192 vdd gnd cell_6t
Xbit_r193_c191 bl_191 br_191 wl_193 vdd gnd cell_6t
Xbit_r194_c191 bl_191 br_191 wl_194 vdd gnd cell_6t
Xbit_r195_c191 bl_191 br_191 wl_195 vdd gnd cell_6t
Xbit_r196_c191 bl_191 br_191 wl_196 vdd gnd cell_6t
Xbit_r197_c191 bl_191 br_191 wl_197 vdd gnd cell_6t
Xbit_r198_c191 bl_191 br_191 wl_198 vdd gnd cell_6t
Xbit_r199_c191 bl_191 br_191 wl_199 vdd gnd cell_6t
Xbit_r200_c191 bl_191 br_191 wl_200 vdd gnd cell_6t
Xbit_r201_c191 bl_191 br_191 wl_201 vdd gnd cell_6t
Xbit_r202_c191 bl_191 br_191 wl_202 vdd gnd cell_6t
Xbit_r203_c191 bl_191 br_191 wl_203 vdd gnd cell_6t
Xbit_r204_c191 bl_191 br_191 wl_204 vdd gnd cell_6t
Xbit_r205_c191 bl_191 br_191 wl_205 vdd gnd cell_6t
Xbit_r206_c191 bl_191 br_191 wl_206 vdd gnd cell_6t
Xbit_r207_c191 bl_191 br_191 wl_207 vdd gnd cell_6t
Xbit_r208_c191 bl_191 br_191 wl_208 vdd gnd cell_6t
Xbit_r209_c191 bl_191 br_191 wl_209 vdd gnd cell_6t
Xbit_r210_c191 bl_191 br_191 wl_210 vdd gnd cell_6t
Xbit_r211_c191 bl_191 br_191 wl_211 vdd gnd cell_6t
Xbit_r212_c191 bl_191 br_191 wl_212 vdd gnd cell_6t
Xbit_r213_c191 bl_191 br_191 wl_213 vdd gnd cell_6t
Xbit_r214_c191 bl_191 br_191 wl_214 vdd gnd cell_6t
Xbit_r215_c191 bl_191 br_191 wl_215 vdd gnd cell_6t
Xbit_r216_c191 bl_191 br_191 wl_216 vdd gnd cell_6t
Xbit_r217_c191 bl_191 br_191 wl_217 vdd gnd cell_6t
Xbit_r218_c191 bl_191 br_191 wl_218 vdd gnd cell_6t
Xbit_r219_c191 bl_191 br_191 wl_219 vdd gnd cell_6t
Xbit_r220_c191 bl_191 br_191 wl_220 vdd gnd cell_6t
Xbit_r221_c191 bl_191 br_191 wl_221 vdd gnd cell_6t
Xbit_r222_c191 bl_191 br_191 wl_222 vdd gnd cell_6t
Xbit_r223_c191 bl_191 br_191 wl_223 vdd gnd cell_6t
Xbit_r224_c191 bl_191 br_191 wl_224 vdd gnd cell_6t
Xbit_r225_c191 bl_191 br_191 wl_225 vdd gnd cell_6t
Xbit_r226_c191 bl_191 br_191 wl_226 vdd gnd cell_6t
Xbit_r227_c191 bl_191 br_191 wl_227 vdd gnd cell_6t
Xbit_r228_c191 bl_191 br_191 wl_228 vdd gnd cell_6t
Xbit_r229_c191 bl_191 br_191 wl_229 vdd gnd cell_6t
Xbit_r230_c191 bl_191 br_191 wl_230 vdd gnd cell_6t
Xbit_r231_c191 bl_191 br_191 wl_231 vdd gnd cell_6t
Xbit_r232_c191 bl_191 br_191 wl_232 vdd gnd cell_6t
Xbit_r233_c191 bl_191 br_191 wl_233 vdd gnd cell_6t
Xbit_r234_c191 bl_191 br_191 wl_234 vdd gnd cell_6t
Xbit_r235_c191 bl_191 br_191 wl_235 vdd gnd cell_6t
Xbit_r236_c191 bl_191 br_191 wl_236 vdd gnd cell_6t
Xbit_r237_c191 bl_191 br_191 wl_237 vdd gnd cell_6t
Xbit_r238_c191 bl_191 br_191 wl_238 vdd gnd cell_6t
Xbit_r239_c191 bl_191 br_191 wl_239 vdd gnd cell_6t
Xbit_r240_c191 bl_191 br_191 wl_240 vdd gnd cell_6t
Xbit_r241_c191 bl_191 br_191 wl_241 vdd gnd cell_6t
Xbit_r242_c191 bl_191 br_191 wl_242 vdd gnd cell_6t
Xbit_r243_c191 bl_191 br_191 wl_243 vdd gnd cell_6t
Xbit_r244_c191 bl_191 br_191 wl_244 vdd gnd cell_6t
Xbit_r245_c191 bl_191 br_191 wl_245 vdd gnd cell_6t
Xbit_r246_c191 bl_191 br_191 wl_246 vdd gnd cell_6t
Xbit_r247_c191 bl_191 br_191 wl_247 vdd gnd cell_6t
Xbit_r248_c191 bl_191 br_191 wl_248 vdd gnd cell_6t
Xbit_r249_c191 bl_191 br_191 wl_249 vdd gnd cell_6t
Xbit_r250_c191 bl_191 br_191 wl_250 vdd gnd cell_6t
Xbit_r251_c191 bl_191 br_191 wl_251 vdd gnd cell_6t
Xbit_r252_c191 bl_191 br_191 wl_252 vdd gnd cell_6t
Xbit_r253_c191 bl_191 br_191 wl_253 vdd gnd cell_6t
Xbit_r254_c191 bl_191 br_191 wl_254 vdd gnd cell_6t
Xbit_r255_c191 bl_191 br_191 wl_255 vdd gnd cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd cell_6t
Xbit_r1_c192 bl_192 br_192 wl_1 vdd gnd cell_6t
Xbit_r2_c192 bl_192 br_192 wl_2 vdd gnd cell_6t
Xbit_r3_c192 bl_192 br_192 wl_3 vdd gnd cell_6t
Xbit_r4_c192 bl_192 br_192 wl_4 vdd gnd cell_6t
Xbit_r5_c192 bl_192 br_192 wl_5 vdd gnd cell_6t
Xbit_r6_c192 bl_192 br_192 wl_6 vdd gnd cell_6t
Xbit_r7_c192 bl_192 br_192 wl_7 vdd gnd cell_6t
Xbit_r8_c192 bl_192 br_192 wl_8 vdd gnd cell_6t
Xbit_r9_c192 bl_192 br_192 wl_9 vdd gnd cell_6t
Xbit_r10_c192 bl_192 br_192 wl_10 vdd gnd cell_6t
Xbit_r11_c192 bl_192 br_192 wl_11 vdd gnd cell_6t
Xbit_r12_c192 bl_192 br_192 wl_12 vdd gnd cell_6t
Xbit_r13_c192 bl_192 br_192 wl_13 vdd gnd cell_6t
Xbit_r14_c192 bl_192 br_192 wl_14 vdd gnd cell_6t
Xbit_r15_c192 bl_192 br_192 wl_15 vdd gnd cell_6t
Xbit_r16_c192 bl_192 br_192 wl_16 vdd gnd cell_6t
Xbit_r17_c192 bl_192 br_192 wl_17 vdd gnd cell_6t
Xbit_r18_c192 bl_192 br_192 wl_18 vdd gnd cell_6t
Xbit_r19_c192 bl_192 br_192 wl_19 vdd gnd cell_6t
Xbit_r20_c192 bl_192 br_192 wl_20 vdd gnd cell_6t
Xbit_r21_c192 bl_192 br_192 wl_21 vdd gnd cell_6t
Xbit_r22_c192 bl_192 br_192 wl_22 vdd gnd cell_6t
Xbit_r23_c192 bl_192 br_192 wl_23 vdd gnd cell_6t
Xbit_r24_c192 bl_192 br_192 wl_24 vdd gnd cell_6t
Xbit_r25_c192 bl_192 br_192 wl_25 vdd gnd cell_6t
Xbit_r26_c192 bl_192 br_192 wl_26 vdd gnd cell_6t
Xbit_r27_c192 bl_192 br_192 wl_27 vdd gnd cell_6t
Xbit_r28_c192 bl_192 br_192 wl_28 vdd gnd cell_6t
Xbit_r29_c192 bl_192 br_192 wl_29 vdd gnd cell_6t
Xbit_r30_c192 bl_192 br_192 wl_30 vdd gnd cell_6t
Xbit_r31_c192 bl_192 br_192 wl_31 vdd gnd cell_6t
Xbit_r32_c192 bl_192 br_192 wl_32 vdd gnd cell_6t
Xbit_r33_c192 bl_192 br_192 wl_33 vdd gnd cell_6t
Xbit_r34_c192 bl_192 br_192 wl_34 vdd gnd cell_6t
Xbit_r35_c192 bl_192 br_192 wl_35 vdd gnd cell_6t
Xbit_r36_c192 bl_192 br_192 wl_36 vdd gnd cell_6t
Xbit_r37_c192 bl_192 br_192 wl_37 vdd gnd cell_6t
Xbit_r38_c192 bl_192 br_192 wl_38 vdd gnd cell_6t
Xbit_r39_c192 bl_192 br_192 wl_39 vdd gnd cell_6t
Xbit_r40_c192 bl_192 br_192 wl_40 vdd gnd cell_6t
Xbit_r41_c192 bl_192 br_192 wl_41 vdd gnd cell_6t
Xbit_r42_c192 bl_192 br_192 wl_42 vdd gnd cell_6t
Xbit_r43_c192 bl_192 br_192 wl_43 vdd gnd cell_6t
Xbit_r44_c192 bl_192 br_192 wl_44 vdd gnd cell_6t
Xbit_r45_c192 bl_192 br_192 wl_45 vdd gnd cell_6t
Xbit_r46_c192 bl_192 br_192 wl_46 vdd gnd cell_6t
Xbit_r47_c192 bl_192 br_192 wl_47 vdd gnd cell_6t
Xbit_r48_c192 bl_192 br_192 wl_48 vdd gnd cell_6t
Xbit_r49_c192 bl_192 br_192 wl_49 vdd gnd cell_6t
Xbit_r50_c192 bl_192 br_192 wl_50 vdd gnd cell_6t
Xbit_r51_c192 bl_192 br_192 wl_51 vdd gnd cell_6t
Xbit_r52_c192 bl_192 br_192 wl_52 vdd gnd cell_6t
Xbit_r53_c192 bl_192 br_192 wl_53 vdd gnd cell_6t
Xbit_r54_c192 bl_192 br_192 wl_54 vdd gnd cell_6t
Xbit_r55_c192 bl_192 br_192 wl_55 vdd gnd cell_6t
Xbit_r56_c192 bl_192 br_192 wl_56 vdd gnd cell_6t
Xbit_r57_c192 bl_192 br_192 wl_57 vdd gnd cell_6t
Xbit_r58_c192 bl_192 br_192 wl_58 vdd gnd cell_6t
Xbit_r59_c192 bl_192 br_192 wl_59 vdd gnd cell_6t
Xbit_r60_c192 bl_192 br_192 wl_60 vdd gnd cell_6t
Xbit_r61_c192 bl_192 br_192 wl_61 vdd gnd cell_6t
Xbit_r62_c192 bl_192 br_192 wl_62 vdd gnd cell_6t
Xbit_r63_c192 bl_192 br_192 wl_63 vdd gnd cell_6t
Xbit_r64_c192 bl_192 br_192 wl_64 vdd gnd cell_6t
Xbit_r65_c192 bl_192 br_192 wl_65 vdd gnd cell_6t
Xbit_r66_c192 bl_192 br_192 wl_66 vdd gnd cell_6t
Xbit_r67_c192 bl_192 br_192 wl_67 vdd gnd cell_6t
Xbit_r68_c192 bl_192 br_192 wl_68 vdd gnd cell_6t
Xbit_r69_c192 bl_192 br_192 wl_69 vdd gnd cell_6t
Xbit_r70_c192 bl_192 br_192 wl_70 vdd gnd cell_6t
Xbit_r71_c192 bl_192 br_192 wl_71 vdd gnd cell_6t
Xbit_r72_c192 bl_192 br_192 wl_72 vdd gnd cell_6t
Xbit_r73_c192 bl_192 br_192 wl_73 vdd gnd cell_6t
Xbit_r74_c192 bl_192 br_192 wl_74 vdd gnd cell_6t
Xbit_r75_c192 bl_192 br_192 wl_75 vdd gnd cell_6t
Xbit_r76_c192 bl_192 br_192 wl_76 vdd gnd cell_6t
Xbit_r77_c192 bl_192 br_192 wl_77 vdd gnd cell_6t
Xbit_r78_c192 bl_192 br_192 wl_78 vdd gnd cell_6t
Xbit_r79_c192 bl_192 br_192 wl_79 vdd gnd cell_6t
Xbit_r80_c192 bl_192 br_192 wl_80 vdd gnd cell_6t
Xbit_r81_c192 bl_192 br_192 wl_81 vdd gnd cell_6t
Xbit_r82_c192 bl_192 br_192 wl_82 vdd gnd cell_6t
Xbit_r83_c192 bl_192 br_192 wl_83 vdd gnd cell_6t
Xbit_r84_c192 bl_192 br_192 wl_84 vdd gnd cell_6t
Xbit_r85_c192 bl_192 br_192 wl_85 vdd gnd cell_6t
Xbit_r86_c192 bl_192 br_192 wl_86 vdd gnd cell_6t
Xbit_r87_c192 bl_192 br_192 wl_87 vdd gnd cell_6t
Xbit_r88_c192 bl_192 br_192 wl_88 vdd gnd cell_6t
Xbit_r89_c192 bl_192 br_192 wl_89 vdd gnd cell_6t
Xbit_r90_c192 bl_192 br_192 wl_90 vdd gnd cell_6t
Xbit_r91_c192 bl_192 br_192 wl_91 vdd gnd cell_6t
Xbit_r92_c192 bl_192 br_192 wl_92 vdd gnd cell_6t
Xbit_r93_c192 bl_192 br_192 wl_93 vdd gnd cell_6t
Xbit_r94_c192 bl_192 br_192 wl_94 vdd gnd cell_6t
Xbit_r95_c192 bl_192 br_192 wl_95 vdd gnd cell_6t
Xbit_r96_c192 bl_192 br_192 wl_96 vdd gnd cell_6t
Xbit_r97_c192 bl_192 br_192 wl_97 vdd gnd cell_6t
Xbit_r98_c192 bl_192 br_192 wl_98 vdd gnd cell_6t
Xbit_r99_c192 bl_192 br_192 wl_99 vdd gnd cell_6t
Xbit_r100_c192 bl_192 br_192 wl_100 vdd gnd cell_6t
Xbit_r101_c192 bl_192 br_192 wl_101 vdd gnd cell_6t
Xbit_r102_c192 bl_192 br_192 wl_102 vdd gnd cell_6t
Xbit_r103_c192 bl_192 br_192 wl_103 vdd gnd cell_6t
Xbit_r104_c192 bl_192 br_192 wl_104 vdd gnd cell_6t
Xbit_r105_c192 bl_192 br_192 wl_105 vdd gnd cell_6t
Xbit_r106_c192 bl_192 br_192 wl_106 vdd gnd cell_6t
Xbit_r107_c192 bl_192 br_192 wl_107 vdd gnd cell_6t
Xbit_r108_c192 bl_192 br_192 wl_108 vdd gnd cell_6t
Xbit_r109_c192 bl_192 br_192 wl_109 vdd gnd cell_6t
Xbit_r110_c192 bl_192 br_192 wl_110 vdd gnd cell_6t
Xbit_r111_c192 bl_192 br_192 wl_111 vdd gnd cell_6t
Xbit_r112_c192 bl_192 br_192 wl_112 vdd gnd cell_6t
Xbit_r113_c192 bl_192 br_192 wl_113 vdd gnd cell_6t
Xbit_r114_c192 bl_192 br_192 wl_114 vdd gnd cell_6t
Xbit_r115_c192 bl_192 br_192 wl_115 vdd gnd cell_6t
Xbit_r116_c192 bl_192 br_192 wl_116 vdd gnd cell_6t
Xbit_r117_c192 bl_192 br_192 wl_117 vdd gnd cell_6t
Xbit_r118_c192 bl_192 br_192 wl_118 vdd gnd cell_6t
Xbit_r119_c192 bl_192 br_192 wl_119 vdd gnd cell_6t
Xbit_r120_c192 bl_192 br_192 wl_120 vdd gnd cell_6t
Xbit_r121_c192 bl_192 br_192 wl_121 vdd gnd cell_6t
Xbit_r122_c192 bl_192 br_192 wl_122 vdd gnd cell_6t
Xbit_r123_c192 bl_192 br_192 wl_123 vdd gnd cell_6t
Xbit_r124_c192 bl_192 br_192 wl_124 vdd gnd cell_6t
Xbit_r125_c192 bl_192 br_192 wl_125 vdd gnd cell_6t
Xbit_r126_c192 bl_192 br_192 wl_126 vdd gnd cell_6t
Xbit_r127_c192 bl_192 br_192 wl_127 vdd gnd cell_6t
Xbit_r128_c192 bl_192 br_192 wl_128 vdd gnd cell_6t
Xbit_r129_c192 bl_192 br_192 wl_129 vdd gnd cell_6t
Xbit_r130_c192 bl_192 br_192 wl_130 vdd gnd cell_6t
Xbit_r131_c192 bl_192 br_192 wl_131 vdd gnd cell_6t
Xbit_r132_c192 bl_192 br_192 wl_132 vdd gnd cell_6t
Xbit_r133_c192 bl_192 br_192 wl_133 vdd gnd cell_6t
Xbit_r134_c192 bl_192 br_192 wl_134 vdd gnd cell_6t
Xbit_r135_c192 bl_192 br_192 wl_135 vdd gnd cell_6t
Xbit_r136_c192 bl_192 br_192 wl_136 vdd gnd cell_6t
Xbit_r137_c192 bl_192 br_192 wl_137 vdd gnd cell_6t
Xbit_r138_c192 bl_192 br_192 wl_138 vdd gnd cell_6t
Xbit_r139_c192 bl_192 br_192 wl_139 vdd gnd cell_6t
Xbit_r140_c192 bl_192 br_192 wl_140 vdd gnd cell_6t
Xbit_r141_c192 bl_192 br_192 wl_141 vdd gnd cell_6t
Xbit_r142_c192 bl_192 br_192 wl_142 vdd gnd cell_6t
Xbit_r143_c192 bl_192 br_192 wl_143 vdd gnd cell_6t
Xbit_r144_c192 bl_192 br_192 wl_144 vdd gnd cell_6t
Xbit_r145_c192 bl_192 br_192 wl_145 vdd gnd cell_6t
Xbit_r146_c192 bl_192 br_192 wl_146 vdd gnd cell_6t
Xbit_r147_c192 bl_192 br_192 wl_147 vdd gnd cell_6t
Xbit_r148_c192 bl_192 br_192 wl_148 vdd gnd cell_6t
Xbit_r149_c192 bl_192 br_192 wl_149 vdd gnd cell_6t
Xbit_r150_c192 bl_192 br_192 wl_150 vdd gnd cell_6t
Xbit_r151_c192 bl_192 br_192 wl_151 vdd gnd cell_6t
Xbit_r152_c192 bl_192 br_192 wl_152 vdd gnd cell_6t
Xbit_r153_c192 bl_192 br_192 wl_153 vdd gnd cell_6t
Xbit_r154_c192 bl_192 br_192 wl_154 vdd gnd cell_6t
Xbit_r155_c192 bl_192 br_192 wl_155 vdd gnd cell_6t
Xbit_r156_c192 bl_192 br_192 wl_156 vdd gnd cell_6t
Xbit_r157_c192 bl_192 br_192 wl_157 vdd gnd cell_6t
Xbit_r158_c192 bl_192 br_192 wl_158 vdd gnd cell_6t
Xbit_r159_c192 bl_192 br_192 wl_159 vdd gnd cell_6t
Xbit_r160_c192 bl_192 br_192 wl_160 vdd gnd cell_6t
Xbit_r161_c192 bl_192 br_192 wl_161 vdd gnd cell_6t
Xbit_r162_c192 bl_192 br_192 wl_162 vdd gnd cell_6t
Xbit_r163_c192 bl_192 br_192 wl_163 vdd gnd cell_6t
Xbit_r164_c192 bl_192 br_192 wl_164 vdd gnd cell_6t
Xbit_r165_c192 bl_192 br_192 wl_165 vdd gnd cell_6t
Xbit_r166_c192 bl_192 br_192 wl_166 vdd gnd cell_6t
Xbit_r167_c192 bl_192 br_192 wl_167 vdd gnd cell_6t
Xbit_r168_c192 bl_192 br_192 wl_168 vdd gnd cell_6t
Xbit_r169_c192 bl_192 br_192 wl_169 vdd gnd cell_6t
Xbit_r170_c192 bl_192 br_192 wl_170 vdd gnd cell_6t
Xbit_r171_c192 bl_192 br_192 wl_171 vdd gnd cell_6t
Xbit_r172_c192 bl_192 br_192 wl_172 vdd gnd cell_6t
Xbit_r173_c192 bl_192 br_192 wl_173 vdd gnd cell_6t
Xbit_r174_c192 bl_192 br_192 wl_174 vdd gnd cell_6t
Xbit_r175_c192 bl_192 br_192 wl_175 vdd gnd cell_6t
Xbit_r176_c192 bl_192 br_192 wl_176 vdd gnd cell_6t
Xbit_r177_c192 bl_192 br_192 wl_177 vdd gnd cell_6t
Xbit_r178_c192 bl_192 br_192 wl_178 vdd gnd cell_6t
Xbit_r179_c192 bl_192 br_192 wl_179 vdd gnd cell_6t
Xbit_r180_c192 bl_192 br_192 wl_180 vdd gnd cell_6t
Xbit_r181_c192 bl_192 br_192 wl_181 vdd gnd cell_6t
Xbit_r182_c192 bl_192 br_192 wl_182 vdd gnd cell_6t
Xbit_r183_c192 bl_192 br_192 wl_183 vdd gnd cell_6t
Xbit_r184_c192 bl_192 br_192 wl_184 vdd gnd cell_6t
Xbit_r185_c192 bl_192 br_192 wl_185 vdd gnd cell_6t
Xbit_r186_c192 bl_192 br_192 wl_186 vdd gnd cell_6t
Xbit_r187_c192 bl_192 br_192 wl_187 vdd gnd cell_6t
Xbit_r188_c192 bl_192 br_192 wl_188 vdd gnd cell_6t
Xbit_r189_c192 bl_192 br_192 wl_189 vdd gnd cell_6t
Xbit_r190_c192 bl_192 br_192 wl_190 vdd gnd cell_6t
Xbit_r191_c192 bl_192 br_192 wl_191 vdd gnd cell_6t
Xbit_r192_c192 bl_192 br_192 wl_192 vdd gnd cell_6t
Xbit_r193_c192 bl_192 br_192 wl_193 vdd gnd cell_6t
Xbit_r194_c192 bl_192 br_192 wl_194 vdd gnd cell_6t
Xbit_r195_c192 bl_192 br_192 wl_195 vdd gnd cell_6t
Xbit_r196_c192 bl_192 br_192 wl_196 vdd gnd cell_6t
Xbit_r197_c192 bl_192 br_192 wl_197 vdd gnd cell_6t
Xbit_r198_c192 bl_192 br_192 wl_198 vdd gnd cell_6t
Xbit_r199_c192 bl_192 br_192 wl_199 vdd gnd cell_6t
Xbit_r200_c192 bl_192 br_192 wl_200 vdd gnd cell_6t
Xbit_r201_c192 bl_192 br_192 wl_201 vdd gnd cell_6t
Xbit_r202_c192 bl_192 br_192 wl_202 vdd gnd cell_6t
Xbit_r203_c192 bl_192 br_192 wl_203 vdd gnd cell_6t
Xbit_r204_c192 bl_192 br_192 wl_204 vdd gnd cell_6t
Xbit_r205_c192 bl_192 br_192 wl_205 vdd gnd cell_6t
Xbit_r206_c192 bl_192 br_192 wl_206 vdd gnd cell_6t
Xbit_r207_c192 bl_192 br_192 wl_207 vdd gnd cell_6t
Xbit_r208_c192 bl_192 br_192 wl_208 vdd gnd cell_6t
Xbit_r209_c192 bl_192 br_192 wl_209 vdd gnd cell_6t
Xbit_r210_c192 bl_192 br_192 wl_210 vdd gnd cell_6t
Xbit_r211_c192 bl_192 br_192 wl_211 vdd gnd cell_6t
Xbit_r212_c192 bl_192 br_192 wl_212 vdd gnd cell_6t
Xbit_r213_c192 bl_192 br_192 wl_213 vdd gnd cell_6t
Xbit_r214_c192 bl_192 br_192 wl_214 vdd gnd cell_6t
Xbit_r215_c192 bl_192 br_192 wl_215 vdd gnd cell_6t
Xbit_r216_c192 bl_192 br_192 wl_216 vdd gnd cell_6t
Xbit_r217_c192 bl_192 br_192 wl_217 vdd gnd cell_6t
Xbit_r218_c192 bl_192 br_192 wl_218 vdd gnd cell_6t
Xbit_r219_c192 bl_192 br_192 wl_219 vdd gnd cell_6t
Xbit_r220_c192 bl_192 br_192 wl_220 vdd gnd cell_6t
Xbit_r221_c192 bl_192 br_192 wl_221 vdd gnd cell_6t
Xbit_r222_c192 bl_192 br_192 wl_222 vdd gnd cell_6t
Xbit_r223_c192 bl_192 br_192 wl_223 vdd gnd cell_6t
Xbit_r224_c192 bl_192 br_192 wl_224 vdd gnd cell_6t
Xbit_r225_c192 bl_192 br_192 wl_225 vdd gnd cell_6t
Xbit_r226_c192 bl_192 br_192 wl_226 vdd gnd cell_6t
Xbit_r227_c192 bl_192 br_192 wl_227 vdd gnd cell_6t
Xbit_r228_c192 bl_192 br_192 wl_228 vdd gnd cell_6t
Xbit_r229_c192 bl_192 br_192 wl_229 vdd gnd cell_6t
Xbit_r230_c192 bl_192 br_192 wl_230 vdd gnd cell_6t
Xbit_r231_c192 bl_192 br_192 wl_231 vdd gnd cell_6t
Xbit_r232_c192 bl_192 br_192 wl_232 vdd gnd cell_6t
Xbit_r233_c192 bl_192 br_192 wl_233 vdd gnd cell_6t
Xbit_r234_c192 bl_192 br_192 wl_234 vdd gnd cell_6t
Xbit_r235_c192 bl_192 br_192 wl_235 vdd gnd cell_6t
Xbit_r236_c192 bl_192 br_192 wl_236 vdd gnd cell_6t
Xbit_r237_c192 bl_192 br_192 wl_237 vdd gnd cell_6t
Xbit_r238_c192 bl_192 br_192 wl_238 vdd gnd cell_6t
Xbit_r239_c192 bl_192 br_192 wl_239 vdd gnd cell_6t
Xbit_r240_c192 bl_192 br_192 wl_240 vdd gnd cell_6t
Xbit_r241_c192 bl_192 br_192 wl_241 vdd gnd cell_6t
Xbit_r242_c192 bl_192 br_192 wl_242 vdd gnd cell_6t
Xbit_r243_c192 bl_192 br_192 wl_243 vdd gnd cell_6t
Xbit_r244_c192 bl_192 br_192 wl_244 vdd gnd cell_6t
Xbit_r245_c192 bl_192 br_192 wl_245 vdd gnd cell_6t
Xbit_r246_c192 bl_192 br_192 wl_246 vdd gnd cell_6t
Xbit_r247_c192 bl_192 br_192 wl_247 vdd gnd cell_6t
Xbit_r248_c192 bl_192 br_192 wl_248 vdd gnd cell_6t
Xbit_r249_c192 bl_192 br_192 wl_249 vdd gnd cell_6t
Xbit_r250_c192 bl_192 br_192 wl_250 vdd gnd cell_6t
Xbit_r251_c192 bl_192 br_192 wl_251 vdd gnd cell_6t
Xbit_r252_c192 bl_192 br_192 wl_252 vdd gnd cell_6t
Xbit_r253_c192 bl_192 br_192 wl_253 vdd gnd cell_6t
Xbit_r254_c192 bl_192 br_192 wl_254 vdd gnd cell_6t
Xbit_r255_c192 bl_192 br_192 wl_255 vdd gnd cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd cell_6t
Xbit_r1_c193 bl_193 br_193 wl_1 vdd gnd cell_6t
Xbit_r2_c193 bl_193 br_193 wl_2 vdd gnd cell_6t
Xbit_r3_c193 bl_193 br_193 wl_3 vdd gnd cell_6t
Xbit_r4_c193 bl_193 br_193 wl_4 vdd gnd cell_6t
Xbit_r5_c193 bl_193 br_193 wl_5 vdd gnd cell_6t
Xbit_r6_c193 bl_193 br_193 wl_6 vdd gnd cell_6t
Xbit_r7_c193 bl_193 br_193 wl_7 vdd gnd cell_6t
Xbit_r8_c193 bl_193 br_193 wl_8 vdd gnd cell_6t
Xbit_r9_c193 bl_193 br_193 wl_9 vdd gnd cell_6t
Xbit_r10_c193 bl_193 br_193 wl_10 vdd gnd cell_6t
Xbit_r11_c193 bl_193 br_193 wl_11 vdd gnd cell_6t
Xbit_r12_c193 bl_193 br_193 wl_12 vdd gnd cell_6t
Xbit_r13_c193 bl_193 br_193 wl_13 vdd gnd cell_6t
Xbit_r14_c193 bl_193 br_193 wl_14 vdd gnd cell_6t
Xbit_r15_c193 bl_193 br_193 wl_15 vdd gnd cell_6t
Xbit_r16_c193 bl_193 br_193 wl_16 vdd gnd cell_6t
Xbit_r17_c193 bl_193 br_193 wl_17 vdd gnd cell_6t
Xbit_r18_c193 bl_193 br_193 wl_18 vdd gnd cell_6t
Xbit_r19_c193 bl_193 br_193 wl_19 vdd gnd cell_6t
Xbit_r20_c193 bl_193 br_193 wl_20 vdd gnd cell_6t
Xbit_r21_c193 bl_193 br_193 wl_21 vdd gnd cell_6t
Xbit_r22_c193 bl_193 br_193 wl_22 vdd gnd cell_6t
Xbit_r23_c193 bl_193 br_193 wl_23 vdd gnd cell_6t
Xbit_r24_c193 bl_193 br_193 wl_24 vdd gnd cell_6t
Xbit_r25_c193 bl_193 br_193 wl_25 vdd gnd cell_6t
Xbit_r26_c193 bl_193 br_193 wl_26 vdd gnd cell_6t
Xbit_r27_c193 bl_193 br_193 wl_27 vdd gnd cell_6t
Xbit_r28_c193 bl_193 br_193 wl_28 vdd gnd cell_6t
Xbit_r29_c193 bl_193 br_193 wl_29 vdd gnd cell_6t
Xbit_r30_c193 bl_193 br_193 wl_30 vdd gnd cell_6t
Xbit_r31_c193 bl_193 br_193 wl_31 vdd gnd cell_6t
Xbit_r32_c193 bl_193 br_193 wl_32 vdd gnd cell_6t
Xbit_r33_c193 bl_193 br_193 wl_33 vdd gnd cell_6t
Xbit_r34_c193 bl_193 br_193 wl_34 vdd gnd cell_6t
Xbit_r35_c193 bl_193 br_193 wl_35 vdd gnd cell_6t
Xbit_r36_c193 bl_193 br_193 wl_36 vdd gnd cell_6t
Xbit_r37_c193 bl_193 br_193 wl_37 vdd gnd cell_6t
Xbit_r38_c193 bl_193 br_193 wl_38 vdd gnd cell_6t
Xbit_r39_c193 bl_193 br_193 wl_39 vdd gnd cell_6t
Xbit_r40_c193 bl_193 br_193 wl_40 vdd gnd cell_6t
Xbit_r41_c193 bl_193 br_193 wl_41 vdd gnd cell_6t
Xbit_r42_c193 bl_193 br_193 wl_42 vdd gnd cell_6t
Xbit_r43_c193 bl_193 br_193 wl_43 vdd gnd cell_6t
Xbit_r44_c193 bl_193 br_193 wl_44 vdd gnd cell_6t
Xbit_r45_c193 bl_193 br_193 wl_45 vdd gnd cell_6t
Xbit_r46_c193 bl_193 br_193 wl_46 vdd gnd cell_6t
Xbit_r47_c193 bl_193 br_193 wl_47 vdd gnd cell_6t
Xbit_r48_c193 bl_193 br_193 wl_48 vdd gnd cell_6t
Xbit_r49_c193 bl_193 br_193 wl_49 vdd gnd cell_6t
Xbit_r50_c193 bl_193 br_193 wl_50 vdd gnd cell_6t
Xbit_r51_c193 bl_193 br_193 wl_51 vdd gnd cell_6t
Xbit_r52_c193 bl_193 br_193 wl_52 vdd gnd cell_6t
Xbit_r53_c193 bl_193 br_193 wl_53 vdd gnd cell_6t
Xbit_r54_c193 bl_193 br_193 wl_54 vdd gnd cell_6t
Xbit_r55_c193 bl_193 br_193 wl_55 vdd gnd cell_6t
Xbit_r56_c193 bl_193 br_193 wl_56 vdd gnd cell_6t
Xbit_r57_c193 bl_193 br_193 wl_57 vdd gnd cell_6t
Xbit_r58_c193 bl_193 br_193 wl_58 vdd gnd cell_6t
Xbit_r59_c193 bl_193 br_193 wl_59 vdd gnd cell_6t
Xbit_r60_c193 bl_193 br_193 wl_60 vdd gnd cell_6t
Xbit_r61_c193 bl_193 br_193 wl_61 vdd gnd cell_6t
Xbit_r62_c193 bl_193 br_193 wl_62 vdd gnd cell_6t
Xbit_r63_c193 bl_193 br_193 wl_63 vdd gnd cell_6t
Xbit_r64_c193 bl_193 br_193 wl_64 vdd gnd cell_6t
Xbit_r65_c193 bl_193 br_193 wl_65 vdd gnd cell_6t
Xbit_r66_c193 bl_193 br_193 wl_66 vdd gnd cell_6t
Xbit_r67_c193 bl_193 br_193 wl_67 vdd gnd cell_6t
Xbit_r68_c193 bl_193 br_193 wl_68 vdd gnd cell_6t
Xbit_r69_c193 bl_193 br_193 wl_69 vdd gnd cell_6t
Xbit_r70_c193 bl_193 br_193 wl_70 vdd gnd cell_6t
Xbit_r71_c193 bl_193 br_193 wl_71 vdd gnd cell_6t
Xbit_r72_c193 bl_193 br_193 wl_72 vdd gnd cell_6t
Xbit_r73_c193 bl_193 br_193 wl_73 vdd gnd cell_6t
Xbit_r74_c193 bl_193 br_193 wl_74 vdd gnd cell_6t
Xbit_r75_c193 bl_193 br_193 wl_75 vdd gnd cell_6t
Xbit_r76_c193 bl_193 br_193 wl_76 vdd gnd cell_6t
Xbit_r77_c193 bl_193 br_193 wl_77 vdd gnd cell_6t
Xbit_r78_c193 bl_193 br_193 wl_78 vdd gnd cell_6t
Xbit_r79_c193 bl_193 br_193 wl_79 vdd gnd cell_6t
Xbit_r80_c193 bl_193 br_193 wl_80 vdd gnd cell_6t
Xbit_r81_c193 bl_193 br_193 wl_81 vdd gnd cell_6t
Xbit_r82_c193 bl_193 br_193 wl_82 vdd gnd cell_6t
Xbit_r83_c193 bl_193 br_193 wl_83 vdd gnd cell_6t
Xbit_r84_c193 bl_193 br_193 wl_84 vdd gnd cell_6t
Xbit_r85_c193 bl_193 br_193 wl_85 vdd gnd cell_6t
Xbit_r86_c193 bl_193 br_193 wl_86 vdd gnd cell_6t
Xbit_r87_c193 bl_193 br_193 wl_87 vdd gnd cell_6t
Xbit_r88_c193 bl_193 br_193 wl_88 vdd gnd cell_6t
Xbit_r89_c193 bl_193 br_193 wl_89 vdd gnd cell_6t
Xbit_r90_c193 bl_193 br_193 wl_90 vdd gnd cell_6t
Xbit_r91_c193 bl_193 br_193 wl_91 vdd gnd cell_6t
Xbit_r92_c193 bl_193 br_193 wl_92 vdd gnd cell_6t
Xbit_r93_c193 bl_193 br_193 wl_93 vdd gnd cell_6t
Xbit_r94_c193 bl_193 br_193 wl_94 vdd gnd cell_6t
Xbit_r95_c193 bl_193 br_193 wl_95 vdd gnd cell_6t
Xbit_r96_c193 bl_193 br_193 wl_96 vdd gnd cell_6t
Xbit_r97_c193 bl_193 br_193 wl_97 vdd gnd cell_6t
Xbit_r98_c193 bl_193 br_193 wl_98 vdd gnd cell_6t
Xbit_r99_c193 bl_193 br_193 wl_99 vdd gnd cell_6t
Xbit_r100_c193 bl_193 br_193 wl_100 vdd gnd cell_6t
Xbit_r101_c193 bl_193 br_193 wl_101 vdd gnd cell_6t
Xbit_r102_c193 bl_193 br_193 wl_102 vdd gnd cell_6t
Xbit_r103_c193 bl_193 br_193 wl_103 vdd gnd cell_6t
Xbit_r104_c193 bl_193 br_193 wl_104 vdd gnd cell_6t
Xbit_r105_c193 bl_193 br_193 wl_105 vdd gnd cell_6t
Xbit_r106_c193 bl_193 br_193 wl_106 vdd gnd cell_6t
Xbit_r107_c193 bl_193 br_193 wl_107 vdd gnd cell_6t
Xbit_r108_c193 bl_193 br_193 wl_108 vdd gnd cell_6t
Xbit_r109_c193 bl_193 br_193 wl_109 vdd gnd cell_6t
Xbit_r110_c193 bl_193 br_193 wl_110 vdd gnd cell_6t
Xbit_r111_c193 bl_193 br_193 wl_111 vdd gnd cell_6t
Xbit_r112_c193 bl_193 br_193 wl_112 vdd gnd cell_6t
Xbit_r113_c193 bl_193 br_193 wl_113 vdd gnd cell_6t
Xbit_r114_c193 bl_193 br_193 wl_114 vdd gnd cell_6t
Xbit_r115_c193 bl_193 br_193 wl_115 vdd gnd cell_6t
Xbit_r116_c193 bl_193 br_193 wl_116 vdd gnd cell_6t
Xbit_r117_c193 bl_193 br_193 wl_117 vdd gnd cell_6t
Xbit_r118_c193 bl_193 br_193 wl_118 vdd gnd cell_6t
Xbit_r119_c193 bl_193 br_193 wl_119 vdd gnd cell_6t
Xbit_r120_c193 bl_193 br_193 wl_120 vdd gnd cell_6t
Xbit_r121_c193 bl_193 br_193 wl_121 vdd gnd cell_6t
Xbit_r122_c193 bl_193 br_193 wl_122 vdd gnd cell_6t
Xbit_r123_c193 bl_193 br_193 wl_123 vdd gnd cell_6t
Xbit_r124_c193 bl_193 br_193 wl_124 vdd gnd cell_6t
Xbit_r125_c193 bl_193 br_193 wl_125 vdd gnd cell_6t
Xbit_r126_c193 bl_193 br_193 wl_126 vdd gnd cell_6t
Xbit_r127_c193 bl_193 br_193 wl_127 vdd gnd cell_6t
Xbit_r128_c193 bl_193 br_193 wl_128 vdd gnd cell_6t
Xbit_r129_c193 bl_193 br_193 wl_129 vdd gnd cell_6t
Xbit_r130_c193 bl_193 br_193 wl_130 vdd gnd cell_6t
Xbit_r131_c193 bl_193 br_193 wl_131 vdd gnd cell_6t
Xbit_r132_c193 bl_193 br_193 wl_132 vdd gnd cell_6t
Xbit_r133_c193 bl_193 br_193 wl_133 vdd gnd cell_6t
Xbit_r134_c193 bl_193 br_193 wl_134 vdd gnd cell_6t
Xbit_r135_c193 bl_193 br_193 wl_135 vdd gnd cell_6t
Xbit_r136_c193 bl_193 br_193 wl_136 vdd gnd cell_6t
Xbit_r137_c193 bl_193 br_193 wl_137 vdd gnd cell_6t
Xbit_r138_c193 bl_193 br_193 wl_138 vdd gnd cell_6t
Xbit_r139_c193 bl_193 br_193 wl_139 vdd gnd cell_6t
Xbit_r140_c193 bl_193 br_193 wl_140 vdd gnd cell_6t
Xbit_r141_c193 bl_193 br_193 wl_141 vdd gnd cell_6t
Xbit_r142_c193 bl_193 br_193 wl_142 vdd gnd cell_6t
Xbit_r143_c193 bl_193 br_193 wl_143 vdd gnd cell_6t
Xbit_r144_c193 bl_193 br_193 wl_144 vdd gnd cell_6t
Xbit_r145_c193 bl_193 br_193 wl_145 vdd gnd cell_6t
Xbit_r146_c193 bl_193 br_193 wl_146 vdd gnd cell_6t
Xbit_r147_c193 bl_193 br_193 wl_147 vdd gnd cell_6t
Xbit_r148_c193 bl_193 br_193 wl_148 vdd gnd cell_6t
Xbit_r149_c193 bl_193 br_193 wl_149 vdd gnd cell_6t
Xbit_r150_c193 bl_193 br_193 wl_150 vdd gnd cell_6t
Xbit_r151_c193 bl_193 br_193 wl_151 vdd gnd cell_6t
Xbit_r152_c193 bl_193 br_193 wl_152 vdd gnd cell_6t
Xbit_r153_c193 bl_193 br_193 wl_153 vdd gnd cell_6t
Xbit_r154_c193 bl_193 br_193 wl_154 vdd gnd cell_6t
Xbit_r155_c193 bl_193 br_193 wl_155 vdd gnd cell_6t
Xbit_r156_c193 bl_193 br_193 wl_156 vdd gnd cell_6t
Xbit_r157_c193 bl_193 br_193 wl_157 vdd gnd cell_6t
Xbit_r158_c193 bl_193 br_193 wl_158 vdd gnd cell_6t
Xbit_r159_c193 bl_193 br_193 wl_159 vdd gnd cell_6t
Xbit_r160_c193 bl_193 br_193 wl_160 vdd gnd cell_6t
Xbit_r161_c193 bl_193 br_193 wl_161 vdd gnd cell_6t
Xbit_r162_c193 bl_193 br_193 wl_162 vdd gnd cell_6t
Xbit_r163_c193 bl_193 br_193 wl_163 vdd gnd cell_6t
Xbit_r164_c193 bl_193 br_193 wl_164 vdd gnd cell_6t
Xbit_r165_c193 bl_193 br_193 wl_165 vdd gnd cell_6t
Xbit_r166_c193 bl_193 br_193 wl_166 vdd gnd cell_6t
Xbit_r167_c193 bl_193 br_193 wl_167 vdd gnd cell_6t
Xbit_r168_c193 bl_193 br_193 wl_168 vdd gnd cell_6t
Xbit_r169_c193 bl_193 br_193 wl_169 vdd gnd cell_6t
Xbit_r170_c193 bl_193 br_193 wl_170 vdd gnd cell_6t
Xbit_r171_c193 bl_193 br_193 wl_171 vdd gnd cell_6t
Xbit_r172_c193 bl_193 br_193 wl_172 vdd gnd cell_6t
Xbit_r173_c193 bl_193 br_193 wl_173 vdd gnd cell_6t
Xbit_r174_c193 bl_193 br_193 wl_174 vdd gnd cell_6t
Xbit_r175_c193 bl_193 br_193 wl_175 vdd gnd cell_6t
Xbit_r176_c193 bl_193 br_193 wl_176 vdd gnd cell_6t
Xbit_r177_c193 bl_193 br_193 wl_177 vdd gnd cell_6t
Xbit_r178_c193 bl_193 br_193 wl_178 vdd gnd cell_6t
Xbit_r179_c193 bl_193 br_193 wl_179 vdd gnd cell_6t
Xbit_r180_c193 bl_193 br_193 wl_180 vdd gnd cell_6t
Xbit_r181_c193 bl_193 br_193 wl_181 vdd gnd cell_6t
Xbit_r182_c193 bl_193 br_193 wl_182 vdd gnd cell_6t
Xbit_r183_c193 bl_193 br_193 wl_183 vdd gnd cell_6t
Xbit_r184_c193 bl_193 br_193 wl_184 vdd gnd cell_6t
Xbit_r185_c193 bl_193 br_193 wl_185 vdd gnd cell_6t
Xbit_r186_c193 bl_193 br_193 wl_186 vdd gnd cell_6t
Xbit_r187_c193 bl_193 br_193 wl_187 vdd gnd cell_6t
Xbit_r188_c193 bl_193 br_193 wl_188 vdd gnd cell_6t
Xbit_r189_c193 bl_193 br_193 wl_189 vdd gnd cell_6t
Xbit_r190_c193 bl_193 br_193 wl_190 vdd gnd cell_6t
Xbit_r191_c193 bl_193 br_193 wl_191 vdd gnd cell_6t
Xbit_r192_c193 bl_193 br_193 wl_192 vdd gnd cell_6t
Xbit_r193_c193 bl_193 br_193 wl_193 vdd gnd cell_6t
Xbit_r194_c193 bl_193 br_193 wl_194 vdd gnd cell_6t
Xbit_r195_c193 bl_193 br_193 wl_195 vdd gnd cell_6t
Xbit_r196_c193 bl_193 br_193 wl_196 vdd gnd cell_6t
Xbit_r197_c193 bl_193 br_193 wl_197 vdd gnd cell_6t
Xbit_r198_c193 bl_193 br_193 wl_198 vdd gnd cell_6t
Xbit_r199_c193 bl_193 br_193 wl_199 vdd gnd cell_6t
Xbit_r200_c193 bl_193 br_193 wl_200 vdd gnd cell_6t
Xbit_r201_c193 bl_193 br_193 wl_201 vdd gnd cell_6t
Xbit_r202_c193 bl_193 br_193 wl_202 vdd gnd cell_6t
Xbit_r203_c193 bl_193 br_193 wl_203 vdd gnd cell_6t
Xbit_r204_c193 bl_193 br_193 wl_204 vdd gnd cell_6t
Xbit_r205_c193 bl_193 br_193 wl_205 vdd gnd cell_6t
Xbit_r206_c193 bl_193 br_193 wl_206 vdd gnd cell_6t
Xbit_r207_c193 bl_193 br_193 wl_207 vdd gnd cell_6t
Xbit_r208_c193 bl_193 br_193 wl_208 vdd gnd cell_6t
Xbit_r209_c193 bl_193 br_193 wl_209 vdd gnd cell_6t
Xbit_r210_c193 bl_193 br_193 wl_210 vdd gnd cell_6t
Xbit_r211_c193 bl_193 br_193 wl_211 vdd gnd cell_6t
Xbit_r212_c193 bl_193 br_193 wl_212 vdd gnd cell_6t
Xbit_r213_c193 bl_193 br_193 wl_213 vdd gnd cell_6t
Xbit_r214_c193 bl_193 br_193 wl_214 vdd gnd cell_6t
Xbit_r215_c193 bl_193 br_193 wl_215 vdd gnd cell_6t
Xbit_r216_c193 bl_193 br_193 wl_216 vdd gnd cell_6t
Xbit_r217_c193 bl_193 br_193 wl_217 vdd gnd cell_6t
Xbit_r218_c193 bl_193 br_193 wl_218 vdd gnd cell_6t
Xbit_r219_c193 bl_193 br_193 wl_219 vdd gnd cell_6t
Xbit_r220_c193 bl_193 br_193 wl_220 vdd gnd cell_6t
Xbit_r221_c193 bl_193 br_193 wl_221 vdd gnd cell_6t
Xbit_r222_c193 bl_193 br_193 wl_222 vdd gnd cell_6t
Xbit_r223_c193 bl_193 br_193 wl_223 vdd gnd cell_6t
Xbit_r224_c193 bl_193 br_193 wl_224 vdd gnd cell_6t
Xbit_r225_c193 bl_193 br_193 wl_225 vdd gnd cell_6t
Xbit_r226_c193 bl_193 br_193 wl_226 vdd gnd cell_6t
Xbit_r227_c193 bl_193 br_193 wl_227 vdd gnd cell_6t
Xbit_r228_c193 bl_193 br_193 wl_228 vdd gnd cell_6t
Xbit_r229_c193 bl_193 br_193 wl_229 vdd gnd cell_6t
Xbit_r230_c193 bl_193 br_193 wl_230 vdd gnd cell_6t
Xbit_r231_c193 bl_193 br_193 wl_231 vdd gnd cell_6t
Xbit_r232_c193 bl_193 br_193 wl_232 vdd gnd cell_6t
Xbit_r233_c193 bl_193 br_193 wl_233 vdd gnd cell_6t
Xbit_r234_c193 bl_193 br_193 wl_234 vdd gnd cell_6t
Xbit_r235_c193 bl_193 br_193 wl_235 vdd gnd cell_6t
Xbit_r236_c193 bl_193 br_193 wl_236 vdd gnd cell_6t
Xbit_r237_c193 bl_193 br_193 wl_237 vdd gnd cell_6t
Xbit_r238_c193 bl_193 br_193 wl_238 vdd gnd cell_6t
Xbit_r239_c193 bl_193 br_193 wl_239 vdd gnd cell_6t
Xbit_r240_c193 bl_193 br_193 wl_240 vdd gnd cell_6t
Xbit_r241_c193 bl_193 br_193 wl_241 vdd gnd cell_6t
Xbit_r242_c193 bl_193 br_193 wl_242 vdd gnd cell_6t
Xbit_r243_c193 bl_193 br_193 wl_243 vdd gnd cell_6t
Xbit_r244_c193 bl_193 br_193 wl_244 vdd gnd cell_6t
Xbit_r245_c193 bl_193 br_193 wl_245 vdd gnd cell_6t
Xbit_r246_c193 bl_193 br_193 wl_246 vdd gnd cell_6t
Xbit_r247_c193 bl_193 br_193 wl_247 vdd gnd cell_6t
Xbit_r248_c193 bl_193 br_193 wl_248 vdd gnd cell_6t
Xbit_r249_c193 bl_193 br_193 wl_249 vdd gnd cell_6t
Xbit_r250_c193 bl_193 br_193 wl_250 vdd gnd cell_6t
Xbit_r251_c193 bl_193 br_193 wl_251 vdd gnd cell_6t
Xbit_r252_c193 bl_193 br_193 wl_252 vdd gnd cell_6t
Xbit_r253_c193 bl_193 br_193 wl_253 vdd gnd cell_6t
Xbit_r254_c193 bl_193 br_193 wl_254 vdd gnd cell_6t
Xbit_r255_c193 bl_193 br_193 wl_255 vdd gnd cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd cell_6t
Xbit_r1_c194 bl_194 br_194 wl_1 vdd gnd cell_6t
Xbit_r2_c194 bl_194 br_194 wl_2 vdd gnd cell_6t
Xbit_r3_c194 bl_194 br_194 wl_3 vdd gnd cell_6t
Xbit_r4_c194 bl_194 br_194 wl_4 vdd gnd cell_6t
Xbit_r5_c194 bl_194 br_194 wl_5 vdd gnd cell_6t
Xbit_r6_c194 bl_194 br_194 wl_6 vdd gnd cell_6t
Xbit_r7_c194 bl_194 br_194 wl_7 vdd gnd cell_6t
Xbit_r8_c194 bl_194 br_194 wl_8 vdd gnd cell_6t
Xbit_r9_c194 bl_194 br_194 wl_9 vdd gnd cell_6t
Xbit_r10_c194 bl_194 br_194 wl_10 vdd gnd cell_6t
Xbit_r11_c194 bl_194 br_194 wl_11 vdd gnd cell_6t
Xbit_r12_c194 bl_194 br_194 wl_12 vdd gnd cell_6t
Xbit_r13_c194 bl_194 br_194 wl_13 vdd gnd cell_6t
Xbit_r14_c194 bl_194 br_194 wl_14 vdd gnd cell_6t
Xbit_r15_c194 bl_194 br_194 wl_15 vdd gnd cell_6t
Xbit_r16_c194 bl_194 br_194 wl_16 vdd gnd cell_6t
Xbit_r17_c194 bl_194 br_194 wl_17 vdd gnd cell_6t
Xbit_r18_c194 bl_194 br_194 wl_18 vdd gnd cell_6t
Xbit_r19_c194 bl_194 br_194 wl_19 vdd gnd cell_6t
Xbit_r20_c194 bl_194 br_194 wl_20 vdd gnd cell_6t
Xbit_r21_c194 bl_194 br_194 wl_21 vdd gnd cell_6t
Xbit_r22_c194 bl_194 br_194 wl_22 vdd gnd cell_6t
Xbit_r23_c194 bl_194 br_194 wl_23 vdd gnd cell_6t
Xbit_r24_c194 bl_194 br_194 wl_24 vdd gnd cell_6t
Xbit_r25_c194 bl_194 br_194 wl_25 vdd gnd cell_6t
Xbit_r26_c194 bl_194 br_194 wl_26 vdd gnd cell_6t
Xbit_r27_c194 bl_194 br_194 wl_27 vdd gnd cell_6t
Xbit_r28_c194 bl_194 br_194 wl_28 vdd gnd cell_6t
Xbit_r29_c194 bl_194 br_194 wl_29 vdd gnd cell_6t
Xbit_r30_c194 bl_194 br_194 wl_30 vdd gnd cell_6t
Xbit_r31_c194 bl_194 br_194 wl_31 vdd gnd cell_6t
Xbit_r32_c194 bl_194 br_194 wl_32 vdd gnd cell_6t
Xbit_r33_c194 bl_194 br_194 wl_33 vdd gnd cell_6t
Xbit_r34_c194 bl_194 br_194 wl_34 vdd gnd cell_6t
Xbit_r35_c194 bl_194 br_194 wl_35 vdd gnd cell_6t
Xbit_r36_c194 bl_194 br_194 wl_36 vdd gnd cell_6t
Xbit_r37_c194 bl_194 br_194 wl_37 vdd gnd cell_6t
Xbit_r38_c194 bl_194 br_194 wl_38 vdd gnd cell_6t
Xbit_r39_c194 bl_194 br_194 wl_39 vdd gnd cell_6t
Xbit_r40_c194 bl_194 br_194 wl_40 vdd gnd cell_6t
Xbit_r41_c194 bl_194 br_194 wl_41 vdd gnd cell_6t
Xbit_r42_c194 bl_194 br_194 wl_42 vdd gnd cell_6t
Xbit_r43_c194 bl_194 br_194 wl_43 vdd gnd cell_6t
Xbit_r44_c194 bl_194 br_194 wl_44 vdd gnd cell_6t
Xbit_r45_c194 bl_194 br_194 wl_45 vdd gnd cell_6t
Xbit_r46_c194 bl_194 br_194 wl_46 vdd gnd cell_6t
Xbit_r47_c194 bl_194 br_194 wl_47 vdd gnd cell_6t
Xbit_r48_c194 bl_194 br_194 wl_48 vdd gnd cell_6t
Xbit_r49_c194 bl_194 br_194 wl_49 vdd gnd cell_6t
Xbit_r50_c194 bl_194 br_194 wl_50 vdd gnd cell_6t
Xbit_r51_c194 bl_194 br_194 wl_51 vdd gnd cell_6t
Xbit_r52_c194 bl_194 br_194 wl_52 vdd gnd cell_6t
Xbit_r53_c194 bl_194 br_194 wl_53 vdd gnd cell_6t
Xbit_r54_c194 bl_194 br_194 wl_54 vdd gnd cell_6t
Xbit_r55_c194 bl_194 br_194 wl_55 vdd gnd cell_6t
Xbit_r56_c194 bl_194 br_194 wl_56 vdd gnd cell_6t
Xbit_r57_c194 bl_194 br_194 wl_57 vdd gnd cell_6t
Xbit_r58_c194 bl_194 br_194 wl_58 vdd gnd cell_6t
Xbit_r59_c194 bl_194 br_194 wl_59 vdd gnd cell_6t
Xbit_r60_c194 bl_194 br_194 wl_60 vdd gnd cell_6t
Xbit_r61_c194 bl_194 br_194 wl_61 vdd gnd cell_6t
Xbit_r62_c194 bl_194 br_194 wl_62 vdd gnd cell_6t
Xbit_r63_c194 bl_194 br_194 wl_63 vdd gnd cell_6t
Xbit_r64_c194 bl_194 br_194 wl_64 vdd gnd cell_6t
Xbit_r65_c194 bl_194 br_194 wl_65 vdd gnd cell_6t
Xbit_r66_c194 bl_194 br_194 wl_66 vdd gnd cell_6t
Xbit_r67_c194 bl_194 br_194 wl_67 vdd gnd cell_6t
Xbit_r68_c194 bl_194 br_194 wl_68 vdd gnd cell_6t
Xbit_r69_c194 bl_194 br_194 wl_69 vdd gnd cell_6t
Xbit_r70_c194 bl_194 br_194 wl_70 vdd gnd cell_6t
Xbit_r71_c194 bl_194 br_194 wl_71 vdd gnd cell_6t
Xbit_r72_c194 bl_194 br_194 wl_72 vdd gnd cell_6t
Xbit_r73_c194 bl_194 br_194 wl_73 vdd gnd cell_6t
Xbit_r74_c194 bl_194 br_194 wl_74 vdd gnd cell_6t
Xbit_r75_c194 bl_194 br_194 wl_75 vdd gnd cell_6t
Xbit_r76_c194 bl_194 br_194 wl_76 vdd gnd cell_6t
Xbit_r77_c194 bl_194 br_194 wl_77 vdd gnd cell_6t
Xbit_r78_c194 bl_194 br_194 wl_78 vdd gnd cell_6t
Xbit_r79_c194 bl_194 br_194 wl_79 vdd gnd cell_6t
Xbit_r80_c194 bl_194 br_194 wl_80 vdd gnd cell_6t
Xbit_r81_c194 bl_194 br_194 wl_81 vdd gnd cell_6t
Xbit_r82_c194 bl_194 br_194 wl_82 vdd gnd cell_6t
Xbit_r83_c194 bl_194 br_194 wl_83 vdd gnd cell_6t
Xbit_r84_c194 bl_194 br_194 wl_84 vdd gnd cell_6t
Xbit_r85_c194 bl_194 br_194 wl_85 vdd gnd cell_6t
Xbit_r86_c194 bl_194 br_194 wl_86 vdd gnd cell_6t
Xbit_r87_c194 bl_194 br_194 wl_87 vdd gnd cell_6t
Xbit_r88_c194 bl_194 br_194 wl_88 vdd gnd cell_6t
Xbit_r89_c194 bl_194 br_194 wl_89 vdd gnd cell_6t
Xbit_r90_c194 bl_194 br_194 wl_90 vdd gnd cell_6t
Xbit_r91_c194 bl_194 br_194 wl_91 vdd gnd cell_6t
Xbit_r92_c194 bl_194 br_194 wl_92 vdd gnd cell_6t
Xbit_r93_c194 bl_194 br_194 wl_93 vdd gnd cell_6t
Xbit_r94_c194 bl_194 br_194 wl_94 vdd gnd cell_6t
Xbit_r95_c194 bl_194 br_194 wl_95 vdd gnd cell_6t
Xbit_r96_c194 bl_194 br_194 wl_96 vdd gnd cell_6t
Xbit_r97_c194 bl_194 br_194 wl_97 vdd gnd cell_6t
Xbit_r98_c194 bl_194 br_194 wl_98 vdd gnd cell_6t
Xbit_r99_c194 bl_194 br_194 wl_99 vdd gnd cell_6t
Xbit_r100_c194 bl_194 br_194 wl_100 vdd gnd cell_6t
Xbit_r101_c194 bl_194 br_194 wl_101 vdd gnd cell_6t
Xbit_r102_c194 bl_194 br_194 wl_102 vdd gnd cell_6t
Xbit_r103_c194 bl_194 br_194 wl_103 vdd gnd cell_6t
Xbit_r104_c194 bl_194 br_194 wl_104 vdd gnd cell_6t
Xbit_r105_c194 bl_194 br_194 wl_105 vdd gnd cell_6t
Xbit_r106_c194 bl_194 br_194 wl_106 vdd gnd cell_6t
Xbit_r107_c194 bl_194 br_194 wl_107 vdd gnd cell_6t
Xbit_r108_c194 bl_194 br_194 wl_108 vdd gnd cell_6t
Xbit_r109_c194 bl_194 br_194 wl_109 vdd gnd cell_6t
Xbit_r110_c194 bl_194 br_194 wl_110 vdd gnd cell_6t
Xbit_r111_c194 bl_194 br_194 wl_111 vdd gnd cell_6t
Xbit_r112_c194 bl_194 br_194 wl_112 vdd gnd cell_6t
Xbit_r113_c194 bl_194 br_194 wl_113 vdd gnd cell_6t
Xbit_r114_c194 bl_194 br_194 wl_114 vdd gnd cell_6t
Xbit_r115_c194 bl_194 br_194 wl_115 vdd gnd cell_6t
Xbit_r116_c194 bl_194 br_194 wl_116 vdd gnd cell_6t
Xbit_r117_c194 bl_194 br_194 wl_117 vdd gnd cell_6t
Xbit_r118_c194 bl_194 br_194 wl_118 vdd gnd cell_6t
Xbit_r119_c194 bl_194 br_194 wl_119 vdd gnd cell_6t
Xbit_r120_c194 bl_194 br_194 wl_120 vdd gnd cell_6t
Xbit_r121_c194 bl_194 br_194 wl_121 vdd gnd cell_6t
Xbit_r122_c194 bl_194 br_194 wl_122 vdd gnd cell_6t
Xbit_r123_c194 bl_194 br_194 wl_123 vdd gnd cell_6t
Xbit_r124_c194 bl_194 br_194 wl_124 vdd gnd cell_6t
Xbit_r125_c194 bl_194 br_194 wl_125 vdd gnd cell_6t
Xbit_r126_c194 bl_194 br_194 wl_126 vdd gnd cell_6t
Xbit_r127_c194 bl_194 br_194 wl_127 vdd gnd cell_6t
Xbit_r128_c194 bl_194 br_194 wl_128 vdd gnd cell_6t
Xbit_r129_c194 bl_194 br_194 wl_129 vdd gnd cell_6t
Xbit_r130_c194 bl_194 br_194 wl_130 vdd gnd cell_6t
Xbit_r131_c194 bl_194 br_194 wl_131 vdd gnd cell_6t
Xbit_r132_c194 bl_194 br_194 wl_132 vdd gnd cell_6t
Xbit_r133_c194 bl_194 br_194 wl_133 vdd gnd cell_6t
Xbit_r134_c194 bl_194 br_194 wl_134 vdd gnd cell_6t
Xbit_r135_c194 bl_194 br_194 wl_135 vdd gnd cell_6t
Xbit_r136_c194 bl_194 br_194 wl_136 vdd gnd cell_6t
Xbit_r137_c194 bl_194 br_194 wl_137 vdd gnd cell_6t
Xbit_r138_c194 bl_194 br_194 wl_138 vdd gnd cell_6t
Xbit_r139_c194 bl_194 br_194 wl_139 vdd gnd cell_6t
Xbit_r140_c194 bl_194 br_194 wl_140 vdd gnd cell_6t
Xbit_r141_c194 bl_194 br_194 wl_141 vdd gnd cell_6t
Xbit_r142_c194 bl_194 br_194 wl_142 vdd gnd cell_6t
Xbit_r143_c194 bl_194 br_194 wl_143 vdd gnd cell_6t
Xbit_r144_c194 bl_194 br_194 wl_144 vdd gnd cell_6t
Xbit_r145_c194 bl_194 br_194 wl_145 vdd gnd cell_6t
Xbit_r146_c194 bl_194 br_194 wl_146 vdd gnd cell_6t
Xbit_r147_c194 bl_194 br_194 wl_147 vdd gnd cell_6t
Xbit_r148_c194 bl_194 br_194 wl_148 vdd gnd cell_6t
Xbit_r149_c194 bl_194 br_194 wl_149 vdd gnd cell_6t
Xbit_r150_c194 bl_194 br_194 wl_150 vdd gnd cell_6t
Xbit_r151_c194 bl_194 br_194 wl_151 vdd gnd cell_6t
Xbit_r152_c194 bl_194 br_194 wl_152 vdd gnd cell_6t
Xbit_r153_c194 bl_194 br_194 wl_153 vdd gnd cell_6t
Xbit_r154_c194 bl_194 br_194 wl_154 vdd gnd cell_6t
Xbit_r155_c194 bl_194 br_194 wl_155 vdd gnd cell_6t
Xbit_r156_c194 bl_194 br_194 wl_156 vdd gnd cell_6t
Xbit_r157_c194 bl_194 br_194 wl_157 vdd gnd cell_6t
Xbit_r158_c194 bl_194 br_194 wl_158 vdd gnd cell_6t
Xbit_r159_c194 bl_194 br_194 wl_159 vdd gnd cell_6t
Xbit_r160_c194 bl_194 br_194 wl_160 vdd gnd cell_6t
Xbit_r161_c194 bl_194 br_194 wl_161 vdd gnd cell_6t
Xbit_r162_c194 bl_194 br_194 wl_162 vdd gnd cell_6t
Xbit_r163_c194 bl_194 br_194 wl_163 vdd gnd cell_6t
Xbit_r164_c194 bl_194 br_194 wl_164 vdd gnd cell_6t
Xbit_r165_c194 bl_194 br_194 wl_165 vdd gnd cell_6t
Xbit_r166_c194 bl_194 br_194 wl_166 vdd gnd cell_6t
Xbit_r167_c194 bl_194 br_194 wl_167 vdd gnd cell_6t
Xbit_r168_c194 bl_194 br_194 wl_168 vdd gnd cell_6t
Xbit_r169_c194 bl_194 br_194 wl_169 vdd gnd cell_6t
Xbit_r170_c194 bl_194 br_194 wl_170 vdd gnd cell_6t
Xbit_r171_c194 bl_194 br_194 wl_171 vdd gnd cell_6t
Xbit_r172_c194 bl_194 br_194 wl_172 vdd gnd cell_6t
Xbit_r173_c194 bl_194 br_194 wl_173 vdd gnd cell_6t
Xbit_r174_c194 bl_194 br_194 wl_174 vdd gnd cell_6t
Xbit_r175_c194 bl_194 br_194 wl_175 vdd gnd cell_6t
Xbit_r176_c194 bl_194 br_194 wl_176 vdd gnd cell_6t
Xbit_r177_c194 bl_194 br_194 wl_177 vdd gnd cell_6t
Xbit_r178_c194 bl_194 br_194 wl_178 vdd gnd cell_6t
Xbit_r179_c194 bl_194 br_194 wl_179 vdd gnd cell_6t
Xbit_r180_c194 bl_194 br_194 wl_180 vdd gnd cell_6t
Xbit_r181_c194 bl_194 br_194 wl_181 vdd gnd cell_6t
Xbit_r182_c194 bl_194 br_194 wl_182 vdd gnd cell_6t
Xbit_r183_c194 bl_194 br_194 wl_183 vdd gnd cell_6t
Xbit_r184_c194 bl_194 br_194 wl_184 vdd gnd cell_6t
Xbit_r185_c194 bl_194 br_194 wl_185 vdd gnd cell_6t
Xbit_r186_c194 bl_194 br_194 wl_186 vdd gnd cell_6t
Xbit_r187_c194 bl_194 br_194 wl_187 vdd gnd cell_6t
Xbit_r188_c194 bl_194 br_194 wl_188 vdd gnd cell_6t
Xbit_r189_c194 bl_194 br_194 wl_189 vdd gnd cell_6t
Xbit_r190_c194 bl_194 br_194 wl_190 vdd gnd cell_6t
Xbit_r191_c194 bl_194 br_194 wl_191 vdd gnd cell_6t
Xbit_r192_c194 bl_194 br_194 wl_192 vdd gnd cell_6t
Xbit_r193_c194 bl_194 br_194 wl_193 vdd gnd cell_6t
Xbit_r194_c194 bl_194 br_194 wl_194 vdd gnd cell_6t
Xbit_r195_c194 bl_194 br_194 wl_195 vdd gnd cell_6t
Xbit_r196_c194 bl_194 br_194 wl_196 vdd gnd cell_6t
Xbit_r197_c194 bl_194 br_194 wl_197 vdd gnd cell_6t
Xbit_r198_c194 bl_194 br_194 wl_198 vdd gnd cell_6t
Xbit_r199_c194 bl_194 br_194 wl_199 vdd gnd cell_6t
Xbit_r200_c194 bl_194 br_194 wl_200 vdd gnd cell_6t
Xbit_r201_c194 bl_194 br_194 wl_201 vdd gnd cell_6t
Xbit_r202_c194 bl_194 br_194 wl_202 vdd gnd cell_6t
Xbit_r203_c194 bl_194 br_194 wl_203 vdd gnd cell_6t
Xbit_r204_c194 bl_194 br_194 wl_204 vdd gnd cell_6t
Xbit_r205_c194 bl_194 br_194 wl_205 vdd gnd cell_6t
Xbit_r206_c194 bl_194 br_194 wl_206 vdd gnd cell_6t
Xbit_r207_c194 bl_194 br_194 wl_207 vdd gnd cell_6t
Xbit_r208_c194 bl_194 br_194 wl_208 vdd gnd cell_6t
Xbit_r209_c194 bl_194 br_194 wl_209 vdd gnd cell_6t
Xbit_r210_c194 bl_194 br_194 wl_210 vdd gnd cell_6t
Xbit_r211_c194 bl_194 br_194 wl_211 vdd gnd cell_6t
Xbit_r212_c194 bl_194 br_194 wl_212 vdd gnd cell_6t
Xbit_r213_c194 bl_194 br_194 wl_213 vdd gnd cell_6t
Xbit_r214_c194 bl_194 br_194 wl_214 vdd gnd cell_6t
Xbit_r215_c194 bl_194 br_194 wl_215 vdd gnd cell_6t
Xbit_r216_c194 bl_194 br_194 wl_216 vdd gnd cell_6t
Xbit_r217_c194 bl_194 br_194 wl_217 vdd gnd cell_6t
Xbit_r218_c194 bl_194 br_194 wl_218 vdd gnd cell_6t
Xbit_r219_c194 bl_194 br_194 wl_219 vdd gnd cell_6t
Xbit_r220_c194 bl_194 br_194 wl_220 vdd gnd cell_6t
Xbit_r221_c194 bl_194 br_194 wl_221 vdd gnd cell_6t
Xbit_r222_c194 bl_194 br_194 wl_222 vdd gnd cell_6t
Xbit_r223_c194 bl_194 br_194 wl_223 vdd gnd cell_6t
Xbit_r224_c194 bl_194 br_194 wl_224 vdd gnd cell_6t
Xbit_r225_c194 bl_194 br_194 wl_225 vdd gnd cell_6t
Xbit_r226_c194 bl_194 br_194 wl_226 vdd gnd cell_6t
Xbit_r227_c194 bl_194 br_194 wl_227 vdd gnd cell_6t
Xbit_r228_c194 bl_194 br_194 wl_228 vdd gnd cell_6t
Xbit_r229_c194 bl_194 br_194 wl_229 vdd gnd cell_6t
Xbit_r230_c194 bl_194 br_194 wl_230 vdd gnd cell_6t
Xbit_r231_c194 bl_194 br_194 wl_231 vdd gnd cell_6t
Xbit_r232_c194 bl_194 br_194 wl_232 vdd gnd cell_6t
Xbit_r233_c194 bl_194 br_194 wl_233 vdd gnd cell_6t
Xbit_r234_c194 bl_194 br_194 wl_234 vdd gnd cell_6t
Xbit_r235_c194 bl_194 br_194 wl_235 vdd gnd cell_6t
Xbit_r236_c194 bl_194 br_194 wl_236 vdd gnd cell_6t
Xbit_r237_c194 bl_194 br_194 wl_237 vdd gnd cell_6t
Xbit_r238_c194 bl_194 br_194 wl_238 vdd gnd cell_6t
Xbit_r239_c194 bl_194 br_194 wl_239 vdd gnd cell_6t
Xbit_r240_c194 bl_194 br_194 wl_240 vdd gnd cell_6t
Xbit_r241_c194 bl_194 br_194 wl_241 vdd gnd cell_6t
Xbit_r242_c194 bl_194 br_194 wl_242 vdd gnd cell_6t
Xbit_r243_c194 bl_194 br_194 wl_243 vdd gnd cell_6t
Xbit_r244_c194 bl_194 br_194 wl_244 vdd gnd cell_6t
Xbit_r245_c194 bl_194 br_194 wl_245 vdd gnd cell_6t
Xbit_r246_c194 bl_194 br_194 wl_246 vdd gnd cell_6t
Xbit_r247_c194 bl_194 br_194 wl_247 vdd gnd cell_6t
Xbit_r248_c194 bl_194 br_194 wl_248 vdd gnd cell_6t
Xbit_r249_c194 bl_194 br_194 wl_249 vdd gnd cell_6t
Xbit_r250_c194 bl_194 br_194 wl_250 vdd gnd cell_6t
Xbit_r251_c194 bl_194 br_194 wl_251 vdd gnd cell_6t
Xbit_r252_c194 bl_194 br_194 wl_252 vdd gnd cell_6t
Xbit_r253_c194 bl_194 br_194 wl_253 vdd gnd cell_6t
Xbit_r254_c194 bl_194 br_194 wl_254 vdd gnd cell_6t
Xbit_r255_c194 bl_194 br_194 wl_255 vdd gnd cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd cell_6t
Xbit_r1_c195 bl_195 br_195 wl_1 vdd gnd cell_6t
Xbit_r2_c195 bl_195 br_195 wl_2 vdd gnd cell_6t
Xbit_r3_c195 bl_195 br_195 wl_3 vdd gnd cell_6t
Xbit_r4_c195 bl_195 br_195 wl_4 vdd gnd cell_6t
Xbit_r5_c195 bl_195 br_195 wl_5 vdd gnd cell_6t
Xbit_r6_c195 bl_195 br_195 wl_6 vdd gnd cell_6t
Xbit_r7_c195 bl_195 br_195 wl_7 vdd gnd cell_6t
Xbit_r8_c195 bl_195 br_195 wl_8 vdd gnd cell_6t
Xbit_r9_c195 bl_195 br_195 wl_9 vdd gnd cell_6t
Xbit_r10_c195 bl_195 br_195 wl_10 vdd gnd cell_6t
Xbit_r11_c195 bl_195 br_195 wl_11 vdd gnd cell_6t
Xbit_r12_c195 bl_195 br_195 wl_12 vdd gnd cell_6t
Xbit_r13_c195 bl_195 br_195 wl_13 vdd gnd cell_6t
Xbit_r14_c195 bl_195 br_195 wl_14 vdd gnd cell_6t
Xbit_r15_c195 bl_195 br_195 wl_15 vdd gnd cell_6t
Xbit_r16_c195 bl_195 br_195 wl_16 vdd gnd cell_6t
Xbit_r17_c195 bl_195 br_195 wl_17 vdd gnd cell_6t
Xbit_r18_c195 bl_195 br_195 wl_18 vdd gnd cell_6t
Xbit_r19_c195 bl_195 br_195 wl_19 vdd gnd cell_6t
Xbit_r20_c195 bl_195 br_195 wl_20 vdd gnd cell_6t
Xbit_r21_c195 bl_195 br_195 wl_21 vdd gnd cell_6t
Xbit_r22_c195 bl_195 br_195 wl_22 vdd gnd cell_6t
Xbit_r23_c195 bl_195 br_195 wl_23 vdd gnd cell_6t
Xbit_r24_c195 bl_195 br_195 wl_24 vdd gnd cell_6t
Xbit_r25_c195 bl_195 br_195 wl_25 vdd gnd cell_6t
Xbit_r26_c195 bl_195 br_195 wl_26 vdd gnd cell_6t
Xbit_r27_c195 bl_195 br_195 wl_27 vdd gnd cell_6t
Xbit_r28_c195 bl_195 br_195 wl_28 vdd gnd cell_6t
Xbit_r29_c195 bl_195 br_195 wl_29 vdd gnd cell_6t
Xbit_r30_c195 bl_195 br_195 wl_30 vdd gnd cell_6t
Xbit_r31_c195 bl_195 br_195 wl_31 vdd gnd cell_6t
Xbit_r32_c195 bl_195 br_195 wl_32 vdd gnd cell_6t
Xbit_r33_c195 bl_195 br_195 wl_33 vdd gnd cell_6t
Xbit_r34_c195 bl_195 br_195 wl_34 vdd gnd cell_6t
Xbit_r35_c195 bl_195 br_195 wl_35 vdd gnd cell_6t
Xbit_r36_c195 bl_195 br_195 wl_36 vdd gnd cell_6t
Xbit_r37_c195 bl_195 br_195 wl_37 vdd gnd cell_6t
Xbit_r38_c195 bl_195 br_195 wl_38 vdd gnd cell_6t
Xbit_r39_c195 bl_195 br_195 wl_39 vdd gnd cell_6t
Xbit_r40_c195 bl_195 br_195 wl_40 vdd gnd cell_6t
Xbit_r41_c195 bl_195 br_195 wl_41 vdd gnd cell_6t
Xbit_r42_c195 bl_195 br_195 wl_42 vdd gnd cell_6t
Xbit_r43_c195 bl_195 br_195 wl_43 vdd gnd cell_6t
Xbit_r44_c195 bl_195 br_195 wl_44 vdd gnd cell_6t
Xbit_r45_c195 bl_195 br_195 wl_45 vdd gnd cell_6t
Xbit_r46_c195 bl_195 br_195 wl_46 vdd gnd cell_6t
Xbit_r47_c195 bl_195 br_195 wl_47 vdd gnd cell_6t
Xbit_r48_c195 bl_195 br_195 wl_48 vdd gnd cell_6t
Xbit_r49_c195 bl_195 br_195 wl_49 vdd gnd cell_6t
Xbit_r50_c195 bl_195 br_195 wl_50 vdd gnd cell_6t
Xbit_r51_c195 bl_195 br_195 wl_51 vdd gnd cell_6t
Xbit_r52_c195 bl_195 br_195 wl_52 vdd gnd cell_6t
Xbit_r53_c195 bl_195 br_195 wl_53 vdd gnd cell_6t
Xbit_r54_c195 bl_195 br_195 wl_54 vdd gnd cell_6t
Xbit_r55_c195 bl_195 br_195 wl_55 vdd gnd cell_6t
Xbit_r56_c195 bl_195 br_195 wl_56 vdd gnd cell_6t
Xbit_r57_c195 bl_195 br_195 wl_57 vdd gnd cell_6t
Xbit_r58_c195 bl_195 br_195 wl_58 vdd gnd cell_6t
Xbit_r59_c195 bl_195 br_195 wl_59 vdd gnd cell_6t
Xbit_r60_c195 bl_195 br_195 wl_60 vdd gnd cell_6t
Xbit_r61_c195 bl_195 br_195 wl_61 vdd gnd cell_6t
Xbit_r62_c195 bl_195 br_195 wl_62 vdd gnd cell_6t
Xbit_r63_c195 bl_195 br_195 wl_63 vdd gnd cell_6t
Xbit_r64_c195 bl_195 br_195 wl_64 vdd gnd cell_6t
Xbit_r65_c195 bl_195 br_195 wl_65 vdd gnd cell_6t
Xbit_r66_c195 bl_195 br_195 wl_66 vdd gnd cell_6t
Xbit_r67_c195 bl_195 br_195 wl_67 vdd gnd cell_6t
Xbit_r68_c195 bl_195 br_195 wl_68 vdd gnd cell_6t
Xbit_r69_c195 bl_195 br_195 wl_69 vdd gnd cell_6t
Xbit_r70_c195 bl_195 br_195 wl_70 vdd gnd cell_6t
Xbit_r71_c195 bl_195 br_195 wl_71 vdd gnd cell_6t
Xbit_r72_c195 bl_195 br_195 wl_72 vdd gnd cell_6t
Xbit_r73_c195 bl_195 br_195 wl_73 vdd gnd cell_6t
Xbit_r74_c195 bl_195 br_195 wl_74 vdd gnd cell_6t
Xbit_r75_c195 bl_195 br_195 wl_75 vdd gnd cell_6t
Xbit_r76_c195 bl_195 br_195 wl_76 vdd gnd cell_6t
Xbit_r77_c195 bl_195 br_195 wl_77 vdd gnd cell_6t
Xbit_r78_c195 bl_195 br_195 wl_78 vdd gnd cell_6t
Xbit_r79_c195 bl_195 br_195 wl_79 vdd gnd cell_6t
Xbit_r80_c195 bl_195 br_195 wl_80 vdd gnd cell_6t
Xbit_r81_c195 bl_195 br_195 wl_81 vdd gnd cell_6t
Xbit_r82_c195 bl_195 br_195 wl_82 vdd gnd cell_6t
Xbit_r83_c195 bl_195 br_195 wl_83 vdd gnd cell_6t
Xbit_r84_c195 bl_195 br_195 wl_84 vdd gnd cell_6t
Xbit_r85_c195 bl_195 br_195 wl_85 vdd gnd cell_6t
Xbit_r86_c195 bl_195 br_195 wl_86 vdd gnd cell_6t
Xbit_r87_c195 bl_195 br_195 wl_87 vdd gnd cell_6t
Xbit_r88_c195 bl_195 br_195 wl_88 vdd gnd cell_6t
Xbit_r89_c195 bl_195 br_195 wl_89 vdd gnd cell_6t
Xbit_r90_c195 bl_195 br_195 wl_90 vdd gnd cell_6t
Xbit_r91_c195 bl_195 br_195 wl_91 vdd gnd cell_6t
Xbit_r92_c195 bl_195 br_195 wl_92 vdd gnd cell_6t
Xbit_r93_c195 bl_195 br_195 wl_93 vdd gnd cell_6t
Xbit_r94_c195 bl_195 br_195 wl_94 vdd gnd cell_6t
Xbit_r95_c195 bl_195 br_195 wl_95 vdd gnd cell_6t
Xbit_r96_c195 bl_195 br_195 wl_96 vdd gnd cell_6t
Xbit_r97_c195 bl_195 br_195 wl_97 vdd gnd cell_6t
Xbit_r98_c195 bl_195 br_195 wl_98 vdd gnd cell_6t
Xbit_r99_c195 bl_195 br_195 wl_99 vdd gnd cell_6t
Xbit_r100_c195 bl_195 br_195 wl_100 vdd gnd cell_6t
Xbit_r101_c195 bl_195 br_195 wl_101 vdd gnd cell_6t
Xbit_r102_c195 bl_195 br_195 wl_102 vdd gnd cell_6t
Xbit_r103_c195 bl_195 br_195 wl_103 vdd gnd cell_6t
Xbit_r104_c195 bl_195 br_195 wl_104 vdd gnd cell_6t
Xbit_r105_c195 bl_195 br_195 wl_105 vdd gnd cell_6t
Xbit_r106_c195 bl_195 br_195 wl_106 vdd gnd cell_6t
Xbit_r107_c195 bl_195 br_195 wl_107 vdd gnd cell_6t
Xbit_r108_c195 bl_195 br_195 wl_108 vdd gnd cell_6t
Xbit_r109_c195 bl_195 br_195 wl_109 vdd gnd cell_6t
Xbit_r110_c195 bl_195 br_195 wl_110 vdd gnd cell_6t
Xbit_r111_c195 bl_195 br_195 wl_111 vdd gnd cell_6t
Xbit_r112_c195 bl_195 br_195 wl_112 vdd gnd cell_6t
Xbit_r113_c195 bl_195 br_195 wl_113 vdd gnd cell_6t
Xbit_r114_c195 bl_195 br_195 wl_114 vdd gnd cell_6t
Xbit_r115_c195 bl_195 br_195 wl_115 vdd gnd cell_6t
Xbit_r116_c195 bl_195 br_195 wl_116 vdd gnd cell_6t
Xbit_r117_c195 bl_195 br_195 wl_117 vdd gnd cell_6t
Xbit_r118_c195 bl_195 br_195 wl_118 vdd gnd cell_6t
Xbit_r119_c195 bl_195 br_195 wl_119 vdd gnd cell_6t
Xbit_r120_c195 bl_195 br_195 wl_120 vdd gnd cell_6t
Xbit_r121_c195 bl_195 br_195 wl_121 vdd gnd cell_6t
Xbit_r122_c195 bl_195 br_195 wl_122 vdd gnd cell_6t
Xbit_r123_c195 bl_195 br_195 wl_123 vdd gnd cell_6t
Xbit_r124_c195 bl_195 br_195 wl_124 vdd gnd cell_6t
Xbit_r125_c195 bl_195 br_195 wl_125 vdd gnd cell_6t
Xbit_r126_c195 bl_195 br_195 wl_126 vdd gnd cell_6t
Xbit_r127_c195 bl_195 br_195 wl_127 vdd gnd cell_6t
Xbit_r128_c195 bl_195 br_195 wl_128 vdd gnd cell_6t
Xbit_r129_c195 bl_195 br_195 wl_129 vdd gnd cell_6t
Xbit_r130_c195 bl_195 br_195 wl_130 vdd gnd cell_6t
Xbit_r131_c195 bl_195 br_195 wl_131 vdd gnd cell_6t
Xbit_r132_c195 bl_195 br_195 wl_132 vdd gnd cell_6t
Xbit_r133_c195 bl_195 br_195 wl_133 vdd gnd cell_6t
Xbit_r134_c195 bl_195 br_195 wl_134 vdd gnd cell_6t
Xbit_r135_c195 bl_195 br_195 wl_135 vdd gnd cell_6t
Xbit_r136_c195 bl_195 br_195 wl_136 vdd gnd cell_6t
Xbit_r137_c195 bl_195 br_195 wl_137 vdd gnd cell_6t
Xbit_r138_c195 bl_195 br_195 wl_138 vdd gnd cell_6t
Xbit_r139_c195 bl_195 br_195 wl_139 vdd gnd cell_6t
Xbit_r140_c195 bl_195 br_195 wl_140 vdd gnd cell_6t
Xbit_r141_c195 bl_195 br_195 wl_141 vdd gnd cell_6t
Xbit_r142_c195 bl_195 br_195 wl_142 vdd gnd cell_6t
Xbit_r143_c195 bl_195 br_195 wl_143 vdd gnd cell_6t
Xbit_r144_c195 bl_195 br_195 wl_144 vdd gnd cell_6t
Xbit_r145_c195 bl_195 br_195 wl_145 vdd gnd cell_6t
Xbit_r146_c195 bl_195 br_195 wl_146 vdd gnd cell_6t
Xbit_r147_c195 bl_195 br_195 wl_147 vdd gnd cell_6t
Xbit_r148_c195 bl_195 br_195 wl_148 vdd gnd cell_6t
Xbit_r149_c195 bl_195 br_195 wl_149 vdd gnd cell_6t
Xbit_r150_c195 bl_195 br_195 wl_150 vdd gnd cell_6t
Xbit_r151_c195 bl_195 br_195 wl_151 vdd gnd cell_6t
Xbit_r152_c195 bl_195 br_195 wl_152 vdd gnd cell_6t
Xbit_r153_c195 bl_195 br_195 wl_153 vdd gnd cell_6t
Xbit_r154_c195 bl_195 br_195 wl_154 vdd gnd cell_6t
Xbit_r155_c195 bl_195 br_195 wl_155 vdd gnd cell_6t
Xbit_r156_c195 bl_195 br_195 wl_156 vdd gnd cell_6t
Xbit_r157_c195 bl_195 br_195 wl_157 vdd gnd cell_6t
Xbit_r158_c195 bl_195 br_195 wl_158 vdd gnd cell_6t
Xbit_r159_c195 bl_195 br_195 wl_159 vdd gnd cell_6t
Xbit_r160_c195 bl_195 br_195 wl_160 vdd gnd cell_6t
Xbit_r161_c195 bl_195 br_195 wl_161 vdd gnd cell_6t
Xbit_r162_c195 bl_195 br_195 wl_162 vdd gnd cell_6t
Xbit_r163_c195 bl_195 br_195 wl_163 vdd gnd cell_6t
Xbit_r164_c195 bl_195 br_195 wl_164 vdd gnd cell_6t
Xbit_r165_c195 bl_195 br_195 wl_165 vdd gnd cell_6t
Xbit_r166_c195 bl_195 br_195 wl_166 vdd gnd cell_6t
Xbit_r167_c195 bl_195 br_195 wl_167 vdd gnd cell_6t
Xbit_r168_c195 bl_195 br_195 wl_168 vdd gnd cell_6t
Xbit_r169_c195 bl_195 br_195 wl_169 vdd gnd cell_6t
Xbit_r170_c195 bl_195 br_195 wl_170 vdd gnd cell_6t
Xbit_r171_c195 bl_195 br_195 wl_171 vdd gnd cell_6t
Xbit_r172_c195 bl_195 br_195 wl_172 vdd gnd cell_6t
Xbit_r173_c195 bl_195 br_195 wl_173 vdd gnd cell_6t
Xbit_r174_c195 bl_195 br_195 wl_174 vdd gnd cell_6t
Xbit_r175_c195 bl_195 br_195 wl_175 vdd gnd cell_6t
Xbit_r176_c195 bl_195 br_195 wl_176 vdd gnd cell_6t
Xbit_r177_c195 bl_195 br_195 wl_177 vdd gnd cell_6t
Xbit_r178_c195 bl_195 br_195 wl_178 vdd gnd cell_6t
Xbit_r179_c195 bl_195 br_195 wl_179 vdd gnd cell_6t
Xbit_r180_c195 bl_195 br_195 wl_180 vdd gnd cell_6t
Xbit_r181_c195 bl_195 br_195 wl_181 vdd gnd cell_6t
Xbit_r182_c195 bl_195 br_195 wl_182 vdd gnd cell_6t
Xbit_r183_c195 bl_195 br_195 wl_183 vdd gnd cell_6t
Xbit_r184_c195 bl_195 br_195 wl_184 vdd gnd cell_6t
Xbit_r185_c195 bl_195 br_195 wl_185 vdd gnd cell_6t
Xbit_r186_c195 bl_195 br_195 wl_186 vdd gnd cell_6t
Xbit_r187_c195 bl_195 br_195 wl_187 vdd gnd cell_6t
Xbit_r188_c195 bl_195 br_195 wl_188 vdd gnd cell_6t
Xbit_r189_c195 bl_195 br_195 wl_189 vdd gnd cell_6t
Xbit_r190_c195 bl_195 br_195 wl_190 vdd gnd cell_6t
Xbit_r191_c195 bl_195 br_195 wl_191 vdd gnd cell_6t
Xbit_r192_c195 bl_195 br_195 wl_192 vdd gnd cell_6t
Xbit_r193_c195 bl_195 br_195 wl_193 vdd gnd cell_6t
Xbit_r194_c195 bl_195 br_195 wl_194 vdd gnd cell_6t
Xbit_r195_c195 bl_195 br_195 wl_195 vdd gnd cell_6t
Xbit_r196_c195 bl_195 br_195 wl_196 vdd gnd cell_6t
Xbit_r197_c195 bl_195 br_195 wl_197 vdd gnd cell_6t
Xbit_r198_c195 bl_195 br_195 wl_198 vdd gnd cell_6t
Xbit_r199_c195 bl_195 br_195 wl_199 vdd gnd cell_6t
Xbit_r200_c195 bl_195 br_195 wl_200 vdd gnd cell_6t
Xbit_r201_c195 bl_195 br_195 wl_201 vdd gnd cell_6t
Xbit_r202_c195 bl_195 br_195 wl_202 vdd gnd cell_6t
Xbit_r203_c195 bl_195 br_195 wl_203 vdd gnd cell_6t
Xbit_r204_c195 bl_195 br_195 wl_204 vdd gnd cell_6t
Xbit_r205_c195 bl_195 br_195 wl_205 vdd gnd cell_6t
Xbit_r206_c195 bl_195 br_195 wl_206 vdd gnd cell_6t
Xbit_r207_c195 bl_195 br_195 wl_207 vdd gnd cell_6t
Xbit_r208_c195 bl_195 br_195 wl_208 vdd gnd cell_6t
Xbit_r209_c195 bl_195 br_195 wl_209 vdd gnd cell_6t
Xbit_r210_c195 bl_195 br_195 wl_210 vdd gnd cell_6t
Xbit_r211_c195 bl_195 br_195 wl_211 vdd gnd cell_6t
Xbit_r212_c195 bl_195 br_195 wl_212 vdd gnd cell_6t
Xbit_r213_c195 bl_195 br_195 wl_213 vdd gnd cell_6t
Xbit_r214_c195 bl_195 br_195 wl_214 vdd gnd cell_6t
Xbit_r215_c195 bl_195 br_195 wl_215 vdd gnd cell_6t
Xbit_r216_c195 bl_195 br_195 wl_216 vdd gnd cell_6t
Xbit_r217_c195 bl_195 br_195 wl_217 vdd gnd cell_6t
Xbit_r218_c195 bl_195 br_195 wl_218 vdd gnd cell_6t
Xbit_r219_c195 bl_195 br_195 wl_219 vdd gnd cell_6t
Xbit_r220_c195 bl_195 br_195 wl_220 vdd gnd cell_6t
Xbit_r221_c195 bl_195 br_195 wl_221 vdd gnd cell_6t
Xbit_r222_c195 bl_195 br_195 wl_222 vdd gnd cell_6t
Xbit_r223_c195 bl_195 br_195 wl_223 vdd gnd cell_6t
Xbit_r224_c195 bl_195 br_195 wl_224 vdd gnd cell_6t
Xbit_r225_c195 bl_195 br_195 wl_225 vdd gnd cell_6t
Xbit_r226_c195 bl_195 br_195 wl_226 vdd gnd cell_6t
Xbit_r227_c195 bl_195 br_195 wl_227 vdd gnd cell_6t
Xbit_r228_c195 bl_195 br_195 wl_228 vdd gnd cell_6t
Xbit_r229_c195 bl_195 br_195 wl_229 vdd gnd cell_6t
Xbit_r230_c195 bl_195 br_195 wl_230 vdd gnd cell_6t
Xbit_r231_c195 bl_195 br_195 wl_231 vdd gnd cell_6t
Xbit_r232_c195 bl_195 br_195 wl_232 vdd gnd cell_6t
Xbit_r233_c195 bl_195 br_195 wl_233 vdd gnd cell_6t
Xbit_r234_c195 bl_195 br_195 wl_234 vdd gnd cell_6t
Xbit_r235_c195 bl_195 br_195 wl_235 vdd gnd cell_6t
Xbit_r236_c195 bl_195 br_195 wl_236 vdd gnd cell_6t
Xbit_r237_c195 bl_195 br_195 wl_237 vdd gnd cell_6t
Xbit_r238_c195 bl_195 br_195 wl_238 vdd gnd cell_6t
Xbit_r239_c195 bl_195 br_195 wl_239 vdd gnd cell_6t
Xbit_r240_c195 bl_195 br_195 wl_240 vdd gnd cell_6t
Xbit_r241_c195 bl_195 br_195 wl_241 vdd gnd cell_6t
Xbit_r242_c195 bl_195 br_195 wl_242 vdd gnd cell_6t
Xbit_r243_c195 bl_195 br_195 wl_243 vdd gnd cell_6t
Xbit_r244_c195 bl_195 br_195 wl_244 vdd gnd cell_6t
Xbit_r245_c195 bl_195 br_195 wl_245 vdd gnd cell_6t
Xbit_r246_c195 bl_195 br_195 wl_246 vdd gnd cell_6t
Xbit_r247_c195 bl_195 br_195 wl_247 vdd gnd cell_6t
Xbit_r248_c195 bl_195 br_195 wl_248 vdd gnd cell_6t
Xbit_r249_c195 bl_195 br_195 wl_249 vdd gnd cell_6t
Xbit_r250_c195 bl_195 br_195 wl_250 vdd gnd cell_6t
Xbit_r251_c195 bl_195 br_195 wl_251 vdd gnd cell_6t
Xbit_r252_c195 bl_195 br_195 wl_252 vdd gnd cell_6t
Xbit_r253_c195 bl_195 br_195 wl_253 vdd gnd cell_6t
Xbit_r254_c195 bl_195 br_195 wl_254 vdd gnd cell_6t
Xbit_r255_c195 bl_195 br_195 wl_255 vdd gnd cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd cell_6t
Xbit_r1_c196 bl_196 br_196 wl_1 vdd gnd cell_6t
Xbit_r2_c196 bl_196 br_196 wl_2 vdd gnd cell_6t
Xbit_r3_c196 bl_196 br_196 wl_3 vdd gnd cell_6t
Xbit_r4_c196 bl_196 br_196 wl_4 vdd gnd cell_6t
Xbit_r5_c196 bl_196 br_196 wl_5 vdd gnd cell_6t
Xbit_r6_c196 bl_196 br_196 wl_6 vdd gnd cell_6t
Xbit_r7_c196 bl_196 br_196 wl_7 vdd gnd cell_6t
Xbit_r8_c196 bl_196 br_196 wl_8 vdd gnd cell_6t
Xbit_r9_c196 bl_196 br_196 wl_9 vdd gnd cell_6t
Xbit_r10_c196 bl_196 br_196 wl_10 vdd gnd cell_6t
Xbit_r11_c196 bl_196 br_196 wl_11 vdd gnd cell_6t
Xbit_r12_c196 bl_196 br_196 wl_12 vdd gnd cell_6t
Xbit_r13_c196 bl_196 br_196 wl_13 vdd gnd cell_6t
Xbit_r14_c196 bl_196 br_196 wl_14 vdd gnd cell_6t
Xbit_r15_c196 bl_196 br_196 wl_15 vdd gnd cell_6t
Xbit_r16_c196 bl_196 br_196 wl_16 vdd gnd cell_6t
Xbit_r17_c196 bl_196 br_196 wl_17 vdd gnd cell_6t
Xbit_r18_c196 bl_196 br_196 wl_18 vdd gnd cell_6t
Xbit_r19_c196 bl_196 br_196 wl_19 vdd gnd cell_6t
Xbit_r20_c196 bl_196 br_196 wl_20 vdd gnd cell_6t
Xbit_r21_c196 bl_196 br_196 wl_21 vdd gnd cell_6t
Xbit_r22_c196 bl_196 br_196 wl_22 vdd gnd cell_6t
Xbit_r23_c196 bl_196 br_196 wl_23 vdd gnd cell_6t
Xbit_r24_c196 bl_196 br_196 wl_24 vdd gnd cell_6t
Xbit_r25_c196 bl_196 br_196 wl_25 vdd gnd cell_6t
Xbit_r26_c196 bl_196 br_196 wl_26 vdd gnd cell_6t
Xbit_r27_c196 bl_196 br_196 wl_27 vdd gnd cell_6t
Xbit_r28_c196 bl_196 br_196 wl_28 vdd gnd cell_6t
Xbit_r29_c196 bl_196 br_196 wl_29 vdd gnd cell_6t
Xbit_r30_c196 bl_196 br_196 wl_30 vdd gnd cell_6t
Xbit_r31_c196 bl_196 br_196 wl_31 vdd gnd cell_6t
Xbit_r32_c196 bl_196 br_196 wl_32 vdd gnd cell_6t
Xbit_r33_c196 bl_196 br_196 wl_33 vdd gnd cell_6t
Xbit_r34_c196 bl_196 br_196 wl_34 vdd gnd cell_6t
Xbit_r35_c196 bl_196 br_196 wl_35 vdd gnd cell_6t
Xbit_r36_c196 bl_196 br_196 wl_36 vdd gnd cell_6t
Xbit_r37_c196 bl_196 br_196 wl_37 vdd gnd cell_6t
Xbit_r38_c196 bl_196 br_196 wl_38 vdd gnd cell_6t
Xbit_r39_c196 bl_196 br_196 wl_39 vdd gnd cell_6t
Xbit_r40_c196 bl_196 br_196 wl_40 vdd gnd cell_6t
Xbit_r41_c196 bl_196 br_196 wl_41 vdd gnd cell_6t
Xbit_r42_c196 bl_196 br_196 wl_42 vdd gnd cell_6t
Xbit_r43_c196 bl_196 br_196 wl_43 vdd gnd cell_6t
Xbit_r44_c196 bl_196 br_196 wl_44 vdd gnd cell_6t
Xbit_r45_c196 bl_196 br_196 wl_45 vdd gnd cell_6t
Xbit_r46_c196 bl_196 br_196 wl_46 vdd gnd cell_6t
Xbit_r47_c196 bl_196 br_196 wl_47 vdd gnd cell_6t
Xbit_r48_c196 bl_196 br_196 wl_48 vdd gnd cell_6t
Xbit_r49_c196 bl_196 br_196 wl_49 vdd gnd cell_6t
Xbit_r50_c196 bl_196 br_196 wl_50 vdd gnd cell_6t
Xbit_r51_c196 bl_196 br_196 wl_51 vdd gnd cell_6t
Xbit_r52_c196 bl_196 br_196 wl_52 vdd gnd cell_6t
Xbit_r53_c196 bl_196 br_196 wl_53 vdd gnd cell_6t
Xbit_r54_c196 bl_196 br_196 wl_54 vdd gnd cell_6t
Xbit_r55_c196 bl_196 br_196 wl_55 vdd gnd cell_6t
Xbit_r56_c196 bl_196 br_196 wl_56 vdd gnd cell_6t
Xbit_r57_c196 bl_196 br_196 wl_57 vdd gnd cell_6t
Xbit_r58_c196 bl_196 br_196 wl_58 vdd gnd cell_6t
Xbit_r59_c196 bl_196 br_196 wl_59 vdd gnd cell_6t
Xbit_r60_c196 bl_196 br_196 wl_60 vdd gnd cell_6t
Xbit_r61_c196 bl_196 br_196 wl_61 vdd gnd cell_6t
Xbit_r62_c196 bl_196 br_196 wl_62 vdd gnd cell_6t
Xbit_r63_c196 bl_196 br_196 wl_63 vdd gnd cell_6t
Xbit_r64_c196 bl_196 br_196 wl_64 vdd gnd cell_6t
Xbit_r65_c196 bl_196 br_196 wl_65 vdd gnd cell_6t
Xbit_r66_c196 bl_196 br_196 wl_66 vdd gnd cell_6t
Xbit_r67_c196 bl_196 br_196 wl_67 vdd gnd cell_6t
Xbit_r68_c196 bl_196 br_196 wl_68 vdd gnd cell_6t
Xbit_r69_c196 bl_196 br_196 wl_69 vdd gnd cell_6t
Xbit_r70_c196 bl_196 br_196 wl_70 vdd gnd cell_6t
Xbit_r71_c196 bl_196 br_196 wl_71 vdd gnd cell_6t
Xbit_r72_c196 bl_196 br_196 wl_72 vdd gnd cell_6t
Xbit_r73_c196 bl_196 br_196 wl_73 vdd gnd cell_6t
Xbit_r74_c196 bl_196 br_196 wl_74 vdd gnd cell_6t
Xbit_r75_c196 bl_196 br_196 wl_75 vdd gnd cell_6t
Xbit_r76_c196 bl_196 br_196 wl_76 vdd gnd cell_6t
Xbit_r77_c196 bl_196 br_196 wl_77 vdd gnd cell_6t
Xbit_r78_c196 bl_196 br_196 wl_78 vdd gnd cell_6t
Xbit_r79_c196 bl_196 br_196 wl_79 vdd gnd cell_6t
Xbit_r80_c196 bl_196 br_196 wl_80 vdd gnd cell_6t
Xbit_r81_c196 bl_196 br_196 wl_81 vdd gnd cell_6t
Xbit_r82_c196 bl_196 br_196 wl_82 vdd gnd cell_6t
Xbit_r83_c196 bl_196 br_196 wl_83 vdd gnd cell_6t
Xbit_r84_c196 bl_196 br_196 wl_84 vdd gnd cell_6t
Xbit_r85_c196 bl_196 br_196 wl_85 vdd gnd cell_6t
Xbit_r86_c196 bl_196 br_196 wl_86 vdd gnd cell_6t
Xbit_r87_c196 bl_196 br_196 wl_87 vdd gnd cell_6t
Xbit_r88_c196 bl_196 br_196 wl_88 vdd gnd cell_6t
Xbit_r89_c196 bl_196 br_196 wl_89 vdd gnd cell_6t
Xbit_r90_c196 bl_196 br_196 wl_90 vdd gnd cell_6t
Xbit_r91_c196 bl_196 br_196 wl_91 vdd gnd cell_6t
Xbit_r92_c196 bl_196 br_196 wl_92 vdd gnd cell_6t
Xbit_r93_c196 bl_196 br_196 wl_93 vdd gnd cell_6t
Xbit_r94_c196 bl_196 br_196 wl_94 vdd gnd cell_6t
Xbit_r95_c196 bl_196 br_196 wl_95 vdd gnd cell_6t
Xbit_r96_c196 bl_196 br_196 wl_96 vdd gnd cell_6t
Xbit_r97_c196 bl_196 br_196 wl_97 vdd gnd cell_6t
Xbit_r98_c196 bl_196 br_196 wl_98 vdd gnd cell_6t
Xbit_r99_c196 bl_196 br_196 wl_99 vdd gnd cell_6t
Xbit_r100_c196 bl_196 br_196 wl_100 vdd gnd cell_6t
Xbit_r101_c196 bl_196 br_196 wl_101 vdd gnd cell_6t
Xbit_r102_c196 bl_196 br_196 wl_102 vdd gnd cell_6t
Xbit_r103_c196 bl_196 br_196 wl_103 vdd gnd cell_6t
Xbit_r104_c196 bl_196 br_196 wl_104 vdd gnd cell_6t
Xbit_r105_c196 bl_196 br_196 wl_105 vdd gnd cell_6t
Xbit_r106_c196 bl_196 br_196 wl_106 vdd gnd cell_6t
Xbit_r107_c196 bl_196 br_196 wl_107 vdd gnd cell_6t
Xbit_r108_c196 bl_196 br_196 wl_108 vdd gnd cell_6t
Xbit_r109_c196 bl_196 br_196 wl_109 vdd gnd cell_6t
Xbit_r110_c196 bl_196 br_196 wl_110 vdd gnd cell_6t
Xbit_r111_c196 bl_196 br_196 wl_111 vdd gnd cell_6t
Xbit_r112_c196 bl_196 br_196 wl_112 vdd gnd cell_6t
Xbit_r113_c196 bl_196 br_196 wl_113 vdd gnd cell_6t
Xbit_r114_c196 bl_196 br_196 wl_114 vdd gnd cell_6t
Xbit_r115_c196 bl_196 br_196 wl_115 vdd gnd cell_6t
Xbit_r116_c196 bl_196 br_196 wl_116 vdd gnd cell_6t
Xbit_r117_c196 bl_196 br_196 wl_117 vdd gnd cell_6t
Xbit_r118_c196 bl_196 br_196 wl_118 vdd gnd cell_6t
Xbit_r119_c196 bl_196 br_196 wl_119 vdd gnd cell_6t
Xbit_r120_c196 bl_196 br_196 wl_120 vdd gnd cell_6t
Xbit_r121_c196 bl_196 br_196 wl_121 vdd gnd cell_6t
Xbit_r122_c196 bl_196 br_196 wl_122 vdd gnd cell_6t
Xbit_r123_c196 bl_196 br_196 wl_123 vdd gnd cell_6t
Xbit_r124_c196 bl_196 br_196 wl_124 vdd gnd cell_6t
Xbit_r125_c196 bl_196 br_196 wl_125 vdd gnd cell_6t
Xbit_r126_c196 bl_196 br_196 wl_126 vdd gnd cell_6t
Xbit_r127_c196 bl_196 br_196 wl_127 vdd gnd cell_6t
Xbit_r128_c196 bl_196 br_196 wl_128 vdd gnd cell_6t
Xbit_r129_c196 bl_196 br_196 wl_129 vdd gnd cell_6t
Xbit_r130_c196 bl_196 br_196 wl_130 vdd gnd cell_6t
Xbit_r131_c196 bl_196 br_196 wl_131 vdd gnd cell_6t
Xbit_r132_c196 bl_196 br_196 wl_132 vdd gnd cell_6t
Xbit_r133_c196 bl_196 br_196 wl_133 vdd gnd cell_6t
Xbit_r134_c196 bl_196 br_196 wl_134 vdd gnd cell_6t
Xbit_r135_c196 bl_196 br_196 wl_135 vdd gnd cell_6t
Xbit_r136_c196 bl_196 br_196 wl_136 vdd gnd cell_6t
Xbit_r137_c196 bl_196 br_196 wl_137 vdd gnd cell_6t
Xbit_r138_c196 bl_196 br_196 wl_138 vdd gnd cell_6t
Xbit_r139_c196 bl_196 br_196 wl_139 vdd gnd cell_6t
Xbit_r140_c196 bl_196 br_196 wl_140 vdd gnd cell_6t
Xbit_r141_c196 bl_196 br_196 wl_141 vdd gnd cell_6t
Xbit_r142_c196 bl_196 br_196 wl_142 vdd gnd cell_6t
Xbit_r143_c196 bl_196 br_196 wl_143 vdd gnd cell_6t
Xbit_r144_c196 bl_196 br_196 wl_144 vdd gnd cell_6t
Xbit_r145_c196 bl_196 br_196 wl_145 vdd gnd cell_6t
Xbit_r146_c196 bl_196 br_196 wl_146 vdd gnd cell_6t
Xbit_r147_c196 bl_196 br_196 wl_147 vdd gnd cell_6t
Xbit_r148_c196 bl_196 br_196 wl_148 vdd gnd cell_6t
Xbit_r149_c196 bl_196 br_196 wl_149 vdd gnd cell_6t
Xbit_r150_c196 bl_196 br_196 wl_150 vdd gnd cell_6t
Xbit_r151_c196 bl_196 br_196 wl_151 vdd gnd cell_6t
Xbit_r152_c196 bl_196 br_196 wl_152 vdd gnd cell_6t
Xbit_r153_c196 bl_196 br_196 wl_153 vdd gnd cell_6t
Xbit_r154_c196 bl_196 br_196 wl_154 vdd gnd cell_6t
Xbit_r155_c196 bl_196 br_196 wl_155 vdd gnd cell_6t
Xbit_r156_c196 bl_196 br_196 wl_156 vdd gnd cell_6t
Xbit_r157_c196 bl_196 br_196 wl_157 vdd gnd cell_6t
Xbit_r158_c196 bl_196 br_196 wl_158 vdd gnd cell_6t
Xbit_r159_c196 bl_196 br_196 wl_159 vdd gnd cell_6t
Xbit_r160_c196 bl_196 br_196 wl_160 vdd gnd cell_6t
Xbit_r161_c196 bl_196 br_196 wl_161 vdd gnd cell_6t
Xbit_r162_c196 bl_196 br_196 wl_162 vdd gnd cell_6t
Xbit_r163_c196 bl_196 br_196 wl_163 vdd gnd cell_6t
Xbit_r164_c196 bl_196 br_196 wl_164 vdd gnd cell_6t
Xbit_r165_c196 bl_196 br_196 wl_165 vdd gnd cell_6t
Xbit_r166_c196 bl_196 br_196 wl_166 vdd gnd cell_6t
Xbit_r167_c196 bl_196 br_196 wl_167 vdd gnd cell_6t
Xbit_r168_c196 bl_196 br_196 wl_168 vdd gnd cell_6t
Xbit_r169_c196 bl_196 br_196 wl_169 vdd gnd cell_6t
Xbit_r170_c196 bl_196 br_196 wl_170 vdd gnd cell_6t
Xbit_r171_c196 bl_196 br_196 wl_171 vdd gnd cell_6t
Xbit_r172_c196 bl_196 br_196 wl_172 vdd gnd cell_6t
Xbit_r173_c196 bl_196 br_196 wl_173 vdd gnd cell_6t
Xbit_r174_c196 bl_196 br_196 wl_174 vdd gnd cell_6t
Xbit_r175_c196 bl_196 br_196 wl_175 vdd gnd cell_6t
Xbit_r176_c196 bl_196 br_196 wl_176 vdd gnd cell_6t
Xbit_r177_c196 bl_196 br_196 wl_177 vdd gnd cell_6t
Xbit_r178_c196 bl_196 br_196 wl_178 vdd gnd cell_6t
Xbit_r179_c196 bl_196 br_196 wl_179 vdd gnd cell_6t
Xbit_r180_c196 bl_196 br_196 wl_180 vdd gnd cell_6t
Xbit_r181_c196 bl_196 br_196 wl_181 vdd gnd cell_6t
Xbit_r182_c196 bl_196 br_196 wl_182 vdd gnd cell_6t
Xbit_r183_c196 bl_196 br_196 wl_183 vdd gnd cell_6t
Xbit_r184_c196 bl_196 br_196 wl_184 vdd gnd cell_6t
Xbit_r185_c196 bl_196 br_196 wl_185 vdd gnd cell_6t
Xbit_r186_c196 bl_196 br_196 wl_186 vdd gnd cell_6t
Xbit_r187_c196 bl_196 br_196 wl_187 vdd gnd cell_6t
Xbit_r188_c196 bl_196 br_196 wl_188 vdd gnd cell_6t
Xbit_r189_c196 bl_196 br_196 wl_189 vdd gnd cell_6t
Xbit_r190_c196 bl_196 br_196 wl_190 vdd gnd cell_6t
Xbit_r191_c196 bl_196 br_196 wl_191 vdd gnd cell_6t
Xbit_r192_c196 bl_196 br_196 wl_192 vdd gnd cell_6t
Xbit_r193_c196 bl_196 br_196 wl_193 vdd gnd cell_6t
Xbit_r194_c196 bl_196 br_196 wl_194 vdd gnd cell_6t
Xbit_r195_c196 bl_196 br_196 wl_195 vdd gnd cell_6t
Xbit_r196_c196 bl_196 br_196 wl_196 vdd gnd cell_6t
Xbit_r197_c196 bl_196 br_196 wl_197 vdd gnd cell_6t
Xbit_r198_c196 bl_196 br_196 wl_198 vdd gnd cell_6t
Xbit_r199_c196 bl_196 br_196 wl_199 vdd gnd cell_6t
Xbit_r200_c196 bl_196 br_196 wl_200 vdd gnd cell_6t
Xbit_r201_c196 bl_196 br_196 wl_201 vdd gnd cell_6t
Xbit_r202_c196 bl_196 br_196 wl_202 vdd gnd cell_6t
Xbit_r203_c196 bl_196 br_196 wl_203 vdd gnd cell_6t
Xbit_r204_c196 bl_196 br_196 wl_204 vdd gnd cell_6t
Xbit_r205_c196 bl_196 br_196 wl_205 vdd gnd cell_6t
Xbit_r206_c196 bl_196 br_196 wl_206 vdd gnd cell_6t
Xbit_r207_c196 bl_196 br_196 wl_207 vdd gnd cell_6t
Xbit_r208_c196 bl_196 br_196 wl_208 vdd gnd cell_6t
Xbit_r209_c196 bl_196 br_196 wl_209 vdd gnd cell_6t
Xbit_r210_c196 bl_196 br_196 wl_210 vdd gnd cell_6t
Xbit_r211_c196 bl_196 br_196 wl_211 vdd gnd cell_6t
Xbit_r212_c196 bl_196 br_196 wl_212 vdd gnd cell_6t
Xbit_r213_c196 bl_196 br_196 wl_213 vdd gnd cell_6t
Xbit_r214_c196 bl_196 br_196 wl_214 vdd gnd cell_6t
Xbit_r215_c196 bl_196 br_196 wl_215 vdd gnd cell_6t
Xbit_r216_c196 bl_196 br_196 wl_216 vdd gnd cell_6t
Xbit_r217_c196 bl_196 br_196 wl_217 vdd gnd cell_6t
Xbit_r218_c196 bl_196 br_196 wl_218 vdd gnd cell_6t
Xbit_r219_c196 bl_196 br_196 wl_219 vdd gnd cell_6t
Xbit_r220_c196 bl_196 br_196 wl_220 vdd gnd cell_6t
Xbit_r221_c196 bl_196 br_196 wl_221 vdd gnd cell_6t
Xbit_r222_c196 bl_196 br_196 wl_222 vdd gnd cell_6t
Xbit_r223_c196 bl_196 br_196 wl_223 vdd gnd cell_6t
Xbit_r224_c196 bl_196 br_196 wl_224 vdd gnd cell_6t
Xbit_r225_c196 bl_196 br_196 wl_225 vdd gnd cell_6t
Xbit_r226_c196 bl_196 br_196 wl_226 vdd gnd cell_6t
Xbit_r227_c196 bl_196 br_196 wl_227 vdd gnd cell_6t
Xbit_r228_c196 bl_196 br_196 wl_228 vdd gnd cell_6t
Xbit_r229_c196 bl_196 br_196 wl_229 vdd gnd cell_6t
Xbit_r230_c196 bl_196 br_196 wl_230 vdd gnd cell_6t
Xbit_r231_c196 bl_196 br_196 wl_231 vdd gnd cell_6t
Xbit_r232_c196 bl_196 br_196 wl_232 vdd gnd cell_6t
Xbit_r233_c196 bl_196 br_196 wl_233 vdd gnd cell_6t
Xbit_r234_c196 bl_196 br_196 wl_234 vdd gnd cell_6t
Xbit_r235_c196 bl_196 br_196 wl_235 vdd gnd cell_6t
Xbit_r236_c196 bl_196 br_196 wl_236 vdd gnd cell_6t
Xbit_r237_c196 bl_196 br_196 wl_237 vdd gnd cell_6t
Xbit_r238_c196 bl_196 br_196 wl_238 vdd gnd cell_6t
Xbit_r239_c196 bl_196 br_196 wl_239 vdd gnd cell_6t
Xbit_r240_c196 bl_196 br_196 wl_240 vdd gnd cell_6t
Xbit_r241_c196 bl_196 br_196 wl_241 vdd gnd cell_6t
Xbit_r242_c196 bl_196 br_196 wl_242 vdd gnd cell_6t
Xbit_r243_c196 bl_196 br_196 wl_243 vdd gnd cell_6t
Xbit_r244_c196 bl_196 br_196 wl_244 vdd gnd cell_6t
Xbit_r245_c196 bl_196 br_196 wl_245 vdd gnd cell_6t
Xbit_r246_c196 bl_196 br_196 wl_246 vdd gnd cell_6t
Xbit_r247_c196 bl_196 br_196 wl_247 vdd gnd cell_6t
Xbit_r248_c196 bl_196 br_196 wl_248 vdd gnd cell_6t
Xbit_r249_c196 bl_196 br_196 wl_249 vdd gnd cell_6t
Xbit_r250_c196 bl_196 br_196 wl_250 vdd gnd cell_6t
Xbit_r251_c196 bl_196 br_196 wl_251 vdd gnd cell_6t
Xbit_r252_c196 bl_196 br_196 wl_252 vdd gnd cell_6t
Xbit_r253_c196 bl_196 br_196 wl_253 vdd gnd cell_6t
Xbit_r254_c196 bl_196 br_196 wl_254 vdd gnd cell_6t
Xbit_r255_c196 bl_196 br_196 wl_255 vdd gnd cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd cell_6t
Xbit_r1_c197 bl_197 br_197 wl_1 vdd gnd cell_6t
Xbit_r2_c197 bl_197 br_197 wl_2 vdd gnd cell_6t
Xbit_r3_c197 bl_197 br_197 wl_3 vdd gnd cell_6t
Xbit_r4_c197 bl_197 br_197 wl_4 vdd gnd cell_6t
Xbit_r5_c197 bl_197 br_197 wl_5 vdd gnd cell_6t
Xbit_r6_c197 bl_197 br_197 wl_6 vdd gnd cell_6t
Xbit_r7_c197 bl_197 br_197 wl_7 vdd gnd cell_6t
Xbit_r8_c197 bl_197 br_197 wl_8 vdd gnd cell_6t
Xbit_r9_c197 bl_197 br_197 wl_9 vdd gnd cell_6t
Xbit_r10_c197 bl_197 br_197 wl_10 vdd gnd cell_6t
Xbit_r11_c197 bl_197 br_197 wl_11 vdd gnd cell_6t
Xbit_r12_c197 bl_197 br_197 wl_12 vdd gnd cell_6t
Xbit_r13_c197 bl_197 br_197 wl_13 vdd gnd cell_6t
Xbit_r14_c197 bl_197 br_197 wl_14 vdd gnd cell_6t
Xbit_r15_c197 bl_197 br_197 wl_15 vdd gnd cell_6t
Xbit_r16_c197 bl_197 br_197 wl_16 vdd gnd cell_6t
Xbit_r17_c197 bl_197 br_197 wl_17 vdd gnd cell_6t
Xbit_r18_c197 bl_197 br_197 wl_18 vdd gnd cell_6t
Xbit_r19_c197 bl_197 br_197 wl_19 vdd gnd cell_6t
Xbit_r20_c197 bl_197 br_197 wl_20 vdd gnd cell_6t
Xbit_r21_c197 bl_197 br_197 wl_21 vdd gnd cell_6t
Xbit_r22_c197 bl_197 br_197 wl_22 vdd gnd cell_6t
Xbit_r23_c197 bl_197 br_197 wl_23 vdd gnd cell_6t
Xbit_r24_c197 bl_197 br_197 wl_24 vdd gnd cell_6t
Xbit_r25_c197 bl_197 br_197 wl_25 vdd gnd cell_6t
Xbit_r26_c197 bl_197 br_197 wl_26 vdd gnd cell_6t
Xbit_r27_c197 bl_197 br_197 wl_27 vdd gnd cell_6t
Xbit_r28_c197 bl_197 br_197 wl_28 vdd gnd cell_6t
Xbit_r29_c197 bl_197 br_197 wl_29 vdd gnd cell_6t
Xbit_r30_c197 bl_197 br_197 wl_30 vdd gnd cell_6t
Xbit_r31_c197 bl_197 br_197 wl_31 vdd gnd cell_6t
Xbit_r32_c197 bl_197 br_197 wl_32 vdd gnd cell_6t
Xbit_r33_c197 bl_197 br_197 wl_33 vdd gnd cell_6t
Xbit_r34_c197 bl_197 br_197 wl_34 vdd gnd cell_6t
Xbit_r35_c197 bl_197 br_197 wl_35 vdd gnd cell_6t
Xbit_r36_c197 bl_197 br_197 wl_36 vdd gnd cell_6t
Xbit_r37_c197 bl_197 br_197 wl_37 vdd gnd cell_6t
Xbit_r38_c197 bl_197 br_197 wl_38 vdd gnd cell_6t
Xbit_r39_c197 bl_197 br_197 wl_39 vdd gnd cell_6t
Xbit_r40_c197 bl_197 br_197 wl_40 vdd gnd cell_6t
Xbit_r41_c197 bl_197 br_197 wl_41 vdd gnd cell_6t
Xbit_r42_c197 bl_197 br_197 wl_42 vdd gnd cell_6t
Xbit_r43_c197 bl_197 br_197 wl_43 vdd gnd cell_6t
Xbit_r44_c197 bl_197 br_197 wl_44 vdd gnd cell_6t
Xbit_r45_c197 bl_197 br_197 wl_45 vdd gnd cell_6t
Xbit_r46_c197 bl_197 br_197 wl_46 vdd gnd cell_6t
Xbit_r47_c197 bl_197 br_197 wl_47 vdd gnd cell_6t
Xbit_r48_c197 bl_197 br_197 wl_48 vdd gnd cell_6t
Xbit_r49_c197 bl_197 br_197 wl_49 vdd gnd cell_6t
Xbit_r50_c197 bl_197 br_197 wl_50 vdd gnd cell_6t
Xbit_r51_c197 bl_197 br_197 wl_51 vdd gnd cell_6t
Xbit_r52_c197 bl_197 br_197 wl_52 vdd gnd cell_6t
Xbit_r53_c197 bl_197 br_197 wl_53 vdd gnd cell_6t
Xbit_r54_c197 bl_197 br_197 wl_54 vdd gnd cell_6t
Xbit_r55_c197 bl_197 br_197 wl_55 vdd gnd cell_6t
Xbit_r56_c197 bl_197 br_197 wl_56 vdd gnd cell_6t
Xbit_r57_c197 bl_197 br_197 wl_57 vdd gnd cell_6t
Xbit_r58_c197 bl_197 br_197 wl_58 vdd gnd cell_6t
Xbit_r59_c197 bl_197 br_197 wl_59 vdd gnd cell_6t
Xbit_r60_c197 bl_197 br_197 wl_60 vdd gnd cell_6t
Xbit_r61_c197 bl_197 br_197 wl_61 vdd gnd cell_6t
Xbit_r62_c197 bl_197 br_197 wl_62 vdd gnd cell_6t
Xbit_r63_c197 bl_197 br_197 wl_63 vdd gnd cell_6t
Xbit_r64_c197 bl_197 br_197 wl_64 vdd gnd cell_6t
Xbit_r65_c197 bl_197 br_197 wl_65 vdd gnd cell_6t
Xbit_r66_c197 bl_197 br_197 wl_66 vdd gnd cell_6t
Xbit_r67_c197 bl_197 br_197 wl_67 vdd gnd cell_6t
Xbit_r68_c197 bl_197 br_197 wl_68 vdd gnd cell_6t
Xbit_r69_c197 bl_197 br_197 wl_69 vdd gnd cell_6t
Xbit_r70_c197 bl_197 br_197 wl_70 vdd gnd cell_6t
Xbit_r71_c197 bl_197 br_197 wl_71 vdd gnd cell_6t
Xbit_r72_c197 bl_197 br_197 wl_72 vdd gnd cell_6t
Xbit_r73_c197 bl_197 br_197 wl_73 vdd gnd cell_6t
Xbit_r74_c197 bl_197 br_197 wl_74 vdd gnd cell_6t
Xbit_r75_c197 bl_197 br_197 wl_75 vdd gnd cell_6t
Xbit_r76_c197 bl_197 br_197 wl_76 vdd gnd cell_6t
Xbit_r77_c197 bl_197 br_197 wl_77 vdd gnd cell_6t
Xbit_r78_c197 bl_197 br_197 wl_78 vdd gnd cell_6t
Xbit_r79_c197 bl_197 br_197 wl_79 vdd gnd cell_6t
Xbit_r80_c197 bl_197 br_197 wl_80 vdd gnd cell_6t
Xbit_r81_c197 bl_197 br_197 wl_81 vdd gnd cell_6t
Xbit_r82_c197 bl_197 br_197 wl_82 vdd gnd cell_6t
Xbit_r83_c197 bl_197 br_197 wl_83 vdd gnd cell_6t
Xbit_r84_c197 bl_197 br_197 wl_84 vdd gnd cell_6t
Xbit_r85_c197 bl_197 br_197 wl_85 vdd gnd cell_6t
Xbit_r86_c197 bl_197 br_197 wl_86 vdd gnd cell_6t
Xbit_r87_c197 bl_197 br_197 wl_87 vdd gnd cell_6t
Xbit_r88_c197 bl_197 br_197 wl_88 vdd gnd cell_6t
Xbit_r89_c197 bl_197 br_197 wl_89 vdd gnd cell_6t
Xbit_r90_c197 bl_197 br_197 wl_90 vdd gnd cell_6t
Xbit_r91_c197 bl_197 br_197 wl_91 vdd gnd cell_6t
Xbit_r92_c197 bl_197 br_197 wl_92 vdd gnd cell_6t
Xbit_r93_c197 bl_197 br_197 wl_93 vdd gnd cell_6t
Xbit_r94_c197 bl_197 br_197 wl_94 vdd gnd cell_6t
Xbit_r95_c197 bl_197 br_197 wl_95 vdd gnd cell_6t
Xbit_r96_c197 bl_197 br_197 wl_96 vdd gnd cell_6t
Xbit_r97_c197 bl_197 br_197 wl_97 vdd gnd cell_6t
Xbit_r98_c197 bl_197 br_197 wl_98 vdd gnd cell_6t
Xbit_r99_c197 bl_197 br_197 wl_99 vdd gnd cell_6t
Xbit_r100_c197 bl_197 br_197 wl_100 vdd gnd cell_6t
Xbit_r101_c197 bl_197 br_197 wl_101 vdd gnd cell_6t
Xbit_r102_c197 bl_197 br_197 wl_102 vdd gnd cell_6t
Xbit_r103_c197 bl_197 br_197 wl_103 vdd gnd cell_6t
Xbit_r104_c197 bl_197 br_197 wl_104 vdd gnd cell_6t
Xbit_r105_c197 bl_197 br_197 wl_105 vdd gnd cell_6t
Xbit_r106_c197 bl_197 br_197 wl_106 vdd gnd cell_6t
Xbit_r107_c197 bl_197 br_197 wl_107 vdd gnd cell_6t
Xbit_r108_c197 bl_197 br_197 wl_108 vdd gnd cell_6t
Xbit_r109_c197 bl_197 br_197 wl_109 vdd gnd cell_6t
Xbit_r110_c197 bl_197 br_197 wl_110 vdd gnd cell_6t
Xbit_r111_c197 bl_197 br_197 wl_111 vdd gnd cell_6t
Xbit_r112_c197 bl_197 br_197 wl_112 vdd gnd cell_6t
Xbit_r113_c197 bl_197 br_197 wl_113 vdd gnd cell_6t
Xbit_r114_c197 bl_197 br_197 wl_114 vdd gnd cell_6t
Xbit_r115_c197 bl_197 br_197 wl_115 vdd gnd cell_6t
Xbit_r116_c197 bl_197 br_197 wl_116 vdd gnd cell_6t
Xbit_r117_c197 bl_197 br_197 wl_117 vdd gnd cell_6t
Xbit_r118_c197 bl_197 br_197 wl_118 vdd gnd cell_6t
Xbit_r119_c197 bl_197 br_197 wl_119 vdd gnd cell_6t
Xbit_r120_c197 bl_197 br_197 wl_120 vdd gnd cell_6t
Xbit_r121_c197 bl_197 br_197 wl_121 vdd gnd cell_6t
Xbit_r122_c197 bl_197 br_197 wl_122 vdd gnd cell_6t
Xbit_r123_c197 bl_197 br_197 wl_123 vdd gnd cell_6t
Xbit_r124_c197 bl_197 br_197 wl_124 vdd gnd cell_6t
Xbit_r125_c197 bl_197 br_197 wl_125 vdd gnd cell_6t
Xbit_r126_c197 bl_197 br_197 wl_126 vdd gnd cell_6t
Xbit_r127_c197 bl_197 br_197 wl_127 vdd gnd cell_6t
Xbit_r128_c197 bl_197 br_197 wl_128 vdd gnd cell_6t
Xbit_r129_c197 bl_197 br_197 wl_129 vdd gnd cell_6t
Xbit_r130_c197 bl_197 br_197 wl_130 vdd gnd cell_6t
Xbit_r131_c197 bl_197 br_197 wl_131 vdd gnd cell_6t
Xbit_r132_c197 bl_197 br_197 wl_132 vdd gnd cell_6t
Xbit_r133_c197 bl_197 br_197 wl_133 vdd gnd cell_6t
Xbit_r134_c197 bl_197 br_197 wl_134 vdd gnd cell_6t
Xbit_r135_c197 bl_197 br_197 wl_135 vdd gnd cell_6t
Xbit_r136_c197 bl_197 br_197 wl_136 vdd gnd cell_6t
Xbit_r137_c197 bl_197 br_197 wl_137 vdd gnd cell_6t
Xbit_r138_c197 bl_197 br_197 wl_138 vdd gnd cell_6t
Xbit_r139_c197 bl_197 br_197 wl_139 vdd gnd cell_6t
Xbit_r140_c197 bl_197 br_197 wl_140 vdd gnd cell_6t
Xbit_r141_c197 bl_197 br_197 wl_141 vdd gnd cell_6t
Xbit_r142_c197 bl_197 br_197 wl_142 vdd gnd cell_6t
Xbit_r143_c197 bl_197 br_197 wl_143 vdd gnd cell_6t
Xbit_r144_c197 bl_197 br_197 wl_144 vdd gnd cell_6t
Xbit_r145_c197 bl_197 br_197 wl_145 vdd gnd cell_6t
Xbit_r146_c197 bl_197 br_197 wl_146 vdd gnd cell_6t
Xbit_r147_c197 bl_197 br_197 wl_147 vdd gnd cell_6t
Xbit_r148_c197 bl_197 br_197 wl_148 vdd gnd cell_6t
Xbit_r149_c197 bl_197 br_197 wl_149 vdd gnd cell_6t
Xbit_r150_c197 bl_197 br_197 wl_150 vdd gnd cell_6t
Xbit_r151_c197 bl_197 br_197 wl_151 vdd gnd cell_6t
Xbit_r152_c197 bl_197 br_197 wl_152 vdd gnd cell_6t
Xbit_r153_c197 bl_197 br_197 wl_153 vdd gnd cell_6t
Xbit_r154_c197 bl_197 br_197 wl_154 vdd gnd cell_6t
Xbit_r155_c197 bl_197 br_197 wl_155 vdd gnd cell_6t
Xbit_r156_c197 bl_197 br_197 wl_156 vdd gnd cell_6t
Xbit_r157_c197 bl_197 br_197 wl_157 vdd gnd cell_6t
Xbit_r158_c197 bl_197 br_197 wl_158 vdd gnd cell_6t
Xbit_r159_c197 bl_197 br_197 wl_159 vdd gnd cell_6t
Xbit_r160_c197 bl_197 br_197 wl_160 vdd gnd cell_6t
Xbit_r161_c197 bl_197 br_197 wl_161 vdd gnd cell_6t
Xbit_r162_c197 bl_197 br_197 wl_162 vdd gnd cell_6t
Xbit_r163_c197 bl_197 br_197 wl_163 vdd gnd cell_6t
Xbit_r164_c197 bl_197 br_197 wl_164 vdd gnd cell_6t
Xbit_r165_c197 bl_197 br_197 wl_165 vdd gnd cell_6t
Xbit_r166_c197 bl_197 br_197 wl_166 vdd gnd cell_6t
Xbit_r167_c197 bl_197 br_197 wl_167 vdd gnd cell_6t
Xbit_r168_c197 bl_197 br_197 wl_168 vdd gnd cell_6t
Xbit_r169_c197 bl_197 br_197 wl_169 vdd gnd cell_6t
Xbit_r170_c197 bl_197 br_197 wl_170 vdd gnd cell_6t
Xbit_r171_c197 bl_197 br_197 wl_171 vdd gnd cell_6t
Xbit_r172_c197 bl_197 br_197 wl_172 vdd gnd cell_6t
Xbit_r173_c197 bl_197 br_197 wl_173 vdd gnd cell_6t
Xbit_r174_c197 bl_197 br_197 wl_174 vdd gnd cell_6t
Xbit_r175_c197 bl_197 br_197 wl_175 vdd gnd cell_6t
Xbit_r176_c197 bl_197 br_197 wl_176 vdd gnd cell_6t
Xbit_r177_c197 bl_197 br_197 wl_177 vdd gnd cell_6t
Xbit_r178_c197 bl_197 br_197 wl_178 vdd gnd cell_6t
Xbit_r179_c197 bl_197 br_197 wl_179 vdd gnd cell_6t
Xbit_r180_c197 bl_197 br_197 wl_180 vdd gnd cell_6t
Xbit_r181_c197 bl_197 br_197 wl_181 vdd gnd cell_6t
Xbit_r182_c197 bl_197 br_197 wl_182 vdd gnd cell_6t
Xbit_r183_c197 bl_197 br_197 wl_183 vdd gnd cell_6t
Xbit_r184_c197 bl_197 br_197 wl_184 vdd gnd cell_6t
Xbit_r185_c197 bl_197 br_197 wl_185 vdd gnd cell_6t
Xbit_r186_c197 bl_197 br_197 wl_186 vdd gnd cell_6t
Xbit_r187_c197 bl_197 br_197 wl_187 vdd gnd cell_6t
Xbit_r188_c197 bl_197 br_197 wl_188 vdd gnd cell_6t
Xbit_r189_c197 bl_197 br_197 wl_189 vdd gnd cell_6t
Xbit_r190_c197 bl_197 br_197 wl_190 vdd gnd cell_6t
Xbit_r191_c197 bl_197 br_197 wl_191 vdd gnd cell_6t
Xbit_r192_c197 bl_197 br_197 wl_192 vdd gnd cell_6t
Xbit_r193_c197 bl_197 br_197 wl_193 vdd gnd cell_6t
Xbit_r194_c197 bl_197 br_197 wl_194 vdd gnd cell_6t
Xbit_r195_c197 bl_197 br_197 wl_195 vdd gnd cell_6t
Xbit_r196_c197 bl_197 br_197 wl_196 vdd gnd cell_6t
Xbit_r197_c197 bl_197 br_197 wl_197 vdd gnd cell_6t
Xbit_r198_c197 bl_197 br_197 wl_198 vdd gnd cell_6t
Xbit_r199_c197 bl_197 br_197 wl_199 vdd gnd cell_6t
Xbit_r200_c197 bl_197 br_197 wl_200 vdd gnd cell_6t
Xbit_r201_c197 bl_197 br_197 wl_201 vdd gnd cell_6t
Xbit_r202_c197 bl_197 br_197 wl_202 vdd gnd cell_6t
Xbit_r203_c197 bl_197 br_197 wl_203 vdd gnd cell_6t
Xbit_r204_c197 bl_197 br_197 wl_204 vdd gnd cell_6t
Xbit_r205_c197 bl_197 br_197 wl_205 vdd gnd cell_6t
Xbit_r206_c197 bl_197 br_197 wl_206 vdd gnd cell_6t
Xbit_r207_c197 bl_197 br_197 wl_207 vdd gnd cell_6t
Xbit_r208_c197 bl_197 br_197 wl_208 vdd gnd cell_6t
Xbit_r209_c197 bl_197 br_197 wl_209 vdd gnd cell_6t
Xbit_r210_c197 bl_197 br_197 wl_210 vdd gnd cell_6t
Xbit_r211_c197 bl_197 br_197 wl_211 vdd gnd cell_6t
Xbit_r212_c197 bl_197 br_197 wl_212 vdd gnd cell_6t
Xbit_r213_c197 bl_197 br_197 wl_213 vdd gnd cell_6t
Xbit_r214_c197 bl_197 br_197 wl_214 vdd gnd cell_6t
Xbit_r215_c197 bl_197 br_197 wl_215 vdd gnd cell_6t
Xbit_r216_c197 bl_197 br_197 wl_216 vdd gnd cell_6t
Xbit_r217_c197 bl_197 br_197 wl_217 vdd gnd cell_6t
Xbit_r218_c197 bl_197 br_197 wl_218 vdd gnd cell_6t
Xbit_r219_c197 bl_197 br_197 wl_219 vdd gnd cell_6t
Xbit_r220_c197 bl_197 br_197 wl_220 vdd gnd cell_6t
Xbit_r221_c197 bl_197 br_197 wl_221 vdd gnd cell_6t
Xbit_r222_c197 bl_197 br_197 wl_222 vdd gnd cell_6t
Xbit_r223_c197 bl_197 br_197 wl_223 vdd gnd cell_6t
Xbit_r224_c197 bl_197 br_197 wl_224 vdd gnd cell_6t
Xbit_r225_c197 bl_197 br_197 wl_225 vdd gnd cell_6t
Xbit_r226_c197 bl_197 br_197 wl_226 vdd gnd cell_6t
Xbit_r227_c197 bl_197 br_197 wl_227 vdd gnd cell_6t
Xbit_r228_c197 bl_197 br_197 wl_228 vdd gnd cell_6t
Xbit_r229_c197 bl_197 br_197 wl_229 vdd gnd cell_6t
Xbit_r230_c197 bl_197 br_197 wl_230 vdd gnd cell_6t
Xbit_r231_c197 bl_197 br_197 wl_231 vdd gnd cell_6t
Xbit_r232_c197 bl_197 br_197 wl_232 vdd gnd cell_6t
Xbit_r233_c197 bl_197 br_197 wl_233 vdd gnd cell_6t
Xbit_r234_c197 bl_197 br_197 wl_234 vdd gnd cell_6t
Xbit_r235_c197 bl_197 br_197 wl_235 vdd gnd cell_6t
Xbit_r236_c197 bl_197 br_197 wl_236 vdd gnd cell_6t
Xbit_r237_c197 bl_197 br_197 wl_237 vdd gnd cell_6t
Xbit_r238_c197 bl_197 br_197 wl_238 vdd gnd cell_6t
Xbit_r239_c197 bl_197 br_197 wl_239 vdd gnd cell_6t
Xbit_r240_c197 bl_197 br_197 wl_240 vdd gnd cell_6t
Xbit_r241_c197 bl_197 br_197 wl_241 vdd gnd cell_6t
Xbit_r242_c197 bl_197 br_197 wl_242 vdd gnd cell_6t
Xbit_r243_c197 bl_197 br_197 wl_243 vdd gnd cell_6t
Xbit_r244_c197 bl_197 br_197 wl_244 vdd gnd cell_6t
Xbit_r245_c197 bl_197 br_197 wl_245 vdd gnd cell_6t
Xbit_r246_c197 bl_197 br_197 wl_246 vdd gnd cell_6t
Xbit_r247_c197 bl_197 br_197 wl_247 vdd gnd cell_6t
Xbit_r248_c197 bl_197 br_197 wl_248 vdd gnd cell_6t
Xbit_r249_c197 bl_197 br_197 wl_249 vdd gnd cell_6t
Xbit_r250_c197 bl_197 br_197 wl_250 vdd gnd cell_6t
Xbit_r251_c197 bl_197 br_197 wl_251 vdd gnd cell_6t
Xbit_r252_c197 bl_197 br_197 wl_252 vdd gnd cell_6t
Xbit_r253_c197 bl_197 br_197 wl_253 vdd gnd cell_6t
Xbit_r254_c197 bl_197 br_197 wl_254 vdd gnd cell_6t
Xbit_r255_c197 bl_197 br_197 wl_255 vdd gnd cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd cell_6t
Xbit_r1_c198 bl_198 br_198 wl_1 vdd gnd cell_6t
Xbit_r2_c198 bl_198 br_198 wl_2 vdd gnd cell_6t
Xbit_r3_c198 bl_198 br_198 wl_3 vdd gnd cell_6t
Xbit_r4_c198 bl_198 br_198 wl_4 vdd gnd cell_6t
Xbit_r5_c198 bl_198 br_198 wl_5 vdd gnd cell_6t
Xbit_r6_c198 bl_198 br_198 wl_6 vdd gnd cell_6t
Xbit_r7_c198 bl_198 br_198 wl_7 vdd gnd cell_6t
Xbit_r8_c198 bl_198 br_198 wl_8 vdd gnd cell_6t
Xbit_r9_c198 bl_198 br_198 wl_9 vdd gnd cell_6t
Xbit_r10_c198 bl_198 br_198 wl_10 vdd gnd cell_6t
Xbit_r11_c198 bl_198 br_198 wl_11 vdd gnd cell_6t
Xbit_r12_c198 bl_198 br_198 wl_12 vdd gnd cell_6t
Xbit_r13_c198 bl_198 br_198 wl_13 vdd gnd cell_6t
Xbit_r14_c198 bl_198 br_198 wl_14 vdd gnd cell_6t
Xbit_r15_c198 bl_198 br_198 wl_15 vdd gnd cell_6t
Xbit_r16_c198 bl_198 br_198 wl_16 vdd gnd cell_6t
Xbit_r17_c198 bl_198 br_198 wl_17 vdd gnd cell_6t
Xbit_r18_c198 bl_198 br_198 wl_18 vdd gnd cell_6t
Xbit_r19_c198 bl_198 br_198 wl_19 vdd gnd cell_6t
Xbit_r20_c198 bl_198 br_198 wl_20 vdd gnd cell_6t
Xbit_r21_c198 bl_198 br_198 wl_21 vdd gnd cell_6t
Xbit_r22_c198 bl_198 br_198 wl_22 vdd gnd cell_6t
Xbit_r23_c198 bl_198 br_198 wl_23 vdd gnd cell_6t
Xbit_r24_c198 bl_198 br_198 wl_24 vdd gnd cell_6t
Xbit_r25_c198 bl_198 br_198 wl_25 vdd gnd cell_6t
Xbit_r26_c198 bl_198 br_198 wl_26 vdd gnd cell_6t
Xbit_r27_c198 bl_198 br_198 wl_27 vdd gnd cell_6t
Xbit_r28_c198 bl_198 br_198 wl_28 vdd gnd cell_6t
Xbit_r29_c198 bl_198 br_198 wl_29 vdd gnd cell_6t
Xbit_r30_c198 bl_198 br_198 wl_30 vdd gnd cell_6t
Xbit_r31_c198 bl_198 br_198 wl_31 vdd gnd cell_6t
Xbit_r32_c198 bl_198 br_198 wl_32 vdd gnd cell_6t
Xbit_r33_c198 bl_198 br_198 wl_33 vdd gnd cell_6t
Xbit_r34_c198 bl_198 br_198 wl_34 vdd gnd cell_6t
Xbit_r35_c198 bl_198 br_198 wl_35 vdd gnd cell_6t
Xbit_r36_c198 bl_198 br_198 wl_36 vdd gnd cell_6t
Xbit_r37_c198 bl_198 br_198 wl_37 vdd gnd cell_6t
Xbit_r38_c198 bl_198 br_198 wl_38 vdd gnd cell_6t
Xbit_r39_c198 bl_198 br_198 wl_39 vdd gnd cell_6t
Xbit_r40_c198 bl_198 br_198 wl_40 vdd gnd cell_6t
Xbit_r41_c198 bl_198 br_198 wl_41 vdd gnd cell_6t
Xbit_r42_c198 bl_198 br_198 wl_42 vdd gnd cell_6t
Xbit_r43_c198 bl_198 br_198 wl_43 vdd gnd cell_6t
Xbit_r44_c198 bl_198 br_198 wl_44 vdd gnd cell_6t
Xbit_r45_c198 bl_198 br_198 wl_45 vdd gnd cell_6t
Xbit_r46_c198 bl_198 br_198 wl_46 vdd gnd cell_6t
Xbit_r47_c198 bl_198 br_198 wl_47 vdd gnd cell_6t
Xbit_r48_c198 bl_198 br_198 wl_48 vdd gnd cell_6t
Xbit_r49_c198 bl_198 br_198 wl_49 vdd gnd cell_6t
Xbit_r50_c198 bl_198 br_198 wl_50 vdd gnd cell_6t
Xbit_r51_c198 bl_198 br_198 wl_51 vdd gnd cell_6t
Xbit_r52_c198 bl_198 br_198 wl_52 vdd gnd cell_6t
Xbit_r53_c198 bl_198 br_198 wl_53 vdd gnd cell_6t
Xbit_r54_c198 bl_198 br_198 wl_54 vdd gnd cell_6t
Xbit_r55_c198 bl_198 br_198 wl_55 vdd gnd cell_6t
Xbit_r56_c198 bl_198 br_198 wl_56 vdd gnd cell_6t
Xbit_r57_c198 bl_198 br_198 wl_57 vdd gnd cell_6t
Xbit_r58_c198 bl_198 br_198 wl_58 vdd gnd cell_6t
Xbit_r59_c198 bl_198 br_198 wl_59 vdd gnd cell_6t
Xbit_r60_c198 bl_198 br_198 wl_60 vdd gnd cell_6t
Xbit_r61_c198 bl_198 br_198 wl_61 vdd gnd cell_6t
Xbit_r62_c198 bl_198 br_198 wl_62 vdd gnd cell_6t
Xbit_r63_c198 bl_198 br_198 wl_63 vdd gnd cell_6t
Xbit_r64_c198 bl_198 br_198 wl_64 vdd gnd cell_6t
Xbit_r65_c198 bl_198 br_198 wl_65 vdd gnd cell_6t
Xbit_r66_c198 bl_198 br_198 wl_66 vdd gnd cell_6t
Xbit_r67_c198 bl_198 br_198 wl_67 vdd gnd cell_6t
Xbit_r68_c198 bl_198 br_198 wl_68 vdd gnd cell_6t
Xbit_r69_c198 bl_198 br_198 wl_69 vdd gnd cell_6t
Xbit_r70_c198 bl_198 br_198 wl_70 vdd gnd cell_6t
Xbit_r71_c198 bl_198 br_198 wl_71 vdd gnd cell_6t
Xbit_r72_c198 bl_198 br_198 wl_72 vdd gnd cell_6t
Xbit_r73_c198 bl_198 br_198 wl_73 vdd gnd cell_6t
Xbit_r74_c198 bl_198 br_198 wl_74 vdd gnd cell_6t
Xbit_r75_c198 bl_198 br_198 wl_75 vdd gnd cell_6t
Xbit_r76_c198 bl_198 br_198 wl_76 vdd gnd cell_6t
Xbit_r77_c198 bl_198 br_198 wl_77 vdd gnd cell_6t
Xbit_r78_c198 bl_198 br_198 wl_78 vdd gnd cell_6t
Xbit_r79_c198 bl_198 br_198 wl_79 vdd gnd cell_6t
Xbit_r80_c198 bl_198 br_198 wl_80 vdd gnd cell_6t
Xbit_r81_c198 bl_198 br_198 wl_81 vdd gnd cell_6t
Xbit_r82_c198 bl_198 br_198 wl_82 vdd gnd cell_6t
Xbit_r83_c198 bl_198 br_198 wl_83 vdd gnd cell_6t
Xbit_r84_c198 bl_198 br_198 wl_84 vdd gnd cell_6t
Xbit_r85_c198 bl_198 br_198 wl_85 vdd gnd cell_6t
Xbit_r86_c198 bl_198 br_198 wl_86 vdd gnd cell_6t
Xbit_r87_c198 bl_198 br_198 wl_87 vdd gnd cell_6t
Xbit_r88_c198 bl_198 br_198 wl_88 vdd gnd cell_6t
Xbit_r89_c198 bl_198 br_198 wl_89 vdd gnd cell_6t
Xbit_r90_c198 bl_198 br_198 wl_90 vdd gnd cell_6t
Xbit_r91_c198 bl_198 br_198 wl_91 vdd gnd cell_6t
Xbit_r92_c198 bl_198 br_198 wl_92 vdd gnd cell_6t
Xbit_r93_c198 bl_198 br_198 wl_93 vdd gnd cell_6t
Xbit_r94_c198 bl_198 br_198 wl_94 vdd gnd cell_6t
Xbit_r95_c198 bl_198 br_198 wl_95 vdd gnd cell_6t
Xbit_r96_c198 bl_198 br_198 wl_96 vdd gnd cell_6t
Xbit_r97_c198 bl_198 br_198 wl_97 vdd gnd cell_6t
Xbit_r98_c198 bl_198 br_198 wl_98 vdd gnd cell_6t
Xbit_r99_c198 bl_198 br_198 wl_99 vdd gnd cell_6t
Xbit_r100_c198 bl_198 br_198 wl_100 vdd gnd cell_6t
Xbit_r101_c198 bl_198 br_198 wl_101 vdd gnd cell_6t
Xbit_r102_c198 bl_198 br_198 wl_102 vdd gnd cell_6t
Xbit_r103_c198 bl_198 br_198 wl_103 vdd gnd cell_6t
Xbit_r104_c198 bl_198 br_198 wl_104 vdd gnd cell_6t
Xbit_r105_c198 bl_198 br_198 wl_105 vdd gnd cell_6t
Xbit_r106_c198 bl_198 br_198 wl_106 vdd gnd cell_6t
Xbit_r107_c198 bl_198 br_198 wl_107 vdd gnd cell_6t
Xbit_r108_c198 bl_198 br_198 wl_108 vdd gnd cell_6t
Xbit_r109_c198 bl_198 br_198 wl_109 vdd gnd cell_6t
Xbit_r110_c198 bl_198 br_198 wl_110 vdd gnd cell_6t
Xbit_r111_c198 bl_198 br_198 wl_111 vdd gnd cell_6t
Xbit_r112_c198 bl_198 br_198 wl_112 vdd gnd cell_6t
Xbit_r113_c198 bl_198 br_198 wl_113 vdd gnd cell_6t
Xbit_r114_c198 bl_198 br_198 wl_114 vdd gnd cell_6t
Xbit_r115_c198 bl_198 br_198 wl_115 vdd gnd cell_6t
Xbit_r116_c198 bl_198 br_198 wl_116 vdd gnd cell_6t
Xbit_r117_c198 bl_198 br_198 wl_117 vdd gnd cell_6t
Xbit_r118_c198 bl_198 br_198 wl_118 vdd gnd cell_6t
Xbit_r119_c198 bl_198 br_198 wl_119 vdd gnd cell_6t
Xbit_r120_c198 bl_198 br_198 wl_120 vdd gnd cell_6t
Xbit_r121_c198 bl_198 br_198 wl_121 vdd gnd cell_6t
Xbit_r122_c198 bl_198 br_198 wl_122 vdd gnd cell_6t
Xbit_r123_c198 bl_198 br_198 wl_123 vdd gnd cell_6t
Xbit_r124_c198 bl_198 br_198 wl_124 vdd gnd cell_6t
Xbit_r125_c198 bl_198 br_198 wl_125 vdd gnd cell_6t
Xbit_r126_c198 bl_198 br_198 wl_126 vdd gnd cell_6t
Xbit_r127_c198 bl_198 br_198 wl_127 vdd gnd cell_6t
Xbit_r128_c198 bl_198 br_198 wl_128 vdd gnd cell_6t
Xbit_r129_c198 bl_198 br_198 wl_129 vdd gnd cell_6t
Xbit_r130_c198 bl_198 br_198 wl_130 vdd gnd cell_6t
Xbit_r131_c198 bl_198 br_198 wl_131 vdd gnd cell_6t
Xbit_r132_c198 bl_198 br_198 wl_132 vdd gnd cell_6t
Xbit_r133_c198 bl_198 br_198 wl_133 vdd gnd cell_6t
Xbit_r134_c198 bl_198 br_198 wl_134 vdd gnd cell_6t
Xbit_r135_c198 bl_198 br_198 wl_135 vdd gnd cell_6t
Xbit_r136_c198 bl_198 br_198 wl_136 vdd gnd cell_6t
Xbit_r137_c198 bl_198 br_198 wl_137 vdd gnd cell_6t
Xbit_r138_c198 bl_198 br_198 wl_138 vdd gnd cell_6t
Xbit_r139_c198 bl_198 br_198 wl_139 vdd gnd cell_6t
Xbit_r140_c198 bl_198 br_198 wl_140 vdd gnd cell_6t
Xbit_r141_c198 bl_198 br_198 wl_141 vdd gnd cell_6t
Xbit_r142_c198 bl_198 br_198 wl_142 vdd gnd cell_6t
Xbit_r143_c198 bl_198 br_198 wl_143 vdd gnd cell_6t
Xbit_r144_c198 bl_198 br_198 wl_144 vdd gnd cell_6t
Xbit_r145_c198 bl_198 br_198 wl_145 vdd gnd cell_6t
Xbit_r146_c198 bl_198 br_198 wl_146 vdd gnd cell_6t
Xbit_r147_c198 bl_198 br_198 wl_147 vdd gnd cell_6t
Xbit_r148_c198 bl_198 br_198 wl_148 vdd gnd cell_6t
Xbit_r149_c198 bl_198 br_198 wl_149 vdd gnd cell_6t
Xbit_r150_c198 bl_198 br_198 wl_150 vdd gnd cell_6t
Xbit_r151_c198 bl_198 br_198 wl_151 vdd gnd cell_6t
Xbit_r152_c198 bl_198 br_198 wl_152 vdd gnd cell_6t
Xbit_r153_c198 bl_198 br_198 wl_153 vdd gnd cell_6t
Xbit_r154_c198 bl_198 br_198 wl_154 vdd gnd cell_6t
Xbit_r155_c198 bl_198 br_198 wl_155 vdd gnd cell_6t
Xbit_r156_c198 bl_198 br_198 wl_156 vdd gnd cell_6t
Xbit_r157_c198 bl_198 br_198 wl_157 vdd gnd cell_6t
Xbit_r158_c198 bl_198 br_198 wl_158 vdd gnd cell_6t
Xbit_r159_c198 bl_198 br_198 wl_159 vdd gnd cell_6t
Xbit_r160_c198 bl_198 br_198 wl_160 vdd gnd cell_6t
Xbit_r161_c198 bl_198 br_198 wl_161 vdd gnd cell_6t
Xbit_r162_c198 bl_198 br_198 wl_162 vdd gnd cell_6t
Xbit_r163_c198 bl_198 br_198 wl_163 vdd gnd cell_6t
Xbit_r164_c198 bl_198 br_198 wl_164 vdd gnd cell_6t
Xbit_r165_c198 bl_198 br_198 wl_165 vdd gnd cell_6t
Xbit_r166_c198 bl_198 br_198 wl_166 vdd gnd cell_6t
Xbit_r167_c198 bl_198 br_198 wl_167 vdd gnd cell_6t
Xbit_r168_c198 bl_198 br_198 wl_168 vdd gnd cell_6t
Xbit_r169_c198 bl_198 br_198 wl_169 vdd gnd cell_6t
Xbit_r170_c198 bl_198 br_198 wl_170 vdd gnd cell_6t
Xbit_r171_c198 bl_198 br_198 wl_171 vdd gnd cell_6t
Xbit_r172_c198 bl_198 br_198 wl_172 vdd gnd cell_6t
Xbit_r173_c198 bl_198 br_198 wl_173 vdd gnd cell_6t
Xbit_r174_c198 bl_198 br_198 wl_174 vdd gnd cell_6t
Xbit_r175_c198 bl_198 br_198 wl_175 vdd gnd cell_6t
Xbit_r176_c198 bl_198 br_198 wl_176 vdd gnd cell_6t
Xbit_r177_c198 bl_198 br_198 wl_177 vdd gnd cell_6t
Xbit_r178_c198 bl_198 br_198 wl_178 vdd gnd cell_6t
Xbit_r179_c198 bl_198 br_198 wl_179 vdd gnd cell_6t
Xbit_r180_c198 bl_198 br_198 wl_180 vdd gnd cell_6t
Xbit_r181_c198 bl_198 br_198 wl_181 vdd gnd cell_6t
Xbit_r182_c198 bl_198 br_198 wl_182 vdd gnd cell_6t
Xbit_r183_c198 bl_198 br_198 wl_183 vdd gnd cell_6t
Xbit_r184_c198 bl_198 br_198 wl_184 vdd gnd cell_6t
Xbit_r185_c198 bl_198 br_198 wl_185 vdd gnd cell_6t
Xbit_r186_c198 bl_198 br_198 wl_186 vdd gnd cell_6t
Xbit_r187_c198 bl_198 br_198 wl_187 vdd gnd cell_6t
Xbit_r188_c198 bl_198 br_198 wl_188 vdd gnd cell_6t
Xbit_r189_c198 bl_198 br_198 wl_189 vdd gnd cell_6t
Xbit_r190_c198 bl_198 br_198 wl_190 vdd gnd cell_6t
Xbit_r191_c198 bl_198 br_198 wl_191 vdd gnd cell_6t
Xbit_r192_c198 bl_198 br_198 wl_192 vdd gnd cell_6t
Xbit_r193_c198 bl_198 br_198 wl_193 vdd gnd cell_6t
Xbit_r194_c198 bl_198 br_198 wl_194 vdd gnd cell_6t
Xbit_r195_c198 bl_198 br_198 wl_195 vdd gnd cell_6t
Xbit_r196_c198 bl_198 br_198 wl_196 vdd gnd cell_6t
Xbit_r197_c198 bl_198 br_198 wl_197 vdd gnd cell_6t
Xbit_r198_c198 bl_198 br_198 wl_198 vdd gnd cell_6t
Xbit_r199_c198 bl_198 br_198 wl_199 vdd gnd cell_6t
Xbit_r200_c198 bl_198 br_198 wl_200 vdd gnd cell_6t
Xbit_r201_c198 bl_198 br_198 wl_201 vdd gnd cell_6t
Xbit_r202_c198 bl_198 br_198 wl_202 vdd gnd cell_6t
Xbit_r203_c198 bl_198 br_198 wl_203 vdd gnd cell_6t
Xbit_r204_c198 bl_198 br_198 wl_204 vdd gnd cell_6t
Xbit_r205_c198 bl_198 br_198 wl_205 vdd gnd cell_6t
Xbit_r206_c198 bl_198 br_198 wl_206 vdd gnd cell_6t
Xbit_r207_c198 bl_198 br_198 wl_207 vdd gnd cell_6t
Xbit_r208_c198 bl_198 br_198 wl_208 vdd gnd cell_6t
Xbit_r209_c198 bl_198 br_198 wl_209 vdd gnd cell_6t
Xbit_r210_c198 bl_198 br_198 wl_210 vdd gnd cell_6t
Xbit_r211_c198 bl_198 br_198 wl_211 vdd gnd cell_6t
Xbit_r212_c198 bl_198 br_198 wl_212 vdd gnd cell_6t
Xbit_r213_c198 bl_198 br_198 wl_213 vdd gnd cell_6t
Xbit_r214_c198 bl_198 br_198 wl_214 vdd gnd cell_6t
Xbit_r215_c198 bl_198 br_198 wl_215 vdd gnd cell_6t
Xbit_r216_c198 bl_198 br_198 wl_216 vdd gnd cell_6t
Xbit_r217_c198 bl_198 br_198 wl_217 vdd gnd cell_6t
Xbit_r218_c198 bl_198 br_198 wl_218 vdd gnd cell_6t
Xbit_r219_c198 bl_198 br_198 wl_219 vdd gnd cell_6t
Xbit_r220_c198 bl_198 br_198 wl_220 vdd gnd cell_6t
Xbit_r221_c198 bl_198 br_198 wl_221 vdd gnd cell_6t
Xbit_r222_c198 bl_198 br_198 wl_222 vdd gnd cell_6t
Xbit_r223_c198 bl_198 br_198 wl_223 vdd gnd cell_6t
Xbit_r224_c198 bl_198 br_198 wl_224 vdd gnd cell_6t
Xbit_r225_c198 bl_198 br_198 wl_225 vdd gnd cell_6t
Xbit_r226_c198 bl_198 br_198 wl_226 vdd gnd cell_6t
Xbit_r227_c198 bl_198 br_198 wl_227 vdd gnd cell_6t
Xbit_r228_c198 bl_198 br_198 wl_228 vdd gnd cell_6t
Xbit_r229_c198 bl_198 br_198 wl_229 vdd gnd cell_6t
Xbit_r230_c198 bl_198 br_198 wl_230 vdd gnd cell_6t
Xbit_r231_c198 bl_198 br_198 wl_231 vdd gnd cell_6t
Xbit_r232_c198 bl_198 br_198 wl_232 vdd gnd cell_6t
Xbit_r233_c198 bl_198 br_198 wl_233 vdd gnd cell_6t
Xbit_r234_c198 bl_198 br_198 wl_234 vdd gnd cell_6t
Xbit_r235_c198 bl_198 br_198 wl_235 vdd gnd cell_6t
Xbit_r236_c198 bl_198 br_198 wl_236 vdd gnd cell_6t
Xbit_r237_c198 bl_198 br_198 wl_237 vdd gnd cell_6t
Xbit_r238_c198 bl_198 br_198 wl_238 vdd gnd cell_6t
Xbit_r239_c198 bl_198 br_198 wl_239 vdd gnd cell_6t
Xbit_r240_c198 bl_198 br_198 wl_240 vdd gnd cell_6t
Xbit_r241_c198 bl_198 br_198 wl_241 vdd gnd cell_6t
Xbit_r242_c198 bl_198 br_198 wl_242 vdd gnd cell_6t
Xbit_r243_c198 bl_198 br_198 wl_243 vdd gnd cell_6t
Xbit_r244_c198 bl_198 br_198 wl_244 vdd gnd cell_6t
Xbit_r245_c198 bl_198 br_198 wl_245 vdd gnd cell_6t
Xbit_r246_c198 bl_198 br_198 wl_246 vdd gnd cell_6t
Xbit_r247_c198 bl_198 br_198 wl_247 vdd gnd cell_6t
Xbit_r248_c198 bl_198 br_198 wl_248 vdd gnd cell_6t
Xbit_r249_c198 bl_198 br_198 wl_249 vdd gnd cell_6t
Xbit_r250_c198 bl_198 br_198 wl_250 vdd gnd cell_6t
Xbit_r251_c198 bl_198 br_198 wl_251 vdd gnd cell_6t
Xbit_r252_c198 bl_198 br_198 wl_252 vdd gnd cell_6t
Xbit_r253_c198 bl_198 br_198 wl_253 vdd gnd cell_6t
Xbit_r254_c198 bl_198 br_198 wl_254 vdd gnd cell_6t
Xbit_r255_c198 bl_198 br_198 wl_255 vdd gnd cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd cell_6t
Xbit_r1_c199 bl_199 br_199 wl_1 vdd gnd cell_6t
Xbit_r2_c199 bl_199 br_199 wl_2 vdd gnd cell_6t
Xbit_r3_c199 bl_199 br_199 wl_3 vdd gnd cell_6t
Xbit_r4_c199 bl_199 br_199 wl_4 vdd gnd cell_6t
Xbit_r5_c199 bl_199 br_199 wl_5 vdd gnd cell_6t
Xbit_r6_c199 bl_199 br_199 wl_6 vdd gnd cell_6t
Xbit_r7_c199 bl_199 br_199 wl_7 vdd gnd cell_6t
Xbit_r8_c199 bl_199 br_199 wl_8 vdd gnd cell_6t
Xbit_r9_c199 bl_199 br_199 wl_9 vdd gnd cell_6t
Xbit_r10_c199 bl_199 br_199 wl_10 vdd gnd cell_6t
Xbit_r11_c199 bl_199 br_199 wl_11 vdd gnd cell_6t
Xbit_r12_c199 bl_199 br_199 wl_12 vdd gnd cell_6t
Xbit_r13_c199 bl_199 br_199 wl_13 vdd gnd cell_6t
Xbit_r14_c199 bl_199 br_199 wl_14 vdd gnd cell_6t
Xbit_r15_c199 bl_199 br_199 wl_15 vdd gnd cell_6t
Xbit_r16_c199 bl_199 br_199 wl_16 vdd gnd cell_6t
Xbit_r17_c199 bl_199 br_199 wl_17 vdd gnd cell_6t
Xbit_r18_c199 bl_199 br_199 wl_18 vdd gnd cell_6t
Xbit_r19_c199 bl_199 br_199 wl_19 vdd gnd cell_6t
Xbit_r20_c199 bl_199 br_199 wl_20 vdd gnd cell_6t
Xbit_r21_c199 bl_199 br_199 wl_21 vdd gnd cell_6t
Xbit_r22_c199 bl_199 br_199 wl_22 vdd gnd cell_6t
Xbit_r23_c199 bl_199 br_199 wl_23 vdd gnd cell_6t
Xbit_r24_c199 bl_199 br_199 wl_24 vdd gnd cell_6t
Xbit_r25_c199 bl_199 br_199 wl_25 vdd gnd cell_6t
Xbit_r26_c199 bl_199 br_199 wl_26 vdd gnd cell_6t
Xbit_r27_c199 bl_199 br_199 wl_27 vdd gnd cell_6t
Xbit_r28_c199 bl_199 br_199 wl_28 vdd gnd cell_6t
Xbit_r29_c199 bl_199 br_199 wl_29 vdd gnd cell_6t
Xbit_r30_c199 bl_199 br_199 wl_30 vdd gnd cell_6t
Xbit_r31_c199 bl_199 br_199 wl_31 vdd gnd cell_6t
Xbit_r32_c199 bl_199 br_199 wl_32 vdd gnd cell_6t
Xbit_r33_c199 bl_199 br_199 wl_33 vdd gnd cell_6t
Xbit_r34_c199 bl_199 br_199 wl_34 vdd gnd cell_6t
Xbit_r35_c199 bl_199 br_199 wl_35 vdd gnd cell_6t
Xbit_r36_c199 bl_199 br_199 wl_36 vdd gnd cell_6t
Xbit_r37_c199 bl_199 br_199 wl_37 vdd gnd cell_6t
Xbit_r38_c199 bl_199 br_199 wl_38 vdd gnd cell_6t
Xbit_r39_c199 bl_199 br_199 wl_39 vdd gnd cell_6t
Xbit_r40_c199 bl_199 br_199 wl_40 vdd gnd cell_6t
Xbit_r41_c199 bl_199 br_199 wl_41 vdd gnd cell_6t
Xbit_r42_c199 bl_199 br_199 wl_42 vdd gnd cell_6t
Xbit_r43_c199 bl_199 br_199 wl_43 vdd gnd cell_6t
Xbit_r44_c199 bl_199 br_199 wl_44 vdd gnd cell_6t
Xbit_r45_c199 bl_199 br_199 wl_45 vdd gnd cell_6t
Xbit_r46_c199 bl_199 br_199 wl_46 vdd gnd cell_6t
Xbit_r47_c199 bl_199 br_199 wl_47 vdd gnd cell_6t
Xbit_r48_c199 bl_199 br_199 wl_48 vdd gnd cell_6t
Xbit_r49_c199 bl_199 br_199 wl_49 vdd gnd cell_6t
Xbit_r50_c199 bl_199 br_199 wl_50 vdd gnd cell_6t
Xbit_r51_c199 bl_199 br_199 wl_51 vdd gnd cell_6t
Xbit_r52_c199 bl_199 br_199 wl_52 vdd gnd cell_6t
Xbit_r53_c199 bl_199 br_199 wl_53 vdd gnd cell_6t
Xbit_r54_c199 bl_199 br_199 wl_54 vdd gnd cell_6t
Xbit_r55_c199 bl_199 br_199 wl_55 vdd gnd cell_6t
Xbit_r56_c199 bl_199 br_199 wl_56 vdd gnd cell_6t
Xbit_r57_c199 bl_199 br_199 wl_57 vdd gnd cell_6t
Xbit_r58_c199 bl_199 br_199 wl_58 vdd gnd cell_6t
Xbit_r59_c199 bl_199 br_199 wl_59 vdd gnd cell_6t
Xbit_r60_c199 bl_199 br_199 wl_60 vdd gnd cell_6t
Xbit_r61_c199 bl_199 br_199 wl_61 vdd gnd cell_6t
Xbit_r62_c199 bl_199 br_199 wl_62 vdd gnd cell_6t
Xbit_r63_c199 bl_199 br_199 wl_63 vdd gnd cell_6t
Xbit_r64_c199 bl_199 br_199 wl_64 vdd gnd cell_6t
Xbit_r65_c199 bl_199 br_199 wl_65 vdd gnd cell_6t
Xbit_r66_c199 bl_199 br_199 wl_66 vdd gnd cell_6t
Xbit_r67_c199 bl_199 br_199 wl_67 vdd gnd cell_6t
Xbit_r68_c199 bl_199 br_199 wl_68 vdd gnd cell_6t
Xbit_r69_c199 bl_199 br_199 wl_69 vdd gnd cell_6t
Xbit_r70_c199 bl_199 br_199 wl_70 vdd gnd cell_6t
Xbit_r71_c199 bl_199 br_199 wl_71 vdd gnd cell_6t
Xbit_r72_c199 bl_199 br_199 wl_72 vdd gnd cell_6t
Xbit_r73_c199 bl_199 br_199 wl_73 vdd gnd cell_6t
Xbit_r74_c199 bl_199 br_199 wl_74 vdd gnd cell_6t
Xbit_r75_c199 bl_199 br_199 wl_75 vdd gnd cell_6t
Xbit_r76_c199 bl_199 br_199 wl_76 vdd gnd cell_6t
Xbit_r77_c199 bl_199 br_199 wl_77 vdd gnd cell_6t
Xbit_r78_c199 bl_199 br_199 wl_78 vdd gnd cell_6t
Xbit_r79_c199 bl_199 br_199 wl_79 vdd gnd cell_6t
Xbit_r80_c199 bl_199 br_199 wl_80 vdd gnd cell_6t
Xbit_r81_c199 bl_199 br_199 wl_81 vdd gnd cell_6t
Xbit_r82_c199 bl_199 br_199 wl_82 vdd gnd cell_6t
Xbit_r83_c199 bl_199 br_199 wl_83 vdd gnd cell_6t
Xbit_r84_c199 bl_199 br_199 wl_84 vdd gnd cell_6t
Xbit_r85_c199 bl_199 br_199 wl_85 vdd gnd cell_6t
Xbit_r86_c199 bl_199 br_199 wl_86 vdd gnd cell_6t
Xbit_r87_c199 bl_199 br_199 wl_87 vdd gnd cell_6t
Xbit_r88_c199 bl_199 br_199 wl_88 vdd gnd cell_6t
Xbit_r89_c199 bl_199 br_199 wl_89 vdd gnd cell_6t
Xbit_r90_c199 bl_199 br_199 wl_90 vdd gnd cell_6t
Xbit_r91_c199 bl_199 br_199 wl_91 vdd gnd cell_6t
Xbit_r92_c199 bl_199 br_199 wl_92 vdd gnd cell_6t
Xbit_r93_c199 bl_199 br_199 wl_93 vdd gnd cell_6t
Xbit_r94_c199 bl_199 br_199 wl_94 vdd gnd cell_6t
Xbit_r95_c199 bl_199 br_199 wl_95 vdd gnd cell_6t
Xbit_r96_c199 bl_199 br_199 wl_96 vdd gnd cell_6t
Xbit_r97_c199 bl_199 br_199 wl_97 vdd gnd cell_6t
Xbit_r98_c199 bl_199 br_199 wl_98 vdd gnd cell_6t
Xbit_r99_c199 bl_199 br_199 wl_99 vdd gnd cell_6t
Xbit_r100_c199 bl_199 br_199 wl_100 vdd gnd cell_6t
Xbit_r101_c199 bl_199 br_199 wl_101 vdd gnd cell_6t
Xbit_r102_c199 bl_199 br_199 wl_102 vdd gnd cell_6t
Xbit_r103_c199 bl_199 br_199 wl_103 vdd gnd cell_6t
Xbit_r104_c199 bl_199 br_199 wl_104 vdd gnd cell_6t
Xbit_r105_c199 bl_199 br_199 wl_105 vdd gnd cell_6t
Xbit_r106_c199 bl_199 br_199 wl_106 vdd gnd cell_6t
Xbit_r107_c199 bl_199 br_199 wl_107 vdd gnd cell_6t
Xbit_r108_c199 bl_199 br_199 wl_108 vdd gnd cell_6t
Xbit_r109_c199 bl_199 br_199 wl_109 vdd gnd cell_6t
Xbit_r110_c199 bl_199 br_199 wl_110 vdd gnd cell_6t
Xbit_r111_c199 bl_199 br_199 wl_111 vdd gnd cell_6t
Xbit_r112_c199 bl_199 br_199 wl_112 vdd gnd cell_6t
Xbit_r113_c199 bl_199 br_199 wl_113 vdd gnd cell_6t
Xbit_r114_c199 bl_199 br_199 wl_114 vdd gnd cell_6t
Xbit_r115_c199 bl_199 br_199 wl_115 vdd gnd cell_6t
Xbit_r116_c199 bl_199 br_199 wl_116 vdd gnd cell_6t
Xbit_r117_c199 bl_199 br_199 wl_117 vdd gnd cell_6t
Xbit_r118_c199 bl_199 br_199 wl_118 vdd gnd cell_6t
Xbit_r119_c199 bl_199 br_199 wl_119 vdd gnd cell_6t
Xbit_r120_c199 bl_199 br_199 wl_120 vdd gnd cell_6t
Xbit_r121_c199 bl_199 br_199 wl_121 vdd gnd cell_6t
Xbit_r122_c199 bl_199 br_199 wl_122 vdd gnd cell_6t
Xbit_r123_c199 bl_199 br_199 wl_123 vdd gnd cell_6t
Xbit_r124_c199 bl_199 br_199 wl_124 vdd gnd cell_6t
Xbit_r125_c199 bl_199 br_199 wl_125 vdd gnd cell_6t
Xbit_r126_c199 bl_199 br_199 wl_126 vdd gnd cell_6t
Xbit_r127_c199 bl_199 br_199 wl_127 vdd gnd cell_6t
Xbit_r128_c199 bl_199 br_199 wl_128 vdd gnd cell_6t
Xbit_r129_c199 bl_199 br_199 wl_129 vdd gnd cell_6t
Xbit_r130_c199 bl_199 br_199 wl_130 vdd gnd cell_6t
Xbit_r131_c199 bl_199 br_199 wl_131 vdd gnd cell_6t
Xbit_r132_c199 bl_199 br_199 wl_132 vdd gnd cell_6t
Xbit_r133_c199 bl_199 br_199 wl_133 vdd gnd cell_6t
Xbit_r134_c199 bl_199 br_199 wl_134 vdd gnd cell_6t
Xbit_r135_c199 bl_199 br_199 wl_135 vdd gnd cell_6t
Xbit_r136_c199 bl_199 br_199 wl_136 vdd gnd cell_6t
Xbit_r137_c199 bl_199 br_199 wl_137 vdd gnd cell_6t
Xbit_r138_c199 bl_199 br_199 wl_138 vdd gnd cell_6t
Xbit_r139_c199 bl_199 br_199 wl_139 vdd gnd cell_6t
Xbit_r140_c199 bl_199 br_199 wl_140 vdd gnd cell_6t
Xbit_r141_c199 bl_199 br_199 wl_141 vdd gnd cell_6t
Xbit_r142_c199 bl_199 br_199 wl_142 vdd gnd cell_6t
Xbit_r143_c199 bl_199 br_199 wl_143 vdd gnd cell_6t
Xbit_r144_c199 bl_199 br_199 wl_144 vdd gnd cell_6t
Xbit_r145_c199 bl_199 br_199 wl_145 vdd gnd cell_6t
Xbit_r146_c199 bl_199 br_199 wl_146 vdd gnd cell_6t
Xbit_r147_c199 bl_199 br_199 wl_147 vdd gnd cell_6t
Xbit_r148_c199 bl_199 br_199 wl_148 vdd gnd cell_6t
Xbit_r149_c199 bl_199 br_199 wl_149 vdd gnd cell_6t
Xbit_r150_c199 bl_199 br_199 wl_150 vdd gnd cell_6t
Xbit_r151_c199 bl_199 br_199 wl_151 vdd gnd cell_6t
Xbit_r152_c199 bl_199 br_199 wl_152 vdd gnd cell_6t
Xbit_r153_c199 bl_199 br_199 wl_153 vdd gnd cell_6t
Xbit_r154_c199 bl_199 br_199 wl_154 vdd gnd cell_6t
Xbit_r155_c199 bl_199 br_199 wl_155 vdd gnd cell_6t
Xbit_r156_c199 bl_199 br_199 wl_156 vdd gnd cell_6t
Xbit_r157_c199 bl_199 br_199 wl_157 vdd gnd cell_6t
Xbit_r158_c199 bl_199 br_199 wl_158 vdd gnd cell_6t
Xbit_r159_c199 bl_199 br_199 wl_159 vdd gnd cell_6t
Xbit_r160_c199 bl_199 br_199 wl_160 vdd gnd cell_6t
Xbit_r161_c199 bl_199 br_199 wl_161 vdd gnd cell_6t
Xbit_r162_c199 bl_199 br_199 wl_162 vdd gnd cell_6t
Xbit_r163_c199 bl_199 br_199 wl_163 vdd gnd cell_6t
Xbit_r164_c199 bl_199 br_199 wl_164 vdd gnd cell_6t
Xbit_r165_c199 bl_199 br_199 wl_165 vdd gnd cell_6t
Xbit_r166_c199 bl_199 br_199 wl_166 vdd gnd cell_6t
Xbit_r167_c199 bl_199 br_199 wl_167 vdd gnd cell_6t
Xbit_r168_c199 bl_199 br_199 wl_168 vdd gnd cell_6t
Xbit_r169_c199 bl_199 br_199 wl_169 vdd gnd cell_6t
Xbit_r170_c199 bl_199 br_199 wl_170 vdd gnd cell_6t
Xbit_r171_c199 bl_199 br_199 wl_171 vdd gnd cell_6t
Xbit_r172_c199 bl_199 br_199 wl_172 vdd gnd cell_6t
Xbit_r173_c199 bl_199 br_199 wl_173 vdd gnd cell_6t
Xbit_r174_c199 bl_199 br_199 wl_174 vdd gnd cell_6t
Xbit_r175_c199 bl_199 br_199 wl_175 vdd gnd cell_6t
Xbit_r176_c199 bl_199 br_199 wl_176 vdd gnd cell_6t
Xbit_r177_c199 bl_199 br_199 wl_177 vdd gnd cell_6t
Xbit_r178_c199 bl_199 br_199 wl_178 vdd gnd cell_6t
Xbit_r179_c199 bl_199 br_199 wl_179 vdd gnd cell_6t
Xbit_r180_c199 bl_199 br_199 wl_180 vdd gnd cell_6t
Xbit_r181_c199 bl_199 br_199 wl_181 vdd gnd cell_6t
Xbit_r182_c199 bl_199 br_199 wl_182 vdd gnd cell_6t
Xbit_r183_c199 bl_199 br_199 wl_183 vdd gnd cell_6t
Xbit_r184_c199 bl_199 br_199 wl_184 vdd gnd cell_6t
Xbit_r185_c199 bl_199 br_199 wl_185 vdd gnd cell_6t
Xbit_r186_c199 bl_199 br_199 wl_186 vdd gnd cell_6t
Xbit_r187_c199 bl_199 br_199 wl_187 vdd gnd cell_6t
Xbit_r188_c199 bl_199 br_199 wl_188 vdd gnd cell_6t
Xbit_r189_c199 bl_199 br_199 wl_189 vdd gnd cell_6t
Xbit_r190_c199 bl_199 br_199 wl_190 vdd gnd cell_6t
Xbit_r191_c199 bl_199 br_199 wl_191 vdd gnd cell_6t
Xbit_r192_c199 bl_199 br_199 wl_192 vdd gnd cell_6t
Xbit_r193_c199 bl_199 br_199 wl_193 vdd gnd cell_6t
Xbit_r194_c199 bl_199 br_199 wl_194 vdd gnd cell_6t
Xbit_r195_c199 bl_199 br_199 wl_195 vdd gnd cell_6t
Xbit_r196_c199 bl_199 br_199 wl_196 vdd gnd cell_6t
Xbit_r197_c199 bl_199 br_199 wl_197 vdd gnd cell_6t
Xbit_r198_c199 bl_199 br_199 wl_198 vdd gnd cell_6t
Xbit_r199_c199 bl_199 br_199 wl_199 vdd gnd cell_6t
Xbit_r200_c199 bl_199 br_199 wl_200 vdd gnd cell_6t
Xbit_r201_c199 bl_199 br_199 wl_201 vdd gnd cell_6t
Xbit_r202_c199 bl_199 br_199 wl_202 vdd gnd cell_6t
Xbit_r203_c199 bl_199 br_199 wl_203 vdd gnd cell_6t
Xbit_r204_c199 bl_199 br_199 wl_204 vdd gnd cell_6t
Xbit_r205_c199 bl_199 br_199 wl_205 vdd gnd cell_6t
Xbit_r206_c199 bl_199 br_199 wl_206 vdd gnd cell_6t
Xbit_r207_c199 bl_199 br_199 wl_207 vdd gnd cell_6t
Xbit_r208_c199 bl_199 br_199 wl_208 vdd gnd cell_6t
Xbit_r209_c199 bl_199 br_199 wl_209 vdd gnd cell_6t
Xbit_r210_c199 bl_199 br_199 wl_210 vdd gnd cell_6t
Xbit_r211_c199 bl_199 br_199 wl_211 vdd gnd cell_6t
Xbit_r212_c199 bl_199 br_199 wl_212 vdd gnd cell_6t
Xbit_r213_c199 bl_199 br_199 wl_213 vdd gnd cell_6t
Xbit_r214_c199 bl_199 br_199 wl_214 vdd gnd cell_6t
Xbit_r215_c199 bl_199 br_199 wl_215 vdd gnd cell_6t
Xbit_r216_c199 bl_199 br_199 wl_216 vdd gnd cell_6t
Xbit_r217_c199 bl_199 br_199 wl_217 vdd gnd cell_6t
Xbit_r218_c199 bl_199 br_199 wl_218 vdd gnd cell_6t
Xbit_r219_c199 bl_199 br_199 wl_219 vdd gnd cell_6t
Xbit_r220_c199 bl_199 br_199 wl_220 vdd gnd cell_6t
Xbit_r221_c199 bl_199 br_199 wl_221 vdd gnd cell_6t
Xbit_r222_c199 bl_199 br_199 wl_222 vdd gnd cell_6t
Xbit_r223_c199 bl_199 br_199 wl_223 vdd gnd cell_6t
Xbit_r224_c199 bl_199 br_199 wl_224 vdd gnd cell_6t
Xbit_r225_c199 bl_199 br_199 wl_225 vdd gnd cell_6t
Xbit_r226_c199 bl_199 br_199 wl_226 vdd gnd cell_6t
Xbit_r227_c199 bl_199 br_199 wl_227 vdd gnd cell_6t
Xbit_r228_c199 bl_199 br_199 wl_228 vdd gnd cell_6t
Xbit_r229_c199 bl_199 br_199 wl_229 vdd gnd cell_6t
Xbit_r230_c199 bl_199 br_199 wl_230 vdd gnd cell_6t
Xbit_r231_c199 bl_199 br_199 wl_231 vdd gnd cell_6t
Xbit_r232_c199 bl_199 br_199 wl_232 vdd gnd cell_6t
Xbit_r233_c199 bl_199 br_199 wl_233 vdd gnd cell_6t
Xbit_r234_c199 bl_199 br_199 wl_234 vdd gnd cell_6t
Xbit_r235_c199 bl_199 br_199 wl_235 vdd gnd cell_6t
Xbit_r236_c199 bl_199 br_199 wl_236 vdd gnd cell_6t
Xbit_r237_c199 bl_199 br_199 wl_237 vdd gnd cell_6t
Xbit_r238_c199 bl_199 br_199 wl_238 vdd gnd cell_6t
Xbit_r239_c199 bl_199 br_199 wl_239 vdd gnd cell_6t
Xbit_r240_c199 bl_199 br_199 wl_240 vdd gnd cell_6t
Xbit_r241_c199 bl_199 br_199 wl_241 vdd gnd cell_6t
Xbit_r242_c199 bl_199 br_199 wl_242 vdd gnd cell_6t
Xbit_r243_c199 bl_199 br_199 wl_243 vdd gnd cell_6t
Xbit_r244_c199 bl_199 br_199 wl_244 vdd gnd cell_6t
Xbit_r245_c199 bl_199 br_199 wl_245 vdd gnd cell_6t
Xbit_r246_c199 bl_199 br_199 wl_246 vdd gnd cell_6t
Xbit_r247_c199 bl_199 br_199 wl_247 vdd gnd cell_6t
Xbit_r248_c199 bl_199 br_199 wl_248 vdd gnd cell_6t
Xbit_r249_c199 bl_199 br_199 wl_249 vdd gnd cell_6t
Xbit_r250_c199 bl_199 br_199 wl_250 vdd gnd cell_6t
Xbit_r251_c199 bl_199 br_199 wl_251 vdd gnd cell_6t
Xbit_r252_c199 bl_199 br_199 wl_252 vdd gnd cell_6t
Xbit_r253_c199 bl_199 br_199 wl_253 vdd gnd cell_6t
Xbit_r254_c199 bl_199 br_199 wl_254 vdd gnd cell_6t
Xbit_r255_c199 bl_199 br_199 wl_255 vdd gnd cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd cell_6t
Xbit_r1_c200 bl_200 br_200 wl_1 vdd gnd cell_6t
Xbit_r2_c200 bl_200 br_200 wl_2 vdd gnd cell_6t
Xbit_r3_c200 bl_200 br_200 wl_3 vdd gnd cell_6t
Xbit_r4_c200 bl_200 br_200 wl_4 vdd gnd cell_6t
Xbit_r5_c200 bl_200 br_200 wl_5 vdd gnd cell_6t
Xbit_r6_c200 bl_200 br_200 wl_6 vdd gnd cell_6t
Xbit_r7_c200 bl_200 br_200 wl_7 vdd gnd cell_6t
Xbit_r8_c200 bl_200 br_200 wl_8 vdd gnd cell_6t
Xbit_r9_c200 bl_200 br_200 wl_9 vdd gnd cell_6t
Xbit_r10_c200 bl_200 br_200 wl_10 vdd gnd cell_6t
Xbit_r11_c200 bl_200 br_200 wl_11 vdd gnd cell_6t
Xbit_r12_c200 bl_200 br_200 wl_12 vdd gnd cell_6t
Xbit_r13_c200 bl_200 br_200 wl_13 vdd gnd cell_6t
Xbit_r14_c200 bl_200 br_200 wl_14 vdd gnd cell_6t
Xbit_r15_c200 bl_200 br_200 wl_15 vdd gnd cell_6t
Xbit_r16_c200 bl_200 br_200 wl_16 vdd gnd cell_6t
Xbit_r17_c200 bl_200 br_200 wl_17 vdd gnd cell_6t
Xbit_r18_c200 bl_200 br_200 wl_18 vdd gnd cell_6t
Xbit_r19_c200 bl_200 br_200 wl_19 vdd gnd cell_6t
Xbit_r20_c200 bl_200 br_200 wl_20 vdd gnd cell_6t
Xbit_r21_c200 bl_200 br_200 wl_21 vdd gnd cell_6t
Xbit_r22_c200 bl_200 br_200 wl_22 vdd gnd cell_6t
Xbit_r23_c200 bl_200 br_200 wl_23 vdd gnd cell_6t
Xbit_r24_c200 bl_200 br_200 wl_24 vdd gnd cell_6t
Xbit_r25_c200 bl_200 br_200 wl_25 vdd gnd cell_6t
Xbit_r26_c200 bl_200 br_200 wl_26 vdd gnd cell_6t
Xbit_r27_c200 bl_200 br_200 wl_27 vdd gnd cell_6t
Xbit_r28_c200 bl_200 br_200 wl_28 vdd gnd cell_6t
Xbit_r29_c200 bl_200 br_200 wl_29 vdd gnd cell_6t
Xbit_r30_c200 bl_200 br_200 wl_30 vdd gnd cell_6t
Xbit_r31_c200 bl_200 br_200 wl_31 vdd gnd cell_6t
Xbit_r32_c200 bl_200 br_200 wl_32 vdd gnd cell_6t
Xbit_r33_c200 bl_200 br_200 wl_33 vdd gnd cell_6t
Xbit_r34_c200 bl_200 br_200 wl_34 vdd gnd cell_6t
Xbit_r35_c200 bl_200 br_200 wl_35 vdd gnd cell_6t
Xbit_r36_c200 bl_200 br_200 wl_36 vdd gnd cell_6t
Xbit_r37_c200 bl_200 br_200 wl_37 vdd gnd cell_6t
Xbit_r38_c200 bl_200 br_200 wl_38 vdd gnd cell_6t
Xbit_r39_c200 bl_200 br_200 wl_39 vdd gnd cell_6t
Xbit_r40_c200 bl_200 br_200 wl_40 vdd gnd cell_6t
Xbit_r41_c200 bl_200 br_200 wl_41 vdd gnd cell_6t
Xbit_r42_c200 bl_200 br_200 wl_42 vdd gnd cell_6t
Xbit_r43_c200 bl_200 br_200 wl_43 vdd gnd cell_6t
Xbit_r44_c200 bl_200 br_200 wl_44 vdd gnd cell_6t
Xbit_r45_c200 bl_200 br_200 wl_45 vdd gnd cell_6t
Xbit_r46_c200 bl_200 br_200 wl_46 vdd gnd cell_6t
Xbit_r47_c200 bl_200 br_200 wl_47 vdd gnd cell_6t
Xbit_r48_c200 bl_200 br_200 wl_48 vdd gnd cell_6t
Xbit_r49_c200 bl_200 br_200 wl_49 vdd gnd cell_6t
Xbit_r50_c200 bl_200 br_200 wl_50 vdd gnd cell_6t
Xbit_r51_c200 bl_200 br_200 wl_51 vdd gnd cell_6t
Xbit_r52_c200 bl_200 br_200 wl_52 vdd gnd cell_6t
Xbit_r53_c200 bl_200 br_200 wl_53 vdd gnd cell_6t
Xbit_r54_c200 bl_200 br_200 wl_54 vdd gnd cell_6t
Xbit_r55_c200 bl_200 br_200 wl_55 vdd gnd cell_6t
Xbit_r56_c200 bl_200 br_200 wl_56 vdd gnd cell_6t
Xbit_r57_c200 bl_200 br_200 wl_57 vdd gnd cell_6t
Xbit_r58_c200 bl_200 br_200 wl_58 vdd gnd cell_6t
Xbit_r59_c200 bl_200 br_200 wl_59 vdd gnd cell_6t
Xbit_r60_c200 bl_200 br_200 wl_60 vdd gnd cell_6t
Xbit_r61_c200 bl_200 br_200 wl_61 vdd gnd cell_6t
Xbit_r62_c200 bl_200 br_200 wl_62 vdd gnd cell_6t
Xbit_r63_c200 bl_200 br_200 wl_63 vdd gnd cell_6t
Xbit_r64_c200 bl_200 br_200 wl_64 vdd gnd cell_6t
Xbit_r65_c200 bl_200 br_200 wl_65 vdd gnd cell_6t
Xbit_r66_c200 bl_200 br_200 wl_66 vdd gnd cell_6t
Xbit_r67_c200 bl_200 br_200 wl_67 vdd gnd cell_6t
Xbit_r68_c200 bl_200 br_200 wl_68 vdd gnd cell_6t
Xbit_r69_c200 bl_200 br_200 wl_69 vdd gnd cell_6t
Xbit_r70_c200 bl_200 br_200 wl_70 vdd gnd cell_6t
Xbit_r71_c200 bl_200 br_200 wl_71 vdd gnd cell_6t
Xbit_r72_c200 bl_200 br_200 wl_72 vdd gnd cell_6t
Xbit_r73_c200 bl_200 br_200 wl_73 vdd gnd cell_6t
Xbit_r74_c200 bl_200 br_200 wl_74 vdd gnd cell_6t
Xbit_r75_c200 bl_200 br_200 wl_75 vdd gnd cell_6t
Xbit_r76_c200 bl_200 br_200 wl_76 vdd gnd cell_6t
Xbit_r77_c200 bl_200 br_200 wl_77 vdd gnd cell_6t
Xbit_r78_c200 bl_200 br_200 wl_78 vdd gnd cell_6t
Xbit_r79_c200 bl_200 br_200 wl_79 vdd gnd cell_6t
Xbit_r80_c200 bl_200 br_200 wl_80 vdd gnd cell_6t
Xbit_r81_c200 bl_200 br_200 wl_81 vdd gnd cell_6t
Xbit_r82_c200 bl_200 br_200 wl_82 vdd gnd cell_6t
Xbit_r83_c200 bl_200 br_200 wl_83 vdd gnd cell_6t
Xbit_r84_c200 bl_200 br_200 wl_84 vdd gnd cell_6t
Xbit_r85_c200 bl_200 br_200 wl_85 vdd gnd cell_6t
Xbit_r86_c200 bl_200 br_200 wl_86 vdd gnd cell_6t
Xbit_r87_c200 bl_200 br_200 wl_87 vdd gnd cell_6t
Xbit_r88_c200 bl_200 br_200 wl_88 vdd gnd cell_6t
Xbit_r89_c200 bl_200 br_200 wl_89 vdd gnd cell_6t
Xbit_r90_c200 bl_200 br_200 wl_90 vdd gnd cell_6t
Xbit_r91_c200 bl_200 br_200 wl_91 vdd gnd cell_6t
Xbit_r92_c200 bl_200 br_200 wl_92 vdd gnd cell_6t
Xbit_r93_c200 bl_200 br_200 wl_93 vdd gnd cell_6t
Xbit_r94_c200 bl_200 br_200 wl_94 vdd gnd cell_6t
Xbit_r95_c200 bl_200 br_200 wl_95 vdd gnd cell_6t
Xbit_r96_c200 bl_200 br_200 wl_96 vdd gnd cell_6t
Xbit_r97_c200 bl_200 br_200 wl_97 vdd gnd cell_6t
Xbit_r98_c200 bl_200 br_200 wl_98 vdd gnd cell_6t
Xbit_r99_c200 bl_200 br_200 wl_99 vdd gnd cell_6t
Xbit_r100_c200 bl_200 br_200 wl_100 vdd gnd cell_6t
Xbit_r101_c200 bl_200 br_200 wl_101 vdd gnd cell_6t
Xbit_r102_c200 bl_200 br_200 wl_102 vdd gnd cell_6t
Xbit_r103_c200 bl_200 br_200 wl_103 vdd gnd cell_6t
Xbit_r104_c200 bl_200 br_200 wl_104 vdd gnd cell_6t
Xbit_r105_c200 bl_200 br_200 wl_105 vdd gnd cell_6t
Xbit_r106_c200 bl_200 br_200 wl_106 vdd gnd cell_6t
Xbit_r107_c200 bl_200 br_200 wl_107 vdd gnd cell_6t
Xbit_r108_c200 bl_200 br_200 wl_108 vdd gnd cell_6t
Xbit_r109_c200 bl_200 br_200 wl_109 vdd gnd cell_6t
Xbit_r110_c200 bl_200 br_200 wl_110 vdd gnd cell_6t
Xbit_r111_c200 bl_200 br_200 wl_111 vdd gnd cell_6t
Xbit_r112_c200 bl_200 br_200 wl_112 vdd gnd cell_6t
Xbit_r113_c200 bl_200 br_200 wl_113 vdd gnd cell_6t
Xbit_r114_c200 bl_200 br_200 wl_114 vdd gnd cell_6t
Xbit_r115_c200 bl_200 br_200 wl_115 vdd gnd cell_6t
Xbit_r116_c200 bl_200 br_200 wl_116 vdd gnd cell_6t
Xbit_r117_c200 bl_200 br_200 wl_117 vdd gnd cell_6t
Xbit_r118_c200 bl_200 br_200 wl_118 vdd gnd cell_6t
Xbit_r119_c200 bl_200 br_200 wl_119 vdd gnd cell_6t
Xbit_r120_c200 bl_200 br_200 wl_120 vdd gnd cell_6t
Xbit_r121_c200 bl_200 br_200 wl_121 vdd gnd cell_6t
Xbit_r122_c200 bl_200 br_200 wl_122 vdd gnd cell_6t
Xbit_r123_c200 bl_200 br_200 wl_123 vdd gnd cell_6t
Xbit_r124_c200 bl_200 br_200 wl_124 vdd gnd cell_6t
Xbit_r125_c200 bl_200 br_200 wl_125 vdd gnd cell_6t
Xbit_r126_c200 bl_200 br_200 wl_126 vdd gnd cell_6t
Xbit_r127_c200 bl_200 br_200 wl_127 vdd gnd cell_6t
Xbit_r128_c200 bl_200 br_200 wl_128 vdd gnd cell_6t
Xbit_r129_c200 bl_200 br_200 wl_129 vdd gnd cell_6t
Xbit_r130_c200 bl_200 br_200 wl_130 vdd gnd cell_6t
Xbit_r131_c200 bl_200 br_200 wl_131 vdd gnd cell_6t
Xbit_r132_c200 bl_200 br_200 wl_132 vdd gnd cell_6t
Xbit_r133_c200 bl_200 br_200 wl_133 vdd gnd cell_6t
Xbit_r134_c200 bl_200 br_200 wl_134 vdd gnd cell_6t
Xbit_r135_c200 bl_200 br_200 wl_135 vdd gnd cell_6t
Xbit_r136_c200 bl_200 br_200 wl_136 vdd gnd cell_6t
Xbit_r137_c200 bl_200 br_200 wl_137 vdd gnd cell_6t
Xbit_r138_c200 bl_200 br_200 wl_138 vdd gnd cell_6t
Xbit_r139_c200 bl_200 br_200 wl_139 vdd gnd cell_6t
Xbit_r140_c200 bl_200 br_200 wl_140 vdd gnd cell_6t
Xbit_r141_c200 bl_200 br_200 wl_141 vdd gnd cell_6t
Xbit_r142_c200 bl_200 br_200 wl_142 vdd gnd cell_6t
Xbit_r143_c200 bl_200 br_200 wl_143 vdd gnd cell_6t
Xbit_r144_c200 bl_200 br_200 wl_144 vdd gnd cell_6t
Xbit_r145_c200 bl_200 br_200 wl_145 vdd gnd cell_6t
Xbit_r146_c200 bl_200 br_200 wl_146 vdd gnd cell_6t
Xbit_r147_c200 bl_200 br_200 wl_147 vdd gnd cell_6t
Xbit_r148_c200 bl_200 br_200 wl_148 vdd gnd cell_6t
Xbit_r149_c200 bl_200 br_200 wl_149 vdd gnd cell_6t
Xbit_r150_c200 bl_200 br_200 wl_150 vdd gnd cell_6t
Xbit_r151_c200 bl_200 br_200 wl_151 vdd gnd cell_6t
Xbit_r152_c200 bl_200 br_200 wl_152 vdd gnd cell_6t
Xbit_r153_c200 bl_200 br_200 wl_153 vdd gnd cell_6t
Xbit_r154_c200 bl_200 br_200 wl_154 vdd gnd cell_6t
Xbit_r155_c200 bl_200 br_200 wl_155 vdd gnd cell_6t
Xbit_r156_c200 bl_200 br_200 wl_156 vdd gnd cell_6t
Xbit_r157_c200 bl_200 br_200 wl_157 vdd gnd cell_6t
Xbit_r158_c200 bl_200 br_200 wl_158 vdd gnd cell_6t
Xbit_r159_c200 bl_200 br_200 wl_159 vdd gnd cell_6t
Xbit_r160_c200 bl_200 br_200 wl_160 vdd gnd cell_6t
Xbit_r161_c200 bl_200 br_200 wl_161 vdd gnd cell_6t
Xbit_r162_c200 bl_200 br_200 wl_162 vdd gnd cell_6t
Xbit_r163_c200 bl_200 br_200 wl_163 vdd gnd cell_6t
Xbit_r164_c200 bl_200 br_200 wl_164 vdd gnd cell_6t
Xbit_r165_c200 bl_200 br_200 wl_165 vdd gnd cell_6t
Xbit_r166_c200 bl_200 br_200 wl_166 vdd gnd cell_6t
Xbit_r167_c200 bl_200 br_200 wl_167 vdd gnd cell_6t
Xbit_r168_c200 bl_200 br_200 wl_168 vdd gnd cell_6t
Xbit_r169_c200 bl_200 br_200 wl_169 vdd gnd cell_6t
Xbit_r170_c200 bl_200 br_200 wl_170 vdd gnd cell_6t
Xbit_r171_c200 bl_200 br_200 wl_171 vdd gnd cell_6t
Xbit_r172_c200 bl_200 br_200 wl_172 vdd gnd cell_6t
Xbit_r173_c200 bl_200 br_200 wl_173 vdd gnd cell_6t
Xbit_r174_c200 bl_200 br_200 wl_174 vdd gnd cell_6t
Xbit_r175_c200 bl_200 br_200 wl_175 vdd gnd cell_6t
Xbit_r176_c200 bl_200 br_200 wl_176 vdd gnd cell_6t
Xbit_r177_c200 bl_200 br_200 wl_177 vdd gnd cell_6t
Xbit_r178_c200 bl_200 br_200 wl_178 vdd gnd cell_6t
Xbit_r179_c200 bl_200 br_200 wl_179 vdd gnd cell_6t
Xbit_r180_c200 bl_200 br_200 wl_180 vdd gnd cell_6t
Xbit_r181_c200 bl_200 br_200 wl_181 vdd gnd cell_6t
Xbit_r182_c200 bl_200 br_200 wl_182 vdd gnd cell_6t
Xbit_r183_c200 bl_200 br_200 wl_183 vdd gnd cell_6t
Xbit_r184_c200 bl_200 br_200 wl_184 vdd gnd cell_6t
Xbit_r185_c200 bl_200 br_200 wl_185 vdd gnd cell_6t
Xbit_r186_c200 bl_200 br_200 wl_186 vdd gnd cell_6t
Xbit_r187_c200 bl_200 br_200 wl_187 vdd gnd cell_6t
Xbit_r188_c200 bl_200 br_200 wl_188 vdd gnd cell_6t
Xbit_r189_c200 bl_200 br_200 wl_189 vdd gnd cell_6t
Xbit_r190_c200 bl_200 br_200 wl_190 vdd gnd cell_6t
Xbit_r191_c200 bl_200 br_200 wl_191 vdd gnd cell_6t
Xbit_r192_c200 bl_200 br_200 wl_192 vdd gnd cell_6t
Xbit_r193_c200 bl_200 br_200 wl_193 vdd gnd cell_6t
Xbit_r194_c200 bl_200 br_200 wl_194 vdd gnd cell_6t
Xbit_r195_c200 bl_200 br_200 wl_195 vdd gnd cell_6t
Xbit_r196_c200 bl_200 br_200 wl_196 vdd gnd cell_6t
Xbit_r197_c200 bl_200 br_200 wl_197 vdd gnd cell_6t
Xbit_r198_c200 bl_200 br_200 wl_198 vdd gnd cell_6t
Xbit_r199_c200 bl_200 br_200 wl_199 vdd gnd cell_6t
Xbit_r200_c200 bl_200 br_200 wl_200 vdd gnd cell_6t
Xbit_r201_c200 bl_200 br_200 wl_201 vdd gnd cell_6t
Xbit_r202_c200 bl_200 br_200 wl_202 vdd gnd cell_6t
Xbit_r203_c200 bl_200 br_200 wl_203 vdd gnd cell_6t
Xbit_r204_c200 bl_200 br_200 wl_204 vdd gnd cell_6t
Xbit_r205_c200 bl_200 br_200 wl_205 vdd gnd cell_6t
Xbit_r206_c200 bl_200 br_200 wl_206 vdd gnd cell_6t
Xbit_r207_c200 bl_200 br_200 wl_207 vdd gnd cell_6t
Xbit_r208_c200 bl_200 br_200 wl_208 vdd gnd cell_6t
Xbit_r209_c200 bl_200 br_200 wl_209 vdd gnd cell_6t
Xbit_r210_c200 bl_200 br_200 wl_210 vdd gnd cell_6t
Xbit_r211_c200 bl_200 br_200 wl_211 vdd gnd cell_6t
Xbit_r212_c200 bl_200 br_200 wl_212 vdd gnd cell_6t
Xbit_r213_c200 bl_200 br_200 wl_213 vdd gnd cell_6t
Xbit_r214_c200 bl_200 br_200 wl_214 vdd gnd cell_6t
Xbit_r215_c200 bl_200 br_200 wl_215 vdd gnd cell_6t
Xbit_r216_c200 bl_200 br_200 wl_216 vdd gnd cell_6t
Xbit_r217_c200 bl_200 br_200 wl_217 vdd gnd cell_6t
Xbit_r218_c200 bl_200 br_200 wl_218 vdd gnd cell_6t
Xbit_r219_c200 bl_200 br_200 wl_219 vdd gnd cell_6t
Xbit_r220_c200 bl_200 br_200 wl_220 vdd gnd cell_6t
Xbit_r221_c200 bl_200 br_200 wl_221 vdd gnd cell_6t
Xbit_r222_c200 bl_200 br_200 wl_222 vdd gnd cell_6t
Xbit_r223_c200 bl_200 br_200 wl_223 vdd gnd cell_6t
Xbit_r224_c200 bl_200 br_200 wl_224 vdd gnd cell_6t
Xbit_r225_c200 bl_200 br_200 wl_225 vdd gnd cell_6t
Xbit_r226_c200 bl_200 br_200 wl_226 vdd gnd cell_6t
Xbit_r227_c200 bl_200 br_200 wl_227 vdd gnd cell_6t
Xbit_r228_c200 bl_200 br_200 wl_228 vdd gnd cell_6t
Xbit_r229_c200 bl_200 br_200 wl_229 vdd gnd cell_6t
Xbit_r230_c200 bl_200 br_200 wl_230 vdd gnd cell_6t
Xbit_r231_c200 bl_200 br_200 wl_231 vdd gnd cell_6t
Xbit_r232_c200 bl_200 br_200 wl_232 vdd gnd cell_6t
Xbit_r233_c200 bl_200 br_200 wl_233 vdd gnd cell_6t
Xbit_r234_c200 bl_200 br_200 wl_234 vdd gnd cell_6t
Xbit_r235_c200 bl_200 br_200 wl_235 vdd gnd cell_6t
Xbit_r236_c200 bl_200 br_200 wl_236 vdd gnd cell_6t
Xbit_r237_c200 bl_200 br_200 wl_237 vdd gnd cell_6t
Xbit_r238_c200 bl_200 br_200 wl_238 vdd gnd cell_6t
Xbit_r239_c200 bl_200 br_200 wl_239 vdd gnd cell_6t
Xbit_r240_c200 bl_200 br_200 wl_240 vdd gnd cell_6t
Xbit_r241_c200 bl_200 br_200 wl_241 vdd gnd cell_6t
Xbit_r242_c200 bl_200 br_200 wl_242 vdd gnd cell_6t
Xbit_r243_c200 bl_200 br_200 wl_243 vdd gnd cell_6t
Xbit_r244_c200 bl_200 br_200 wl_244 vdd gnd cell_6t
Xbit_r245_c200 bl_200 br_200 wl_245 vdd gnd cell_6t
Xbit_r246_c200 bl_200 br_200 wl_246 vdd gnd cell_6t
Xbit_r247_c200 bl_200 br_200 wl_247 vdd gnd cell_6t
Xbit_r248_c200 bl_200 br_200 wl_248 vdd gnd cell_6t
Xbit_r249_c200 bl_200 br_200 wl_249 vdd gnd cell_6t
Xbit_r250_c200 bl_200 br_200 wl_250 vdd gnd cell_6t
Xbit_r251_c200 bl_200 br_200 wl_251 vdd gnd cell_6t
Xbit_r252_c200 bl_200 br_200 wl_252 vdd gnd cell_6t
Xbit_r253_c200 bl_200 br_200 wl_253 vdd gnd cell_6t
Xbit_r254_c200 bl_200 br_200 wl_254 vdd gnd cell_6t
Xbit_r255_c200 bl_200 br_200 wl_255 vdd gnd cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd cell_6t
Xbit_r1_c201 bl_201 br_201 wl_1 vdd gnd cell_6t
Xbit_r2_c201 bl_201 br_201 wl_2 vdd gnd cell_6t
Xbit_r3_c201 bl_201 br_201 wl_3 vdd gnd cell_6t
Xbit_r4_c201 bl_201 br_201 wl_4 vdd gnd cell_6t
Xbit_r5_c201 bl_201 br_201 wl_5 vdd gnd cell_6t
Xbit_r6_c201 bl_201 br_201 wl_6 vdd gnd cell_6t
Xbit_r7_c201 bl_201 br_201 wl_7 vdd gnd cell_6t
Xbit_r8_c201 bl_201 br_201 wl_8 vdd gnd cell_6t
Xbit_r9_c201 bl_201 br_201 wl_9 vdd gnd cell_6t
Xbit_r10_c201 bl_201 br_201 wl_10 vdd gnd cell_6t
Xbit_r11_c201 bl_201 br_201 wl_11 vdd gnd cell_6t
Xbit_r12_c201 bl_201 br_201 wl_12 vdd gnd cell_6t
Xbit_r13_c201 bl_201 br_201 wl_13 vdd gnd cell_6t
Xbit_r14_c201 bl_201 br_201 wl_14 vdd gnd cell_6t
Xbit_r15_c201 bl_201 br_201 wl_15 vdd gnd cell_6t
Xbit_r16_c201 bl_201 br_201 wl_16 vdd gnd cell_6t
Xbit_r17_c201 bl_201 br_201 wl_17 vdd gnd cell_6t
Xbit_r18_c201 bl_201 br_201 wl_18 vdd gnd cell_6t
Xbit_r19_c201 bl_201 br_201 wl_19 vdd gnd cell_6t
Xbit_r20_c201 bl_201 br_201 wl_20 vdd gnd cell_6t
Xbit_r21_c201 bl_201 br_201 wl_21 vdd gnd cell_6t
Xbit_r22_c201 bl_201 br_201 wl_22 vdd gnd cell_6t
Xbit_r23_c201 bl_201 br_201 wl_23 vdd gnd cell_6t
Xbit_r24_c201 bl_201 br_201 wl_24 vdd gnd cell_6t
Xbit_r25_c201 bl_201 br_201 wl_25 vdd gnd cell_6t
Xbit_r26_c201 bl_201 br_201 wl_26 vdd gnd cell_6t
Xbit_r27_c201 bl_201 br_201 wl_27 vdd gnd cell_6t
Xbit_r28_c201 bl_201 br_201 wl_28 vdd gnd cell_6t
Xbit_r29_c201 bl_201 br_201 wl_29 vdd gnd cell_6t
Xbit_r30_c201 bl_201 br_201 wl_30 vdd gnd cell_6t
Xbit_r31_c201 bl_201 br_201 wl_31 vdd gnd cell_6t
Xbit_r32_c201 bl_201 br_201 wl_32 vdd gnd cell_6t
Xbit_r33_c201 bl_201 br_201 wl_33 vdd gnd cell_6t
Xbit_r34_c201 bl_201 br_201 wl_34 vdd gnd cell_6t
Xbit_r35_c201 bl_201 br_201 wl_35 vdd gnd cell_6t
Xbit_r36_c201 bl_201 br_201 wl_36 vdd gnd cell_6t
Xbit_r37_c201 bl_201 br_201 wl_37 vdd gnd cell_6t
Xbit_r38_c201 bl_201 br_201 wl_38 vdd gnd cell_6t
Xbit_r39_c201 bl_201 br_201 wl_39 vdd gnd cell_6t
Xbit_r40_c201 bl_201 br_201 wl_40 vdd gnd cell_6t
Xbit_r41_c201 bl_201 br_201 wl_41 vdd gnd cell_6t
Xbit_r42_c201 bl_201 br_201 wl_42 vdd gnd cell_6t
Xbit_r43_c201 bl_201 br_201 wl_43 vdd gnd cell_6t
Xbit_r44_c201 bl_201 br_201 wl_44 vdd gnd cell_6t
Xbit_r45_c201 bl_201 br_201 wl_45 vdd gnd cell_6t
Xbit_r46_c201 bl_201 br_201 wl_46 vdd gnd cell_6t
Xbit_r47_c201 bl_201 br_201 wl_47 vdd gnd cell_6t
Xbit_r48_c201 bl_201 br_201 wl_48 vdd gnd cell_6t
Xbit_r49_c201 bl_201 br_201 wl_49 vdd gnd cell_6t
Xbit_r50_c201 bl_201 br_201 wl_50 vdd gnd cell_6t
Xbit_r51_c201 bl_201 br_201 wl_51 vdd gnd cell_6t
Xbit_r52_c201 bl_201 br_201 wl_52 vdd gnd cell_6t
Xbit_r53_c201 bl_201 br_201 wl_53 vdd gnd cell_6t
Xbit_r54_c201 bl_201 br_201 wl_54 vdd gnd cell_6t
Xbit_r55_c201 bl_201 br_201 wl_55 vdd gnd cell_6t
Xbit_r56_c201 bl_201 br_201 wl_56 vdd gnd cell_6t
Xbit_r57_c201 bl_201 br_201 wl_57 vdd gnd cell_6t
Xbit_r58_c201 bl_201 br_201 wl_58 vdd gnd cell_6t
Xbit_r59_c201 bl_201 br_201 wl_59 vdd gnd cell_6t
Xbit_r60_c201 bl_201 br_201 wl_60 vdd gnd cell_6t
Xbit_r61_c201 bl_201 br_201 wl_61 vdd gnd cell_6t
Xbit_r62_c201 bl_201 br_201 wl_62 vdd gnd cell_6t
Xbit_r63_c201 bl_201 br_201 wl_63 vdd gnd cell_6t
Xbit_r64_c201 bl_201 br_201 wl_64 vdd gnd cell_6t
Xbit_r65_c201 bl_201 br_201 wl_65 vdd gnd cell_6t
Xbit_r66_c201 bl_201 br_201 wl_66 vdd gnd cell_6t
Xbit_r67_c201 bl_201 br_201 wl_67 vdd gnd cell_6t
Xbit_r68_c201 bl_201 br_201 wl_68 vdd gnd cell_6t
Xbit_r69_c201 bl_201 br_201 wl_69 vdd gnd cell_6t
Xbit_r70_c201 bl_201 br_201 wl_70 vdd gnd cell_6t
Xbit_r71_c201 bl_201 br_201 wl_71 vdd gnd cell_6t
Xbit_r72_c201 bl_201 br_201 wl_72 vdd gnd cell_6t
Xbit_r73_c201 bl_201 br_201 wl_73 vdd gnd cell_6t
Xbit_r74_c201 bl_201 br_201 wl_74 vdd gnd cell_6t
Xbit_r75_c201 bl_201 br_201 wl_75 vdd gnd cell_6t
Xbit_r76_c201 bl_201 br_201 wl_76 vdd gnd cell_6t
Xbit_r77_c201 bl_201 br_201 wl_77 vdd gnd cell_6t
Xbit_r78_c201 bl_201 br_201 wl_78 vdd gnd cell_6t
Xbit_r79_c201 bl_201 br_201 wl_79 vdd gnd cell_6t
Xbit_r80_c201 bl_201 br_201 wl_80 vdd gnd cell_6t
Xbit_r81_c201 bl_201 br_201 wl_81 vdd gnd cell_6t
Xbit_r82_c201 bl_201 br_201 wl_82 vdd gnd cell_6t
Xbit_r83_c201 bl_201 br_201 wl_83 vdd gnd cell_6t
Xbit_r84_c201 bl_201 br_201 wl_84 vdd gnd cell_6t
Xbit_r85_c201 bl_201 br_201 wl_85 vdd gnd cell_6t
Xbit_r86_c201 bl_201 br_201 wl_86 vdd gnd cell_6t
Xbit_r87_c201 bl_201 br_201 wl_87 vdd gnd cell_6t
Xbit_r88_c201 bl_201 br_201 wl_88 vdd gnd cell_6t
Xbit_r89_c201 bl_201 br_201 wl_89 vdd gnd cell_6t
Xbit_r90_c201 bl_201 br_201 wl_90 vdd gnd cell_6t
Xbit_r91_c201 bl_201 br_201 wl_91 vdd gnd cell_6t
Xbit_r92_c201 bl_201 br_201 wl_92 vdd gnd cell_6t
Xbit_r93_c201 bl_201 br_201 wl_93 vdd gnd cell_6t
Xbit_r94_c201 bl_201 br_201 wl_94 vdd gnd cell_6t
Xbit_r95_c201 bl_201 br_201 wl_95 vdd gnd cell_6t
Xbit_r96_c201 bl_201 br_201 wl_96 vdd gnd cell_6t
Xbit_r97_c201 bl_201 br_201 wl_97 vdd gnd cell_6t
Xbit_r98_c201 bl_201 br_201 wl_98 vdd gnd cell_6t
Xbit_r99_c201 bl_201 br_201 wl_99 vdd gnd cell_6t
Xbit_r100_c201 bl_201 br_201 wl_100 vdd gnd cell_6t
Xbit_r101_c201 bl_201 br_201 wl_101 vdd gnd cell_6t
Xbit_r102_c201 bl_201 br_201 wl_102 vdd gnd cell_6t
Xbit_r103_c201 bl_201 br_201 wl_103 vdd gnd cell_6t
Xbit_r104_c201 bl_201 br_201 wl_104 vdd gnd cell_6t
Xbit_r105_c201 bl_201 br_201 wl_105 vdd gnd cell_6t
Xbit_r106_c201 bl_201 br_201 wl_106 vdd gnd cell_6t
Xbit_r107_c201 bl_201 br_201 wl_107 vdd gnd cell_6t
Xbit_r108_c201 bl_201 br_201 wl_108 vdd gnd cell_6t
Xbit_r109_c201 bl_201 br_201 wl_109 vdd gnd cell_6t
Xbit_r110_c201 bl_201 br_201 wl_110 vdd gnd cell_6t
Xbit_r111_c201 bl_201 br_201 wl_111 vdd gnd cell_6t
Xbit_r112_c201 bl_201 br_201 wl_112 vdd gnd cell_6t
Xbit_r113_c201 bl_201 br_201 wl_113 vdd gnd cell_6t
Xbit_r114_c201 bl_201 br_201 wl_114 vdd gnd cell_6t
Xbit_r115_c201 bl_201 br_201 wl_115 vdd gnd cell_6t
Xbit_r116_c201 bl_201 br_201 wl_116 vdd gnd cell_6t
Xbit_r117_c201 bl_201 br_201 wl_117 vdd gnd cell_6t
Xbit_r118_c201 bl_201 br_201 wl_118 vdd gnd cell_6t
Xbit_r119_c201 bl_201 br_201 wl_119 vdd gnd cell_6t
Xbit_r120_c201 bl_201 br_201 wl_120 vdd gnd cell_6t
Xbit_r121_c201 bl_201 br_201 wl_121 vdd gnd cell_6t
Xbit_r122_c201 bl_201 br_201 wl_122 vdd gnd cell_6t
Xbit_r123_c201 bl_201 br_201 wl_123 vdd gnd cell_6t
Xbit_r124_c201 bl_201 br_201 wl_124 vdd gnd cell_6t
Xbit_r125_c201 bl_201 br_201 wl_125 vdd gnd cell_6t
Xbit_r126_c201 bl_201 br_201 wl_126 vdd gnd cell_6t
Xbit_r127_c201 bl_201 br_201 wl_127 vdd gnd cell_6t
Xbit_r128_c201 bl_201 br_201 wl_128 vdd gnd cell_6t
Xbit_r129_c201 bl_201 br_201 wl_129 vdd gnd cell_6t
Xbit_r130_c201 bl_201 br_201 wl_130 vdd gnd cell_6t
Xbit_r131_c201 bl_201 br_201 wl_131 vdd gnd cell_6t
Xbit_r132_c201 bl_201 br_201 wl_132 vdd gnd cell_6t
Xbit_r133_c201 bl_201 br_201 wl_133 vdd gnd cell_6t
Xbit_r134_c201 bl_201 br_201 wl_134 vdd gnd cell_6t
Xbit_r135_c201 bl_201 br_201 wl_135 vdd gnd cell_6t
Xbit_r136_c201 bl_201 br_201 wl_136 vdd gnd cell_6t
Xbit_r137_c201 bl_201 br_201 wl_137 vdd gnd cell_6t
Xbit_r138_c201 bl_201 br_201 wl_138 vdd gnd cell_6t
Xbit_r139_c201 bl_201 br_201 wl_139 vdd gnd cell_6t
Xbit_r140_c201 bl_201 br_201 wl_140 vdd gnd cell_6t
Xbit_r141_c201 bl_201 br_201 wl_141 vdd gnd cell_6t
Xbit_r142_c201 bl_201 br_201 wl_142 vdd gnd cell_6t
Xbit_r143_c201 bl_201 br_201 wl_143 vdd gnd cell_6t
Xbit_r144_c201 bl_201 br_201 wl_144 vdd gnd cell_6t
Xbit_r145_c201 bl_201 br_201 wl_145 vdd gnd cell_6t
Xbit_r146_c201 bl_201 br_201 wl_146 vdd gnd cell_6t
Xbit_r147_c201 bl_201 br_201 wl_147 vdd gnd cell_6t
Xbit_r148_c201 bl_201 br_201 wl_148 vdd gnd cell_6t
Xbit_r149_c201 bl_201 br_201 wl_149 vdd gnd cell_6t
Xbit_r150_c201 bl_201 br_201 wl_150 vdd gnd cell_6t
Xbit_r151_c201 bl_201 br_201 wl_151 vdd gnd cell_6t
Xbit_r152_c201 bl_201 br_201 wl_152 vdd gnd cell_6t
Xbit_r153_c201 bl_201 br_201 wl_153 vdd gnd cell_6t
Xbit_r154_c201 bl_201 br_201 wl_154 vdd gnd cell_6t
Xbit_r155_c201 bl_201 br_201 wl_155 vdd gnd cell_6t
Xbit_r156_c201 bl_201 br_201 wl_156 vdd gnd cell_6t
Xbit_r157_c201 bl_201 br_201 wl_157 vdd gnd cell_6t
Xbit_r158_c201 bl_201 br_201 wl_158 vdd gnd cell_6t
Xbit_r159_c201 bl_201 br_201 wl_159 vdd gnd cell_6t
Xbit_r160_c201 bl_201 br_201 wl_160 vdd gnd cell_6t
Xbit_r161_c201 bl_201 br_201 wl_161 vdd gnd cell_6t
Xbit_r162_c201 bl_201 br_201 wl_162 vdd gnd cell_6t
Xbit_r163_c201 bl_201 br_201 wl_163 vdd gnd cell_6t
Xbit_r164_c201 bl_201 br_201 wl_164 vdd gnd cell_6t
Xbit_r165_c201 bl_201 br_201 wl_165 vdd gnd cell_6t
Xbit_r166_c201 bl_201 br_201 wl_166 vdd gnd cell_6t
Xbit_r167_c201 bl_201 br_201 wl_167 vdd gnd cell_6t
Xbit_r168_c201 bl_201 br_201 wl_168 vdd gnd cell_6t
Xbit_r169_c201 bl_201 br_201 wl_169 vdd gnd cell_6t
Xbit_r170_c201 bl_201 br_201 wl_170 vdd gnd cell_6t
Xbit_r171_c201 bl_201 br_201 wl_171 vdd gnd cell_6t
Xbit_r172_c201 bl_201 br_201 wl_172 vdd gnd cell_6t
Xbit_r173_c201 bl_201 br_201 wl_173 vdd gnd cell_6t
Xbit_r174_c201 bl_201 br_201 wl_174 vdd gnd cell_6t
Xbit_r175_c201 bl_201 br_201 wl_175 vdd gnd cell_6t
Xbit_r176_c201 bl_201 br_201 wl_176 vdd gnd cell_6t
Xbit_r177_c201 bl_201 br_201 wl_177 vdd gnd cell_6t
Xbit_r178_c201 bl_201 br_201 wl_178 vdd gnd cell_6t
Xbit_r179_c201 bl_201 br_201 wl_179 vdd gnd cell_6t
Xbit_r180_c201 bl_201 br_201 wl_180 vdd gnd cell_6t
Xbit_r181_c201 bl_201 br_201 wl_181 vdd gnd cell_6t
Xbit_r182_c201 bl_201 br_201 wl_182 vdd gnd cell_6t
Xbit_r183_c201 bl_201 br_201 wl_183 vdd gnd cell_6t
Xbit_r184_c201 bl_201 br_201 wl_184 vdd gnd cell_6t
Xbit_r185_c201 bl_201 br_201 wl_185 vdd gnd cell_6t
Xbit_r186_c201 bl_201 br_201 wl_186 vdd gnd cell_6t
Xbit_r187_c201 bl_201 br_201 wl_187 vdd gnd cell_6t
Xbit_r188_c201 bl_201 br_201 wl_188 vdd gnd cell_6t
Xbit_r189_c201 bl_201 br_201 wl_189 vdd gnd cell_6t
Xbit_r190_c201 bl_201 br_201 wl_190 vdd gnd cell_6t
Xbit_r191_c201 bl_201 br_201 wl_191 vdd gnd cell_6t
Xbit_r192_c201 bl_201 br_201 wl_192 vdd gnd cell_6t
Xbit_r193_c201 bl_201 br_201 wl_193 vdd gnd cell_6t
Xbit_r194_c201 bl_201 br_201 wl_194 vdd gnd cell_6t
Xbit_r195_c201 bl_201 br_201 wl_195 vdd gnd cell_6t
Xbit_r196_c201 bl_201 br_201 wl_196 vdd gnd cell_6t
Xbit_r197_c201 bl_201 br_201 wl_197 vdd gnd cell_6t
Xbit_r198_c201 bl_201 br_201 wl_198 vdd gnd cell_6t
Xbit_r199_c201 bl_201 br_201 wl_199 vdd gnd cell_6t
Xbit_r200_c201 bl_201 br_201 wl_200 vdd gnd cell_6t
Xbit_r201_c201 bl_201 br_201 wl_201 vdd gnd cell_6t
Xbit_r202_c201 bl_201 br_201 wl_202 vdd gnd cell_6t
Xbit_r203_c201 bl_201 br_201 wl_203 vdd gnd cell_6t
Xbit_r204_c201 bl_201 br_201 wl_204 vdd gnd cell_6t
Xbit_r205_c201 bl_201 br_201 wl_205 vdd gnd cell_6t
Xbit_r206_c201 bl_201 br_201 wl_206 vdd gnd cell_6t
Xbit_r207_c201 bl_201 br_201 wl_207 vdd gnd cell_6t
Xbit_r208_c201 bl_201 br_201 wl_208 vdd gnd cell_6t
Xbit_r209_c201 bl_201 br_201 wl_209 vdd gnd cell_6t
Xbit_r210_c201 bl_201 br_201 wl_210 vdd gnd cell_6t
Xbit_r211_c201 bl_201 br_201 wl_211 vdd gnd cell_6t
Xbit_r212_c201 bl_201 br_201 wl_212 vdd gnd cell_6t
Xbit_r213_c201 bl_201 br_201 wl_213 vdd gnd cell_6t
Xbit_r214_c201 bl_201 br_201 wl_214 vdd gnd cell_6t
Xbit_r215_c201 bl_201 br_201 wl_215 vdd gnd cell_6t
Xbit_r216_c201 bl_201 br_201 wl_216 vdd gnd cell_6t
Xbit_r217_c201 bl_201 br_201 wl_217 vdd gnd cell_6t
Xbit_r218_c201 bl_201 br_201 wl_218 vdd gnd cell_6t
Xbit_r219_c201 bl_201 br_201 wl_219 vdd gnd cell_6t
Xbit_r220_c201 bl_201 br_201 wl_220 vdd gnd cell_6t
Xbit_r221_c201 bl_201 br_201 wl_221 vdd gnd cell_6t
Xbit_r222_c201 bl_201 br_201 wl_222 vdd gnd cell_6t
Xbit_r223_c201 bl_201 br_201 wl_223 vdd gnd cell_6t
Xbit_r224_c201 bl_201 br_201 wl_224 vdd gnd cell_6t
Xbit_r225_c201 bl_201 br_201 wl_225 vdd gnd cell_6t
Xbit_r226_c201 bl_201 br_201 wl_226 vdd gnd cell_6t
Xbit_r227_c201 bl_201 br_201 wl_227 vdd gnd cell_6t
Xbit_r228_c201 bl_201 br_201 wl_228 vdd gnd cell_6t
Xbit_r229_c201 bl_201 br_201 wl_229 vdd gnd cell_6t
Xbit_r230_c201 bl_201 br_201 wl_230 vdd gnd cell_6t
Xbit_r231_c201 bl_201 br_201 wl_231 vdd gnd cell_6t
Xbit_r232_c201 bl_201 br_201 wl_232 vdd gnd cell_6t
Xbit_r233_c201 bl_201 br_201 wl_233 vdd gnd cell_6t
Xbit_r234_c201 bl_201 br_201 wl_234 vdd gnd cell_6t
Xbit_r235_c201 bl_201 br_201 wl_235 vdd gnd cell_6t
Xbit_r236_c201 bl_201 br_201 wl_236 vdd gnd cell_6t
Xbit_r237_c201 bl_201 br_201 wl_237 vdd gnd cell_6t
Xbit_r238_c201 bl_201 br_201 wl_238 vdd gnd cell_6t
Xbit_r239_c201 bl_201 br_201 wl_239 vdd gnd cell_6t
Xbit_r240_c201 bl_201 br_201 wl_240 vdd gnd cell_6t
Xbit_r241_c201 bl_201 br_201 wl_241 vdd gnd cell_6t
Xbit_r242_c201 bl_201 br_201 wl_242 vdd gnd cell_6t
Xbit_r243_c201 bl_201 br_201 wl_243 vdd gnd cell_6t
Xbit_r244_c201 bl_201 br_201 wl_244 vdd gnd cell_6t
Xbit_r245_c201 bl_201 br_201 wl_245 vdd gnd cell_6t
Xbit_r246_c201 bl_201 br_201 wl_246 vdd gnd cell_6t
Xbit_r247_c201 bl_201 br_201 wl_247 vdd gnd cell_6t
Xbit_r248_c201 bl_201 br_201 wl_248 vdd gnd cell_6t
Xbit_r249_c201 bl_201 br_201 wl_249 vdd gnd cell_6t
Xbit_r250_c201 bl_201 br_201 wl_250 vdd gnd cell_6t
Xbit_r251_c201 bl_201 br_201 wl_251 vdd gnd cell_6t
Xbit_r252_c201 bl_201 br_201 wl_252 vdd gnd cell_6t
Xbit_r253_c201 bl_201 br_201 wl_253 vdd gnd cell_6t
Xbit_r254_c201 bl_201 br_201 wl_254 vdd gnd cell_6t
Xbit_r255_c201 bl_201 br_201 wl_255 vdd gnd cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd cell_6t
Xbit_r1_c202 bl_202 br_202 wl_1 vdd gnd cell_6t
Xbit_r2_c202 bl_202 br_202 wl_2 vdd gnd cell_6t
Xbit_r3_c202 bl_202 br_202 wl_3 vdd gnd cell_6t
Xbit_r4_c202 bl_202 br_202 wl_4 vdd gnd cell_6t
Xbit_r5_c202 bl_202 br_202 wl_5 vdd gnd cell_6t
Xbit_r6_c202 bl_202 br_202 wl_6 vdd gnd cell_6t
Xbit_r7_c202 bl_202 br_202 wl_7 vdd gnd cell_6t
Xbit_r8_c202 bl_202 br_202 wl_8 vdd gnd cell_6t
Xbit_r9_c202 bl_202 br_202 wl_9 vdd gnd cell_6t
Xbit_r10_c202 bl_202 br_202 wl_10 vdd gnd cell_6t
Xbit_r11_c202 bl_202 br_202 wl_11 vdd gnd cell_6t
Xbit_r12_c202 bl_202 br_202 wl_12 vdd gnd cell_6t
Xbit_r13_c202 bl_202 br_202 wl_13 vdd gnd cell_6t
Xbit_r14_c202 bl_202 br_202 wl_14 vdd gnd cell_6t
Xbit_r15_c202 bl_202 br_202 wl_15 vdd gnd cell_6t
Xbit_r16_c202 bl_202 br_202 wl_16 vdd gnd cell_6t
Xbit_r17_c202 bl_202 br_202 wl_17 vdd gnd cell_6t
Xbit_r18_c202 bl_202 br_202 wl_18 vdd gnd cell_6t
Xbit_r19_c202 bl_202 br_202 wl_19 vdd gnd cell_6t
Xbit_r20_c202 bl_202 br_202 wl_20 vdd gnd cell_6t
Xbit_r21_c202 bl_202 br_202 wl_21 vdd gnd cell_6t
Xbit_r22_c202 bl_202 br_202 wl_22 vdd gnd cell_6t
Xbit_r23_c202 bl_202 br_202 wl_23 vdd gnd cell_6t
Xbit_r24_c202 bl_202 br_202 wl_24 vdd gnd cell_6t
Xbit_r25_c202 bl_202 br_202 wl_25 vdd gnd cell_6t
Xbit_r26_c202 bl_202 br_202 wl_26 vdd gnd cell_6t
Xbit_r27_c202 bl_202 br_202 wl_27 vdd gnd cell_6t
Xbit_r28_c202 bl_202 br_202 wl_28 vdd gnd cell_6t
Xbit_r29_c202 bl_202 br_202 wl_29 vdd gnd cell_6t
Xbit_r30_c202 bl_202 br_202 wl_30 vdd gnd cell_6t
Xbit_r31_c202 bl_202 br_202 wl_31 vdd gnd cell_6t
Xbit_r32_c202 bl_202 br_202 wl_32 vdd gnd cell_6t
Xbit_r33_c202 bl_202 br_202 wl_33 vdd gnd cell_6t
Xbit_r34_c202 bl_202 br_202 wl_34 vdd gnd cell_6t
Xbit_r35_c202 bl_202 br_202 wl_35 vdd gnd cell_6t
Xbit_r36_c202 bl_202 br_202 wl_36 vdd gnd cell_6t
Xbit_r37_c202 bl_202 br_202 wl_37 vdd gnd cell_6t
Xbit_r38_c202 bl_202 br_202 wl_38 vdd gnd cell_6t
Xbit_r39_c202 bl_202 br_202 wl_39 vdd gnd cell_6t
Xbit_r40_c202 bl_202 br_202 wl_40 vdd gnd cell_6t
Xbit_r41_c202 bl_202 br_202 wl_41 vdd gnd cell_6t
Xbit_r42_c202 bl_202 br_202 wl_42 vdd gnd cell_6t
Xbit_r43_c202 bl_202 br_202 wl_43 vdd gnd cell_6t
Xbit_r44_c202 bl_202 br_202 wl_44 vdd gnd cell_6t
Xbit_r45_c202 bl_202 br_202 wl_45 vdd gnd cell_6t
Xbit_r46_c202 bl_202 br_202 wl_46 vdd gnd cell_6t
Xbit_r47_c202 bl_202 br_202 wl_47 vdd gnd cell_6t
Xbit_r48_c202 bl_202 br_202 wl_48 vdd gnd cell_6t
Xbit_r49_c202 bl_202 br_202 wl_49 vdd gnd cell_6t
Xbit_r50_c202 bl_202 br_202 wl_50 vdd gnd cell_6t
Xbit_r51_c202 bl_202 br_202 wl_51 vdd gnd cell_6t
Xbit_r52_c202 bl_202 br_202 wl_52 vdd gnd cell_6t
Xbit_r53_c202 bl_202 br_202 wl_53 vdd gnd cell_6t
Xbit_r54_c202 bl_202 br_202 wl_54 vdd gnd cell_6t
Xbit_r55_c202 bl_202 br_202 wl_55 vdd gnd cell_6t
Xbit_r56_c202 bl_202 br_202 wl_56 vdd gnd cell_6t
Xbit_r57_c202 bl_202 br_202 wl_57 vdd gnd cell_6t
Xbit_r58_c202 bl_202 br_202 wl_58 vdd gnd cell_6t
Xbit_r59_c202 bl_202 br_202 wl_59 vdd gnd cell_6t
Xbit_r60_c202 bl_202 br_202 wl_60 vdd gnd cell_6t
Xbit_r61_c202 bl_202 br_202 wl_61 vdd gnd cell_6t
Xbit_r62_c202 bl_202 br_202 wl_62 vdd gnd cell_6t
Xbit_r63_c202 bl_202 br_202 wl_63 vdd gnd cell_6t
Xbit_r64_c202 bl_202 br_202 wl_64 vdd gnd cell_6t
Xbit_r65_c202 bl_202 br_202 wl_65 vdd gnd cell_6t
Xbit_r66_c202 bl_202 br_202 wl_66 vdd gnd cell_6t
Xbit_r67_c202 bl_202 br_202 wl_67 vdd gnd cell_6t
Xbit_r68_c202 bl_202 br_202 wl_68 vdd gnd cell_6t
Xbit_r69_c202 bl_202 br_202 wl_69 vdd gnd cell_6t
Xbit_r70_c202 bl_202 br_202 wl_70 vdd gnd cell_6t
Xbit_r71_c202 bl_202 br_202 wl_71 vdd gnd cell_6t
Xbit_r72_c202 bl_202 br_202 wl_72 vdd gnd cell_6t
Xbit_r73_c202 bl_202 br_202 wl_73 vdd gnd cell_6t
Xbit_r74_c202 bl_202 br_202 wl_74 vdd gnd cell_6t
Xbit_r75_c202 bl_202 br_202 wl_75 vdd gnd cell_6t
Xbit_r76_c202 bl_202 br_202 wl_76 vdd gnd cell_6t
Xbit_r77_c202 bl_202 br_202 wl_77 vdd gnd cell_6t
Xbit_r78_c202 bl_202 br_202 wl_78 vdd gnd cell_6t
Xbit_r79_c202 bl_202 br_202 wl_79 vdd gnd cell_6t
Xbit_r80_c202 bl_202 br_202 wl_80 vdd gnd cell_6t
Xbit_r81_c202 bl_202 br_202 wl_81 vdd gnd cell_6t
Xbit_r82_c202 bl_202 br_202 wl_82 vdd gnd cell_6t
Xbit_r83_c202 bl_202 br_202 wl_83 vdd gnd cell_6t
Xbit_r84_c202 bl_202 br_202 wl_84 vdd gnd cell_6t
Xbit_r85_c202 bl_202 br_202 wl_85 vdd gnd cell_6t
Xbit_r86_c202 bl_202 br_202 wl_86 vdd gnd cell_6t
Xbit_r87_c202 bl_202 br_202 wl_87 vdd gnd cell_6t
Xbit_r88_c202 bl_202 br_202 wl_88 vdd gnd cell_6t
Xbit_r89_c202 bl_202 br_202 wl_89 vdd gnd cell_6t
Xbit_r90_c202 bl_202 br_202 wl_90 vdd gnd cell_6t
Xbit_r91_c202 bl_202 br_202 wl_91 vdd gnd cell_6t
Xbit_r92_c202 bl_202 br_202 wl_92 vdd gnd cell_6t
Xbit_r93_c202 bl_202 br_202 wl_93 vdd gnd cell_6t
Xbit_r94_c202 bl_202 br_202 wl_94 vdd gnd cell_6t
Xbit_r95_c202 bl_202 br_202 wl_95 vdd gnd cell_6t
Xbit_r96_c202 bl_202 br_202 wl_96 vdd gnd cell_6t
Xbit_r97_c202 bl_202 br_202 wl_97 vdd gnd cell_6t
Xbit_r98_c202 bl_202 br_202 wl_98 vdd gnd cell_6t
Xbit_r99_c202 bl_202 br_202 wl_99 vdd gnd cell_6t
Xbit_r100_c202 bl_202 br_202 wl_100 vdd gnd cell_6t
Xbit_r101_c202 bl_202 br_202 wl_101 vdd gnd cell_6t
Xbit_r102_c202 bl_202 br_202 wl_102 vdd gnd cell_6t
Xbit_r103_c202 bl_202 br_202 wl_103 vdd gnd cell_6t
Xbit_r104_c202 bl_202 br_202 wl_104 vdd gnd cell_6t
Xbit_r105_c202 bl_202 br_202 wl_105 vdd gnd cell_6t
Xbit_r106_c202 bl_202 br_202 wl_106 vdd gnd cell_6t
Xbit_r107_c202 bl_202 br_202 wl_107 vdd gnd cell_6t
Xbit_r108_c202 bl_202 br_202 wl_108 vdd gnd cell_6t
Xbit_r109_c202 bl_202 br_202 wl_109 vdd gnd cell_6t
Xbit_r110_c202 bl_202 br_202 wl_110 vdd gnd cell_6t
Xbit_r111_c202 bl_202 br_202 wl_111 vdd gnd cell_6t
Xbit_r112_c202 bl_202 br_202 wl_112 vdd gnd cell_6t
Xbit_r113_c202 bl_202 br_202 wl_113 vdd gnd cell_6t
Xbit_r114_c202 bl_202 br_202 wl_114 vdd gnd cell_6t
Xbit_r115_c202 bl_202 br_202 wl_115 vdd gnd cell_6t
Xbit_r116_c202 bl_202 br_202 wl_116 vdd gnd cell_6t
Xbit_r117_c202 bl_202 br_202 wl_117 vdd gnd cell_6t
Xbit_r118_c202 bl_202 br_202 wl_118 vdd gnd cell_6t
Xbit_r119_c202 bl_202 br_202 wl_119 vdd gnd cell_6t
Xbit_r120_c202 bl_202 br_202 wl_120 vdd gnd cell_6t
Xbit_r121_c202 bl_202 br_202 wl_121 vdd gnd cell_6t
Xbit_r122_c202 bl_202 br_202 wl_122 vdd gnd cell_6t
Xbit_r123_c202 bl_202 br_202 wl_123 vdd gnd cell_6t
Xbit_r124_c202 bl_202 br_202 wl_124 vdd gnd cell_6t
Xbit_r125_c202 bl_202 br_202 wl_125 vdd gnd cell_6t
Xbit_r126_c202 bl_202 br_202 wl_126 vdd gnd cell_6t
Xbit_r127_c202 bl_202 br_202 wl_127 vdd gnd cell_6t
Xbit_r128_c202 bl_202 br_202 wl_128 vdd gnd cell_6t
Xbit_r129_c202 bl_202 br_202 wl_129 vdd gnd cell_6t
Xbit_r130_c202 bl_202 br_202 wl_130 vdd gnd cell_6t
Xbit_r131_c202 bl_202 br_202 wl_131 vdd gnd cell_6t
Xbit_r132_c202 bl_202 br_202 wl_132 vdd gnd cell_6t
Xbit_r133_c202 bl_202 br_202 wl_133 vdd gnd cell_6t
Xbit_r134_c202 bl_202 br_202 wl_134 vdd gnd cell_6t
Xbit_r135_c202 bl_202 br_202 wl_135 vdd gnd cell_6t
Xbit_r136_c202 bl_202 br_202 wl_136 vdd gnd cell_6t
Xbit_r137_c202 bl_202 br_202 wl_137 vdd gnd cell_6t
Xbit_r138_c202 bl_202 br_202 wl_138 vdd gnd cell_6t
Xbit_r139_c202 bl_202 br_202 wl_139 vdd gnd cell_6t
Xbit_r140_c202 bl_202 br_202 wl_140 vdd gnd cell_6t
Xbit_r141_c202 bl_202 br_202 wl_141 vdd gnd cell_6t
Xbit_r142_c202 bl_202 br_202 wl_142 vdd gnd cell_6t
Xbit_r143_c202 bl_202 br_202 wl_143 vdd gnd cell_6t
Xbit_r144_c202 bl_202 br_202 wl_144 vdd gnd cell_6t
Xbit_r145_c202 bl_202 br_202 wl_145 vdd gnd cell_6t
Xbit_r146_c202 bl_202 br_202 wl_146 vdd gnd cell_6t
Xbit_r147_c202 bl_202 br_202 wl_147 vdd gnd cell_6t
Xbit_r148_c202 bl_202 br_202 wl_148 vdd gnd cell_6t
Xbit_r149_c202 bl_202 br_202 wl_149 vdd gnd cell_6t
Xbit_r150_c202 bl_202 br_202 wl_150 vdd gnd cell_6t
Xbit_r151_c202 bl_202 br_202 wl_151 vdd gnd cell_6t
Xbit_r152_c202 bl_202 br_202 wl_152 vdd gnd cell_6t
Xbit_r153_c202 bl_202 br_202 wl_153 vdd gnd cell_6t
Xbit_r154_c202 bl_202 br_202 wl_154 vdd gnd cell_6t
Xbit_r155_c202 bl_202 br_202 wl_155 vdd gnd cell_6t
Xbit_r156_c202 bl_202 br_202 wl_156 vdd gnd cell_6t
Xbit_r157_c202 bl_202 br_202 wl_157 vdd gnd cell_6t
Xbit_r158_c202 bl_202 br_202 wl_158 vdd gnd cell_6t
Xbit_r159_c202 bl_202 br_202 wl_159 vdd gnd cell_6t
Xbit_r160_c202 bl_202 br_202 wl_160 vdd gnd cell_6t
Xbit_r161_c202 bl_202 br_202 wl_161 vdd gnd cell_6t
Xbit_r162_c202 bl_202 br_202 wl_162 vdd gnd cell_6t
Xbit_r163_c202 bl_202 br_202 wl_163 vdd gnd cell_6t
Xbit_r164_c202 bl_202 br_202 wl_164 vdd gnd cell_6t
Xbit_r165_c202 bl_202 br_202 wl_165 vdd gnd cell_6t
Xbit_r166_c202 bl_202 br_202 wl_166 vdd gnd cell_6t
Xbit_r167_c202 bl_202 br_202 wl_167 vdd gnd cell_6t
Xbit_r168_c202 bl_202 br_202 wl_168 vdd gnd cell_6t
Xbit_r169_c202 bl_202 br_202 wl_169 vdd gnd cell_6t
Xbit_r170_c202 bl_202 br_202 wl_170 vdd gnd cell_6t
Xbit_r171_c202 bl_202 br_202 wl_171 vdd gnd cell_6t
Xbit_r172_c202 bl_202 br_202 wl_172 vdd gnd cell_6t
Xbit_r173_c202 bl_202 br_202 wl_173 vdd gnd cell_6t
Xbit_r174_c202 bl_202 br_202 wl_174 vdd gnd cell_6t
Xbit_r175_c202 bl_202 br_202 wl_175 vdd gnd cell_6t
Xbit_r176_c202 bl_202 br_202 wl_176 vdd gnd cell_6t
Xbit_r177_c202 bl_202 br_202 wl_177 vdd gnd cell_6t
Xbit_r178_c202 bl_202 br_202 wl_178 vdd gnd cell_6t
Xbit_r179_c202 bl_202 br_202 wl_179 vdd gnd cell_6t
Xbit_r180_c202 bl_202 br_202 wl_180 vdd gnd cell_6t
Xbit_r181_c202 bl_202 br_202 wl_181 vdd gnd cell_6t
Xbit_r182_c202 bl_202 br_202 wl_182 vdd gnd cell_6t
Xbit_r183_c202 bl_202 br_202 wl_183 vdd gnd cell_6t
Xbit_r184_c202 bl_202 br_202 wl_184 vdd gnd cell_6t
Xbit_r185_c202 bl_202 br_202 wl_185 vdd gnd cell_6t
Xbit_r186_c202 bl_202 br_202 wl_186 vdd gnd cell_6t
Xbit_r187_c202 bl_202 br_202 wl_187 vdd gnd cell_6t
Xbit_r188_c202 bl_202 br_202 wl_188 vdd gnd cell_6t
Xbit_r189_c202 bl_202 br_202 wl_189 vdd gnd cell_6t
Xbit_r190_c202 bl_202 br_202 wl_190 vdd gnd cell_6t
Xbit_r191_c202 bl_202 br_202 wl_191 vdd gnd cell_6t
Xbit_r192_c202 bl_202 br_202 wl_192 vdd gnd cell_6t
Xbit_r193_c202 bl_202 br_202 wl_193 vdd gnd cell_6t
Xbit_r194_c202 bl_202 br_202 wl_194 vdd gnd cell_6t
Xbit_r195_c202 bl_202 br_202 wl_195 vdd gnd cell_6t
Xbit_r196_c202 bl_202 br_202 wl_196 vdd gnd cell_6t
Xbit_r197_c202 bl_202 br_202 wl_197 vdd gnd cell_6t
Xbit_r198_c202 bl_202 br_202 wl_198 vdd gnd cell_6t
Xbit_r199_c202 bl_202 br_202 wl_199 vdd gnd cell_6t
Xbit_r200_c202 bl_202 br_202 wl_200 vdd gnd cell_6t
Xbit_r201_c202 bl_202 br_202 wl_201 vdd gnd cell_6t
Xbit_r202_c202 bl_202 br_202 wl_202 vdd gnd cell_6t
Xbit_r203_c202 bl_202 br_202 wl_203 vdd gnd cell_6t
Xbit_r204_c202 bl_202 br_202 wl_204 vdd gnd cell_6t
Xbit_r205_c202 bl_202 br_202 wl_205 vdd gnd cell_6t
Xbit_r206_c202 bl_202 br_202 wl_206 vdd gnd cell_6t
Xbit_r207_c202 bl_202 br_202 wl_207 vdd gnd cell_6t
Xbit_r208_c202 bl_202 br_202 wl_208 vdd gnd cell_6t
Xbit_r209_c202 bl_202 br_202 wl_209 vdd gnd cell_6t
Xbit_r210_c202 bl_202 br_202 wl_210 vdd gnd cell_6t
Xbit_r211_c202 bl_202 br_202 wl_211 vdd gnd cell_6t
Xbit_r212_c202 bl_202 br_202 wl_212 vdd gnd cell_6t
Xbit_r213_c202 bl_202 br_202 wl_213 vdd gnd cell_6t
Xbit_r214_c202 bl_202 br_202 wl_214 vdd gnd cell_6t
Xbit_r215_c202 bl_202 br_202 wl_215 vdd gnd cell_6t
Xbit_r216_c202 bl_202 br_202 wl_216 vdd gnd cell_6t
Xbit_r217_c202 bl_202 br_202 wl_217 vdd gnd cell_6t
Xbit_r218_c202 bl_202 br_202 wl_218 vdd gnd cell_6t
Xbit_r219_c202 bl_202 br_202 wl_219 vdd gnd cell_6t
Xbit_r220_c202 bl_202 br_202 wl_220 vdd gnd cell_6t
Xbit_r221_c202 bl_202 br_202 wl_221 vdd gnd cell_6t
Xbit_r222_c202 bl_202 br_202 wl_222 vdd gnd cell_6t
Xbit_r223_c202 bl_202 br_202 wl_223 vdd gnd cell_6t
Xbit_r224_c202 bl_202 br_202 wl_224 vdd gnd cell_6t
Xbit_r225_c202 bl_202 br_202 wl_225 vdd gnd cell_6t
Xbit_r226_c202 bl_202 br_202 wl_226 vdd gnd cell_6t
Xbit_r227_c202 bl_202 br_202 wl_227 vdd gnd cell_6t
Xbit_r228_c202 bl_202 br_202 wl_228 vdd gnd cell_6t
Xbit_r229_c202 bl_202 br_202 wl_229 vdd gnd cell_6t
Xbit_r230_c202 bl_202 br_202 wl_230 vdd gnd cell_6t
Xbit_r231_c202 bl_202 br_202 wl_231 vdd gnd cell_6t
Xbit_r232_c202 bl_202 br_202 wl_232 vdd gnd cell_6t
Xbit_r233_c202 bl_202 br_202 wl_233 vdd gnd cell_6t
Xbit_r234_c202 bl_202 br_202 wl_234 vdd gnd cell_6t
Xbit_r235_c202 bl_202 br_202 wl_235 vdd gnd cell_6t
Xbit_r236_c202 bl_202 br_202 wl_236 vdd gnd cell_6t
Xbit_r237_c202 bl_202 br_202 wl_237 vdd gnd cell_6t
Xbit_r238_c202 bl_202 br_202 wl_238 vdd gnd cell_6t
Xbit_r239_c202 bl_202 br_202 wl_239 vdd gnd cell_6t
Xbit_r240_c202 bl_202 br_202 wl_240 vdd gnd cell_6t
Xbit_r241_c202 bl_202 br_202 wl_241 vdd gnd cell_6t
Xbit_r242_c202 bl_202 br_202 wl_242 vdd gnd cell_6t
Xbit_r243_c202 bl_202 br_202 wl_243 vdd gnd cell_6t
Xbit_r244_c202 bl_202 br_202 wl_244 vdd gnd cell_6t
Xbit_r245_c202 bl_202 br_202 wl_245 vdd gnd cell_6t
Xbit_r246_c202 bl_202 br_202 wl_246 vdd gnd cell_6t
Xbit_r247_c202 bl_202 br_202 wl_247 vdd gnd cell_6t
Xbit_r248_c202 bl_202 br_202 wl_248 vdd gnd cell_6t
Xbit_r249_c202 bl_202 br_202 wl_249 vdd gnd cell_6t
Xbit_r250_c202 bl_202 br_202 wl_250 vdd gnd cell_6t
Xbit_r251_c202 bl_202 br_202 wl_251 vdd gnd cell_6t
Xbit_r252_c202 bl_202 br_202 wl_252 vdd gnd cell_6t
Xbit_r253_c202 bl_202 br_202 wl_253 vdd gnd cell_6t
Xbit_r254_c202 bl_202 br_202 wl_254 vdd gnd cell_6t
Xbit_r255_c202 bl_202 br_202 wl_255 vdd gnd cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd cell_6t
Xbit_r1_c203 bl_203 br_203 wl_1 vdd gnd cell_6t
Xbit_r2_c203 bl_203 br_203 wl_2 vdd gnd cell_6t
Xbit_r3_c203 bl_203 br_203 wl_3 vdd gnd cell_6t
Xbit_r4_c203 bl_203 br_203 wl_4 vdd gnd cell_6t
Xbit_r5_c203 bl_203 br_203 wl_5 vdd gnd cell_6t
Xbit_r6_c203 bl_203 br_203 wl_6 vdd gnd cell_6t
Xbit_r7_c203 bl_203 br_203 wl_7 vdd gnd cell_6t
Xbit_r8_c203 bl_203 br_203 wl_8 vdd gnd cell_6t
Xbit_r9_c203 bl_203 br_203 wl_9 vdd gnd cell_6t
Xbit_r10_c203 bl_203 br_203 wl_10 vdd gnd cell_6t
Xbit_r11_c203 bl_203 br_203 wl_11 vdd gnd cell_6t
Xbit_r12_c203 bl_203 br_203 wl_12 vdd gnd cell_6t
Xbit_r13_c203 bl_203 br_203 wl_13 vdd gnd cell_6t
Xbit_r14_c203 bl_203 br_203 wl_14 vdd gnd cell_6t
Xbit_r15_c203 bl_203 br_203 wl_15 vdd gnd cell_6t
Xbit_r16_c203 bl_203 br_203 wl_16 vdd gnd cell_6t
Xbit_r17_c203 bl_203 br_203 wl_17 vdd gnd cell_6t
Xbit_r18_c203 bl_203 br_203 wl_18 vdd gnd cell_6t
Xbit_r19_c203 bl_203 br_203 wl_19 vdd gnd cell_6t
Xbit_r20_c203 bl_203 br_203 wl_20 vdd gnd cell_6t
Xbit_r21_c203 bl_203 br_203 wl_21 vdd gnd cell_6t
Xbit_r22_c203 bl_203 br_203 wl_22 vdd gnd cell_6t
Xbit_r23_c203 bl_203 br_203 wl_23 vdd gnd cell_6t
Xbit_r24_c203 bl_203 br_203 wl_24 vdd gnd cell_6t
Xbit_r25_c203 bl_203 br_203 wl_25 vdd gnd cell_6t
Xbit_r26_c203 bl_203 br_203 wl_26 vdd gnd cell_6t
Xbit_r27_c203 bl_203 br_203 wl_27 vdd gnd cell_6t
Xbit_r28_c203 bl_203 br_203 wl_28 vdd gnd cell_6t
Xbit_r29_c203 bl_203 br_203 wl_29 vdd gnd cell_6t
Xbit_r30_c203 bl_203 br_203 wl_30 vdd gnd cell_6t
Xbit_r31_c203 bl_203 br_203 wl_31 vdd gnd cell_6t
Xbit_r32_c203 bl_203 br_203 wl_32 vdd gnd cell_6t
Xbit_r33_c203 bl_203 br_203 wl_33 vdd gnd cell_6t
Xbit_r34_c203 bl_203 br_203 wl_34 vdd gnd cell_6t
Xbit_r35_c203 bl_203 br_203 wl_35 vdd gnd cell_6t
Xbit_r36_c203 bl_203 br_203 wl_36 vdd gnd cell_6t
Xbit_r37_c203 bl_203 br_203 wl_37 vdd gnd cell_6t
Xbit_r38_c203 bl_203 br_203 wl_38 vdd gnd cell_6t
Xbit_r39_c203 bl_203 br_203 wl_39 vdd gnd cell_6t
Xbit_r40_c203 bl_203 br_203 wl_40 vdd gnd cell_6t
Xbit_r41_c203 bl_203 br_203 wl_41 vdd gnd cell_6t
Xbit_r42_c203 bl_203 br_203 wl_42 vdd gnd cell_6t
Xbit_r43_c203 bl_203 br_203 wl_43 vdd gnd cell_6t
Xbit_r44_c203 bl_203 br_203 wl_44 vdd gnd cell_6t
Xbit_r45_c203 bl_203 br_203 wl_45 vdd gnd cell_6t
Xbit_r46_c203 bl_203 br_203 wl_46 vdd gnd cell_6t
Xbit_r47_c203 bl_203 br_203 wl_47 vdd gnd cell_6t
Xbit_r48_c203 bl_203 br_203 wl_48 vdd gnd cell_6t
Xbit_r49_c203 bl_203 br_203 wl_49 vdd gnd cell_6t
Xbit_r50_c203 bl_203 br_203 wl_50 vdd gnd cell_6t
Xbit_r51_c203 bl_203 br_203 wl_51 vdd gnd cell_6t
Xbit_r52_c203 bl_203 br_203 wl_52 vdd gnd cell_6t
Xbit_r53_c203 bl_203 br_203 wl_53 vdd gnd cell_6t
Xbit_r54_c203 bl_203 br_203 wl_54 vdd gnd cell_6t
Xbit_r55_c203 bl_203 br_203 wl_55 vdd gnd cell_6t
Xbit_r56_c203 bl_203 br_203 wl_56 vdd gnd cell_6t
Xbit_r57_c203 bl_203 br_203 wl_57 vdd gnd cell_6t
Xbit_r58_c203 bl_203 br_203 wl_58 vdd gnd cell_6t
Xbit_r59_c203 bl_203 br_203 wl_59 vdd gnd cell_6t
Xbit_r60_c203 bl_203 br_203 wl_60 vdd gnd cell_6t
Xbit_r61_c203 bl_203 br_203 wl_61 vdd gnd cell_6t
Xbit_r62_c203 bl_203 br_203 wl_62 vdd gnd cell_6t
Xbit_r63_c203 bl_203 br_203 wl_63 vdd gnd cell_6t
Xbit_r64_c203 bl_203 br_203 wl_64 vdd gnd cell_6t
Xbit_r65_c203 bl_203 br_203 wl_65 vdd gnd cell_6t
Xbit_r66_c203 bl_203 br_203 wl_66 vdd gnd cell_6t
Xbit_r67_c203 bl_203 br_203 wl_67 vdd gnd cell_6t
Xbit_r68_c203 bl_203 br_203 wl_68 vdd gnd cell_6t
Xbit_r69_c203 bl_203 br_203 wl_69 vdd gnd cell_6t
Xbit_r70_c203 bl_203 br_203 wl_70 vdd gnd cell_6t
Xbit_r71_c203 bl_203 br_203 wl_71 vdd gnd cell_6t
Xbit_r72_c203 bl_203 br_203 wl_72 vdd gnd cell_6t
Xbit_r73_c203 bl_203 br_203 wl_73 vdd gnd cell_6t
Xbit_r74_c203 bl_203 br_203 wl_74 vdd gnd cell_6t
Xbit_r75_c203 bl_203 br_203 wl_75 vdd gnd cell_6t
Xbit_r76_c203 bl_203 br_203 wl_76 vdd gnd cell_6t
Xbit_r77_c203 bl_203 br_203 wl_77 vdd gnd cell_6t
Xbit_r78_c203 bl_203 br_203 wl_78 vdd gnd cell_6t
Xbit_r79_c203 bl_203 br_203 wl_79 vdd gnd cell_6t
Xbit_r80_c203 bl_203 br_203 wl_80 vdd gnd cell_6t
Xbit_r81_c203 bl_203 br_203 wl_81 vdd gnd cell_6t
Xbit_r82_c203 bl_203 br_203 wl_82 vdd gnd cell_6t
Xbit_r83_c203 bl_203 br_203 wl_83 vdd gnd cell_6t
Xbit_r84_c203 bl_203 br_203 wl_84 vdd gnd cell_6t
Xbit_r85_c203 bl_203 br_203 wl_85 vdd gnd cell_6t
Xbit_r86_c203 bl_203 br_203 wl_86 vdd gnd cell_6t
Xbit_r87_c203 bl_203 br_203 wl_87 vdd gnd cell_6t
Xbit_r88_c203 bl_203 br_203 wl_88 vdd gnd cell_6t
Xbit_r89_c203 bl_203 br_203 wl_89 vdd gnd cell_6t
Xbit_r90_c203 bl_203 br_203 wl_90 vdd gnd cell_6t
Xbit_r91_c203 bl_203 br_203 wl_91 vdd gnd cell_6t
Xbit_r92_c203 bl_203 br_203 wl_92 vdd gnd cell_6t
Xbit_r93_c203 bl_203 br_203 wl_93 vdd gnd cell_6t
Xbit_r94_c203 bl_203 br_203 wl_94 vdd gnd cell_6t
Xbit_r95_c203 bl_203 br_203 wl_95 vdd gnd cell_6t
Xbit_r96_c203 bl_203 br_203 wl_96 vdd gnd cell_6t
Xbit_r97_c203 bl_203 br_203 wl_97 vdd gnd cell_6t
Xbit_r98_c203 bl_203 br_203 wl_98 vdd gnd cell_6t
Xbit_r99_c203 bl_203 br_203 wl_99 vdd gnd cell_6t
Xbit_r100_c203 bl_203 br_203 wl_100 vdd gnd cell_6t
Xbit_r101_c203 bl_203 br_203 wl_101 vdd gnd cell_6t
Xbit_r102_c203 bl_203 br_203 wl_102 vdd gnd cell_6t
Xbit_r103_c203 bl_203 br_203 wl_103 vdd gnd cell_6t
Xbit_r104_c203 bl_203 br_203 wl_104 vdd gnd cell_6t
Xbit_r105_c203 bl_203 br_203 wl_105 vdd gnd cell_6t
Xbit_r106_c203 bl_203 br_203 wl_106 vdd gnd cell_6t
Xbit_r107_c203 bl_203 br_203 wl_107 vdd gnd cell_6t
Xbit_r108_c203 bl_203 br_203 wl_108 vdd gnd cell_6t
Xbit_r109_c203 bl_203 br_203 wl_109 vdd gnd cell_6t
Xbit_r110_c203 bl_203 br_203 wl_110 vdd gnd cell_6t
Xbit_r111_c203 bl_203 br_203 wl_111 vdd gnd cell_6t
Xbit_r112_c203 bl_203 br_203 wl_112 vdd gnd cell_6t
Xbit_r113_c203 bl_203 br_203 wl_113 vdd gnd cell_6t
Xbit_r114_c203 bl_203 br_203 wl_114 vdd gnd cell_6t
Xbit_r115_c203 bl_203 br_203 wl_115 vdd gnd cell_6t
Xbit_r116_c203 bl_203 br_203 wl_116 vdd gnd cell_6t
Xbit_r117_c203 bl_203 br_203 wl_117 vdd gnd cell_6t
Xbit_r118_c203 bl_203 br_203 wl_118 vdd gnd cell_6t
Xbit_r119_c203 bl_203 br_203 wl_119 vdd gnd cell_6t
Xbit_r120_c203 bl_203 br_203 wl_120 vdd gnd cell_6t
Xbit_r121_c203 bl_203 br_203 wl_121 vdd gnd cell_6t
Xbit_r122_c203 bl_203 br_203 wl_122 vdd gnd cell_6t
Xbit_r123_c203 bl_203 br_203 wl_123 vdd gnd cell_6t
Xbit_r124_c203 bl_203 br_203 wl_124 vdd gnd cell_6t
Xbit_r125_c203 bl_203 br_203 wl_125 vdd gnd cell_6t
Xbit_r126_c203 bl_203 br_203 wl_126 vdd gnd cell_6t
Xbit_r127_c203 bl_203 br_203 wl_127 vdd gnd cell_6t
Xbit_r128_c203 bl_203 br_203 wl_128 vdd gnd cell_6t
Xbit_r129_c203 bl_203 br_203 wl_129 vdd gnd cell_6t
Xbit_r130_c203 bl_203 br_203 wl_130 vdd gnd cell_6t
Xbit_r131_c203 bl_203 br_203 wl_131 vdd gnd cell_6t
Xbit_r132_c203 bl_203 br_203 wl_132 vdd gnd cell_6t
Xbit_r133_c203 bl_203 br_203 wl_133 vdd gnd cell_6t
Xbit_r134_c203 bl_203 br_203 wl_134 vdd gnd cell_6t
Xbit_r135_c203 bl_203 br_203 wl_135 vdd gnd cell_6t
Xbit_r136_c203 bl_203 br_203 wl_136 vdd gnd cell_6t
Xbit_r137_c203 bl_203 br_203 wl_137 vdd gnd cell_6t
Xbit_r138_c203 bl_203 br_203 wl_138 vdd gnd cell_6t
Xbit_r139_c203 bl_203 br_203 wl_139 vdd gnd cell_6t
Xbit_r140_c203 bl_203 br_203 wl_140 vdd gnd cell_6t
Xbit_r141_c203 bl_203 br_203 wl_141 vdd gnd cell_6t
Xbit_r142_c203 bl_203 br_203 wl_142 vdd gnd cell_6t
Xbit_r143_c203 bl_203 br_203 wl_143 vdd gnd cell_6t
Xbit_r144_c203 bl_203 br_203 wl_144 vdd gnd cell_6t
Xbit_r145_c203 bl_203 br_203 wl_145 vdd gnd cell_6t
Xbit_r146_c203 bl_203 br_203 wl_146 vdd gnd cell_6t
Xbit_r147_c203 bl_203 br_203 wl_147 vdd gnd cell_6t
Xbit_r148_c203 bl_203 br_203 wl_148 vdd gnd cell_6t
Xbit_r149_c203 bl_203 br_203 wl_149 vdd gnd cell_6t
Xbit_r150_c203 bl_203 br_203 wl_150 vdd gnd cell_6t
Xbit_r151_c203 bl_203 br_203 wl_151 vdd gnd cell_6t
Xbit_r152_c203 bl_203 br_203 wl_152 vdd gnd cell_6t
Xbit_r153_c203 bl_203 br_203 wl_153 vdd gnd cell_6t
Xbit_r154_c203 bl_203 br_203 wl_154 vdd gnd cell_6t
Xbit_r155_c203 bl_203 br_203 wl_155 vdd gnd cell_6t
Xbit_r156_c203 bl_203 br_203 wl_156 vdd gnd cell_6t
Xbit_r157_c203 bl_203 br_203 wl_157 vdd gnd cell_6t
Xbit_r158_c203 bl_203 br_203 wl_158 vdd gnd cell_6t
Xbit_r159_c203 bl_203 br_203 wl_159 vdd gnd cell_6t
Xbit_r160_c203 bl_203 br_203 wl_160 vdd gnd cell_6t
Xbit_r161_c203 bl_203 br_203 wl_161 vdd gnd cell_6t
Xbit_r162_c203 bl_203 br_203 wl_162 vdd gnd cell_6t
Xbit_r163_c203 bl_203 br_203 wl_163 vdd gnd cell_6t
Xbit_r164_c203 bl_203 br_203 wl_164 vdd gnd cell_6t
Xbit_r165_c203 bl_203 br_203 wl_165 vdd gnd cell_6t
Xbit_r166_c203 bl_203 br_203 wl_166 vdd gnd cell_6t
Xbit_r167_c203 bl_203 br_203 wl_167 vdd gnd cell_6t
Xbit_r168_c203 bl_203 br_203 wl_168 vdd gnd cell_6t
Xbit_r169_c203 bl_203 br_203 wl_169 vdd gnd cell_6t
Xbit_r170_c203 bl_203 br_203 wl_170 vdd gnd cell_6t
Xbit_r171_c203 bl_203 br_203 wl_171 vdd gnd cell_6t
Xbit_r172_c203 bl_203 br_203 wl_172 vdd gnd cell_6t
Xbit_r173_c203 bl_203 br_203 wl_173 vdd gnd cell_6t
Xbit_r174_c203 bl_203 br_203 wl_174 vdd gnd cell_6t
Xbit_r175_c203 bl_203 br_203 wl_175 vdd gnd cell_6t
Xbit_r176_c203 bl_203 br_203 wl_176 vdd gnd cell_6t
Xbit_r177_c203 bl_203 br_203 wl_177 vdd gnd cell_6t
Xbit_r178_c203 bl_203 br_203 wl_178 vdd gnd cell_6t
Xbit_r179_c203 bl_203 br_203 wl_179 vdd gnd cell_6t
Xbit_r180_c203 bl_203 br_203 wl_180 vdd gnd cell_6t
Xbit_r181_c203 bl_203 br_203 wl_181 vdd gnd cell_6t
Xbit_r182_c203 bl_203 br_203 wl_182 vdd gnd cell_6t
Xbit_r183_c203 bl_203 br_203 wl_183 vdd gnd cell_6t
Xbit_r184_c203 bl_203 br_203 wl_184 vdd gnd cell_6t
Xbit_r185_c203 bl_203 br_203 wl_185 vdd gnd cell_6t
Xbit_r186_c203 bl_203 br_203 wl_186 vdd gnd cell_6t
Xbit_r187_c203 bl_203 br_203 wl_187 vdd gnd cell_6t
Xbit_r188_c203 bl_203 br_203 wl_188 vdd gnd cell_6t
Xbit_r189_c203 bl_203 br_203 wl_189 vdd gnd cell_6t
Xbit_r190_c203 bl_203 br_203 wl_190 vdd gnd cell_6t
Xbit_r191_c203 bl_203 br_203 wl_191 vdd gnd cell_6t
Xbit_r192_c203 bl_203 br_203 wl_192 vdd gnd cell_6t
Xbit_r193_c203 bl_203 br_203 wl_193 vdd gnd cell_6t
Xbit_r194_c203 bl_203 br_203 wl_194 vdd gnd cell_6t
Xbit_r195_c203 bl_203 br_203 wl_195 vdd gnd cell_6t
Xbit_r196_c203 bl_203 br_203 wl_196 vdd gnd cell_6t
Xbit_r197_c203 bl_203 br_203 wl_197 vdd gnd cell_6t
Xbit_r198_c203 bl_203 br_203 wl_198 vdd gnd cell_6t
Xbit_r199_c203 bl_203 br_203 wl_199 vdd gnd cell_6t
Xbit_r200_c203 bl_203 br_203 wl_200 vdd gnd cell_6t
Xbit_r201_c203 bl_203 br_203 wl_201 vdd gnd cell_6t
Xbit_r202_c203 bl_203 br_203 wl_202 vdd gnd cell_6t
Xbit_r203_c203 bl_203 br_203 wl_203 vdd gnd cell_6t
Xbit_r204_c203 bl_203 br_203 wl_204 vdd gnd cell_6t
Xbit_r205_c203 bl_203 br_203 wl_205 vdd gnd cell_6t
Xbit_r206_c203 bl_203 br_203 wl_206 vdd gnd cell_6t
Xbit_r207_c203 bl_203 br_203 wl_207 vdd gnd cell_6t
Xbit_r208_c203 bl_203 br_203 wl_208 vdd gnd cell_6t
Xbit_r209_c203 bl_203 br_203 wl_209 vdd gnd cell_6t
Xbit_r210_c203 bl_203 br_203 wl_210 vdd gnd cell_6t
Xbit_r211_c203 bl_203 br_203 wl_211 vdd gnd cell_6t
Xbit_r212_c203 bl_203 br_203 wl_212 vdd gnd cell_6t
Xbit_r213_c203 bl_203 br_203 wl_213 vdd gnd cell_6t
Xbit_r214_c203 bl_203 br_203 wl_214 vdd gnd cell_6t
Xbit_r215_c203 bl_203 br_203 wl_215 vdd gnd cell_6t
Xbit_r216_c203 bl_203 br_203 wl_216 vdd gnd cell_6t
Xbit_r217_c203 bl_203 br_203 wl_217 vdd gnd cell_6t
Xbit_r218_c203 bl_203 br_203 wl_218 vdd gnd cell_6t
Xbit_r219_c203 bl_203 br_203 wl_219 vdd gnd cell_6t
Xbit_r220_c203 bl_203 br_203 wl_220 vdd gnd cell_6t
Xbit_r221_c203 bl_203 br_203 wl_221 vdd gnd cell_6t
Xbit_r222_c203 bl_203 br_203 wl_222 vdd gnd cell_6t
Xbit_r223_c203 bl_203 br_203 wl_223 vdd gnd cell_6t
Xbit_r224_c203 bl_203 br_203 wl_224 vdd gnd cell_6t
Xbit_r225_c203 bl_203 br_203 wl_225 vdd gnd cell_6t
Xbit_r226_c203 bl_203 br_203 wl_226 vdd gnd cell_6t
Xbit_r227_c203 bl_203 br_203 wl_227 vdd gnd cell_6t
Xbit_r228_c203 bl_203 br_203 wl_228 vdd gnd cell_6t
Xbit_r229_c203 bl_203 br_203 wl_229 vdd gnd cell_6t
Xbit_r230_c203 bl_203 br_203 wl_230 vdd gnd cell_6t
Xbit_r231_c203 bl_203 br_203 wl_231 vdd gnd cell_6t
Xbit_r232_c203 bl_203 br_203 wl_232 vdd gnd cell_6t
Xbit_r233_c203 bl_203 br_203 wl_233 vdd gnd cell_6t
Xbit_r234_c203 bl_203 br_203 wl_234 vdd gnd cell_6t
Xbit_r235_c203 bl_203 br_203 wl_235 vdd gnd cell_6t
Xbit_r236_c203 bl_203 br_203 wl_236 vdd gnd cell_6t
Xbit_r237_c203 bl_203 br_203 wl_237 vdd gnd cell_6t
Xbit_r238_c203 bl_203 br_203 wl_238 vdd gnd cell_6t
Xbit_r239_c203 bl_203 br_203 wl_239 vdd gnd cell_6t
Xbit_r240_c203 bl_203 br_203 wl_240 vdd gnd cell_6t
Xbit_r241_c203 bl_203 br_203 wl_241 vdd gnd cell_6t
Xbit_r242_c203 bl_203 br_203 wl_242 vdd gnd cell_6t
Xbit_r243_c203 bl_203 br_203 wl_243 vdd gnd cell_6t
Xbit_r244_c203 bl_203 br_203 wl_244 vdd gnd cell_6t
Xbit_r245_c203 bl_203 br_203 wl_245 vdd gnd cell_6t
Xbit_r246_c203 bl_203 br_203 wl_246 vdd gnd cell_6t
Xbit_r247_c203 bl_203 br_203 wl_247 vdd gnd cell_6t
Xbit_r248_c203 bl_203 br_203 wl_248 vdd gnd cell_6t
Xbit_r249_c203 bl_203 br_203 wl_249 vdd gnd cell_6t
Xbit_r250_c203 bl_203 br_203 wl_250 vdd gnd cell_6t
Xbit_r251_c203 bl_203 br_203 wl_251 vdd gnd cell_6t
Xbit_r252_c203 bl_203 br_203 wl_252 vdd gnd cell_6t
Xbit_r253_c203 bl_203 br_203 wl_253 vdd gnd cell_6t
Xbit_r254_c203 bl_203 br_203 wl_254 vdd gnd cell_6t
Xbit_r255_c203 bl_203 br_203 wl_255 vdd gnd cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd cell_6t
Xbit_r1_c204 bl_204 br_204 wl_1 vdd gnd cell_6t
Xbit_r2_c204 bl_204 br_204 wl_2 vdd gnd cell_6t
Xbit_r3_c204 bl_204 br_204 wl_3 vdd gnd cell_6t
Xbit_r4_c204 bl_204 br_204 wl_4 vdd gnd cell_6t
Xbit_r5_c204 bl_204 br_204 wl_5 vdd gnd cell_6t
Xbit_r6_c204 bl_204 br_204 wl_6 vdd gnd cell_6t
Xbit_r7_c204 bl_204 br_204 wl_7 vdd gnd cell_6t
Xbit_r8_c204 bl_204 br_204 wl_8 vdd gnd cell_6t
Xbit_r9_c204 bl_204 br_204 wl_9 vdd gnd cell_6t
Xbit_r10_c204 bl_204 br_204 wl_10 vdd gnd cell_6t
Xbit_r11_c204 bl_204 br_204 wl_11 vdd gnd cell_6t
Xbit_r12_c204 bl_204 br_204 wl_12 vdd gnd cell_6t
Xbit_r13_c204 bl_204 br_204 wl_13 vdd gnd cell_6t
Xbit_r14_c204 bl_204 br_204 wl_14 vdd gnd cell_6t
Xbit_r15_c204 bl_204 br_204 wl_15 vdd gnd cell_6t
Xbit_r16_c204 bl_204 br_204 wl_16 vdd gnd cell_6t
Xbit_r17_c204 bl_204 br_204 wl_17 vdd gnd cell_6t
Xbit_r18_c204 bl_204 br_204 wl_18 vdd gnd cell_6t
Xbit_r19_c204 bl_204 br_204 wl_19 vdd gnd cell_6t
Xbit_r20_c204 bl_204 br_204 wl_20 vdd gnd cell_6t
Xbit_r21_c204 bl_204 br_204 wl_21 vdd gnd cell_6t
Xbit_r22_c204 bl_204 br_204 wl_22 vdd gnd cell_6t
Xbit_r23_c204 bl_204 br_204 wl_23 vdd gnd cell_6t
Xbit_r24_c204 bl_204 br_204 wl_24 vdd gnd cell_6t
Xbit_r25_c204 bl_204 br_204 wl_25 vdd gnd cell_6t
Xbit_r26_c204 bl_204 br_204 wl_26 vdd gnd cell_6t
Xbit_r27_c204 bl_204 br_204 wl_27 vdd gnd cell_6t
Xbit_r28_c204 bl_204 br_204 wl_28 vdd gnd cell_6t
Xbit_r29_c204 bl_204 br_204 wl_29 vdd gnd cell_6t
Xbit_r30_c204 bl_204 br_204 wl_30 vdd gnd cell_6t
Xbit_r31_c204 bl_204 br_204 wl_31 vdd gnd cell_6t
Xbit_r32_c204 bl_204 br_204 wl_32 vdd gnd cell_6t
Xbit_r33_c204 bl_204 br_204 wl_33 vdd gnd cell_6t
Xbit_r34_c204 bl_204 br_204 wl_34 vdd gnd cell_6t
Xbit_r35_c204 bl_204 br_204 wl_35 vdd gnd cell_6t
Xbit_r36_c204 bl_204 br_204 wl_36 vdd gnd cell_6t
Xbit_r37_c204 bl_204 br_204 wl_37 vdd gnd cell_6t
Xbit_r38_c204 bl_204 br_204 wl_38 vdd gnd cell_6t
Xbit_r39_c204 bl_204 br_204 wl_39 vdd gnd cell_6t
Xbit_r40_c204 bl_204 br_204 wl_40 vdd gnd cell_6t
Xbit_r41_c204 bl_204 br_204 wl_41 vdd gnd cell_6t
Xbit_r42_c204 bl_204 br_204 wl_42 vdd gnd cell_6t
Xbit_r43_c204 bl_204 br_204 wl_43 vdd gnd cell_6t
Xbit_r44_c204 bl_204 br_204 wl_44 vdd gnd cell_6t
Xbit_r45_c204 bl_204 br_204 wl_45 vdd gnd cell_6t
Xbit_r46_c204 bl_204 br_204 wl_46 vdd gnd cell_6t
Xbit_r47_c204 bl_204 br_204 wl_47 vdd gnd cell_6t
Xbit_r48_c204 bl_204 br_204 wl_48 vdd gnd cell_6t
Xbit_r49_c204 bl_204 br_204 wl_49 vdd gnd cell_6t
Xbit_r50_c204 bl_204 br_204 wl_50 vdd gnd cell_6t
Xbit_r51_c204 bl_204 br_204 wl_51 vdd gnd cell_6t
Xbit_r52_c204 bl_204 br_204 wl_52 vdd gnd cell_6t
Xbit_r53_c204 bl_204 br_204 wl_53 vdd gnd cell_6t
Xbit_r54_c204 bl_204 br_204 wl_54 vdd gnd cell_6t
Xbit_r55_c204 bl_204 br_204 wl_55 vdd gnd cell_6t
Xbit_r56_c204 bl_204 br_204 wl_56 vdd gnd cell_6t
Xbit_r57_c204 bl_204 br_204 wl_57 vdd gnd cell_6t
Xbit_r58_c204 bl_204 br_204 wl_58 vdd gnd cell_6t
Xbit_r59_c204 bl_204 br_204 wl_59 vdd gnd cell_6t
Xbit_r60_c204 bl_204 br_204 wl_60 vdd gnd cell_6t
Xbit_r61_c204 bl_204 br_204 wl_61 vdd gnd cell_6t
Xbit_r62_c204 bl_204 br_204 wl_62 vdd gnd cell_6t
Xbit_r63_c204 bl_204 br_204 wl_63 vdd gnd cell_6t
Xbit_r64_c204 bl_204 br_204 wl_64 vdd gnd cell_6t
Xbit_r65_c204 bl_204 br_204 wl_65 vdd gnd cell_6t
Xbit_r66_c204 bl_204 br_204 wl_66 vdd gnd cell_6t
Xbit_r67_c204 bl_204 br_204 wl_67 vdd gnd cell_6t
Xbit_r68_c204 bl_204 br_204 wl_68 vdd gnd cell_6t
Xbit_r69_c204 bl_204 br_204 wl_69 vdd gnd cell_6t
Xbit_r70_c204 bl_204 br_204 wl_70 vdd gnd cell_6t
Xbit_r71_c204 bl_204 br_204 wl_71 vdd gnd cell_6t
Xbit_r72_c204 bl_204 br_204 wl_72 vdd gnd cell_6t
Xbit_r73_c204 bl_204 br_204 wl_73 vdd gnd cell_6t
Xbit_r74_c204 bl_204 br_204 wl_74 vdd gnd cell_6t
Xbit_r75_c204 bl_204 br_204 wl_75 vdd gnd cell_6t
Xbit_r76_c204 bl_204 br_204 wl_76 vdd gnd cell_6t
Xbit_r77_c204 bl_204 br_204 wl_77 vdd gnd cell_6t
Xbit_r78_c204 bl_204 br_204 wl_78 vdd gnd cell_6t
Xbit_r79_c204 bl_204 br_204 wl_79 vdd gnd cell_6t
Xbit_r80_c204 bl_204 br_204 wl_80 vdd gnd cell_6t
Xbit_r81_c204 bl_204 br_204 wl_81 vdd gnd cell_6t
Xbit_r82_c204 bl_204 br_204 wl_82 vdd gnd cell_6t
Xbit_r83_c204 bl_204 br_204 wl_83 vdd gnd cell_6t
Xbit_r84_c204 bl_204 br_204 wl_84 vdd gnd cell_6t
Xbit_r85_c204 bl_204 br_204 wl_85 vdd gnd cell_6t
Xbit_r86_c204 bl_204 br_204 wl_86 vdd gnd cell_6t
Xbit_r87_c204 bl_204 br_204 wl_87 vdd gnd cell_6t
Xbit_r88_c204 bl_204 br_204 wl_88 vdd gnd cell_6t
Xbit_r89_c204 bl_204 br_204 wl_89 vdd gnd cell_6t
Xbit_r90_c204 bl_204 br_204 wl_90 vdd gnd cell_6t
Xbit_r91_c204 bl_204 br_204 wl_91 vdd gnd cell_6t
Xbit_r92_c204 bl_204 br_204 wl_92 vdd gnd cell_6t
Xbit_r93_c204 bl_204 br_204 wl_93 vdd gnd cell_6t
Xbit_r94_c204 bl_204 br_204 wl_94 vdd gnd cell_6t
Xbit_r95_c204 bl_204 br_204 wl_95 vdd gnd cell_6t
Xbit_r96_c204 bl_204 br_204 wl_96 vdd gnd cell_6t
Xbit_r97_c204 bl_204 br_204 wl_97 vdd gnd cell_6t
Xbit_r98_c204 bl_204 br_204 wl_98 vdd gnd cell_6t
Xbit_r99_c204 bl_204 br_204 wl_99 vdd gnd cell_6t
Xbit_r100_c204 bl_204 br_204 wl_100 vdd gnd cell_6t
Xbit_r101_c204 bl_204 br_204 wl_101 vdd gnd cell_6t
Xbit_r102_c204 bl_204 br_204 wl_102 vdd gnd cell_6t
Xbit_r103_c204 bl_204 br_204 wl_103 vdd gnd cell_6t
Xbit_r104_c204 bl_204 br_204 wl_104 vdd gnd cell_6t
Xbit_r105_c204 bl_204 br_204 wl_105 vdd gnd cell_6t
Xbit_r106_c204 bl_204 br_204 wl_106 vdd gnd cell_6t
Xbit_r107_c204 bl_204 br_204 wl_107 vdd gnd cell_6t
Xbit_r108_c204 bl_204 br_204 wl_108 vdd gnd cell_6t
Xbit_r109_c204 bl_204 br_204 wl_109 vdd gnd cell_6t
Xbit_r110_c204 bl_204 br_204 wl_110 vdd gnd cell_6t
Xbit_r111_c204 bl_204 br_204 wl_111 vdd gnd cell_6t
Xbit_r112_c204 bl_204 br_204 wl_112 vdd gnd cell_6t
Xbit_r113_c204 bl_204 br_204 wl_113 vdd gnd cell_6t
Xbit_r114_c204 bl_204 br_204 wl_114 vdd gnd cell_6t
Xbit_r115_c204 bl_204 br_204 wl_115 vdd gnd cell_6t
Xbit_r116_c204 bl_204 br_204 wl_116 vdd gnd cell_6t
Xbit_r117_c204 bl_204 br_204 wl_117 vdd gnd cell_6t
Xbit_r118_c204 bl_204 br_204 wl_118 vdd gnd cell_6t
Xbit_r119_c204 bl_204 br_204 wl_119 vdd gnd cell_6t
Xbit_r120_c204 bl_204 br_204 wl_120 vdd gnd cell_6t
Xbit_r121_c204 bl_204 br_204 wl_121 vdd gnd cell_6t
Xbit_r122_c204 bl_204 br_204 wl_122 vdd gnd cell_6t
Xbit_r123_c204 bl_204 br_204 wl_123 vdd gnd cell_6t
Xbit_r124_c204 bl_204 br_204 wl_124 vdd gnd cell_6t
Xbit_r125_c204 bl_204 br_204 wl_125 vdd gnd cell_6t
Xbit_r126_c204 bl_204 br_204 wl_126 vdd gnd cell_6t
Xbit_r127_c204 bl_204 br_204 wl_127 vdd gnd cell_6t
Xbit_r128_c204 bl_204 br_204 wl_128 vdd gnd cell_6t
Xbit_r129_c204 bl_204 br_204 wl_129 vdd gnd cell_6t
Xbit_r130_c204 bl_204 br_204 wl_130 vdd gnd cell_6t
Xbit_r131_c204 bl_204 br_204 wl_131 vdd gnd cell_6t
Xbit_r132_c204 bl_204 br_204 wl_132 vdd gnd cell_6t
Xbit_r133_c204 bl_204 br_204 wl_133 vdd gnd cell_6t
Xbit_r134_c204 bl_204 br_204 wl_134 vdd gnd cell_6t
Xbit_r135_c204 bl_204 br_204 wl_135 vdd gnd cell_6t
Xbit_r136_c204 bl_204 br_204 wl_136 vdd gnd cell_6t
Xbit_r137_c204 bl_204 br_204 wl_137 vdd gnd cell_6t
Xbit_r138_c204 bl_204 br_204 wl_138 vdd gnd cell_6t
Xbit_r139_c204 bl_204 br_204 wl_139 vdd gnd cell_6t
Xbit_r140_c204 bl_204 br_204 wl_140 vdd gnd cell_6t
Xbit_r141_c204 bl_204 br_204 wl_141 vdd gnd cell_6t
Xbit_r142_c204 bl_204 br_204 wl_142 vdd gnd cell_6t
Xbit_r143_c204 bl_204 br_204 wl_143 vdd gnd cell_6t
Xbit_r144_c204 bl_204 br_204 wl_144 vdd gnd cell_6t
Xbit_r145_c204 bl_204 br_204 wl_145 vdd gnd cell_6t
Xbit_r146_c204 bl_204 br_204 wl_146 vdd gnd cell_6t
Xbit_r147_c204 bl_204 br_204 wl_147 vdd gnd cell_6t
Xbit_r148_c204 bl_204 br_204 wl_148 vdd gnd cell_6t
Xbit_r149_c204 bl_204 br_204 wl_149 vdd gnd cell_6t
Xbit_r150_c204 bl_204 br_204 wl_150 vdd gnd cell_6t
Xbit_r151_c204 bl_204 br_204 wl_151 vdd gnd cell_6t
Xbit_r152_c204 bl_204 br_204 wl_152 vdd gnd cell_6t
Xbit_r153_c204 bl_204 br_204 wl_153 vdd gnd cell_6t
Xbit_r154_c204 bl_204 br_204 wl_154 vdd gnd cell_6t
Xbit_r155_c204 bl_204 br_204 wl_155 vdd gnd cell_6t
Xbit_r156_c204 bl_204 br_204 wl_156 vdd gnd cell_6t
Xbit_r157_c204 bl_204 br_204 wl_157 vdd gnd cell_6t
Xbit_r158_c204 bl_204 br_204 wl_158 vdd gnd cell_6t
Xbit_r159_c204 bl_204 br_204 wl_159 vdd gnd cell_6t
Xbit_r160_c204 bl_204 br_204 wl_160 vdd gnd cell_6t
Xbit_r161_c204 bl_204 br_204 wl_161 vdd gnd cell_6t
Xbit_r162_c204 bl_204 br_204 wl_162 vdd gnd cell_6t
Xbit_r163_c204 bl_204 br_204 wl_163 vdd gnd cell_6t
Xbit_r164_c204 bl_204 br_204 wl_164 vdd gnd cell_6t
Xbit_r165_c204 bl_204 br_204 wl_165 vdd gnd cell_6t
Xbit_r166_c204 bl_204 br_204 wl_166 vdd gnd cell_6t
Xbit_r167_c204 bl_204 br_204 wl_167 vdd gnd cell_6t
Xbit_r168_c204 bl_204 br_204 wl_168 vdd gnd cell_6t
Xbit_r169_c204 bl_204 br_204 wl_169 vdd gnd cell_6t
Xbit_r170_c204 bl_204 br_204 wl_170 vdd gnd cell_6t
Xbit_r171_c204 bl_204 br_204 wl_171 vdd gnd cell_6t
Xbit_r172_c204 bl_204 br_204 wl_172 vdd gnd cell_6t
Xbit_r173_c204 bl_204 br_204 wl_173 vdd gnd cell_6t
Xbit_r174_c204 bl_204 br_204 wl_174 vdd gnd cell_6t
Xbit_r175_c204 bl_204 br_204 wl_175 vdd gnd cell_6t
Xbit_r176_c204 bl_204 br_204 wl_176 vdd gnd cell_6t
Xbit_r177_c204 bl_204 br_204 wl_177 vdd gnd cell_6t
Xbit_r178_c204 bl_204 br_204 wl_178 vdd gnd cell_6t
Xbit_r179_c204 bl_204 br_204 wl_179 vdd gnd cell_6t
Xbit_r180_c204 bl_204 br_204 wl_180 vdd gnd cell_6t
Xbit_r181_c204 bl_204 br_204 wl_181 vdd gnd cell_6t
Xbit_r182_c204 bl_204 br_204 wl_182 vdd gnd cell_6t
Xbit_r183_c204 bl_204 br_204 wl_183 vdd gnd cell_6t
Xbit_r184_c204 bl_204 br_204 wl_184 vdd gnd cell_6t
Xbit_r185_c204 bl_204 br_204 wl_185 vdd gnd cell_6t
Xbit_r186_c204 bl_204 br_204 wl_186 vdd gnd cell_6t
Xbit_r187_c204 bl_204 br_204 wl_187 vdd gnd cell_6t
Xbit_r188_c204 bl_204 br_204 wl_188 vdd gnd cell_6t
Xbit_r189_c204 bl_204 br_204 wl_189 vdd gnd cell_6t
Xbit_r190_c204 bl_204 br_204 wl_190 vdd gnd cell_6t
Xbit_r191_c204 bl_204 br_204 wl_191 vdd gnd cell_6t
Xbit_r192_c204 bl_204 br_204 wl_192 vdd gnd cell_6t
Xbit_r193_c204 bl_204 br_204 wl_193 vdd gnd cell_6t
Xbit_r194_c204 bl_204 br_204 wl_194 vdd gnd cell_6t
Xbit_r195_c204 bl_204 br_204 wl_195 vdd gnd cell_6t
Xbit_r196_c204 bl_204 br_204 wl_196 vdd gnd cell_6t
Xbit_r197_c204 bl_204 br_204 wl_197 vdd gnd cell_6t
Xbit_r198_c204 bl_204 br_204 wl_198 vdd gnd cell_6t
Xbit_r199_c204 bl_204 br_204 wl_199 vdd gnd cell_6t
Xbit_r200_c204 bl_204 br_204 wl_200 vdd gnd cell_6t
Xbit_r201_c204 bl_204 br_204 wl_201 vdd gnd cell_6t
Xbit_r202_c204 bl_204 br_204 wl_202 vdd gnd cell_6t
Xbit_r203_c204 bl_204 br_204 wl_203 vdd gnd cell_6t
Xbit_r204_c204 bl_204 br_204 wl_204 vdd gnd cell_6t
Xbit_r205_c204 bl_204 br_204 wl_205 vdd gnd cell_6t
Xbit_r206_c204 bl_204 br_204 wl_206 vdd gnd cell_6t
Xbit_r207_c204 bl_204 br_204 wl_207 vdd gnd cell_6t
Xbit_r208_c204 bl_204 br_204 wl_208 vdd gnd cell_6t
Xbit_r209_c204 bl_204 br_204 wl_209 vdd gnd cell_6t
Xbit_r210_c204 bl_204 br_204 wl_210 vdd gnd cell_6t
Xbit_r211_c204 bl_204 br_204 wl_211 vdd gnd cell_6t
Xbit_r212_c204 bl_204 br_204 wl_212 vdd gnd cell_6t
Xbit_r213_c204 bl_204 br_204 wl_213 vdd gnd cell_6t
Xbit_r214_c204 bl_204 br_204 wl_214 vdd gnd cell_6t
Xbit_r215_c204 bl_204 br_204 wl_215 vdd gnd cell_6t
Xbit_r216_c204 bl_204 br_204 wl_216 vdd gnd cell_6t
Xbit_r217_c204 bl_204 br_204 wl_217 vdd gnd cell_6t
Xbit_r218_c204 bl_204 br_204 wl_218 vdd gnd cell_6t
Xbit_r219_c204 bl_204 br_204 wl_219 vdd gnd cell_6t
Xbit_r220_c204 bl_204 br_204 wl_220 vdd gnd cell_6t
Xbit_r221_c204 bl_204 br_204 wl_221 vdd gnd cell_6t
Xbit_r222_c204 bl_204 br_204 wl_222 vdd gnd cell_6t
Xbit_r223_c204 bl_204 br_204 wl_223 vdd gnd cell_6t
Xbit_r224_c204 bl_204 br_204 wl_224 vdd gnd cell_6t
Xbit_r225_c204 bl_204 br_204 wl_225 vdd gnd cell_6t
Xbit_r226_c204 bl_204 br_204 wl_226 vdd gnd cell_6t
Xbit_r227_c204 bl_204 br_204 wl_227 vdd gnd cell_6t
Xbit_r228_c204 bl_204 br_204 wl_228 vdd gnd cell_6t
Xbit_r229_c204 bl_204 br_204 wl_229 vdd gnd cell_6t
Xbit_r230_c204 bl_204 br_204 wl_230 vdd gnd cell_6t
Xbit_r231_c204 bl_204 br_204 wl_231 vdd gnd cell_6t
Xbit_r232_c204 bl_204 br_204 wl_232 vdd gnd cell_6t
Xbit_r233_c204 bl_204 br_204 wl_233 vdd gnd cell_6t
Xbit_r234_c204 bl_204 br_204 wl_234 vdd gnd cell_6t
Xbit_r235_c204 bl_204 br_204 wl_235 vdd gnd cell_6t
Xbit_r236_c204 bl_204 br_204 wl_236 vdd gnd cell_6t
Xbit_r237_c204 bl_204 br_204 wl_237 vdd gnd cell_6t
Xbit_r238_c204 bl_204 br_204 wl_238 vdd gnd cell_6t
Xbit_r239_c204 bl_204 br_204 wl_239 vdd gnd cell_6t
Xbit_r240_c204 bl_204 br_204 wl_240 vdd gnd cell_6t
Xbit_r241_c204 bl_204 br_204 wl_241 vdd gnd cell_6t
Xbit_r242_c204 bl_204 br_204 wl_242 vdd gnd cell_6t
Xbit_r243_c204 bl_204 br_204 wl_243 vdd gnd cell_6t
Xbit_r244_c204 bl_204 br_204 wl_244 vdd gnd cell_6t
Xbit_r245_c204 bl_204 br_204 wl_245 vdd gnd cell_6t
Xbit_r246_c204 bl_204 br_204 wl_246 vdd gnd cell_6t
Xbit_r247_c204 bl_204 br_204 wl_247 vdd gnd cell_6t
Xbit_r248_c204 bl_204 br_204 wl_248 vdd gnd cell_6t
Xbit_r249_c204 bl_204 br_204 wl_249 vdd gnd cell_6t
Xbit_r250_c204 bl_204 br_204 wl_250 vdd gnd cell_6t
Xbit_r251_c204 bl_204 br_204 wl_251 vdd gnd cell_6t
Xbit_r252_c204 bl_204 br_204 wl_252 vdd gnd cell_6t
Xbit_r253_c204 bl_204 br_204 wl_253 vdd gnd cell_6t
Xbit_r254_c204 bl_204 br_204 wl_254 vdd gnd cell_6t
Xbit_r255_c204 bl_204 br_204 wl_255 vdd gnd cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd cell_6t
Xbit_r1_c205 bl_205 br_205 wl_1 vdd gnd cell_6t
Xbit_r2_c205 bl_205 br_205 wl_2 vdd gnd cell_6t
Xbit_r3_c205 bl_205 br_205 wl_3 vdd gnd cell_6t
Xbit_r4_c205 bl_205 br_205 wl_4 vdd gnd cell_6t
Xbit_r5_c205 bl_205 br_205 wl_5 vdd gnd cell_6t
Xbit_r6_c205 bl_205 br_205 wl_6 vdd gnd cell_6t
Xbit_r7_c205 bl_205 br_205 wl_7 vdd gnd cell_6t
Xbit_r8_c205 bl_205 br_205 wl_8 vdd gnd cell_6t
Xbit_r9_c205 bl_205 br_205 wl_9 vdd gnd cell_6t
Xbit_r10_c205 bl_205 br_205 wl_10 vdd gnd cell_6t
Xbit_r11_c205 bl_205 br_205 wl_11 vdd gnd cell_6t
Xbit_r12_c205 bl_205 br_205 wl_12 vdd gnd cell_6t
Xbit_r13_c205 bl_205 br_205 wl_13 vdd gnd cell_6t
Xbit_r14_c205 bl_205 br_205 wl_14 vdd gnd cell_6t
Xbit_r15_c205 bl_205 br_205 wl_15 vdd gnd cell_6t
Xbit_r16_c205 bl_205 br_205 wl_16 vdd gnd cell_6t
Xbit_r17_c205 bl_205 br_205 wl_17 vdd gnd cell_6t
Xbit_r18_c205 bl_205 br_205 wl_18 vdd gnd cell_6t
Xbit_r19_c205 bl_205 br_205 wl_19 vdd gnd cell_6t
Xbit_r20_c205 bl_205 br_205 wl_20 vdd gnd cell_6t
Xbit_r21_c205 bl_205 br_205 wl_21 vdd gnd cell_6t
Xbit_r22_c205 bl_205 br_205 wl_22 vdd gnd cell_6t
Xbit_r23_c205 bl_205 br_205 wl_23 vdd gnd cell_6t
Xbit_r24_c205 bl_205 br_205 wl_24 vdd gnd cell_6t
Xbit_r25_c205 bl_205 br_205 wl_25 vdd gnd cell_6t
Xbit_r26_c205 bl_205 br_205 wl_26 vdd gnd cell_6t
Xbit_r27_c205 bl_205 br_205 wl_27 vdd gnd cell_6t
Xbit_r28_c205 bl_205 br_205 wl_28 vdd gnd cell_6t
Xbit_r29_c205 bl_205 br_205 wl_29 vdd gnd cell_6t
Xbit_r30_c205 bl_205 br_205 wl_30 vdd gnd cell_6t
Xbit_r31_c205 bl_205 br_205 wl_31 vdd gnd cell_6t
Xbit_r32_c205 bl_205 br_205 wl_32 vdd gnd cell_6t
Xbit_r33_c205 bl_205 br_205 wl_33 vdd gnd cell_6t
Xbit_r34_c205 bl_205 br_205 wl_34 vdd gnd cell_6t
Xbit_r35_c205 bl_205 br_205 wl_35 vdd gnd cell_6t
Xbit_r36_c205 bl_205 br_205 wl_36 vdd gnd cell_6t
Xbit_r37_c205 bl_205 br_205 wl_37 vdd gnd cell_6t
Xbit_r38_c205 bl_205 br_205 wl_38 vdd gnd cell_6t
Xbit_r39_c205 bl_205 br_205 wl_39 vdd gnd cell_6t
Xbit_r40_c205 bl_205 br_205 wl_40 vdd gnd cell_6t
Xbit_r41_c205 bl_205 br_205 wl_41 vdd gnd cell_6t
Xbit_r42_c205 bl_205 br_205 wl_42 vdd gnd cell_6t
Xbit_r43_c205 bl_205 br_205 wl_43 vdd gnd cell_6t
Xbit_r44_c205 bl_205 br_205 wl_44 vdd gnd cell_6t
Xbit_r45_c205 bl_205 br_205 wl_45 vdd gnd cell_6t
Xbit_r46_c205 bl_205 br_205 wl_46 vdd gnd cell_6t
Xbit_r47_c205 bl_205 br_205 wl_47 vdd gnd cell_6t
Xbit_r48_c205 bl_205 br_205 wl_48 vdd gnd cell_6t
Xbit_r49_c205 bl_205 br_205 wl_49 vdd gnd cell_6t
Xbit_r50_c205 bl_205 br_205 wl_50 vdd gnd cell_6t
Xbit_r51_c205 bl_205 br_205 wl_51 vdd gnd cell_6t
Xbit_r52_c205 bl_205 br_205 wl_52 vdd gnd cell_6t
Xbit_r53_c205 bl_205 br_205 wl_53 vdd gnd cell_6t
Xbit_r54_c205 bl_205 br_205 wl_54 vdd gnd cell_6t
Xbit_r55_c205 bl_205 br_205 wl_55 vdd gnd cell_6t
Xbit_r56_c205 bl_205 br_205 wl_56 vdd gnd cell_6t
Xbit_r57_c205 bl_205 br_205 wl_57 vdd gnd cell_6t
Xbit_r58_c205 bl_205 br_205 wl_58 vdd gnd cell_6t
Xbit_r59_c205 bl_205 br_205 wl_59 vdd gnd cell_6t
Xbit_r60_c205 bl_205 br_205 wl_60 vdd gnd cell_6t
Xbit_r61_c205 bl_205 br_205 wl_61 vdd gnd cell_6t
Xbit_r62_c205 bl_205 br_205 wl_62 vdd gnd cell_6t
Xbit_r63_c205 bl_205 br_205 wl_63 vdd gnd cell_6t
Xbit_r64_c205 bl_205 br_205 wl_64 vdd gnd cell_6t
Xbit_r65_c205 bl_205 br_205 wl_65 vdd gnd cell_6t
Xbit_r66_c205 bl_205 br_205 wl_66 vdd gnd cell_6t
Xbit_r67_c205 bl_205 br_205 wl_67 vdd gnd cell_6t
Xbit_r68_c205 bl_205 br_205 wl_68 vdd gnd cell_6t
Xbit_r69_c205 bl_205 br_205 wl_69 vdd gnd cell_6t
Xbit_r70_c205 bl_205 br_205 wl_70 vdd gnd cell_6t
Xbit_r71_c205 bl_205 br_205 wl_71 vdd gnd cell_6t
Xbit_r72_c205 bl_205 br_205 wl_72 vdd gnd cell_6t
Xbit_r73_c205 bl_205 br_205 wl_73 vdd gnd cell_6t
Xbit_r74_c205 bl_205 br_205 wl_74 vdd gnd cell_6t
Xbit_r75_c205 bl_205 br_205 wl_75 vdd gnd cell_6t
Xbit_r76_c205 bl_205 br_205 wl_76 vdd gnd cell_6t
Xbit_r77_c205 bl_205 br_205 wl_77 vdd gnd cell_6t
Xbit_r78_c205 bl_205 br_205 wl_78 vdd gnd cell_6t
Xbit_r79_c205 bl_205 br_205 wl_79 vdd gnd cell_6t
Xbit_r80_c205 bl_205 br_205 wl_80 vdd gnd cell_6t
Xbit_r81_c205 bl_205 br_205 wl_81 vdd gnd cell_6t
Xbit_r82_c205 bl_205 br_205 wl_82 vdd gnd cell_6t
Xbit_r83_c205 bl_205 br_205 wl_83 vdd gnd cell_6t
Xbit_r84_c205 bl_205 br_205 wl_84 vdd gnd cell_6t
Xbit_r85_c205 bl_205 br_205 wl_85 vdd gnd cell_6t
Xbit_r86_c205 bl_205 br_205 wl_86 vdd gnd cell_6t
Xbit_r87_c205 bl_205 br_205 wl_87 vdd gnd cell_6t
Xbit_r88_c205 bl_205 br_205 wl_88 vdd gnd cell_6t
Xbit_r89_c205 bl_205 br_205 wl_89 vdd gnd cell_6t
Xbit_r90_c205 bl_205 br_205 wl_90 vdd gnd cell_6t
Xbit_r91_c205 bl_205 br_205 wl_91 vdd gnd cell_6t
Xbit_r92_c205 bl_205 br_205 wl_92 vdd gnd cell_6t
Xbit_r93_c205 bl_205 br_205 wl_93 vdd gnd cell_6t
Xbit_r94_c205 bl_205 br_205 wl_94 vdd gnd cell_6t
Xbit_r95_c205 bl_205 br_205 wl_95 vdd gnd cell_6t
Xbit_r96_c205 bl_205 br_205 wl_96 vdd gnd cell_6t
Xbit_r97_c205 bl_205 br_205 wl_97 vdd gnd cell_6t
Xbit_r98_c205 bl_205 br_205 wl_98 vdd gnd cell_6t
Xbit_r99_c205 bl_205 br_205 wl_99 vdd gnd cell_6t
Xbit_r100_c205 bl_205 br_205 wl_100 vdd gnd cell_6t
Xbit_r101_c205 bl_205 br_205 wl_101 vdd gnd cell_6t
Xbit_r102_c205 bl_205 br_205 wl_102 vdd gnd cell_6t
Xbit_r103_c205 bl_205 br_205 wl_103 vdd gnd cell_6t
Xbit_r104_c205 bl_205 br_205 wl_104 vdd gnd cell_6t
Xbit_r105_c205 bl_205 br_205 wl_105 vdd gnd cell_6t
Xbit_r106_c205 bl_205 br_205 wl_106 vdd gnd cell_6t
Xbit_r107_c205 bl_205 br_205 wl_107 vdd gnd cell_6t
Xbit_r108_c205 bl_205 br_205 wl_108 vdd gnd cell_6t
Xbit_r109_c205 bl_205 br_205 wl_109 vdd gnd cell_6t
Xbit_r110_c205 bl_205 br_205 wl_110 vdd gnd cell_6t
Xbit_r111_c205 bl_205 br_205 wl_111 vdd gnd cell_6t
Xbit_r112_c205 bl_205 br_205 wl_112 vdd gnd cell_6t
Xbit_r113_c205 bl_205 br_205 wl_113 vdd gnd cell_6t
Xbit_r114_c205 bl_205 br_205 wl_114 vdd gnd cell_6t
Xbit_r115_c205 bl_205 br_205 wl_115 vdd gnd cell_6t
Xbit_r116_c205 bl_205 br_205 wl_116 vdd gnd cell_6t
Xbit_r117_c205 bl_205 br_205 wl_117 vdd gnd cell_6t
Xbit_r118_c205 bl_205 br_205 wl_118 vdd gnd cell_6t
Xbit_r119_c205 bl_205 br_205 wl_119 vdd gnd cell_6t
Xbit_r120_c205 bl_205 br_205 wl_120 vdd gnd cell_6t
Xbit_r121_c205 bl_205 br_205 wl_121 vdd gnd cell_6t
Xbit_r122_c205 bl_205 br_205 wl_122 vdd gnd cell_6t
Xbit_r123_c205 bl_205 br_205 wl_123 vdd gnd cell_6t
Xbit_r124_c205 bl_205 br_205 wl_124 vdd gnd cell_6t
Xbit_r125_c205 bl_205 br_205 wl_125 vdd gnd cell_6t
Xbit_r126_c205 bl_205 br_205 wl_126 vdd gnd cell_6t
Xbit_r127_c205 bl_205 br_205 wl_127 vdd gnd cell_6t
Xbit_r128_c205 bl_205 br_205 wl_128 vdd gnd cell_6t
Xbit_r129_c205 bl_205 br_205 wl_129 vdd gnd cell_6t
Xbit_r130_c205 bl_205 br_205 wl_130 vdd gnd cell_6t
Xbit_r131_c205 bl_205 br_205 wl_131 vdd gnd cell_6t
Xbit_r132_c205 bl_205 br_205 wl_132 vdd gnd cell_6t
Xbit_r133_c205 bl_205 br_205 wl_133 vdd gnd cell_6t
Xbit_r134_c205 bl_205 br_205 wl_134 vdd gnd cell_6t
Xbit_r135_c205 bl_205 br_205 wl_135 vdd gnd cell_6t
Xbit_r136_c205 bl_205 br_205 wl_136 vdd gnd cell_6t
Xbit_r137_c205 bl_205 br_205 wl_137 vdd gnd cell_6t
Xbit_r138_c205 bl_205 br_205 wl_138 vdd gnd cell_6t
Xbit_r139_c205 bl_205 br_205 wl_139 vdd gnd cell_6t
Xbit_r140_c205 bl_205 br_205 wl_140 vdd gnd cell_6t
Xbit_r141_c205 bl_205 br_205 wl_141 vdd gnd cell_6t
Xbit_r142_c205 bl_205 br_205 wl_142 vdd gnd cell_6t
Xbit_r143_c205 bl_205 br_205 wl_143 vdd gnd cell_6t
Xbit_r144_c205 bl_205 br_205 wl_144 vdd gnd cell_6t
Xbit_r145_c205 bl_205 br_205 wl_145 vdd gnd cell_6t
Xbit_r146_c205 bl_205 br_205 wl_146 vdd gnd cell_6t
Xbit_r147_c205 bl_205 br_205 wl_147 vdd gnd cell_6t
Xbit_r148_c205 bl_205 br_205 wl_148 vdd gnd cell_6t
Xbit_r149_c205 bl_205 br_205 wl_149 vdd gnd cell_6t
Xbit_r150_c205 bl_205 br_205 wl_150 vdd gnd cell_6t
Xbit_r151_c205 bl_205 br_205 wl_151 vdd gnd cell_6t
Xbit_r152_c205 bl_205 br_205 wl_152 vdd gnd cell_6t
Xbit_r153_c205 bl_205 br_205 wl_153 vdd gnd cell_6t
Xbit_r154_c205 bl_205 br_205 wl_154 vdd gnd cell_6t
Xbit_r155_c205 bl_205 br_205 wl_155 vdd gnd cell_6t
Xbit_r156_c205 bl_205 br_205 wl_156 vdd gnd cell_6t
Xbit_r157_c205 bl_205 br_205 wl_157 vdd gnd cell_6t
Xbit_r158_c205 bl_205 br_205 wl_158 vdd gnd cell_6t
Xbit_r159_c205 bl_205 br_205 wl_159 vdd gnd cell_6t
Xbit_r160_c205 bl_205 br_205 wl_160 vdd gnd cell_6t
Xbit_r161_c205 bl_205 br_205 wl_161 vdd gnd cell_6t
Xbit_r162_c205 bl_205 br_205 wl_162 vdd gnd cell_6t
Xbit_r163_c205 bl_205 br_205 wl_163 vdd gnd cell_6t
Xbit_r164_c205 bl_205 br_205 wl_164 vdd gnd cell_6t
Xbit_r165_c205 bl_205 br_205 wl_165 vdd gnd cell_6t
Xbit_r166_c205 bl_205 br_205 wl_166 vdd gnd cell_6t
Xbit_r167_c205 bl_205 br_205 wl_167 vdd gnd cell_6t
Xbit_r168_c205 bl_205 br_205 wl_168 vdd gnd cell_6t
Xbit_r169_c205 bl_205 br_205 wl_169 vdd gnd cell_6t
Xbit_r170_c205 bl_205 br_205 wl_170 vdd gnd cell_6t
Xbit_r171_c205 bl_205 br_205 wl_171 vdd gnd cell_6t
Xbit_r172_c205 bl_205 br_205 wl_172 vdd gnd cell_6t
Xbit_r173_c205 bl_205 br_205 wl_173 vdd gnd cell_6t
Xbit_r174_c205 bl_205 br_205 wl_174 vdd gnd cell_6t
Xbit_r175_c205 bl_205 br_205 wl_175 vdd gnd cell_6t
Xbit_r176_c205 bl_205 br_205 wl_176 vdd gnd cell_6t
Xbit_r177_c205 bl_205 br_205 wl_177 vdd gnd cell_6t
Xbit_r178_c205 bl_205 br_205 wl_178 vdd gnd cell_6t
Xbit_r179_c205 bl_205 br_205 wl_179 vdd gnd cell_6t
Xbit_r180_c205 bl_205 br_205 wl_180 vdd gnd cell_6t
Xbit_r181_c205 bl_205 br_205 wl_181 vdd gnd cell_6t
Xbit_r182_c205 bl_205 br_205 wl_182 vdd gnd cell_6t
Xbit_r183_c205 bl_205 br_205 wl_183 vdd gnd cell_6t
Xbit_r184_c205 bl_205 br_205 wl_184 vdd gnd cell_6t
Xbit_r185_c205 bl_205 br_205 wl_185 vdd gnd cell_6t
Xbit_r186_c205 bl_205 br_205 wl_186 vdd gnd cell_6t
Xbit_r187_c205 bl_205 br_205 wl_187 vdd gnd cell_6t
Xbit_r188_c205 bl_205 br_205 wl_188 vdd gnd cell_6t
Xbit_r189_c205 bl_205 br_205 wl_189 vdd gnd cell_6t
Xbit_r190_c205 bl_205 br_205 wl_190 vdd gnd cell_6t
Xbit_r191_c205 bl_205 br_205 wl_191 vdd gnd cell_6t
Xbit_r192_c205 bl_205 br_205 wl_192 vdd gnd cell_6t
Xbit_r193_c205 bl_205 br_205 wl_193 vdd gnd cell_6t
Xbit_r194_c205 bl_205 br_205 wl_194 vdd gnd cell_6t
Xbit_r195_c205 bl_205 br_205 wl_195 vdd gnd cell_6t
Xbit_r196_c205 bl_205 br_205 wl_196 vdd gnd cell_6t
Xbit_r197_c205 bl_205 br_205 wl_197 vdd gnd cell_6t
Xbit_r198_c205 bl_205 br_205 wl_198 vdd gnd cell_6t
Xbit_r199_c205 bl_205 br_205 wl_199 vdd gnd cell_6t
Xbit_r200_c205 bl_205 br_205 wl_200 vdd gnd cell_6t
Xbit_r201_c205 bl_205 br_205 wl_201 vdd gnd cell_6t
Xbit_r202_c205 bl_205 br_205 wl_202 vdd gnd cell_6t
Xbit_r203_c205 bl_205 br_205 wl_203 vdd gnd cell_6t
Xbit_r204_c205 bl_205 br_205 wl_204 vdd gnd cell_6t
Xbit_r205_c205 bl_205 br_205 wl_205 vdd gnd cell_6t
Xbit_r206_c205 bl_205 br_205 wl_206 vdd gnd cell_6t
Xbit_r207_c205 bl_205 br_205 wl_207 vdd gnd cell_6t
Xbit_r208_c205 bl_205 br_205 wl_208 vdd gnd cell_6t
Xbit_r209_c205 bl_205 br_205 wl_209 vdd gnd cell_6t
Xbit_r210_c205 bl_205 br_205 wl_210 vdd gnd cell_6t
Xbit_r211_c205 bl_205 br_205 wl_211 vdd gnd cell_6t
Xbit_r212_c205 bl_205 br_205 wl_212 vdd gnd cell_6t
Xbit_r213_c205 bl_205 br_205 wl_213 vdd gnd cell_6t
Xbit_r214_c205 bl_205 br_205 wl_214 vdd gnd cell_6t
Xbit_r215_c205 bl_205 br_205 wl_215 vdd gnd cell_6t
Xbit_r216_c205 bl_205 br_205 wl_216 vdd gnd cell_6t
Xbit_r217_c205 bl_205 br_205 wl_217 vdd gnd cell_6t
Xbit_r218_c205 bl_205 br_205 wl_218 vdd gnd cell_6t
Xbit_r219_c205 bl_205 br_205 wl_219 vdd gnd cell_6t
Xbit_r220_c205 bl_205 br_205 wl_220 vdd gnd cell_6t
Xbit_r221_c205 bl_205 br_205 wl_221 vdd gnd cell_6t
Xbit_r222_c205 bl_205 br_205 wl_222 vdd gnd cell_6t
Xbit_r223_c205 bl_205 br_205 wl_223 vdd gnd cell_6t
Xbit_r224_c205 bl_205 br_205 wl_224 vdd gnd cell_6t
Xbit_r225_c205 bl_205 br_205 wl_225 vdd gnd cell_6t
Xbit_r226_c205 bl_205 br_205 wl_226 vdd gnd cell_6t
Xbit_r227_c205 bl_205 br_205 wl_227 vdd gnd cell_6t
Xbit_r228_c205 bl_205 br_205 wl_228 vdd gnd cell_6t
Xbit_r229_c205 bl_205 br_205 wl_229 vdd gnd cell_6t
Xbit_r230_c205 bl_205 br_205 wl_230 vdd gnd cell_6t
Xbit_r231_c205 bl_205 br_205 wl_231 vdd gnd cell_6t
Xbit_r232_c205 bl_205 br_205 wl_232 vdd gnd cell_6t
Xbit_r233_c205 bl_205 br_205 wl_233 vdd gnd cell_6t
Xbit_r234_c205 bl_205 br_205 wl_234 vdd gnd cell_6t
Xbit_r235_c205 bl_205 br_205 wl_235 vdd gnd cell_6t
Xbit_r236_c205 bl_205 br_205 wl_236 vdd gnd cell_6t
Xbit_r237_c205 bl_205 br_205 wl_237 vdd gnd cell_6t
Xbit_r238_c205 bl_205 br_205 wl_238 vdd gnd cell_6t
Xbit_r239_c205 bl_205 br_205 wl_239 vdd gnd cell_6t
Xbit_r240_c205 bl_205 br_205 wl_240 vdd gnd cell_6t
Xbit_r241_c205 bl_205 br_205 wl_241 vdd gnd cell_6t
Xbit_r242_c205 bl_205 br_205 wl_242 vdd gnd cell_6t
Xbit_r243_c205 bl_205 br_205 wl_243 vdd gnd cell_6t
Xbit_r244_c205 bl_205 br_205 wl_244 vdd gnd cell_6t
Xbit_r245_c205 bl_205 br_205 wl_245 vdd gnd cell_6t
Xbit_r246_c205 bl_205 br_205 wl_246 vdd gnd cell_6t
Xbit_r247_c205 bl_205 br_205 wl_247 vdd gnd cell_6t
Xbit_r248_c205 bl_205 br_205 wl_248 vdd gnd cell_6t
Xbit_r249_c205 bl_205 br_205 wl_249 vdd gnd cell_6t
Xbit_r250_c205 bl_205 br_205 wl_250 vdd gnd cell_6t
Xbit_r251_c205 bl_205 br_205 wl_251 vdd gnd cell_6t
Xbit_r252_c205 bl_205 br_205 wl_252 vdd gnd cell_6t
Xbit_r253_c205 bl_205 br_205 wl_253 vdd gnd cell_6t
Xbit_r254_c205 bl_205 br_205 wl_254 vdd gnd cell_6t
Xbit_r255_c205 bl_205 br_205 wl_255 vdd gnd cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd cell_6t
Xbit_r1_c206 bl_206 br_206 wl_1 vdd gnd cell_6t
Xbit_r2_c206 bl_206 br_206 wl_2 vdd gnd cell_6t
Xbit_r3_c206 bl_206 br_206 wl_3 vdd gnd cell_6t
Xbit_r4_c206 bl_206 br_206 wl_4 vdd gnd cell_6t
Xbit_r5_c206 bl_206 br_206 wl_5 vdd gnd cell_6t
Xbit_r6_c206 bl_206 br_206 wl_6 vdd gnd cell_6t
Xbit_r7_c206 bl_206 br_206 wl_7 vdd gnd cell_6t
Xbit_r8_c206 bl_206 br_206 wl_8 vdd gnd cell_6t
Xbit_r9_c206 bl_206 br_206 wl_9 vdd gnd cell_6t
Xbit_r10_c206 bl_206 br_206 wl_10 vdd gnd cell_6t
Xbit_r11_c206 bl_206 br_206 wl_11 vdd gnd cell_6t
Xbit_r12_c206 bl_206 br_206 wl_12 vdd gnd cell_6t
Xbit_r13_c206 bl_206 br_206 wl_13 vdd gnd cell_6t
Xbit_r14_c206 bl_206 br_206 wl_14 vdd gnd cell_6t
Xbit_r15_c206 bl_206 br_206 wl_15 vdd gnd cell_6t
Xbit_r16_c206 bl_206 br_206 wl_16 vdd gnd cell_6t
Xbit_r17_c206 bl_206 br_206 wl_17 vdd gnd cell_6t
Xbit_r18_c206 bl_206 br_206 wl_18 vdd gnd cell_6t
Xbit_r19_c206 bl_206 br_206 wl_19 vdd gnd cell_6t
Xbit_r20_c206 bl_206 br_206 wl_20 vdd gnd cell_6t
Xbit_r21_c206 bl_206 br_206 wl_21 vdd gnd cell_6t
Xbit_r22_c206 bl_206 br_206 wl_22 vdd gnd cell_6t
Xbit_r23_c206 bl_206 br_206 wl_23 vdd gnd cell_6t
Xbit_r24_c206 bl_206 br_206 wl_24 vdd gnd cell_6t
Xbit_r25_c206 bl_206 br_206 wl_25 vdd gnd cell_6t
Xbit_r26_c206 bl_206 br_206 wl_26 vdd gnd cell_6t
Xbit_r27_c206 bl_206 br_206 wl_27 vdd gnd cell_6t
Xbit_r28_c206 bl_206 br_206 wl_28 vdd gnd cell_6t
Xbit_r29_c206 bl_206 br_206 wl_29 vdd gnd cell_6t
Xbit_r30_c206 bl_206 br_206 wl_30 vdd gnd cell_6t
Xbit_r31_c206 bl_206 br_206 wl_31 vdd gnd cell_6t
Xbit_r32_c206 bl_206 br_206 wl_32 vdd gnd cell_6t
Xbit_r33_c206 bl_206 br_206 wl_33 vdd gnd cell_6t
Xbit_r34_c206 bl_206 br_206 wl_34 vdd gnd cell_6t
Xbit_r35_c206 bl_206 br_206 wl_35 vdd gnd cell_6t
Xbit_r36_c206 bl_206 br_206 wl_36 vdd gnd cell_6t
Xbit_r37_c206 bl_206 br_206 wl_37 vdd gnd cell_6t
Xbit_r38_c206 bl_206 br_206 wl_38 vdd gnd cell_6t
Xbit_r39_c206 bl_206 br_206 wl_39 vdd gnd cell_6t
Xbit_r40_c206 bl_206 br_206 wl_40 vdd gnd cell_6t
Xbit_r41_c206 bl_206 br_206 wl_41 vdd gnd cell_6t
Xbit_r42_c206 bl_206 br_206 wl_42 vdd gnd cell_6t
Xbit_r43_c206 bl_206 br_206 wl_43 vdd gnd cell_6t
Xbit_r44_c206 bl_206 br_206 wl_44 vdd gnd cell_6t
Xbit_r45_c206 bl_206 br_206 wl_45 vdd gnd cell_6t
Xbit_r46_c206 bl_206 br_206 wl_46 vdd gnd cell_6t
Xbit_r47_c206 bl_206 br_206 wl_47 vdd gnd cell_6t
Xbit_r48_c206 bl_206 br_206 wl_48 vdd gnd cell_6t
Xbit_r49_c206 bl_206 br_206 wl_49 vdd gnd cell_6t
Xbit_r50_c206 bl_206 br_206 wl_50 vdd gnd cell_6t
Xbit_r51_c206 bl_206 br_206 wl_51 vdd gnd cell_6t
Xbit_r52_c206 bl_206 br_206 wl_52 vdd gnd cell_6t
Xbit_r53_c206 bl_206 br_206 wl_53 vdd gnd cell_6t
Xbit_r54_c206 bl_206 br_206 wl_54 vdd gnd cell_6t
Xbit_r55_c206 bl_206 br_206 wl_55 vdd gnd cell_6t
Xbit_r56_c206 bl_206 br_206 wl_56 vdd gnd cell_6t
Xbit_r57_c206 bl_206 br_206 wl_57 vdd gnd cell_6t
Xbit_r58_c206 bl_206 br_206 wl_58 vdd gnd cell_6t
Xbit_r59_c206 bl_206 br_206 wl_59 vdd gnd cell_6t
Xbit_r60_c206 bl_206 br_206 wl_60 vdd gnd cell_6t
Xbit_r61_c206 bl_206 br_206 wl_61 vdd gnd cell_6t
Xbit_r62_c206 bl_206 br_206 wl_62 vdd gnd cell_6t
Xbit_r63_c206 bl_206 br_206 wl_63 vdd gnd cell_6t
Xbit_r64_c206 bl_206 br_206 wl_64 vdd gnd cell_6t
Xbit_r65_c206 bl_206 br_206 wl_65 vdd gnd cell_6t
Xbit_r66_c206 bl_206 br_206 wl_66 vdd gnd cell_6t
Xbit_r67_c206 bl_206 br_206 wl_67 vdd gnd cell_6t
Xbit_r68_c206 bl_206 br_206 wl_68 vdd gnd cell_6t
Xbit_r69_c206 bl_206 br_206 wl_69 vdd gnd cell_6t
Xbit_r70_c206 bl_206 br_206 wl_70 vdd gnd cell_6t
Xbit_r71_c206 bl_206 br_206 wl_71 vdd gnd cell_6t
Xbit_r72_c206 bl_206 br_206 wl_72 vdd gnd cell_6t
Xbit_r73_c206 bl_206 br_206 wl_73 vdd gnd cell_6t
Xbit_r74_c206 bl_206 br_206 wl_74 vdd gnd cell_6t
Xbit_r75_c206 bl_206 br_206 wl_75 vdd gnd cell_6t
Xbit_r76_c206 bl_206 br_206 wl_76 vdd gnd cell_6t
Xbit_r77_c206 bl_206 br_206 wl_77 vdd gnd cell_6t
Xbit_r78_c206 bl_206 br_206 wl_78 vdd gnd cell_6t
Xbit_r79_c206 bl_206 br_206 wl_79 vdd gnd cell_6t
Xbit_r80_c206 bl_206 br_206 wl_80 vdd gnd cell_6t
Xbit_r81_c206 bl_206 br_206 wl_81 vdd gnd cell_6t
Xbit_r82_c206 bl_206 br_206 wl_82 vdd gnd cell_6t
Xbit_r83_c206 bl_206 br_206 wl_83 vdd gnd cell_6t
Xbit_r84_c206 bl_206 br_206 wl_84 vdd gnd cell_6t
Xbit_r85_c206 bl_206 br_206 wl_85 vdd gnd cell_6t
Xbit_r86_c206 bl_206 br_206 wl_86 vdd gnd cell_6t
Xbit_r87_c206 bl_206 br_206 wl_87 vdd gnd cell_6t
Xbit_r88_c206 bl_206 br_206 wl_88 vdd gnd cell_6t
Xbit_r89_c206 bl_206 br_206 wl_89 vdd gnd cell_6t
Xbit_r90_c206 bl_206 br_206 wl_90 vdd gnd cell_6t
Xbit_r91_c206 bl_206 br_206 wl_91 vdd gnd cell_6t
Xbit_r92_c206 bl_206 br_206 wl_92 vdd gnd cell_6t
Xbit_r93_c206 bl_206 br_206 wl_93 vdd gnd cell_6t
Xbit_r94_c206 bl_206 br_206 wl_94 vdd gnd cell_6t
Xbit_r95_c206 bl_206 br_206 wl_95 vdd gnd cell_6t
Xbit_r96_c206 bl_206 br_206 wl_96 vdd gnd cell_6t
Xbit_r97_c206 bl_206 br_206 wl_97 vdd gnd cell_6t
Xbit_r98_c206 bl_206 br_206 wl_98 vdd gnd cell_6t
Xbit_r99_c206 bl_206 br_206 wl_99 vdd gnd cell_6t
Xbit_r100_c206 bl_206 br_206 wl_100 vdd gnd cell_6t
Xbit_r101_c206 bl_206 br_206 wl_101 vdd gnd cell_6t
Xbit_r102_c206 bl_206 br_206 wl_102 vdd gnd cell_6t
Xbit_r103_c206 bl_206 br_206 wl_103 vdd gnd cell_6t
Xbit_r104_c206 bl_206 br_206 wl_104 vdd gnd cell_6t
Xbit_r105_c206 bl_206 br_206 wl_105 vdd gnd cell_6t
Xbit_r106_c206 bl_206 br_206 wl_106 vdd gnd cell_6t
Xbit_r107_c206 bl_206 br_206 wl_107 vdd gnd cell_6t
Xbit_r108_c206 bl_206 br_206 wl_108 vdd gnd cell_6t
Xbit_r109_c206 bl_206 br_206 wl_109 vdd gnd cell_6t
Xbit_r110_c206 bl_206 br_206 wl_110 vdd gnd cell_6t
Xbit_r111_c206 bl_206 br_206 wl_111 vdd gnd cell_6t
Xbit_r112_c206 bl_206 br_206 wl_112 vdd gnd cell_6t
Xbit_r113_c206 bl_206 br_206 wl_113 vdd gnd cell_6t
Xbit_r114_c206 bl_206 br_206 wl_114 vdd gnd cell_6t
Xbit_r115_c206 bl_206 br_206 wl_115 vdd gnd cell_6t
Xbit_r116_c206 bl_206 br_206 wl_116 vdd gnd cell_6t
Xbit_r117_c206 bl_206 br_206 wl_117 vdd gnd cell_6t
Xbit_r118_c206 bl_206 br_206 wl_118 vdd gnd cell_6t
Xbit_r119_c206 bl_206 br_206 wl_119 vdd gnd cell_6t
Xbit_r120_c206 bl_206 br_206 wl_120 vdd gnd cell_6t
Xbit_r121_c206 bl_206 br_206 wl_121 vdd gnd cell_6t
Xbit_r122_c206 bl_206 br_206 wl_122 vdd gnd cell_6t
Xbit_r123_c206 bl_206 br_206 wl_123 vdd gnd cell_6t
Xbit_r124_c206 bl_206 br_206 wl_124 vdd gnd cell_6t
Xbit_r125_c206 bl_206 br_206 wl_125 vdd gnd cell_6t
Xbit_r126_c206 bl_206 br_206 wl_126 vdd gnd cell_6t
Xbit_r127_c206 bl_206 br_206 wl_127 vdd gnd cell_6t
Xbit_r128_c206 bl_206 br_206 wl_128 vdd gnd cell_6t
Xbit_r129_c206 bl_206 br_206 wl_129 vdd gnd cell_6t
Xbit_r130_c206 bl_206 br_206 wl_130 vdd gnd cell_6t
Xbit_r131_c206 bl_206 br_206 wl_131 vdd gnd cell_6t
Xbit_r132_c206 bl_206 br_206 wl_132 vdd gnd cell_6t
Xbit_r133_c206 bl_206 br_206 wl_133 vdd gnd cell_6t
Xbit_r134_c206 bl_206 br_206 wl_134 vdd gnd cell_6t
Xbit_r135_c206 bl_206 br_206 wl_135 vdd gnd cell_6t
Xbit_r136_c206 bl_206 br_206 wl_136 vdd gnd cell_6t
Xbit_r137_c206 bl_206 br_206 wl_137 vdd gnd cell_6t
Xbit_r138_c206 bl_206 br_206 wl_138 vdd gnd cell_6t
Xbit_r139_c206 bl_206 br_206 wl_139 vdd gnd cell_6t
Xbit_r140_c206 bl_206 br_206 wl_140 vdd gnd cell_6t
Xbit_r141_c206 bl_206 br_206 wl_141 vdd gnd cell_6t
Xbit_r142_c206 bl_206 br_206 wl_142 vdd gnd cell_6t
Xbit_r143_c206 bl_206 br_206 wl_143 vdd gnd cell_6t
Xbit_r144_c206 bl_206 br_206 wl_144 vdd gnd cell_6t
Xbit_r145_c206 bl_206 br_206 wl_145 vdd gnd cell_6t
Xbit_r146_c206 bl_206 br_206 wl_146 vdd gnd cell_6t
Xbit_r147_c206 bl_206 br_206 wl_147 vdd gnd cell_6t
Xbit_r148_c206 bl_206 br_206 wl_148 vdd gnd cell_6t
Xbit_r149_c206 bl_206 br_206 wl_149 vdd gnd cell_6t
Xbit_r150_c206 bl_206 br_206 wl_150 vdd gnd cell_6t
Xbit_r151_c206 bl_206 br_206 wl_151 vdd gnd cell_6t
Xbit_r152_c206 bl_206 br_206 wl_152 vdd gnd cell_6t
Xbit_r153_c206 bl_206 br_206 wl_153 vdd gnd cell_6t
Xbit_r154_c206 bl_206 br_206 wl_154 vdd gnd cell_6t
Xbit_r155_c206 bl_206 br_206 wl_155 vdd gnd cell_6t
Xbit_r156_c206 bl_206 br_206 wl_156 vdd gnd cell_6t
Xbit_r157_c206 bl_206 br_206 wl_157 vdd gnd cell_6t
Xbit_r158_c206 bl_206 br_206 wl_158 vdd gnd cell_6t
Xbit_r159_c206 bl_206 br_206 wl_159 vdd gnd cell_6t
Xbit_r160_c206 bl_206 br_206 wl_160 vdd gnd cell_6t
Xbit_r161_c206 bl_206 br_206 wl_161 vdd gnd cell_6t
Xbit_r162_c206 bl_206 br_206 wl_162 vdd gnd cell_6t
Xbit_r163_c206 bl_206 br_206 wl_163 vdd gnd cell_6t
Xbit_r164_c206 bl_206 br_206 wl_164 vdd gnd cell_6t
Xbit_r165_c206 bl_206 br_206 wl_165 vdd gnd cell_6t
Xbit_r166_c206 bl_206 br_206 wl_166 vdd gnd cell_6t
Xbit_r167_c206 bl_206 br_206 wl_167 vdd gnd cell_6t
Xbit_r168_c206 bl_206 br_206 wl_168 vdd gnd cell_6t
Xbit_r169_c206 bl_206 br_206 wl_169 vdd gnd cell_6t
Xbit_r170_c206 bl_206 br_206 wl_170 vdd gnd cell_6t
Xbit_r171_c206 bl_206 br_206 wl_171 vdd gnd cell_6t
Xbit_r172_c206 bl_206 br_206 wl_172 vdd gnd cell_6t
Xbit_r173_c206 bl_206 br_206 wl_173 vdd gnd cell_6t
Xbit_r174_c206 bl_206 br_206 wl_174 vdd gnd cell_6t
Xbit_r175_c206 bl_206 br_206 wl_175 vdd gnd cell_6t
Xbit_r176_c206 bl_206 br_206 wl_176 vdd gnd cell_6t
Xbit_r177_c206 bl_206 br_206 wl_177 vdd gnd cell_6t
Xbit_r178_c206 bl_206 br_206 wl_178 vdd gnd cell_6t
Xbit_r179_c206 bl_206 br_206 wl_179 vdd gnd cell_6t
Xbit_r180_c206 bl_206 br_206 wl_180 vdd gnd cell_6t
Xbit_r181_c206 bl_206 br_206 wl_181 vdd gnd cell_6t
Xbit_r182_c206 bl_206 br_206 wl_182 vdd gnd cell_6t
Xbit_r183_c206 bl_206 br_206 wl_183 vdd gnd cell_6t
Xbit_r184_c206 bl_206 br_206 wl_184 vdd gnd cell_6t
Xbit_r185_c206 bl_206 br_206 wl_185 vdd gnd cell_6t
Xbit_r186_c206 bl_206 br_206 wl_186 vdd gnd cell_6t
Xbit_r187_c206 bl_206 br_206 wl_187 vdd gnd cell_6t
Xbit_r188_c206 bl_206 br_206 wl_188 vdd gnd cell_6t
Xbit_r189_c206 bl_206 br_206 wl_189 vdd gnd cell_6t
Xbit_r190_c206 bl_206 br_206 wl_190 vdd gnd cell_6t
Xbit_r191_c206 bl_206 br_206 wl_191 vdd gnd cell_6t
Xbit_r192_c206 bl_206 br_206 wl_192 vdd gnd cell_6t
Xbit_r193_c206 bl_206 br_206 wl_193 vdd gnd cell_6t
Xbit_r194_c206 bl_206 br_206 wl_194 vdd gnd cell_6t
Xbit_r195_c206 bl_206 br_206 wl_195 vdd gnd cell_6t
Xbit_r196_c206 bl_206 br_206 wl_196 vdd gnd cell_6t
Xbit_r197_c206 bl_206 br_206 wl_197 vdd gnd cell_6t
Xbit_r198_c206 bl_206 br_206 wl_198 vdd gnd cell_6t
Xbit_r199_c206 bl_206 br_206 wl_199 vdd gnd cell_6t
Xbit_r200_c206 bl_206 br_206 wl_200 vdd gnd cell_6t
Xbit_r201_c206 bl_206 br_206 wl_201 vdd gnd cell_6t
Xbit_r202_c206 bl_206 br_206 wl_202 vdd gnd cell_6t
Xbit_r203_c206 bl_206 br_206 wl_203 vdd gnd cell_6t
Xbit_r204_c206 bl_206 br_206 wl_204 vdd gnd cell_6t
Xbit_r205_c206 bl_206 br_206 wl_205 vdd gnd cell_6t
Xbit_r206_c206 bl_206 br_206 wl_206 vdd gnd cell_6t
Xbit_r207_c206 bl_206 br_206 wl_207 vdd gnd cell_6t
Xbit_r208_c206 bl_206 br_206 wl_208 vdd gnd cell_6t
Xbit_r209_c206 bl_206 br_206 wl_209 vdd gnd cell_6t
Xbit_r210_c206 bl_206 br_206 wl_210 vdd gnd cell_6t
Xbit_r211_c206 bl_206 br_206 wl_211 vdd gnd cell_6t
Xbit_r212_c206 bl_206 br_206 wl_212 vdd gnd cell_6t
Xbit_r213_c206 bl_206 br_206 wl_213 vdd gnd cell_6t
Xbit_r214_c206 bl_206 br_206 wl_214 vdd gnd cell_6t
Xbit_r215_c206 bl_206 br_206 wl_215 vdd gnd cell_6t
Xbit_r216_c206 bl_206 br_206 wl_216 vdd gnd cell_6t
Xbit_r217_c206 bl_206 br_206 wl_217 vdd gnd cell_6t
Xbit_r218_c206 bl_206 br_206 wl_218 vdd gnd cell_6t
Xbit_r219_c206 bl_206 br_206 wl_219 vdd gnd cell_6t
Xbit_r220_c206 bl_206 br_206 wl_220 vdd gnd cell_6t
Xbit_r221_c206 bl_206 br_206 wl_221 vdd gnd cell_6t
Xbit_r222_c206 bl_206 br_206 wl_222 vdd gnd cell_6t
Xbit_r223_c206 bl_206 br_206 wl_223 vdd gnd cell_6t
Xbit_r224_c206 bl_206 br_206 wl_224 vdd gnd cell_6t
Xbit_r225_c206 bl_206 br_206 wl_225 vdd gnd cell_6t
Xbit_r226_c206 bl_206 br_206 wl_226 vdd gnd cell_6t
Xbit_r227_c206 bl_206 br_206 wl_227 vdd gnd cell_6t
Xbit_r228_c206 bl_206 br_206 wl_228 vdd gnd cell_6t
Xbit_r229_c206 bl_206 br_206 wl_229 vdd gnd cell_6t
Xbit_r230_c206 bl_206 br_206 wl_230 vdd gnd cell_6t
Xbit_r231_c206 bl_206 br_206 wl_231 vdd gnd cell_6t
Xbit_r232_c206 bl_206 br_206 wl_232 vdd gnd cell_6t
Xbit_r233_c206 bl_206 br_206 wl_233 vdd gnd cell_6t
Xbit_r234_c206 bl_206 br_206 wl_234 vdd gnd cell_6t
Xbit_r235_c206 bl_206 br_206 wl_235 vdd gnd cell_6t
Xbit_r236_c206 bl_206 br_206 wl_236 vdd gnd cell_6t
Xbit_r237_c206 bl_206 br_206 wl_237 vdd gnd cell_6t
Xbit_r238_c206 bl_206 br_206 wl_238 vdd gnd cell_6t
Xbit_r239_c206 bl_206 br_206 wl_239 vdd gnd cell_6t
Xbit_r240_c206 bl_206 br_206 wl_240 vdd gnd cell_6t
Xbit_r241_c206 bl_206 br_206 wl_241 vdd gnd cell_6t
Xbit_r242_c206 bl_206 br_206 wl_242 vdd gnd cell_6t
Xbit_r243_c206 bl_206 br_206 wl_243 vdd gnd cell_6t
Xbit_r244_c206 bl_206 br_206 wl_244 vdd gnd cell_6t
Xbit_r245_c206 bl_206 br_206 wl_245 vdd gnd cell_6t
Xbit_r246_c206 bl_206 br_206 wl_246 vdd gnd cell_6t
Xbit_r247_c206 bl_206 br_206 wl_247 vdd gnd cell_6t
Xbit_r248_c206 bl_206 br_206 wl_248 vdd gnd cell_6t
Xbit_r249_c206 bl_206 br_206 wl_249 vdd gnd cell_6t
Xbit_r250_c206 bl_206 br_206 wl_250 vdd gnd cell_6t
Xbit_r251_c206 bl_206 br_206 wl_251 vdd gnd cell_6t
Xbit_r252_c206 bl_206 br_206 wl_252 vdd gnd cell_6t
Xbit_r253_c206 bl_206 br_206 wl_253 vdd gnd cell_6t
Xbit_r254_c206 bl_206 br_206 wl_254 vdd gnd cell_6t
Xbit_r255_c206 bl_206 br_206 wl_255 vdd gnd cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd cell_6t
Xbit_r1_c207 bl_207 br_207 wl_1 vdd gnd cell_6t
Xbit_r2_c207 bl_207 br_207 wl_2 vdd gnd cell_6t
Xbit_r3_c207 bl_207 br_207 wl_3 vdd gnd cell_6t
Xbit_r4_c207 bl_207 br_207 wl_4 vdd gnd cell_6t
Xbit_r5_c207 bl_207 br_207 wl_5 vdd gnd cell_6t
Xbit_r6_c207 bl_207 br_207 wl_6 vdd gnd cell_6t
Xbit_r7_c207 bl_207 br_207 wl_7 vdd gnd cell_6t
Xbit_r8_c207 bl_207 br_207 wl_8 vdd gnd cell_6t
Xbit_r9_c207 bl_207 br_207 wl_9 vdd gnd cell_6t
Xbit_r10_c207 bl_207 br_207 wl_10 vdd gnd cell_6t
Xbit_r11_c207 bl_207 br_207 wl_11 vdd gnd cell_6t
Xbit_r12_c207 bl_207 br_207 wl_12 vdd gnd cell_6t
Xbit_r13_c207 bl_207 br_207 wl_13 vdd gnd cell_6t
Xbit_r14_c207 bl_207 br_207 wl_14 vdd gnd cell_6t
Xbit_r15_c207 bl_207 br_207 wl_15 vdd gnd cell_6t
Xbit_r16_c207 bl_207 br_207 wl_16 vdd gnd cell_6t
Xbit_r17_c207 bl_207 br_207 wl_17 vdd gnd cell_6t
Xbit_r18_c207 bl_207 br_207 wl_18 vdd gnd cell_6t
Xbit_r19_c207 bl_207 br_207 wl_19 vdd gnd cell_6t
Xbit_r20_c207 bl_207 br_207 wl_20 vdd gnd cell_6t
Xbit_r21_c207 bl_207 br_207 wl_21 vdd gnd cell_6t
Xbit_r22_c207 bl_207 br_207 wl_22 vdd gnd cell_6t
Xbit_r23_c207 bl_207 br_207 wl_23 vdd gnd cell_6t
Xbit_r24_c207 bl_207 br_207 wl_24 vdd gnd cell_6t
Xbit_r25_c207 bl_207 br_207 wl_25 vdd gnd cell_6t
Xbit_r26_c207 bl_207 br_207 wl_26 vdd gnd cell_6t
Xbit_r27_c207 bl_207 br_207 wl_27 vdd gnd cell_6t
Xbit_r28_c207 bl_207 br_207 wl_28 vdd gnd cell_6t
Xbit_r29_c207 bl_207 br_207 wl_29 vdd gnd cell_6t
Xbit_r30_c207 bl_207 br_207 wl_30 vdd gnd cell_6t
Xbit_r31_c207 bl_207 br_207 wl_31 vdd gnd cell_6t
Xbit_r32_c207 bl_207 br_207 wl_32 vdd gnd cell_6t
Xbit_r33_c207 bl_207 br_207 wl_33 vdd gnd cell_6t
Xbit_r34_c207 bl_207 br_207 wl_34 vdd gnd cell_6t
Xbit_r35_c207 bl_207 br_207 wl_35 vdd gnd cell_6t
Xbit_r36_c207 bl_207 br_207 wl_36 vdd gnd cell_6t
Xbit_r37_c207 bl_207 br_207 wl_37 vdd gnd cell_6t
Xbit_r38_c207 bl_207 br_207 wl_38 vdd gnd cell_6t
Xbit_r39_c207 bl_207 br_207 wl_39 vdd gnd cell_6t
Xbit_r40_c207 bl_207 br_207 wl_40 vdd gnd cell_6t
Xbit_r41_c207 bl_207 br_207 wl_41 vdd gnd cell_6t
Xbit_r42_c207 bl_207 br_207 wl_42 vdd gnd cell_6t
Xbit_r43_c207 bl_207 br_207 wl_43 vdd gnd cell_6t
Xbit_r44_c207 bl_207 br_207 wl_44 vdd gnd cell_6t
Xbit_r45_c207 bl_207 br_207 wl_45 vdd gnd cell_6t
Xbit_r46_c207 bl_207 br_207 wl_46 vdd gnd cell_6t
Xbit_r47_c207 bl_207 br_207 wl_47 vdd gnd cell_6t
Xbit_r48_c207 bl_207 br_207 wl_48 vdd gnd cell_6t
Xbit_r49_c207 bl_207 br_207 wl_49 vdd gnd cell_6t
Xbit_r50_c207 bl_207 br_207 wl_50 vdd gnd cell_6t
Xbit_r51_c207 bl_207 br_207 wl_51 vdd gnd cell_6t
Xbit_r52_c207 bl_207 br_207 wl_52 vdd gnd cell_6t
Xbit_r53_c207 bl_207 br_207 wl_53 vdd gnd cell_6t
Xbit_r54_c207 bl_207 br_207 wl_54 vdd gnd cell_6t
Xbit_r55_c207 bl_207 br_207 wl_55 vdd gnd cell_6t
Xbit_r56_c207 bl_207 br_207 wl_56 vdd gnd cell_6t
Xbit_r57_c207 bl_207 br_207 wl_57 vdd gnd cell_6t
Xbit_r58_c207 bl_207 br_207 wl_58 vdd gnd cell_6t
Xbit_r59_c207 bl_207 br_207 wl_59 vdd gnd cell_6t
Xbit_r60_c207 bl_207 br_207 wl_60 vdd gnd cell_6t
Xbit_r61_c207 bl_207 br_207 wl_61 vdd gnd cell_6t
Xbit_r62_c207 bl_207 br_207 wl_62 vdd gnd cell_6t
Xbit_r63_c207 bl_207 br_207 wl_63 vdd gnd cell_6t
Xbit_r64_c207 bl_207 br_207 wl_64 vdd gnd cell_6t
Xbit_r65_c207 bl_207 br_207 wl_65 vdd gnd cell_6t
Xbit_r66_c207 bl_207 br_207 wl_66 vdd gnd cell_6t
Xbit_r67_c207 bl_207 br_207 wl_67 vdd gnd cell_6t
Xbit_r68_c207 bl_207 br_207 wl_68 vdd gnd cell_6t
Xbit_r69_c207 bl_207 br_207 wl_69 vdd gnd cell_6t
Xbit_r70_c207 bl_207 br_207 wl_70 vdd gnd cell_6t
Xbit_r71_c207 bl_207 br_207 wl_71 vdd gnd cell_6t
Xbit_r72_c207 bl_207 br_207 wl_72 vdd gnd cell_6t
Xbit_r73_c207 bl_207 br_207 wl_73 vdd gnd cell_6t
Xbit_r74_c207 bl_207 br_207 wl_74 vdd gnd cell_6t
Xbit_r75_c207 bl_207 br_207 wl_75 vdd gnd cell_6t
Xbit_r76_c207 bl_207 br_207 wl_76 vdd gnd cell_6t
Xbit_r77_c207 bl_207 br_207 wl_77 vdd gnd cell_6t
Xbit_r78_c207 bl_207 br_207 wl_78 vdd gnd cell_6t
Xbit_r79_c207 bl_207 br_207 wl_79 vdd gnd cell_6t
Xbit_r80_c207 bl_207 br_207 wl_80 vdd gnd cell_6t
Xbit_r81_c207 bl_207 br_207 wl_81 vdd gnd cell_6t
Xbit_r82_c207 bl_207 br_207 wl_82 vdd gnd cell_6t
Xbit_r83_c207 bl_207 br_207 wl_83 vdd gnd cell_6t
Xbit_r84_c207 bl_207 br_207 wl_84 vdd gnd cell_6t
Xbit_r85_c207 bl_207 br_207 wl_85 vdd gnd cell_6t
Xbit_r86_c207 bl_207 br_207 wl_86 vdd gnd cell_6t
Xbit_r87_c207 bl_207 br_207 wl_87 vdd gnd cell_6t
Xbit_r88_c207 bl_207 br_207 wl_88 vdd gnd cell_6t
Xbit_r89_c207 bl_207 br_207 wl_89 vdd gnd cell_6t
Xbit_r90_c207 bl_207 br_207 wl_90 vdd gnd cell_6t
Xbit_r91_c207 bl_207 br_207 wl_91 vdd gnd cell_6t
Xbit_r92_c207 bl_207 br_207 wl_92 vdd gnd cell_6t
Xbit_r93_c207 bl_207 br_207 wl_93 vdd gnd cell_6t
Xbit_r94_c207 bl_207 br_207 wl_94 vdd gnd cell_6t
Xbit_r95_c207 bl_207 br_207 wl_95 vdd gnd cell_6t
Xbit_r96_c207 bl_207 br_207 wl_96 vdd gnd cell_6t
Xbit_r97_c207 bl_207 br_207 wl_97 vdd gnd cell_6t
Xbit_r98_c207 bl_207 br_207 wl_98 vdd gnd cell_6t
Xbit_r99_c207 bl_207 br_207 wl_99 vdd gnd cell_6t
Xbit_r100_c207 bl_207 br_207 wl_100 vdd gnd cell_6t
Xbit_r101_c207 bl_207 br_207 wl_101 vdd gnd cell_6t
Xbit_r102_c207 bl_207 br_207 wl_102 vdd gnd cell_6t
Xbit_r103_c207 bl_207 br_207 wl_103 vdd gnd cell_6t
Xbit_r104_c207 bl_207 br_207 wl_104 vdd gnd cell_6t
Xbit_r105_c207 bl_207 br_207 wl_105 vdd gnd cell_6t
Xbit_r106_c207 bl_207 br_207 wl_106 vdd gnd cell_6t
Xbit_r107_c207 bl_207 br_207 wl_107 vdd gnd cell_6t
Xbit_r108_c207 bl_207 br_207 wl_108 vdd gnd cell_6t
Xbit_r109_c207 bl_207 br_207 wl_109 vdd gnd cell_6t
Xbit_r110_c207 bl_207 br_207 wl_110 vdd gnd cell_6t
Xbit_r111_c207 bl_207 br_207 wl_111 vdd gnd cell_6t
Xbit_r112_c207 bl_207 br_207 wl_112 vdd gnd cell_6t
Xbit_r113_c207 bl_207 br_207 wl_113 vdd gnd cell_6t
Xbit_r114_c207 bl_207 br_207 wl_114 vdd gnd cell_6t
Xbit_r115_c207 bl_207 br_207 wl_115 vdd gnd cell_6t
Xbit_r116_c207 bl_207 br_207 wl_116 vdd gnd cell_6t
Xbit_r117_c207 bl_207 br_207 wl_117 vdd gnd cell_6t
Xbit_r118_c207 bl_207 br_207 wl_118 vdd gnd cell_6t
Xbit_r119_c207 bl_207 br_207 wl_119 vdd gnd cell_6t
Xbit_r120_c207 bl_207 br_207 wl_120 vdd gnd cell_6t
Xbit_r121_c207 bl_207 br_207 wl_121 vdd gnd cell_6t
Xbit_r122_c207 bl_207 br_207 wl_122 vdd gnd cell_6t
Xbit_r123_c207 bl_207 br_207 wl_123 vdd gnd cell_6t
Xbit_r124_c207 bl_207 br_207 wl_124 vdd gnd cell_6t
Xbit_r125_c207 bl_207 br_207 wl_125 vdd gnd cell_6t
Xbit_r126_c207 bl_207 br_207 wl_126 vdd gnd cell_6t
Xbit_r127_c207 bl_207 br_207 wl_127 vdd gnd cell_6t
Xbit_r128_c207 bl_207 br_207 wl_128 vdd gnd cell_6t
Xbit_r129_c207 bl_207 br_207 wl_129 vdd gnd cell_6t
Xbit_r130_c207 bl_207 br_207 wl_130 vdd gnd cell_6t
Xbit_r131_c207 bl_207 br_207 wl_131 vdd gnd cell_6t
Xbit_r132_c207 bl_207 br_207 wl_132 vdd gnd cell_6t
Xbit_r133_c207 bl_207 br_207 wl_133 vdd gnd cell_6t
Xbit_r134_c207 bl_207 br_207 wl_134 vdd gnd cell_6t
Xbit_r135_c207 bl_207 br_207 wl_135 vdd gnd cell_6t
Xbit_r136_c207 bl_207 br_207 wl_136 vdd gnd cell_6t
Xbit_r137_c207 bl_207 br_207 wl_137 vdd gnd cell_6t
Xbit_r138_c207 bl_207 br_207 wl_138 vdd gnd cell_6t
Xbit_r139_c207 bl_207 br_207 wl_139 vdd gnd cell_6t
Xbit_r140_c207 bl_207 br_207 wl_140 vdd gnd cell_6t
Xbit_r141_c207 bl_207 br_207 wl_141 vdd gnd cell_6t
Xbit_r142_c207 bl_207 br_207 wl_142 vdd gnd cell_6t
Xbit_r143_c207 bl_207 br_207 wl_143 vdd gnd cell_6t
Xbit_r144_c207 bl_207 br_207 wl_144 vdd gnd cell_6t
Xbit_r145_c207 bl_207 br_207 wl_145 vdd gnd cell_6t
Xbit_r146_c207 bl_207 br_207 wl_146 vdd gnd cell_6t
Xbit_r147_c207 bl_207 br_207 wl_147 vdd gnd cell_6t
Xbit_r148_c207 bl_207 br_207 wl_148 vdd gnd cell_6t
Xbit_r149_c207 bl_207 br_207 wl_149 vdd gnd cell_6t
Xbit_r150_c207 bl_207 br_207 wl_150 vdd gnd cell_6t
Xbit_r151_c207 bl_207 br_207 wl_151 vdd gnd cell_6t
Xbit_r152_c207 bl_207 br_207 wl_152 vdd gnd cell_6t
Xbit_r153_c207 bl_207 br_207 wl_153 vdd gnd cell_6t
Xbit_r154_c207 bl_207 br_207 wl_154 vdd gnd cell_6t
Xbit_r155_c207 bl_207 br_207 wl_155 vdd gnd cell_6t
Xbit_r156_c207 bl_207 br_207 wl_156 vdd gnd cell_6t
Xbit_r157_c207 bl_207 br_207 wl_157 vdd gnd cell_6t
Xbit_r158_c207 bl_207 br_207 wl_158 vdd gnd cell_6t
Xbit_r159_c207 bl_207 br_207 wl_159 vdd gnd cell_6t
Xbit_r160_c207 bl_207 br_207 wl_160 vdd gnd cell_6t
Xbit_r161_c207 bl_207 br_207 wl_161 vdd gnd cell_6t
Xbit_r162_c207 bl_207 br_207 wl_162 vdd gnd cell_6t
Xbit_r163_c207 bl_207 br_207 wl_163 vdd gnd cell_6t
Xbit_r164_c207 bl_207 br_207 wl_164 vdd gnd cell_6t
Xbit_r165_c207 bl_207 br_207 wl_165 vdd gnd cell_6t
Xbit_r166_c207 bl_207 br_207 wl_166 vdd gnd cell_6t
Xbit_r167_c207 bl_207 br_207 wl_167 vdd gnd cell_6t
Xbit_r168_c207 bl_207 br_207 wl_168 vdd gnd cell_6t
Xbit_r169_c207 bl_207 br_207 wl_169 vdd gnd cell_6t
Xbit_r170_c207 bl_207 br_207 wl_170 vdd gnd cell_6t
Xbit_r171_c207 bl_207 br_207 wl_171 vdd gnd cell_6t
Xbit_r172_c207 bl_207 br_207 wl_172 vdd gnd cell_6t
Xbit_r173_c207 bl_207 br_207 wl_173 vdd gnd cell_6t
Xbit_r174_c207 bl_207 br_207 wl_174 vdd gnd cell_6t
Xbit_r175_c207 bl_207 br_207 wl_175 vdd gnd cell_6t
Xbit_r176_c207 bl_207 br_207 wl_176 vdd gnd cell_6t
Xbit_r177_c207 bl_207 br_207 wl_177 vdd gnd cell_6t
Xbit_r178_c207 bl_207 br_207 wl_178 vdd gnd cell_6t
Xbit_r179_c207 bl_207 br_207 wl_179 vdd gnd cell_6t
Xbit_r180_c207 bl_207 br_207 wl_180 vdd gnd cell_6t
Xbit_r181_c207 bl_207 br_207 wl_181 vdd gnd cell_6t
Xbit_r182_c207 bl_207 br_207 wl_182 vdd gnd cell_6t
Xbit_r183_c207 bl_207 br_207 wl_183 vdd gnd cell_6t
Xbit_r184_c207 bl_207 br_207 wl_184 vdd gnd cell_6t
Xbit_r185_c207 bl_207 br_207 wl_185 vdd gnd cell_6t
Xbit_r186_c207 bl_207 br_207 wl_186 vdd gnd cell_6t
Xbit_r187_c207 bl_207 br_207 wl_187 vdd gnd cell_6t
Xbit_r188_c207 bl_207 br_207 wl_188 vdd gnd cell_6t
Xbit_r189_c207 bl_207 br_207 wl_189 vdd gnd cell_6t
Xbit_r190_c207 bl_207 br_207 wl_190 vdd gnd cell_6t
Xbit_r191_c207 bl_207 br_207 wl_191 vdd gnd cell_6t
Xbit_r192_c207 bl_207 br_207 wl_192 vdd gnd cell_6t
Xbit_r193_c207 bl_207 br_207 wl_193 vdd gnd cell_6t
Xbit_r194_c207 bl_207 br_207 wl_194 vdd gnd cell_6t
Xbit_r195_c207 bl_207 br_207 wl_195 vdd gnd cell_6t
Xbit_r196_c207 bl_207 br_207 wl_196 vdd gnd cell_6t
Xbit_r197_c207 bl_207 br_207 wl_197 vdd gnd cell_6t
Xbit_r198_c207 bl_207 br_207 wl_198 vdd gnd cell_6t
Xbit_r199_c207 bl_207 br_207 wl_199 vdd gnd cell_6t
Xbit_r200_c207 bl_207 br_207 wl_200 vdd gnd cell_6t
Xbit_r201_c207 bl_207 br_207 wl_201 vdd gnd cell_6t
Xbit_r202_c207 bl_207 br_207 wl_202 vdd gnd cell_6t
Xbit_r203_c207 bl_207 br_207 wl_203 vdd gnd cell_6t
Xbit_r204_c207 bl_207 br_207 wl_204 vdd gnd cell_6t
Xbit_r205_c207 bl_207 br_207 wl_205 vdd gnd cell_6t
Xbit_r206_c207 bl_207 br_207 wl_206 vdd gnd cell_6t
Xbit_r207_c207 bl_207 br_207 wl_207 vdd gnd cell_6t
Xbit_r208_c207 bl_207 br_207 wl_208 vdd gnd cell_6t
Xbit_r209_c207 bl_207 br_207 wl_209 vdd gnd cell_6t
Xbit_r210_c207 bl_207 br_207 wl_210 vdd gnd cell_6t
Xbit_r211_c207 bl_207 br_207 wl_211 vdd gnd cell_6t
Xbit_r212_c207 bl_207 br_207 wl_212 vdd gnd cell_6t
Xbit_r213_c207 bl_207 br_207 wl_213 vdd gnd cell_6t
Xbit_r214_c207 bl_207 br_207 wl_214 vdd gnd cell_6t
Xbit_r215_c207 bl_207 br_207 wl_215 vdd gnd cell_6t
Xbit_r216_c207 bl_207 br_207 wl_216 vdd gnd cell_6t
Xbit_r217_c207 bl_207 br_207 wl_217 vdd gnd cell_6t
Xbit_r218_c207 bl_207 br_207 wl_218 vdd gnd cell_6t
Xbit_r219_c207 bl_207 br_207 wl_219 vdd gnd cell_6t
Xbit_r220_c207 bl_207 br_207 wl_220 vdd gnd cell_6t
Xbit_r221_c207 bl_207 br_207 wl_221 vdd gnd cell_6t
Xbit_r222_c207 bl_207 br_207 wl_222 vdd gnd cell_6t
Xbit_r223_c207 bl_207 br_207 wl_223 vdd gnd cell_6t
Xbit_r224_c207 bl_207 br_207 wl_224 vdd gnd cell_6t
Xbit_r225_c207 bl_207 br_207 wl_225 vdd gnd cell_6t
Xbit_r226_c207 bl_207 br_207 wl_226 vdd gnd cell_6t
Xbit_r227_c207 bl_207 br_207 wl_227 vdd gnd cell_6t
Xbit_r228_c207 bl_207 br_207 wl_228 vdd gnd cell_6t
Xbit_r229_c207 bl_207 br_207 wl_229 vdd gnd cell_6t
Xbit_r230_c207 bl_207 br_207 wl_230 vdd gnd cell_6t
Xbit_r231_c207 bl_207 br_207 wl_231 vdd gnd cell_6t
Xbit_r232_c207 bl_207 br_207 wl_232 vdd gnd cell_6t
Xbit_r233_c207 bl_207 br_207 wl_233 vdd gnd cell_6t
Xbit_r234_c207 bl_207 br_207 wl_234 vdd gnd cell_6t
Xbit_r235_c207 bl_207 br_207 wl_235 vdd gnd cell_6t
Xbit_r236_c207 bl_207 br_207 wl_236 vdd gnd cell_6t
Xbit_r237_c207 bl_207 br_207 wl_237 vdd gnd cell_6t
Xbit_r238_c207 bl_207 br_207 wl_238 vdd gnd cell_6t
Xbit_r239_c207 bl_207 br_207 wl_239 vdd gnd cell_6t
Xbit_r240_c207 bl_207 br_207 wl_240 vdd gnd cell_6t
Xbit_r241_c207 bl_207 br_207 wl_241 vdd gnd cell_6t
Xbit_r242_c207 bl_207 br_207 wl_242 vdd gnd cell_6t
Xbit_r243_c207 bl_207 br_207 wl_243 vdd gnd cell_6t
Xbit_r244_c207 bl_207 br_207 wl_244 vdd gnd cell_6t
Xbit_r245_c207 bl_207 br_207 wl_245 vdd gnd cell_6t
Xbit_r246_c207 bl_207 br_207 wl_246 vdd gnd cell_6t
Xbit_r247_c207 bl_207 br_207 wl_247 vdd gnd cell_6t
Xbit_r248_c207 bl_207 br_207 wl_248 vdd gnd cell_6t
Xbit_r249_c207 bl_207 br_207 wl_249 vdd gnd cell_6t
Xbit_r250_c207 bl_207 br_207 wl_250 vdd gnd cell_6t
Xbit_r251_c207 bl_207 br_207 wl_251 vdd gnd cell_6t
Xbit_r252_c207 bl_207 br_207 wl_252 vdd gnd cell_6t
Xbit_r253_c207 bl_207 br_207 wl_253 vdd gnd cell_6t
Xbit_r254_c207 bl_207 br_207 wl_254 vdd gnd cell_6t
Xbit_r255_c207 bl_207 br_207 wl_255 vdd gnd cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd cell_6t
Xbit_r1_c208 bl_208 br_208 wl_1 vdd gnd cell_6t
Xbit_r2_c208 bl_208 br_208 wl_2 vdd gnd cell_6t
Xbit_r3_c208 bl_208 br_208 wl_3 vdd gnd cell_6t
Xbit_r4_c208 bl_208 br_208 wl_4 vdd gnd cell_6t
Xbit_r5_c208 bl_208 br_208 wl_5 vdd gnd cell_6t
Xbit_r6_c208 bl_208 br_208 wl_6 vdd gnd cell_6t
Xbit_r7_c208 bl_208 br_208 wl_7 vdd gnd cell_6t
Xbit_r8_c208 bl_208 br_208 wl_8 vdd gnd cell_6t
Xbit_r9_c208 bl_208 br_208 wl_9 vdd gnd cell_6t
Xbit_r10_c208 bl_208 br_208 wl_10 vdd gnd cell_6t
Xbit_r11_c208 bl_208 br_208 wl_11 vdd gnd cell_6t
Xbit_r12_c208 bl_208 br_208 wl_12 vdd gnd cell_6t
Xbit_r13_c208 bl_208 br_208 wl_13 vdd gnd cell_6t
Xbit_r14_c208 bl_208 br_208 wl_14 vdd gnd cell_6t
Xbit_r15_c208 bl_208 br_208 wl_15 vdd gnd cell_6t
Xbit_r16_c208 bl_208 br_208 wl_16 vdd gnd cell_6t
Xbit_r17_c208 bl_208 br_208 wl_17 vdd gnd cell_6t
Xbit_r18_c208 bl_208 br_208 wl_18 vdd gnd cell_6t
Xbit_r19_c208 bl_208 br_208 wl_19 vdd gnd cell_6t
Xbit_r20_c208 bl_208 br_208 wl_20 vdd gnd cell_6t
Xbit_r21_c208 bl_208 br_208 wl_21 vdd gnd cell_6t
Xbit_r22_c208 bl_208 br_208 wl_22 vdd gnd cell_6t
Xbit_r23_c208 bl_208 br_208 wl_23 vdd gnd cell_6t
Xbit_r24_c208 bl_208 br_208 wl_24 vdd gnd cell_6t
Xbit_r25_c208 bl_208 br_208 wl_25 vdd gnd cell_6t
Xbit_r26_c208 bl_208 br_208 wl_26 vdd gnd cell_6t
Xbit_r27_c208 bl_208 br_208 wl_27 vdd gnd cell_6t
Xbit_r28_c208 bl_208 br_208 wl_28 vdd gnd cell_6t
Xbit_r29_c208 bl_208 br_208 wl_29 vdd gnd cell_6t
Xbit_r30_c208 bl_208 br_208 wl_30 vdd gnd cell_6t
Xbit_r31_c208 bl_208 br_208 wl_31 vdd gnd cell_6t
Xbit_r32_c208 bl_208 br_208 wl_32 vdd gnd cell_6t
Xbit_r33_c208 bl_208 br_208 wl_33 vdd gnd cell_6t
Xbit_r34_c208 bl_208 br_208 wl_34 vdd gnd cell_6t
Xbit_r35_c208 bl_208 br_208 wl_35 vdd gnd cell_6t
Xbit_r36_c208 bl_208 br_208 wl_36 vdd gnd cell_6t
Xbit_r37_c208 bl_208 br_208 wl_37 vdd gnd cell_6t
Xbit_r38_c208 bl_208 br_208 wl_38 vdd gnd cell_6t
Xbit_r39_c208 bl_208 br_208 wl_39 vdd gnd cell_6t
Xbit_r40_c208 bl_208 br_208 wl_40 vdd gnd cell_6t
Xbit_r41_c208 bl_208 br_208 wl_41 vdd gnd cell_6t
Xbit_r42_c208 bl_208 br_208 wl_42 vdd gnd cell_6t
Xbit_r43_c208 bl_208 br_208 wl_43 vdd gnd cell_6t
Xbit_r44_c208 bl_208 br_208 wl_44 vdd gnd cell_6t
Xbit_r45_c208 bl_208 br_208 wl_45 vdd gnd cell_6t
Xbit_r46_c208 bl_208 br_208 wl_46 vdd gnd cell_6t
Xbit_r47_c208 bl_208 br_208 wl_47 vdd gnd cell_6t
Xbit_r48_c208 bl_208 br_208 wl_48 vdd gnd cell_6t
Xbit_r49_c208 bl_208 br_208 wl_49 vdd gnd cell_6t
Xbit_r50_c208 bl_208 br_208 wl_50 vdd gnd cell_6t
Xbit_r51_c208 bl_208 br_208 wl_51 vdd gnd cell_6t
Xbit_r52_c208 bl_208 br_208 wl_52 vdd gnd cell_6t
Xbit_r53_c208 bl_208 br_208 wl_53 vdd gnd cell_6t
Xbit_r54_c208 bl_208 br_208 wl_54 vdd gnd cell_6t
Xbit_r55_c208 bl_208 br_208 wl_55 vdd gnd cell_6t
Xbit_r56_c208 bl_208 br_208 wl_56 vdd gnd cell_6t
Xbit_r57_c208 bl_208 br_208 wl_57 vdd gnd cell_6t
Xbit_r58_c208 bl_208 br_208 wl_58 vdd gnd cell_6t
Xbit_r59_c208 bl_208 br_208 wl_59 vdd gnd cell_6t
Xbit_r60_c208 bl_208 br_208 wl_60 vdd gnd cell_6t
Xbit_r61_c208 bl_208 br_208 wl_61 vdd gnd cell_6t
Xbit_r62_c208 bl_208 br_208 wl_62 vdd gnd cell_6t
Xbit_r63_c208 bl_208 br_208 wl_63 vdd gnd cell_6t
Xbit_r64_c208 bl_208 br_208 wl_64 vdd gnd cell_6t
Xbit_r65_c208 bl_208 br_208 wl_65 vdd gnd cell_6t
Xbit_r66_c208 bl_208 br_208 wl_66 vdd gnd cell_6t
Xbit_r67_c208 bl_208 br_208 wl_67 vdd gnd cell_6t
Xbit_r68_c208 bl_208 br_208 wl_68 vdd gnd cell_6t
Xbit_r69_c208 bl_208 br_208 wl_69 vdd gnd cell_6t
Xbit_r70_c208 bl_208 br_208 wl_70 vdd gnd cell_6t
Xbit_r71_c208 bl_208 br_208 wl_71 vdd gnd cell_6t
Xbit_r72_c208 bl_208 br_208 wl_72 vdd gnd cell_6t
Xbit_r73_c208 bl_208 br_208 wl_73 vdd gnd cell_6t
Xbit_r74_c208 bl_208 br_208 wl_74 vdd gnd cell_6t
Xbit_r75_c208 bl_208 br_208 wl_75 vdd gnd cell_6t
Xbit_r76_c208 bl_208 br_208 wl_76 vdd gnd cell_6t
Xbit_r77_c208 bl_208 br_208 wl_77 vdd gnd cell_6t
Xbit_r78_c208 bl_208 br_208 wl_78 vdd gnd cell_6t
Xbit_r79_c208 bl_208 br_208 wl_79 vdd gnd cell_6t
Xbit_r80_c208 bl_208 br_208 wl_80 vdd gnd cell_6t
Xbit_r81_c208 bl_208 br_208 wl_81 vdd gnd cell_6t
Xbit_r82_c208 bl_208 br_208 wl_82 vdd gnd cell_6t
Xbit_r83_c208 bl_208 br_208 wl_83 vdd gnd cell_6t
Xbit_r84_c208 bl_208 br_208 wl_84 vdd gnd cell_6t
Xbit_r85_c208 bl_208 br_208 wl_85 vdd gnd cell_6t
Xbit_r86_c208 bl_208 br_208 wl_86 vdd gnd cell_6t
Xbit_r87_c208 bl_208 br_208 wl_87 vdd gnd cell_6t
Xbit_r88_c208 bl_208 br_208 wl_88 vdd gnd cell_6t
Xbit_r89_c208 bl_208 br_208 wl_89 vdd gnd cell_6t
Xbit_r90_c208 bl_208 br_208 wl_90 vdd gnd cell_6t
Xbit_r91_c208 bl_208 br_208 wl_91 vdd gnd cell_6t
Xbit_r92_c208 bl_208 br_208 wl_92 vdd gnd cell_6t
Xbit_r93_c208 bl_208 br_208 wl_93 vdd gnd cell_6t
Xbit_r94_c208 bl_208 br_208 wl_94 vdd gnd cell_6t
Xbit_r95_c208 bl_208 br_208 wl_95 vdd gnd cell_6t
Xbit_r96_c208 bl_208 br_208 wl_96 vdd gnd cell_6t
Xbit_r97_c208 bl_208 br_208 wl_97 vdd gnd cell_6t
Xbit_r98_c208 bl_208 br_208 wl_98 vdd gnd cell_6t
Xbit_r99_c208 bl_208 br_208 wl_99 vdd gnd cell_6t
Xbit_r100_c208 bl_208 br_208 wl_100 vdd gnd cell_6t
Xbit_r101_c208 bl_208 br_208 wl_101 vdd gnd cell_6t
Xbit_r102_c208 bl_208 br_208 wl_102 vdd gnd cell_6t
Xbit_r103_c208 bl_208 br_208 wl_103 vdd gnd cell_6t
Xbit_r104_c208 bl_208 br_208 wl_104 vdd gnd cell_6t
Xbit_r105_c208 bl_208 br_208 wl_105 vdd gnd cell_6t
Xbit_r106_c208 bl_208 br_208 wl_106 vdd gnd cell_6t
Xbit_r107_c208 bl_208 br_208 wl_107 vdd gnd cell_6t
Xbit_r108_c208 bl_208 br_208 wl_108 vdd gnd cell_6t
Xbit_r109_c208 bl_208 br_208 wl_109 vdd gnd cell_6t
Xbit_r110_c208 bl_208 br_208 wl_110 vdd gnd cell_6t
Xbit_r111_c208 bl_208 br_208 wl_111 vdd gnd cell_6t
Xbit_r112_c208 bl_208 br_208 wl_112 vdd gnd cell_6t
Xbit_r113_c208 bl_208 br_208 wl_113 vdd gnd cell_6t
Xbit_r114_c208 bl_208 br_208 wl_114 vdd gnd cell_6t
Xbit_r115_c208 bl_208 br_208 wl_115 vdd gnd cell_6t
Xbit_r116_c208 bl_208 br_208 wl_116 vdd gnd cell_6t
Xbit_r117_c208 bl_208 br_208 wl_117 vdd gnd cell_6t
Xbit_r118_c208 bl_208 br_208 wl_118 vdd gnd cell_6t
Xbit_r119_c208 bl_208 br_208 wl_119 vdd gnd cell_6t
Xbit_r120_c208 bl_208 br_208 wl_120 vdd gnd cell_6t
Xbit_r121_c208 bl_208 br_208 wl_121 vdd gnd cell_6t
Xbit_r122_c208 bl_208 br_208 wl_122 vdd gnd cell_6t
Xbit_r123_c208 bl_208 br_208 wl_123 vdd gnd cell_6t
Xbit_r124_c208 bl_208 br_208 wl_124 vdd gnd cell_6t
Xbit_r125_c208 bl_208 br_208 wl_125 vdd gnd cell_6t
Xbit_r126_c208 bl_208 br_208 wl_126 vdd gnd cell_6t
Xbit_r127_c208 bl_208 br_208 wl_127 vdd gnd cell_6t
Xbit_r128_c208 bl_208 br_208 wl_128 vdd gnd cell_6t
Xbit_r129_c208 bl_208 br_208 wl_129 vdd gnd cell_6t
Xbit_r130_c208 bl_208 br_208 wl_130 vdd gnd cell_6t
Xbit_r131_c208 bl_208 br_208 wl_131 vdd gnd cell_6t
Xbit_r132_c208 bl_208 br_208 wl_132 vdd gnd cell_6t
Xbit_r133_c208 bl_208 br_208 wl_133 vdd gnd cell_6t
Xbit_r134_c208 bl_208 br_208 wl_134 vdd gnd cell_6t
Xbit_r135_c208 bl_208 br_208 wl_135 vdd gnd cell_6t
Xbit_r136_c208 bl_208 br_208 wl_136 vdd gnd cell_6t
Xbit_r137_c208 bl_208 br_208 wl_137 vdd gnd cell_6t
Xbit_r138_c208 bl_208 br_208 wl_138 vdd gnd cell_6t
Xbit_r139_c208 bl_208 br_208 wl_139 vdd gnd cell_6t
Xbit_r140_c208 bl_208 br_208 wl_140 vdd gnd cell_6t
Xbit_r141_c208 bl_208 br_208 wl_141 vdd gnd cell_6t
Xbit_r142_c208 bl_208 br_208 wl_142 vdd gnd cell_6t
Xbit_r143_c208 bl_208 br_208 wl_143 vdd gnd cell_6t
Xbit_r144_c208 bl_208 br_208 wl_144 vdd gnd cell_6t
Xbit_r145_c208 bl_208 br_208 wl_145 vdd gnd cell_6t
Xbit_r146_c208 bl_208 br_208 wl_146 vdd gnd cell_6t
Xbit_r147_c208 bl_208 br_208 wl_147 vdd gnd cell_6t
Xbit_r148_c208 bl_208 br_208 wl_148 vdd gnd cell_6t
Xbit_r149_c208 bl_208 br_208 wl_149 vdd gnd cell_6t
Xbit_r150_c208 bl_208 br_208 wl_150 vdd gnd cell_6t
Xbit_r151_c208 bl_208 br_208 wl_151 vdd gnd cell_6t
Xbit_r152_c208 bl_208 br_208 wl_152 vdd gnd cell_6t
Xbit_r153_c208 bl_208 br_208 wl_153 vdd gnd cell_6t
Xbit_r154_c208 bl_208 br_208 wl_154 vdd gnd cell_6t
Xbit_r155_c208 bl_208 br_208 wl_155 vdd gnd cell_6t
Xbit_r156_c208 bl_208 br_208 wl_156 vdd gnd cell_6t
Xbit_r157_c208 bl_208 br_208 wl_157 vdd gnd cell_6t
Xbit_r158_c208 bl_208 br_208 wl_158 vdd gnd cell_6t
Xbit_r159_c208 bl_208 br_208 wl_159 vdd gnd cell_6t
Xbit_r160_c208 bl_208 br_208 wl_160 vdd gnd cell_6t
Xbit_r161_c208 bl_208 br_208 wl_161 vdd gnd cell_6t
Xbit_r162_c208 bl_208 br_208 wl_162 vdd gnd cell_6t
Xbit_r163_c208 bl_208 br_208 wl_163 vdd gnd cell_6t
Xbit_r164_c208 bl_208 br_208 wl_164 vdd gnd cell_6t
Xbit_r165_c208 bl_208 br_208 wl_165 vdd gnd cell_6t
Xbit_r166_c208 bl_208 br_208 wl_166 vdd gnd cell_6t
Xbit_r167_c208 bl_208 br_208 wl_167 vdd gnd cell_6t
Xbit_r168_c208 bl_208 br_208 wl_168 vdd gnd cell_6t
Xbit_r169_c208 bl_208 br_208 wl_169 vdd gnd cell_6t
Xbit_r170_c208 bl_208 br_208 wl_170 vdd gnd cell_6t
Xbit_r171_c208 bl_208 br_208 wl_171 vdd gnd cell_6t
Xbit_r172_c208 bl_208 br_208 wl_172 vdd gnd cell_6t
Xbit_r173_c208 bl_208 br_208 wl_173 vdd gnd cell_6t
Xbit_r174_c208 bl_208 br_208 wl_174 vdd gnd cell_6t
Xbit_r175_c208 bl_208 br_208 wl_175 vdd gnd cell_6t
Xbit_r176_c208 bl_208 br_208 wl_176 vdd gnd cell_6t
Xbit_r177_c208 bl_208 br_208 wl_177 vdd gnd cell_6t
Xbit_r178_c208 bl_208 br_208 wl_178 vdd gnd cell_6t
Xbit_r179_c208 bl_208 br_208 wl_179 vdd gnd cell_6t
Xbit_r180_c208 bl_208 br_208 wl_180 vdd gnd cell_6t
Xbit_r181_c208 bl_208 br_208 wl_181 vdd gnd cell_6t
Xbit_r182_c208 bl_208 br_208 wl_182 vdd gnd cell_6t
Xbit_r183_c208 bl_208 br_208 wl_183 vdd gnd cell_6t
Xbit_r184_c208 bl_208 br_208 wl_184 vdd gnd cell_6t
Xbit_r185_c208 bl_208 br_208 wl_185 vdd gnd cell_6t
Xbit_r186_c208 bl_208 br_208 wl_186 vdd gnd cell_6t
Xbit_r187_c208 bl_208 br_208 wl_187 vdd gnd cell_6t
Xbit_r188_c208 bl_208 br_208 wl_188 vdd gnd cell_6t
Xbit_r189_c208 bl_208 br_208 wl_189 vdd gnd cell_6t
Xbit_r190_c208 bl_208 br_208 wl_190 vdd gnd cell_6t
Xbit_r191_c208 bl_208 br_208 wl_191 vdd gnd cell_6t
Xbit_r192_c208 bl_208 br_208 wl_192 vdd gnd cell_6t
Xbit_r193_c208 bl_208 br_208 wl_193 vdd gnd cell_6t
Xbit_r194_c208 bl_208 br_208 wl_194 vdd gnd cell_6t
Xbit_r195_c208 bl_208 br_208 wl_195 vdd gnd cell_6t
Xbit_r196_c208 bl_208 br_208 wl_196 vdd gnd cell_6t
Xbit_r197_c208 bl_208 br_208 wl_197 vdd gnd cell_6t
Xbit_r198_c208 bl_208 br_208 wl_198 vdd gnd cell_6t
Xbit_r199_c208 bl_208 br_208 wl_199 vdd gnd cell_6t
Xbit_r200_c208 bl_208 br_208 wl_200 vdd gnd cell_6t
Xbit_r201_c208 bl_208 br_208 wl_201 vdd gnd cell_6t
Xbit_r202_c208 bl_208 br_208 wl_202 vdd gnd cell_6t
Xbit_r203_c208 bl_208 br_208 wl_203 vdd gnd cell_6t
Xbit_r204_c208 bl_208 br_208 wl_204 vdd gnd cell_6t
Xbit_r205_c208 bl_208 br_208 wl_205 vdd gnd cell_6t
Xbit_r206_c208 bl_208 br_208 wl_206 vdd gnd cell_6t
Xbit_r207_c208 bl_208 br_208 wl_207 vdd gnd cell_6t
Xbit_r208_c208 bl_208 br_208 wl_208 vdd gnd cell_6t
Xbit_r209_c208 bl_208 br_208 wl_209 vdd gnd cell_6t
Xbit_r210_c208 bl_208 br_208 wl_210 vdd gnd cell_6t
Xbit_r211_c208 bl_208 br_208 wl_211 vdd gnd cell_6t
Xbit_r212_c208 bl_208 br_208 wl_212 vdd gnd cell_6t
Xbit_r213_c208 bl_208 br_208 wl_213 vdd gnd cell_6t
Xbit_r214_c208 bl_208 br_208 wl_214 vdd gnd cell_6t
Xbit_r215_c208 bl_208 br_208 wl_215 vdd gnd cell_6t
Xbit_r216_c208 bl_208 br_208 wl_216 vdd gnd cell_6t
Xbit_r217_c208 bl_208 br_208 wl_217 vdd gnd cell_6t
Xbit_r218_c208 bl_208 br_208 wl_218 vdd gnd cell_6t
Xbit_r219_c208 bl_208 br_208 wl_219 vdd gnd cell_6t
Xbit_r220_c208 bl_208 br_208 wl_220 vdd gnd cell_6t
Xbit_r221_c208 bl_208 br_208 wl_221 vdd gnd cell_6t
Xbit_r222_c208 bl_208 br_208 wl_222 vdd gnd cell_6t
Xbit_r223_c208 bl_208 br_208 wl_223 vdd gnd cell_6t
Xbit_r224_c208 bl_208 br_208 wl_224 vdd gnd cell_6t
Xbit_r225_c208 bl_208 br_208 wl_225 vdd gnd cell_6t
Xbit_r226_c208 bl_208 br_208 wl_226 vdd gnd cell_6t
Xbit_r227_c208 bl_208 br_208 wl_227 vdd gnd cell_6t
Xbit_r228_c208 bl_208 br_208 wl_228 vdd gnd cell_6t
Xbit_r229_c208 bl_208 br_208 wl_229 vdd gnd cell_6t
Xbit_r230_c208 bl_208 br_208 wl_230 vdd gnd cell_6t
Xbit_r231_c208 bl_208 br_208 wl_231 vdd gnd cell_6t
Xbit_r232_c208 bl_208 br_208 wl_232 vdd gnd cell_6t
Xbit_r233_c208 bl_208 br_208 wl_233 vdd gnd cell_6t
Xbit_r234_c208 bl_208 br_208 wl_234 vdd gnd cell_6t
Xbit_r235_c208 bl_208 br_208 wl_235 vdd gnd cell_6t
Xbit_r236_c208 bl_208 br_208 wl_236 vdd gnd cell_6t
Xbit_r237_c208 bl_208 br_208 wl_237 vdd gnd cell_6t
Xbit_r238_c208 bl_208 br_208 wl_238 vdd gnd cell_6t
Xbit_r239_c208 bl_208 br_208 wl_239 vdd gnd cell_6t
Xbit_r240_c208 bl_208 br_208 wl_240 vdd gnd cell_6t
Xbit_r241_c208 bl_208 br_208 wl_241 vdd gnd cell_6t
Xbit_r242_c208 bl_208 br_208 wl_242 vdd gnd cell_6t
Xbit_r243_c208 bl_208 br_208 wl_243 vdd gnd cell_6t
Xbit_r244_c208 bl_208 br_208 wl_244 vdd gnd cell_6t
Xbit_r245_c208 bl_208 br_208 wl_245 vdd gnd cell_6t
Xbit_r246_c208 bl_208 br_208 wl_246 vdd gnd cell_6t
Xbit_r247_c208 bl_208 br_208 wl_247 vdd gnd cell_6t
Xbit_r248_c208 bl_208 br_208 wl_248 vdd gnd cell_6t
Xbit_r249_c208 bl_208 br_208 wl_249 vdd gnd cell_6t
Xbit_r250_c208 bl_208 br_208 wl_250 vdd gnd cell_6t
Xbit_r251_c208 bl_208 br_208 wl_251 vdd gnd cell_6t
Xbit_r252_c208 bl_208 br_208 wl_252 vdd gnd cell_6t
Xbit_r253_c208 bl_208 br_208 wl_253 vdd gnd cell_6t
Xbit_r254_c208 bl_208 br_208 wl_254 vdd gnd cell_6t
Xbit_r255_c208 bl_208 br_208 wl_255 vdd gnd cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd cell_6t
Xbit_r1_c209 bl_209 br_209 wl_1 vdd gnd cell_6t
Xbit_r2_c209 bl_209 br_209 wl_2 vdd gnd cell_6t
Xbit_r3_c209 bl_209 br_209 wl_3 vdd gnd cell_6t
Xbit_r4_c209 bl_209 br_209 wl_4 vdd gnd cell_6t
Xbit_r5_c209 bl_209 br_209 wl_5 vdd gnd cell_6t
Xbit_r6_c209 bl_209 br_209 wl_6 vdd gnd cell_6t
Xbit_r7_c209 bl_209 br_209 wl_7 vdd gnd cell_6t
Xbit_r8_c209 bl_209 br_209 wl_8 vdd gnd cell_6t
Xbit_r9_c209 bl_209 br_209 wl_9 vdd gnd cell_6t
Xbit_r10_c209 bl_209 br_209 wl_10 vdd gnd cell_6t
Xbit_r11_c209 bl_209 br_209 wl_11 vdd gnd cell_6t
Xbit_r12_c209 bl_209 br_209 wl_12 vdd gnd cell_6t
Xbit_r13_c209 bl_209 br_209 wl_13 vdd gnd cell_6t
Xbit_r14_c209 bl_209 br_209 wl_14 vdd gnd cell_6t
Xbit_r15_c209 bl_209 br_209 wl_15 vdd gnd cell_6t
Xbit_r16_c209 bl_209 br_209 wl_16 vdd gnd cell_6t
Xbit_r17_c209 bl_209 br_209 wl_17 vdd gnd cell_6t
Xbit_r18_c209 bl_209 br_209 wl_18 vdd gnd cell_6t
Xbit_r19_c209 bl_209 br_209 wl_19 vdd gnd cell_6t
Xbit_r20_c209 bl_209 br_209 wl_20 vdd gnd cell_6t
Xbit_r21_c209 bl_209 br_209 wl_21 vdd gnd cell_6t
Xbit_r22_c209 bl_209 br_209 wl_22 vdd gnd cell_6t
Xbit_r23_c209 bl_209 br_209 wl_23 vdd gnd cell_6t
Xbit_r24_c209 bl_209 br_209 wl_24 vdd gnd cell_6t
Xbit_r25_c209 bl_209 br_209 wl_25 vdd gnd cell_6t
Xbit_r26_c209 bl_209 br_209 wl_26 vdd gnd cell_6t
Xbit_r27_c209 bl_209 br_209 wl_27 vdd gnd cell_6t
Xbit_r28_c209 bl_209 br_209 wl_28 vdd gnd cell_6t
Xbit_r29_c209 bl_209 br_209 wl_29 vdd gnd cell_6t
Xbit_r30_c209 bl_209 br_209 wl_30 vdd gnd cell_6t
Xbit_r31_c209 bl_209 br_209 wl_31 vdd gnd cell_6t
Xbit_r32_c209 bl_209 br_209 wl_32 vdd gnd cell_6t
Xbit_r33_c209 bl_209 br_209 wl_33 vdd gnd cell_6t
Xbit_r34_c209 bl_209 br_209 wl_34 vdd gnd cell_6t
Xbit_r35_c209 bl_209 br_209 wl_35 vdd gnd cell_6t
Xbit_r36_c209 bl_209 br_209 wl_36 vdd gnd cell_6t
Xbit_r37_c209 bl_209 br_209 wl_37 vdd gnd cell_6t
Xbit_r38_c209 bl_209 br_209 wl_38 vdd gnd cell_6t
Xbit_r39_c209 bl_209 br_209 wl_39 vdd gnd cell_6t
Xbit_r40_c209 bl_209 br_209 wl_40 vdd gnd cell_6t
Xbit_r41_c209 bl_209 br_209 wl_41 vdd gnd cell_6t
Xbit_r42_c209 bl_209 br_209 wl_42 vdd gnd cell_6t
Xbit_r43_c209 bl_209 br_209 wl_43 vdd gnd cell_6t
Xbit_r44_c209 bl_209 br_209 wl_44 vdd gnd cell_6t
Xbit_r45_c209 bl_209 br_209 wl_45 vdd gnd cell_6t
Xbit_r46_c209 bl_209 br_209 wl_46 vdd gnd cell_6t
Xbit_r47_c209 bl_209 br_209 wl_47 vdd gnd cell_6t
Xbit_r48_c209 bl_209 br_209 wl_48 vdd gnd cell_6t
Xbit_r49_c209 bl_209 br_209 wl_49 vdd gnd cell_6t
Xbit_r50_c209 bl_209 br_209 wl_50 vdd gnd cell_6t
Xbit_r51_c209 bl_209 br_209 wl_51 vdd gnd cell_6t
Xbit_r52_c209 bl_209 br_209 wl_52 vdd gnd cell_6t
Xbit_r53_c209 bl_209 br_209 wl_53 vdd gnd cell_6t
Xbit_r54_c209 bl_209 br_209 wl_54 vdd gnd cell_6t
Xbit_r55_c209 bl_209 br_209 wl_55 vdd gnd cell_6t
Xbit_r56_c209 bl_209 br_209 wl_56 vdd gnd cell_6t
Xbit_r57_c209 bl_209 br_209 wl_57 vdd gnd cell_6t
Xbit_r58_c209 bl_209 br_209 wl_58 vdd gnd cell_6t
Xbit_r59_c209 bl_209 br_209 wl_59 vdd gnd cell_6t
Xbit_r60_c209 bl_209 br_209 wl_60 vdd gnd cell_6t
Xbit_r61_c209 bl_209 br_209 wl_61 vdd gnd cell_6t
Xbit_r62_c209 bl_209 br_209 wl_62 vdd gnd cell_6t
Xbit_r63_c209 bl_209 br_209 wl_63 vdd gnd cell_6t
Xbit_r64_c209 bl_209 br_209 wl_64 vdd gnd cell_6t
Xbit_r65_c209 bl_209 br_209 wl_65 vdd gnd cell_6t
Xbit_r66_c209 bl_209 br_209 wl_66 vdd gnd cell_6t
Xbit_r67_c209 bl_209 br_209 wl_67 vdd gnd cell_6t
Xbit_r68_c209 bl_209 br_209 wl_68 vdd gnd cell_6t
Xbit_r69_c209 bl_209 br_209 wl_69 vdd gnd cell_6t
Xbit_r70_c209 bl_209 br_209 wl_70 vdd gnd cell_6t
Xbit_r71_c209 bl_209 br_209 wl_71 vdd gnd cell_6t
Xbit_r72_c209 bl_209 br_209 wl_72 vdd gnd cell_6t
Xbit_r73_c209 bl_209 br_209 wl_73 vdd gnd cell_6t
Xbit_r74_c209 bl_209 br_209 wl_74 vdd gnd cell_6t
Xbit_r75_c209 bl_209 br_209 wl_75 vdd gnd cell_6t
Xbit_r76_c209 bl_209 br_209 wl_76 vdd gnd cell_6t
Xbit_r77_c209 bl_209 br_209 wl_77 vdd gnd cell_6t
Xbit_r78_c209 bl_209 br_209 wl_78 vdd gnd cell_6t
Xbit_r79_c209 bl_209 br_209 wl_79 vdd gnd cell_6t
Xbit_r80_c209 bl_209 br_209 wl_80 vdd gnd cell_6t
Xbit_r81_c209 bl_209 br_209 wl_81 vdd gnd cell_6t
Xbit_r82_c209 bl_209 br_209 wl_82 vdd gnd cell_6t
Xbit_r83_c209 bl_209 br_209 wl_83 vdd gnd cell_6t
Xbit_r84_c209 bl_209 br_209 wl_84 vdd gnd cell_6t
Xbit_r85_c209 bl_209 br_209 wl_85 vdd gnd cell_6t
Xbit_r86_c209 bl_209 br_209 wl_86 vdd gnd cell_6t
Xbit_r87_c209 bl_209 br_209 wl_87 vdd gnd cell_6t
Xbit_r88_c209 bl_209 br_209 wl_88 vdd gnd cell_6t
Xbit_r89_c209 bl_209 br_209 wl_89 vdd gnd cell_6t
Xbit_r90_c209 bl_209 br_209 wl_90 vdd gnd cell_6t
Xbit_r91_c209 bl_209 br_209 wl_91 vdd gnd cell_6t
Xbit_r92_c209 bl_209 br_209 wl_92 vdd gnd cell_6t
Xbit_r93_c209 bl_209 br_209 wl_93 vdd gnd cell_6t
Xbit_r94_c209 bl_209 br_209 wl_94 vdd gnd cell_6t
Xbit_r95_c209 bl_209 br_209 wl_95 vdd gnd cell_6t
Xbit_r96_c209 bl_209 br_209 wl_96 vdd gnd cell_6t
Xbit_r97_c209 bl_209 br_209 wl_97 vdd gnd cell_6t
Xbit_r98_c209 bl_209 br_209 wl_98 vdd gnd cell_6t
Xbit_r99_c209 bl_209 br_209 wl_99 vdd gnd cell_6t
Xbit_r100_c209 bl_209 br_209 wl_100 vdd gnd cell_6t
Xbit_r101_c209 bl_209 br_209 wl_101 vdd gnd cell_6t
Xbit_r102_c209 bl_209 br_209 wl_102 vdd gnd cell_6t
Xbit_r103_c209 bl_209 br_209 wl_103 vdd gnd cell_6t
Xbit_r104_c209 bl_209 br_209 wl_104 vdd gnd cell_6t
Xbit_r105_c209 bl_209 br_209 wl_105 vdd gnd cell_6t
Xbit_r106_c209 bl_209 br_209 wl_106 vdd gnd cell_6t
Xbit_r107_c209 bl_209 br_209 wl_107 vdd gnd cell_6t
Xbit_r108_c209 bl_209 br_209 wl_108 vdd gnd cell_6t
Xbit_r109_c209 bl_209 br_209 wl_109 vdd gnd cell_6t
Xbit_r110_c209 bl_209 br_209 wl_110 vdd gnd cell_6t
Xbit_r111_c209 bl_209 br_209 wl_111 vdd gnd cell_6t
Xbit_r112_c209 bl_209 br_209 wl_112 vdd gnd cell_6t
Xbit_r113_c209 bl_209 br_209 wl_113 vdd gnd cell_6t
Xbit_r114_c209 bl_209 br_209 wl_114 vdd gnd cell_6t
Xbit_r115_c209 bl_209 br_209 wl_115 vdd gnd cell_6t
Xbit_r116_c209 bl_209 br_209 wl_116 vdd gnd cell_6t
Xbit_r117_c209 bl_209 br_209 wl_117 vdd gnd cell_6t
Xbit_r118_c209 bl_209 br_209 wl_118 vdd gnd cell_6t
Xbit_r119_c209 bl_209 br_209 wl_119 vdd gnd cell_6t
Xbit_r120_c209 bl_209 br_209 wl_120 vdd gnd cell_6t
Xbit_r121_c209 bl_209 br_209 wl_121 vdd gnd cell_6t
Xbit_r122_c209 bl_209 br_209 wl_122 vdd gnd cell_6t
Xbit_r123_c209 bl_209 br_209 wl_123 vdd gnd cell_6t
Xbit_r124_c209 bl_209 br_209 wl_124 vdd gnd cell_6t
Xbit_r125_c209 bl_209 br_209 wl_125 vdd gnd cell_6t
Xbit_r126_c209 bl_209 br_209 wl_126 vdd gnd cell_6t
Xbit_r127_c209 bl_209 br_209 wl_127 vdd gnd cell_6t
Xbit_r128_c209 bl_209 br_209 wl_128 vdd gnd cell_6t
Xbit_r129_c209 bl_209 br_209 wl_129 vdd gnd cell_6t
Xbit_r130_c209 bl_209 br_209 wl_130 vdd gnd cell_6t
Xbit_r131_c209 bl_209 br_209 wl_131 vdd gnd cell_6t
Xbit_r132_c209 bl_209 br_209 wl_132 vdd gnd cell_6t
Xbit_r133_c209 bl_209 br_209 wl_133 vdd gnd cell_6t
Xbit_r134_c209 bl_209 br_209 wl_134 vdd gnd cell_6t
Xbit_r135_c209 bl_209 br_209 wl_135 vdd gnd cell_6t
Xbit_r136_c209 bl_209 br_209 wl_136 vdd gnd cell_6t
Xbit_r137_c209 bl_209 br_209 wl_137 vdd gnd cell_6t
Xbit_r138_c209 bl_209 br_209 wl_138 vdd gnd cell_6t
Xbit_r139_c209 bl_209 br_209 wl_139 vdd gnd cell_6t
Xbit_r140_c209 bl_209 br_209 wl_140 vdd gnd cell_6t
Xbit_r141_c209 bl_209 br_209 wl_141 vdd gnd cell_6t
Xbit_r142_c209 bl_209 br_209 wl_142 vdd gnd cell_6t
Xbit_r143_c209 bl_209 br_209 wl_143 vdd gnd cell_6t
Xbit_r144_c209 bl_209 br_209 wl_144 vdd gnd cell_6t
Xbit_r145_c209 bl_209 br_209 wl_145 vdd gnd cell_6t
Xbit_r146_c209 bl_209 br_209 wl_146 vdd gnd cell_6t
Xbit_r147_c209 bl_209 br_209 wl_147 vdd gnd cell_6t
Xbit_r148_c209 bl_209 br_209 wl_148 vdd gnd cell_6t
Xbit_r149_c209 bl_209 br_209 wl_149 vdd gnd cell_6t
Xbit_r150_c209 bl_209 br_209 wl_150 vdd gnd cell_6t
Xbit_r151_c209 bl_209 br_209 wl_151 vdd gnd cell_6t
Xbit_r152_c209 bl_209 br_209 wl_152 vdd gnd cell_6t
Xbit_r153_c209 bl_209 br_209 wl_153 vdd gnd cell_6t
Xbit_r154_c209 bl_209 br_209 wl_154 vdd gnd cell_6t
Xbit_r155_c209 bl_209 br_209 wl_155 vdd gnd cell_6t
Xbit_r156_c209 bl_209 br_209 wl_156 vdd gnd cell_6t
Xbit_r157_c209 bl_209 br_209 wl_157 vdd gnd cell_6t
Xbit_r158_c209 bl_209 br_209 wl_158 vdd gnd cell_6t
Xbit_r159_c209 bl_209 br_209 wl_159 vdd gnd cell_6t
Xbit_r160_c209 bl_209 br_209 wl_160 vdd gnd cell_6t
Xbit_r161_c209 bl_209 br_209 wl_161 vdd gnd cell_6t
Xbit_r162_c209 bl_209 br_209 wl_162 vdd gnd cell_6t
Xbit_r163_c209 bl_209 br_209 wl_163 vdd gnd cell_6t
Xbit_r164_c209 bl_209 br_209 wl_164 vdd gnd cell_6t
Xbit_r165_c209 bl_209 br_209 wl_165 vdd gnd cell_6t
Xbit_r166_c209 bl_209 br_209 wl_166 vdd gnd cell_6t
Xbit_r167_c209 bl_209 br_209 wl_167 vdd gnd cell_6t
Xbit_r168_c209 bl_209 br_209 wl_168 vdd gnd cell_6t
Xbit_r169_c209 bl_209 br_209 wl_169 vdd gnd cell_6t
Xbit_r170_c209 bl_209 br_209 wl_170 vdd gnd cell_6t
Xbit_r171_c209 bl_209 br_209 wl_171 vdd gnd cell_6t
Xbit_r172_c209 bl_209 br_209 wl_172 vdd gnd cell_6t
Xbit_r173_c209 bl_209 br_209 wl_173 vdd gnd cell_6t
Xbit_r174_c209 bl_209 br_209 wl_174 vdd gnd cell_6t
Xbit_r175_c209 bl_209 br_209 wl_175 vdd gnd cell_6t
Xbit_r176_c209 bl_209 br_209 wl_176 vdd gnd cell_6t
Xbit_r177_c209 bl_209 br_209 wl_177 vdd gnd cell_6t
Xbit_r178_c209 bl_209 br_209 wl_178 vdd gnd cell_6t
Xbit_r179_c209 bl_209 br_209 wl_179 vdd gnd cell_6t
Xbit_r180_c209 bl_209 br_209 wl_180 vdd gnd cell_6t
Xbit_r181_c209 bl_209 br_209 wl_181 vdd gnd cell_6t
Xbit_r182_c209 bl_209 br_209 wl_182 vdd gnd cell_6t
Xbit_r183_c209 bl_209 br_209 wl_183 vdd gnd cell_6t
Xbit_r184_c209 bl_209 br_209 wl_184 vdd gnd cell_6t
Xbit_r185_c209 bl_209 br_209 wl_185 vdd gnd cell_6t
Xbit_r186_c209 bl_209 br_209 wl_186 vdd gnd cell_6t
Xbit_r187_c209 bl_209 br_209 wl_187 vdd gnd cell_6t
Xbit_r188_c209 bl_209 br_209 wl_188 vdd gnd cell_6t
Xbit_r189_c209 bl_209 br_209 wl_189 vdd gnd cell_6t
Xbit_r190_c209 bl_209 br_209 wl_190 vdd gnd cell_6t
Xbit_r191_c209 bl_209 br_209 wl_191 vdd gnd cell_6t
Xbit_r192_c209 bl_209 br_209 wl_192 vdd gnd cell_6t
Xbit_r193_c209 bl_209 br_209 wl_193 vdd gnd cell_6t
Xbit_r194_c209 bl_209 br_209 wl_194 vdd gnd cell_6t
Xbit_r195_c209 bl_209 br_209 wl_195 vdd gnd cell_6t
Xbit_r196_c209 bl_209 br_209 wl_196 vdd gnd cell_6t
Xbit_r197_c209 bl_209 br_209 wl_197 vdd gnd cell_6t
Xbit_r198_c209 bl_209 br_209 wl_198 vdd gnd cell_6t
Xbit_r199_c209 bl_209 br_209 wl_199 vdd gnd cell_6t
Xbit_r200_c209 bl_209 br_209 wl_200 vdd gnd cell_6t
Xbit_r201_c209 bl_209 br_209 wl_201 vdd gnd cell_6t
Xbit_r202_c209 bl_209 br_209 wl_202 vdd gnd cell_6t
Xbit_r203_c209 bl_209 br_209 wl_203 vdd gnd cell_6t
Xbit_r204_c209 bl_209 br_209 wl_204 vdd gnd cell_6t
Xbit_r205_c209 bl_209 br_209 wl_205 vdd gnd cell_6t
Xbit_r206_c209 bl_209 br_209 wl_206 vdd gnd cell_6t
Xbit_r207_c209 bl_209 br_209 wl_207 vdd gnd cell_6t
Xbit_r208_c209 bl_209 br_209 wl_208 vdd gnd cell_6t
Xbit_r209_c209 bl_209 br_209 wl_209 vdd gnd cell_6t
Xbit_r210_c209 bl_209 br_209 wl_210 vdd gnd cell_6t
Xbit_r211_c209 bl_209 br_209 wl_211 vdd gnd cell_6t
Xbit_r212_c209 bl_209 br_209 wl_212 vdd gnd cell_6t
Xbit_r213_c209 bl_209 br_209 wl_213 vdd gnd cell_6t
Xbit_r214_c209 bl_209 br_209 wl_214 vdd gnd cell_6t
Xbit_r215_c209 bl_209 br_209 wl_215 vdd gnd cell_6t
Xbit_r216_c209 bl_209 br_209 wl_216 vdd gnd cell_6t
Xbit_r217_c209 bl_209 br_209 wl_217 vdd gnd cell_6t
Xbit_r218_c209 bl_209 br_209 wl_218 vdd gnd cell_6t
Xbit_r219_c209 bl_209 br_209 wl_219 vdd gnd cell_6t
Xbit_r220_c209 bl_209 br_209 wl_220 vdd gnd cell_6t
Xbit_r221_c209 bl_209 br_209 wl_221 vdd gnd cell_6t
Xbit_r222_c209 bl_209 br_209 wl_222 vdd gnd cell_6t
Xbit_r223_c209 bl_209 br_209 wl_223 vdd gnd cell_6t
Xbit_r224_c209 bl_209 br_209 wl_224 vdd gnd cell_6t
Xbit_r225_c209 bl_209 br_209 wl_225 vdd gnd cell_6t
Xbit_r226_c209 bl_209 br_209 wl_226 vdd gnd cell_6t
Xbit_r227_c209 bl_209 br_209 wl_227 vdd gnd cell_6t
Xbit_r228_c209 bl_209 br_209 wl_228 vdd gnd cell_6t
Xbit_r229_c209 bl_209 br_209 wl_229 vdd gnd cell_6t
Xbit_r230_c209 bl_209 br_209 wl_230 vdd gnd cell_6t
Xbit_r231_c209 bl_209 br_209 wl_231 vdd gnd cell_6t
Xbit_r232_c209 bl_209 br_209 wl_232 vdd gnd cell_6t
Xbit_r233_c209 bl_209 br_209 wl_233 vdd gnd cell_6t
Xbit_r234_c209 bl_209 br_209 wl_234 vdd gnd cell_6t
Xbit_r235_c209 bl_209 br_209 wl_235 vdd gnd cell_6t
Xbit_r236_c209 bl_209 br_209 wl_236 vdd gnd cell_6t
Xbit_r237_c209 bl_209 br_209 wl_237 vdd gnd cell_6t
Xbit_r238_c209 bl_209 br_209 wl_238 vdd gnd cell_6t
Xbit_r239_c209 bl_209 br_209 wl_239 vdd gnd cell_6t
Xbit_r240_c209 bl_209 br_209 wl_240 vdd gnd cell_6t
Xbit_r241_c209 bl_209 br_209 wl_241 vdd gnd cell_6t
Xbit_r242_c209 bl_209 br_209 wl_242 vdd gnd cell_6t
Xbit_r243_c209 bl_209 br_209 wl_243 vdd gnd cell_6t
Xbit_r244_c209 bl_209 br_209 wl_244 vdd gnd cell_6t
Xbit_r245_c209 bl_209 br_209 wl_245 vdd gnd cell_6t
Xbit_r246_c209 bl_209 br_209 wl_246 vdd gnd cell_6t
Xbit_r247_c209 bl_209 br_209 wl_247 vdd gnd cell_6t
Xbit_r248_c209 bl_209 br_209 wl_248 vdd gnd cell_6t
Xbit_r249_c209 bl_209 br_209 wl_249 vdd gnd cell_6t
Xbit_r250_c209 bl_209 br_209 wl_250 vdd gnd cell_6t
Xbit_r251_c209 bl_209 br_209 wl_251 vdd gnd cell_6t
Xbit_r252_c209 bl_209 br_209 wl_252 vdd gnd cell_6t
Xbit_r253_c209 bl_209 br_209 wl_253 vdd gnd cell_6t
Xbit_r254_c209 bl_209 br_209 wl_254 vdd gnd cell_6t
Xbit_r255_c209 bl_209 br_209 wl_255 vdd gnd cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd cell_6t
Xbit_r1_c210 bl_210 br_210 wl_1 vdd gnd cell_6t
Xbit_r2_c210 bl_210 br_210 wl_2 vdd gnd cell_6t
Xbit_r3_c210 bl_210 br_210 wl_3 vdd gnd cell_6t
Xbit_r4_c210 bl_210 br_210 wl_4 vdd gnd cell_6t
Xbit_r5_c210 bl_210 br_210 wl_5 vdd gnd cell_6t
Xbit_r6_c210 bl_210 br_210 wl_6 vdd gnd cell_6t
Xbit_r7_c210 bl_210 br_210 wl_7 vdd gnd cell_6t
Xbit_r8_c210 bl_210 br_210 wl_8 vdd gnd cell_6t
Xbit_r9_c210 bl_210 br_210 wl_9 vdd gnd cell_6t
Xbit_r10_c210 bl_210 br_210 wl_10 vdd gnd cell_6t
Xbit_r11_c210 bl_210 br_210 wl_11 vdd gnd cell_6t
Xbit_r12_c210 bl_210 br_210 wl_12 vdd gnd cell_6t
Xbit_r13_c210 bl_210 br_210 wl_13 vdd gnd cell_6t
Xbit_r14_c210 bl_210 br_210 wl_14 vdd gnd cell_6t
Xbit_r15_c210 bl_210 br_210 wl_15 vdd gnd cell_6t
Xbit_r16_c210 bl_210 br_210 wl_16 vdd gnd cell_6t
Xbit_r17_c210 bl_210 br_210 wl_17 vdd gnd cell_6t
Xbit_r18_c210 bl_210 br_210 wl_18 vdd gnd cell_6t
Xbit_r19_c210 bl_210 br_210 wl_19 vdd gnd cell_6t
Xbit_r20_c210 bl_210 br_210 wl_20 vdd gnd cell_6t
Xbit_r21_c210 bl_210 br_210 wl_21 vdd gnd cell_6t
Xbit_r22_c210 bl_210 br_210 wl_22 vdd gnd cell_6t
Xbit_r23_c210 bl_210 br_210 wl_23 vdd gnd cell_6t
Xbit_r24_c210 bl_210 br_210 wl_24 vdd gnd cell_6t
Xbit_r25_c210 bl_210 br_210 wl_25 vdd gnd cell_6t
Xbit_r26_c210 bl_210 br_210 wl_26 vdd gnd cell_6t
Xbit_r27_c210 bl_210 br_210 wl_27 vdd gnd cell_6t
Xbit_r28_c210 bl_210 br_210 wl_28 vdd gnd cell_6t
Xbit_r29_c210 bl_210 br_210 wl_29 vdd gnd cell_6t
Xbit_r30_c210 bl_210 br_210 wl_30 vdd gnd cell_6t
Xbit_r31_c210 bl_210 br_210 wl_31 vdd gnd cell_6t
Xbit_r32_c210 bl_210 br_210 wl_32 vdd gnd cell_6t
Xbit_r33_c210 bl_210 br_210 wl_33 vdd gnd cell_6t
Xbit_r34_c210 bl_210 br_210 wl_34 vdd gnd cell_6t
Xbit_r35_c210 bl_210 br_210 wl_35 vdd gnd cell_6t
Xbit_r36_c210 bl_210 br_210 wl_36 vdd gnd cell_6t
Xbit_r37_c210 bl_210 br_210 wl_37 vdd gnd cell_6t
Xbit_r38_c210 bl_210 br_210 wl_38 vdd gnd cell_6t
Xbit_r39_c210 bl_210 br_210 wl_39 vdd gnd cell_6t
Xbit_r40_c210 bl_210 br_210 wl_40 vdd gnd cell_6t
Xbit_r41_c210 bl_210 br_210 wl_41 vdd gnd cell_6t
Xbit_r42_c210 bl_210 br_210 wl_42 vdd gnd cell_6t
Xbit_r43_c210 bl_210 br_210 wl_43 vdd gnd cell_6t
Xbit_r44_c210 bl_210 br_210 wl_44 vdd gnd cell_6t
Xbit_r45_c210 bl_210 br_210 wl_45 vdd gnd cell_6t
Xbit_r46_c210 bl_210 br_210 wl_46 vdd gnd cell_6t
Xbit_r47_c210 bl_210 br_210 wl_47 vdd gnd cell_6t
Xbit_r48_c210 bl_210 br_210 wl_48 vdd gnd cell_6t
Xbit_r49_c210 bl_210 br_210 wl_49 vdd gnd cell_6t
Xbit_r50_c210 bl_210 br_210 wl_50 vdd gnd cell_6t
Xbit_r51_c210 bl_210 br_210 wl_51 vdd gnd cell_6t
Xbit_r52_c210 bl_210 br_210 wl_52 vdd gnd cell_6t
Xbit_r53_c210 bl_210 br_210 wl_53 vdd gnd cell_6t
Xbit_r54_c210 bl_210 br_210 wl_54 vdd gnd cell_6t
Xbit_r55_c210 bl_210 br_210 wl_55 vdd gnd cell_6t
Xbit_r56_c210 bl_210 br_210 wl_56 vdd gnd cell_6t
Xbit_r57_c210 bl_210 br_210 wl_57 vdd gnd cell_6t
Xbit_r58_c210 bl_210 br_210 wl_58 vdd gnd cell_6t
Xbit_r59_c210 bl_210 br_210 wl_59 vdd gnd cell_6t
Xbit_r60_c210 bl_210 br_210 wl_60 vdd gnd cell_6t
Xbit_r61_c210 bl_210 br_210 wl_61 vdd gnd cell_6t
Xbit_r62_c210 bl_210 br_210 wl_62 vdd gnd cell_6t
Xbit_r63_c210 bl_210 br_210 wl_63 vdd gnd cell_6t
Xbit_r64_c210 bl_210 br_210 wl_64 vdd gnd cell_6t
Xbit_r65_c210 bl_210 br_210 wl_65 vdd gnd cell_6t
Xbit_r66_c210 bl_210 br_210 wl_66 vdd gnd cell_6t
Xbit_r67_c210 bl_210 br_210 wl_67 vdd gnd cell_6t
Xbit_r68_c210 bl_210 br_210 wl_68 vdd gnd cell_6t
Xbit_r69_c210 bl_210 br_210 wl_69 vdd gnd cell_6t
Xbit_r70_c210 bl_210 br_210 wl_70 vdd gnd cell_6t
Xbit_r71_c210 bl_210 br_210 wl_71 vdd gnd cell_6t
Xbit_r72_c210 bl_210 br_210 wl_72 vdd gnd cell_6t
Xbit_r73_c210 bl_210 br_210 wl_73 vdd gnd cell_6t
Xbit_r74_c210 bl_210 br_210 wl_74 vdd gnd cell_6t
Xbit_r75_c210 bl_210 br_210 wl_75 vdd gnd cell_6t
Xbit_r76_c210 bl_210 br_210 wl_76 vdd gnd cell_6t
Xbit_r77_c210 bl_210 br_210 wl_77 vdd gnd cell_6t
Xbit_r78_c210 bl_210 br_210 wl_78 vdd gnd cell_6t
Xbit_r79_c210 bl_210 br_210 wl_79 vdd gnd cell_6t
Xbit_r80_c210 bl_210 br_210 wl_80 vdd gnd cell_6t
Xbit_r81_c210 bl_210 br_210 wl_81 vdd gnd cell_6t
Xbit_r82_c210 bl_210 br_210 wl_82 vdd gnd cell_6t
Xbit_r83_c210 bl_210 br_210 wl_83 vdd gnd cell_6t
Xbit_r84_c210 bl_210 br_210 wl_84 vdd gnd cell_6t
Xbit_r85_c210 bl_210 br_210 wl_85 vdd gnd cell_6t
Xbit_r86_c210 bl_210 br_210 wl_86 vdd gnd cell_6t
Xbit_r87_c210 bl_210 br_210 wl_87 vdd gnd cell_6t
Xbit_r88_c210 bl_210 br_210 wl_88 vdd gnd cell_6t
Xbit_r89_c210 bl_210 br_210 wl_89 vdd gnd cell_6t
Xbit_r90_c210 bl_210 br_210 wl_90 vdd gnd cell_6t
Xbit_r91_c210 bl_210 br_210 wl_91 vdd gnd cell_6t
Xbit_r92_c210 bl_210 br_210 wl_92 vdd gnd cell_6t
Xbit_r93_c210 bl_210 br_210 wl_93 vdd gnd cell_6t
Xbit_r94_c210 bl_210 br_210 wl_94 vdd gnd cell_6t
Xbit_r95_c210 bl_210 br_210 wl_95 vdd gnd cell_6t
Xbit_r96_c210 bl_210 br_210 wl_96 vdd gnd cell_6t
Xbit_r97_c210 bl_210 br_210 wl_97 vdd gnd cell_6t
Xbit_r98_c210 bl_210 br_210 wl_98 vdd gnd cell_6t
Xbit_r99_c210 bl_210 br_210 wl_99 vdd gnd cell_6t
Xbit_r100_c210 bl_210 br_210 wl_100 vdd gnd cell_6t
Xbit_r101_c210 bl_210 br_210 wl_101 vdd gnd cell_6t
Xbit_r102_c210 bl_210 br_210 wl_102 vdd gnd cell_6t
Xbit_r103_c210 bl_210 br_210 wl_103 vdd gnd cell_6t
Xbit_r104_c210 bl_210 br_210 wl_104 vdd gnd cell_6t
Xbit_r105_c210 bl_210 br_210 wl_105 vdd gnd cell_6t
Xbit_r106_c210 bl_210 br_210 wl_106 vdd gnd cell_6t
Xbit_r107_c210 bl_210 br_210 wl_107 vdd gnd cell_6t
Xbit_r108_c210 bl_210 br_210 wl_108 vdd gnd cell_6t
Xbit_r109_c210 bl_210 br_210 wl_109 vdd gnd cell_6t
Xbit_r110_c210 bl_210 br_210 wl_110 vdd gnd cell_6t
Xbit_r111_c210 bl_210 br_210 wl_111 vdd gnd cell_6t
Xbit_r112_c210 bl_210 br_210 wl_112 vdd gnd cell_6t
Xbit_r113_c210 bl_210 br_210 wl_113 vdd gnd cell_6t
Xbit_r114_c210 bl_210 br_210 wl_114 vdd gnd cell_6t
Xbit_r115_c210 bl_210 br_210 wl_115 vdd gnd cell_6t
Xbit_r116_c210 bl_210 br_210 wl_116 vdd gnd cell_6t
Xbit_r117_c210 bl_210 br_210 wl_117 vdd gnd cell_6t
Xbit_r118_c210 bl_210 br_210 wl_118 vdd gnd cell_6t
Xbit_r119_c210 bl_210 br_210 wl_119 vdd gnd cell_6t
Xbit_r120_c210 bl_210 br_210 wl_120 vdd gnd cell_6t
Xbit_r121_c210 bl_210 br_210 wl_121 vdd gnd cell_6t
Xbit_r122_c210 bl_210 br_210 wl_122 vdd gnd cell_6t
Xbit_r123_c210 bl_210 br_210 wl_123 vdd gnd cell_6t
Xbit_r124_c210 bl_210 br_210 wl_124 vdd gnd cell_6t
Xbit_r125_c210 bl_210 br_210 wl_125 vdd gnd cell_6t
Xbit_r126_c210 bl_210 br_210 wl_126 vdd gnd cell_6t
Xbit_r127_c210 bl_210 br_210 wl_127 vdd gnd cell_6t
Xbit_r128_c210 bl_210 br_210 wl_128 vdd gnd cell_6t
Xbit_r129_c210 bl_210 br_210 wl_129 vdd gnd cell_6t
Xbit_r130_c210 bl_210 br_210 wl_130 vdd gnd cell_6t
Xbit_r131_c210 bl_210 br_210 wl_131 vdd gnd cell_6t
Xbit_r132_c210 bl_210 br_210 wl_132 vdd gnd cell_6t
Xbit_r133_c210 bl_210 br_210 wl_133 vdd gnd cell_6t
Xbit_r134_c210 bl_210 br_210 wl_134 vdd gnd cell_6t
Xbit_r135_c210 bl_210 br_210 wl_135 vdd gnd cell_6t
Xbit_r136_c210 bl_210 br_210 wl_136 vdd gnd cell_6t
Xbit_r137_c210 bl_210 br_210 wl_137 vdd gnd cell_6t
Xbit_r138_c210 bl_210 br_210 wl_138 vdd gnd cell_6t
Xbit_r139_c210 bl_210 br_210 wl_139 vdd gnd cell_6t
Xbit_r140_c210 bl_210 br_210 wl_140 vdd gnd cell_6t
Xbit_r141_c210 bl_210 br_210 wl_141 vdd gnd cell_6t
Xbit_r142_c210 bl_210 br_210 wl_142 vdd gnd cell_6t
Xbit_r143_c210 bl_210 br_210 wl_143 vdd gnd cell_6t
Xbit_r144_c210 bl_210 br_210 wl_144 vdd gnd cell_6t
Xbit_r145_c210 bl_210 br_210 wl_145 vdd gnd cell_6t
Xbit_r146_c210 bl_210 br_210 wl_146 vdd gnd cell_6t
Xbit_r147_c210 bl_210 br_210 wl_147 vdd gnd cell_6t
Xbit_r148_c210 bl_210 br_210 wl_148 vdd gnd cell_6t
Xbit_r149_c210 bl_210 br_210 wl_149 vdd gnd cell_6t
Xbit_r150_c210 bl_210 br_210 wl_150 vdd gnd cell_6t
Xbit_r151_c210 bl_210 br_210 wl_151 vdd gnd cell_6t
Xbit_r152_c210 bl_210 br_210 wl_152 vdd gnd cell_6t
Xbit_r153_c210 bl_210 br_210 wl_153 vdd gnd cell_6t
Xbit_r154_c210 bl_210 br_210 wl_154 vdd gnd cell_6t
Xbit_r155_c210 bl_210 br_210 wl_155 vdd gnd cell_6t
Xbit_r156_c210 bl_210 br_210 wl_156 vdd gnd cell_6t
Xbit_r157_c210 bl_210 br_210 wl_157 vdd gnd cell_6t
Xbit_r158_c210 bl_210 br_210 wl_158 vdd gnd cell_6t
Xbit_r159_c210 bl_210 br_210 wl_159 vdd gnd cell_6t
Xbit_r160_c210 bl_210 br_210 wl_160 vdd gnd cell_6t
Xbit_r161_c210 bl_210 br_210 wl_161 vdd gnd cell_6t
Xbit_r162_c210 bl_210 br_210 wl_162 vdd gnd cell_6t
Xbit_r163_c210 bl_210 br_210 wl_163 vdd gnd cell_6t
Xbit_r164_c210 bl_210 br_210 wl_164 vdd gnd cell_6t
Xbit_r165_c210 bl_210 br_210 wl_165 vdd gnd cell_6t
Xbit_r166_c210 bl_210 br_210 wl_166 vdd gnd cell_6t
Xbit_r167_c210 bl_210 br_210 wl_167 vdd gnd cell_6t
Xbit_r168_c210 bl_210 br_210 wl_168 vdd gnd cell_6t
Xbit_r169_c210 bl_210 br_210 wl_169 vdd gnd cell_6t
Xbit_r170_c210 bl_210 br_210 wl_170 vdd gnd cell_6t
Xbit_r171_c210 bl_210 br_210 wl_171 vdd gnd cell_6t
Xbit_r172_c210 bl_210 br_210 wl_172 vdd gnd cell_6t
Xbit_r173_c210 bl_210 br_210 wl_173 vdd gnd cell_6t
Xbit_r174_c210 bl_210 br_210 wl_174 vdd gnd cell_6t
Xbit_r175_c210 bl_210 br_210 wl_175 vdd gnd cell_6t
Xbit_r176_c210 bl_210 br_210 wl_176 vdd gnd cell_6t
Xbit_r177_c210 bl_210 br_210 wl_177 vdd gnd cell_6t
Xbit_r178_c210 bl_210 br_210 wl_178 vdd gnd cell_6t
Xbit_r179_c210 bl_210 br_210 wl_179 vdd gnd cell_6t
Xbit_r180_c210 bl_210 br_210 wl_180 vdd gnd cell_6t
Xbit_r181_c210 bl_210 br_210 wl_181 vdd gnd cell_6t
Xbit_r182_c210 bl_210 br_210 wl_182 vdd gnd cell_6t
Xbit_r183_c210 bl_210 br_210 wl_183 vdd gnd cell_6t
Xbit_r184_c210 bl_210 br_210 wl_184 vdd gnd cell_6t
Xbit_r185_c210 bl_210 br_210 wl_185 vdd gnd cell_6t
Xbit_r186_c210 bl_210 br_210 wl_186 vdd gnd cell_6t
Xbit_r187_c210 bl_210 br_210 wl_187 vdd gnd cell_6t
Xbit_r188_c210 bl_210 br_210 wl_188 vdd gnd cell_6t
Xbit_r189_c210 bl_210 br_210 wl_189 vdd gnd cell_6t
Xbit_r190_c210 bl_210 br_210 wl_190 vdd gnd cell_6t
Xbit_r191_c210 bl_210 br_210 wl_191 vdd gnd cell_6t
Xbit_r192_c210 bl_210 br_210 wl_192 vdd gnd cell_6t
Xbit_r193_c210 bl_210 br_210 wl_193 vdd gnd cell_6t
Xbit_r194_c210 bl_210 br_210 wl_194 vdd gnd cell_6t
Xbit_r195_c210 bl_210 br_210 wl_195 vdd gnd cell_6t
Xbit_r196_c210 bl_210 br_210 wl_196 vdd gnd cell_6t
Xbit_r197_c210 bl_210 br_210 wl_197 vdd gnd cell_6t
Xbit_r198_c210 bl_210 br_210 wl_198 vdd gnd cell_6t
Xbit_r199_c210 bl_210 br_210 wl_199 vdd gnd cell_6t
Xbit_r200_c210 bl_210 br_210 wl_200 vdd gnd cell_6t
Xbit_r201_c210 bl_210 br_210 wl_201 vdd gnd cell_6t
Xbit_r202_c210 bl_210 br_210 wl_202 vdd gnd cell_6t
Xbit_r203_c210 bl_210 br_210 wl_203 vdd gnd cell_6t
Xbit_r204_c210 bl_210 br_210 wl_204 vdd gnd cell_6t
Xbit_r205_c210 bl_210 br_210 wl_205 vdd gnd cell_6t
Xbit_r206_c210 bl_210 br_210 wl_206 vdd gnd cell_6t
Xbit_r207_c210 bl_210 br_210 wl_207 vdd gnd cell_6t
Xbit_r208_c210 bl_210 br_210 wl_208 vdd gnd cell_6t
Xbit_r209_c210 bl_210 br_210 wl_209 vdd gnd cell_6t
Xbit_r210_c210 bl_210 br_210 wl_210 vdd gnd cell_6t
Xbit_r211_c210 bl_210 br_210 wl_211 vdd gnd cell_6t
Xbit_r212_c210 bl_210 br_210 wl_212 vdd gnd cell_6t
Xbit_r213_c210 bl_210 br_210 wl_213 vdd gnd cell_6t
Xbit_r214_c210 bl_210 br_210 wl_214 vdd gnd cell_6t
Xbit_r215_c210 bl_210 br_210 wl_215 vdd gnd cell_6t
Xbit_r216_c210 bl_210 br_210 wl_216 vdd gnd cell_6t
Xbit_r217_c210 bl_210 br_210 wl_217 vdd gnd cell_6t
Xbit_r218_c210 bl_210 br_210 wl_218 vdd gnd cell_6t
Xbit_r219_c210 bl_210 br_210 wl_219 vdd gnd cell_6t
Xbit_r220_c210 bl_210 br_210 wl_220 vdd gnd cell_6t
Xbit_r221_c210 bl_210 br_210 wl_221 vdd gnd cell_6t
Xbit_r222_c210 bl_210 br_210 wl_222 vdd gnd cell_6t
Xbit_r223_c210 bl_210 br_210 wl_223 vdd gnd cell_6t
Xbit_r224_c210 bl_210 br_210 wl_224 vdd gnd cell_6t
Xbit_r225_c210 bl_210 br_210 wl_225 vdd gnd cell_6t
Xbit_r226_c210 bl_210 br_210 wl_226 vdd gnd cell_6t
Xbit_r227_c210 bl_210 br_210 wl_227 vdd gnd cell_6t
Xbit_r228_c210 bl_210 br_210 wl_228 vdd gnd cell_6t
Xbit_r229_c210 bl_210 br_210 wl_229 vdd gnd cell_6t
Xbit_r230_c210 bl_210 br_210 wl_230 vdd gnd cell_6t
Xbit_r231_c210 bl_210 br_210 wl_231 vdd gnd cell_6t
Xbit_r232_c210 bl_210 br_210 wl_232 vdd gnd cell_6t
Xbit_r233_c210 bl_210 br_210 wl_233 vdd gnd cell_6t
Xbit_r234_c210 bl_210 br_210 wl_234 vdd gnd cell_6t
Xbit_r235_c210 bl_210 br_210 wl_235 vdd gnd cell_6t
Xbit_r236_c210 bl_210 br_210 wl_236 vdd gnd cell_6t
Xbit_r237_c210 bl_210 br_210 wl_237 vdd gnd cell_6t
Xbit_r238_c210 bl_210 br_210 wl_238 vdd gnd cell_6t
Xbit_r239_c210 bl_210 br_210 wl_239 vdd gnd cell_6t
Xbit_r240_c210 bl_210 br_210 wl_240 vdd gnd cell_6t
Xbit_r241_c210 bl_210 br_210 wl_241 vdd gnd cell_6t
Xbit_r242_c210 bl_210 br_210 wl_242 vdd gnd cell_6t
Xbit_r243_c210 bl_210 br_210 wl_243 vdd gnd cell_6t
Xbit_r244_c210 bl_210 br_210 wl_244 vdd gnd cell_6t
Xbit_r245_c210 bl_210 br_210 wl_245 vdd gnd cell_6t
Xbit_r246_c210 bl_210 br_210 wl_246 vdd gnd cell_6t
Xbit_r247_c210 bl_210 br_210 wl_247 vdd gnd cell_6t
Xbit_r248_c210 bl_210 br_210 wl_248 vdd gnd cell_6t
Xbit_r249_c210 bl_210 br_210 wl_249 vdd gnd cell_6t
Xbit_r250_c210 bl_210 br_210 wl_250 vdd gnd cell_6t
Xbit_r251_c210 bl_210 br_210 wl_251 vdd gnd cell_6t
Xbit_r252_c210 bl_210 br_210 wl_252 vdd gnd cell_6t
Xbit_r253_c210 bl_210 br_210 wl_253 vdd gnd cell_6t
Xbit_r254_c210 bl_210 br_210 wl_254 vdd gnd cell_6t
Xbit_r255_c210 bl_210 br_210 wl_255 vdd gnd cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd cell_6t
Xbit_r1_c211 bl_211 br_211 wl_1 vdd gnd cell_6t
Xbit_r2_c211 bl_211 br_211 wl_2 vdd gnd cell_6t
Xbit_r3_c211 bl_211 br_211 wl_3 vdd gnd cell_6t
Xbit_r4_c211 bl_211 br_211 wl_4 vdd gnd cell_6t
Xbit_r5_c211 bl_211 br_211 wl_5 vdd gnd cell_6t
Xbit_r6_c211 bl_211 br_211 wl_6 vdd gnd cell_6t
Xbit_r7_c211 bl_211 br_211 wl_7 vdd gnd cell_6t
Xbit_r8_c211 bl_211 br_211 wl_8 vdd gnd cell_6t
Xbit_r9_c211 bl_211 br_211 wl_9 vdd gnd cell_6t
Xbit_r10_c211 bl_211 br_211 wl_10 vdd gnd cell_6t
Xbit_r11_c211 bl_211 br_211 wl_11 vdd gnd cell_6t
Xbit_r12_c211 bl_211 br_211 wl_12 vdd gnd cell_6t
Xbit_r13_c211 bl_211 br_211 wl_13 vdd gnd cell_6t
Xbit_r14_c211 bl_211 br_211 wl_14 vdd gnd cell_6t
Xbit_r15_c211 bl_211 br_211 wl_15 vdd gnd cell_6t
Xbit_r16_c211 bl_211 br_211 wl_16 vdd gnd cell_6t
Xbit_r17_c211 bl_211 br_211 wl_17 vdd gnd cell_6t
Xbit_r18_c211 bl_211 br_211 wl_18 vdd gnd cell_6t
Xbit_r19_c211 bl_211 br_211 wl_19 vdd gnd cell_6t
Xbit_r20_c211 bl_211 br_211 wl_20 vdd gnd cell_6t
Xbit_r21_c211 bl_211 br_211 wl_21 vdd gnd cell_6t
Xbit_r22_c211 bl_211 br_211 wl_22 vdd gnd cell_6t
Xbit_r23_c211 bl_211 br_211 wl_23 vdd gnd cell_6t
Xbit_r24_c211 bl_211 br_211 wl_24 vdd gnd cell_6t
Xbit_r25_c211 bl_211 br_211 wl_25 vdd gnd cell_6t
Xbit_r26_c211 bl_211 br_211 wl_26 vdd gnd cell_6t
Xbit_r27_c211 bl_211 br_211 wl_27 vdd gnd cell_6t
Xbit_r28_c211 bl_211 br_211 wl_28 vdd gnd cell_6t
Xbit_r29_c211 bl_211 br_211 wl_29 vdd gnd cell_6t
Xbit_r30_c211 bl_211 br_211 wl_30 vdd gnd cell_6t
Xbit_r31_c211 bl_211 br_211 wl_31 vdd gnd cell_6t
Xbit_r32_c211 bl_211 br_211 wl_32 vdd gnd cell_6t
Xbit_r33_c211 bl_211 br_211 wl_33 vdd gnd cell_6t
Xbit_r34_c211 bl_211 br_211 wl_34 vdd gnd cell_6t
Xbit_r35_c211 bl_211 br_211 wl_35 vdd gnd cell_6t
Xbit_r36_c211 bl_211 br_211 wl_36 vdd gnd cell_6t
Xbit_r37_c211 bl_211 br_211 wl_37 vdd gnd cell_6t
Xbit_r38_c211 bl_211 br_211 wl_38 vdd gnd cell_6t
Xbit_r39_c211 bl_211 br_211 wl_39 vdd gnd cell_6t
Xbit_r40_c211 bl_211 br_211 wl_40 vdd gnd cell_6t
Xbit_r41_c211 bl_211 br_211 wl_41 vdd gnd cell_6t
Xbit_r42_c211 bl_211 br_211 wl_42 vdd gnd cell_6t
Xbit_r43_c211 bl_211 br_211 wl_43 vdd gnd cell_6t
Xbit_r44_c211 bl_211 br_211 wl_44 vdd gnd cell_6t
Xbit_r45_c211 bl_211 br_211 wl_45 vdd gnd cell_6t
Xbit_r46_c211 bl_211 br_211 wl_46 vdd gnd cell_6t
Xbit_r47_c211 bl_211 br_211 wl_47 vdd gnd cell_6t
Xbit_r48_c211 bl_211 br_211 wl_48 vdd gnd cell_6t
Xbit_r49_c211 bl_211 br_211 wl_49 vdd gnd cell_6t
Xbit_r50_c211 bl_211 br_211 wl_50 vdd gnd cell_6t
Xbit_r51_c211 bl_211 br_211 wl_51 vdd gnd cell_6t
Xbit_r52_c211 bl_211 br_211 wl_52 vdd gnd cell_6t
Xbit_r53_c211 bl_211 br_211 wl_53 vdd gnd cell_6t
Xbit_r54_c211 bl_211 br_211 wl_54 vdd gnd cell_6t
Xbit_r55_c211 bl_211 br_211 wl_55 vdd gnd cell_6t
Xbit_r56_c211 bl_211 br_211 wl_56 vdd gnd cell_6t
Xbit_r57_c211 bl_211 br_211 wl_57 vdd gnd cell_6t
Xbit_r58_c211 bl_211 br_211 wl_58 vdd gnd cell_6t
Xbit_r59_c211 bl_211 br_211 wl_59 vdd gnd cell_6t
Xbit_r60_c211 bl_211 br_211 wl_60 vdd gnd cell_6t
Xbit_r61_c211 bl_211 br_211 wl_61 vdd gnd cell_6t
Xbit_r62_c211 bl_211 br_211 wl_62 vdd gnd cell_6t
Xbit_r63_c211 bl_211 br_211 wl_63 vdd gnd cell_6t
Xbit_r64_c211 bl_211 br_211 wl_64 vdd gnd cell_6t
Xbit_r65_c211 bl_211 br_211 wl_65 vdd gnd cell_6t
Xbit_r66_c211 bl_211 br_211 wl_66 vdd gnd cell_6t
Xbit_r67_c211 bl_211 br_211 wl_67 vdd gnd cell_6t
Xbit_r68_c211 bl_211 br_211 wl_68 vdd gnd cell_6t
Xbit_r69_c211 bl_211 br_211 wl_69 vdd gnd cell_6t
Xbit_r70_c211 bl_211 br_211 wl_70 vdd gnd cell_6t
Xbit_r71_c211 bl_211 br_211 wl_71 vdd gnd cell_6t
Xbit_r72_c211 bl_211 br_211 wl_72 vdd gnd cell_6t
Xbit_r73_c211 bl_211 br_211 wl_73 vdd gnd cell_6t
Xbit_r74_c211 bl_211 br_211 wl_74 vdd gnd cell_6t
Xbit_r75_c211 bl_211 br_211 wl_75 vdd gnd cell_6t
Xbit_r76_c211 bl_211 br_211 wl_76 vdd gnd cell_6t
Xbit_r77_c211 bl_211 br_211 wl_77 vdd gnd cell_6t
Xbit_r78_c211 bl_211 br_211 wl_78 vdd gnd cell_6t
Xbit_r79_c211 bl_211 br_211 wl_79 vdd gnd cell_6t
Xbit_r80_c211 bl_211 br_211 wl_80 vdd gnd cell_6t
Xbit_r81_c211 bl_211 br_211 wl_81 vdd gnd cell_6t
Xbit_r82_c211 bl_211 br_211 wl_82 vdd gnd cell_6t
Xbit_r83_c211 bl_211 br_211 wl_83 vdd gnd cell_6t
Xbit_r84_c211 bl_211 br_211 wl_84 vdd gnd cell_6t
Xbit_r85_c211 bl_211 br_211 wl_85 vdd gnd cell_6t
Xbit_r86_c211 bl_211 br_211 wl_86 vdd gnd cell_6t
Xbit_r87_c211 bl_211 br_211 wl_87 vdd gnd cell_6t
Xbit_r88_c211 bl_211 br_211 wl_88 vdd gnd cell_6t
Xbit_r89_c211 bl_211 br_211 wl_89 vdd gnd cell_6t
Xbit_r90_c211 bl_211 br_211 wl_90 vdd gnd cell_6t
Xbit_r91_c211 bl_211 br_211 wl_91 vdd gnd cell_6t
Xbit_r92_c211 bl_211 br_211 wl_92 vdd gnd cell_6t
Xbit_r93_c211 bl_211 br_211 wl_93 vdd gnd cell_6t
Xbit_r94_c211 bl_211 br_211 wl_94 vdd gnd cell_6t
Xbit_r95_c211 bl_211 br_211 wl_95 vdd gnd cell_6t
Xbit_r96_c211 bl_211 br_211 wl_96 vdd gnd cell_6t
Xbit_r97_c211 bl_211 br_211 wl_97 vdd gnd cell_6t
Xbit_r98_c211 bl_211 br_211 wl_98 vdd gnd cell_6t
Xbit_r99_c211 bl_211 br_211 wl_99 vdd gnd cell_6t
Xbit_r100_c211 bl_211 br_211 wl_100 vdd gnd cell_6t
Xbit_r101_c211 bl_211 br_211 wl_101 vdd gnd cell_6t
Xbit_r102_c211 bl_211 br_211 wl_102 vdd gnd cell_6t
Xbit_r103_c211 bl_211 br_211 wl_103 vdd gnd cell_6t
Xbit_r104_c211 bl_211 br_211 wl_104 vdd gnd cell_6t
Xbit_r105_c211 bl_211 br_211 wl_105 vdd gnd cell_6t
Xbit_r106_c211 bl_211 br_211 wl_106 vdd gnd cell_6t
Xbit_r107_c211 bl_211 br_211 wl_107 vdd gnd cell_6t
Xbit_r108_c211 bl_211 br_211 wl_108 vdd gnd cell_6t
Xbit_r109_c211 bl_211 br_211 wl_109 vdd gnd cell_6t
Xbit_r110_c211 bl_211 br_211 wl_110 vdd gnd cell_6t
Xbit_r111_c211 bl_211 br_211 wl_111 vdd gnd cell_6t
Xbit_r112_c211 bl_211 br_211 wl_112 vdd gnd cell_6t
Xbit_r113_c211 bl_211 br_211 wl_113 vdd gnd cell_6t
Xbit_r114_c211 bl_211 br_211 wl_114 vdd gnd cell_6t
Xbit_r115_c211 bl_211 br_211 wl_115 vdd gnd cell_6t
Xbit_r116_c211 bl_211 br_211 wl_116 vdd gnd cell_6t
Xbit_r117_c211 bl_211 br_211 wl_117 vdd gnd cell_6t
Xbit_r118_c211 bl_211 br_211 wl_118 vdd gnd cell_6t
Xbit_r119_c211 bl_211 br_211 wl_119 vdd gnd cell_6t
Xbit_r120_c211 bl_211 br_211 wl_120 vdd gnd cell_6t
Xbit_r121_c211 bl_211 br_211 wl_121 vdd gnd cell_6t
Xbit_r122_c211 bl_211 br_211 wl_122 vdd gnd cell_6t
Xbit_r123_c211 bl_211 br_211 wl_123 vdd gnd cell_6t
Xbit_r124_c211 bl_211 br_211 wl_124 vdd gnd cell_6t
Xbit_r125_c211 bl_211 br_211 wl_125 vdd gnd cell_6t
Xbit_r126_c211 bl_211 br_211 wl_126 vdd gnd cell_6t
Xbit_r127_c211 bl_211 br_211 wl_127 vdd gnd cell_6t
Xbit_r128_c211 bl_211 br_211 wl_128 vdd gnd cell_6t
Xbit_r129_c211 bl_211 br_211 wl_129 vdd gnd cell_6t
Xbit_r130_c211 bl_211 br_211 wl_130 vdd gnd cell_6t
Xbit_r131_c211 bl_211 br_211 wl_131 vdd gnd cell_6t
Xbit_r132_c211 bl_211 br_211 wl_132 vdd gnd cell_6t
Xbit_r133_c211 bl_211 br_211 wl_133 vdd gnd cell_6t
Xbit_r134_c211 bl_211 br_211 wl_134 vdd gnd cell_6t
Xbit_r135_c211 bl_211 br_211 wl_135 vdd gnd cell_6t
Xbit_r136_c211 bl_211 br_211 wl_136 vdd gnd cell_6t
Xbit_r137_c211 bl_211 br_211 wl_137 vdd gnd cell_6t
Xbit_r138_c211 bl_211 br_211 wl_138 vdd gnd cell_6t
Xbit_r139_c211 bl_211 br_211 wl_139 vdd gnd cell_6t
Xbit_r140_c211 bl_211 br_211 wl_140 vdd gnd cell_6t
Xbit_r141_c211 bl_211 br_211 wl_141 vdd gnd cell_6t
Xbit_r142_c211 bl_211 br_211 wl_142 vdd gnd cell_6t
Xbit_r143_c211 bl_211 br_211 wl_143 vdd gnd cell_6t
Xbit_r144_c211 bl_211 br_211 wl_144 vdd gnd cell_6t
Xbit_r145_c211 bl_211 br_211 wl_145 vdd gnd cell_6t
Xbit_r146_c211 bl_211 br_211 wl_146 vdd gnd cell_6t
Xbit_r147_c211 bl_211 br_211 wl_147 vdd gnd cell_6t
Xbit_r148_c211 bl_211 br_211 wl_148 vdd gnd cell_6t
Xbit_r149_c211 bl_211 br_211 wl_149 vdd gnd cell_6t
Xbit_r150_c211 bl_211 br_211 wl_150 vdd gnd cell_6t
Xbit_r151_c211 bl_211 br_211 wl_151 vdd gnd cell_6t
Xbit_r152_c211 bl_211 br_211 wl_152 vdd gnd cell_6t
Xbit_r153_c211 bl_211 br_211 wl_153 vdd gnd cell_6t
Xbit_r154_c211 bl_211 br_211 wl_154 vdd gnd cell_6t
Xbit_r155_c211 bl_211 br_211 wl_155 vdd gnd cell_6t
Xbit_r156_c211 bl_211 br_211 wl_156 vdd gnd cell_6t
Xbit_r157_c211 bl_211 br_211 wl_157 vdd gnd cell_6t
Xbit_r158_c211 bl_211 br_211 wl_158 vdd gnd cell_6t
Xbit_r159_c211 bl_211 br_211 wl_159 vdd gnd cell_6t
Xbit_r160_c211 bl_211 br_211 wl_160 vdd gnd cell_6t
Xbit_r161_c211 bl_211 br_211 wl_161 vdd gnd cell_6t
Xbit_r162_c211 bl_211 br_211 wl_162 vdd gnd cell_6t
Xbit_r163_c211 bl_211 br_211 wl_163 vdd gnd cell_6t
Xbit_r164_c211 bl_211 br_211 wl_164 vdd gnd cell_6t
Xbit_r165_c211 bl_211 br_211 wl_165 vdd gnd cell_6t
Xbit_r166_c211 bl_211 br_211 wl_166 vdd gnd cell_6t
Xbit_r167_c211 bl_211 br_211 wl_167 vdd gnd cell_6t
Xbit_r168_c211 bl_211 br_211 wl_168 vdd gnd cell_6t
Xbit_r169_c211 bl_211 br_211 wl_169 vdd gnd cell_6t
Xbit_r170_c211 bl_211 br_211 wl_170 vdd gnd cell_6t
Xbit_r171_c211 bl_211 br_211 wl_171 vdd gnd cell_6t
Xbit_r172_c211 bl_211 br_211 wl_172 vdd gnd cell_6t
Xbit_r173_c211 bl_211 br_211 wl_173 vdd gnd cell_6t
Xbit_r174_c211 bl_211 br_211 wl_174 vdd gnd cell_6t
Xbit_r175_c211 bl_211 br_211 wl_175 vdd gnd cell_6t
Xbit_r176_c211 bl_211 br_211 wl_176 vdd gnd cell_6t
Xbit_r177_c211 bl_211 br_211 wl_177 vdd gnd cell_6t
Xbit_r178_c211 bl_211 br_211 wl_178 vdd gnd cell_6t
Xbit_r179_c211 bl_211 br_211 wl_179 vdd gnd cell_6t
Xbit_r180_c211 bl_211 br_211 wl_180 vdd gnd cell_6t
Xbit_r181_c211 bl_211 br_211 wl_181 vdd gnd cell_6t
Xbit_r182_c211 bl_211 br_211 wl_182 vdd gnd cell_6t
Xbit_r183_c211 bl_211 br_211 wl_183 vdd gnd cell_6t
Xbit_r184_c211 bl_211 br_211 wl_184 vdd gnd cell_6t
Xbit_r185_c211 bl_211 br_211 wl_185 vdd gnd cell_6t
Xbit_r186_c211 bl_211 br_211 wl_186 vdd gnd cell_6t
Xbit_r187_c211 bl_211 br_211 wl_187 vdd gnd cell_6t
Xbit_r188_c211 bl_211 br_211 wl_188 vdd gnd cell_6t
Xbit_r189_c211 bl_211 br_211 wl_189 vdd gnd cell_6t
Xbit_r190_c211 bl_211 br_211 wl_190 vdd gnd cell_6t
Xbit_r191_c211 bl_211 br_211 wl_191 vdd gnd cell_6t
Xbit_r192_c211 bl_211 br_211 wl_192 vdd gnd cell_6t
Xbit_r193_c211 bl_211 br_211 wl_193 vdd gnd cell_6t
Xbit_r194_c211 bl_211 br_211 wl_194 vdd gnd cell_6t
Xbit_r195_c211 bl_211 br_211 wl_195 vdd gnd cell_6t
Xbit_r196_c211 bl_211 br_211 wl_196 vdd gnd cell_6t
Xbit_r197_c211 bl_211 br_211 wl_197 vdd gnd cell_6t
Xbit_r198_c211 bl_211 br_211 wl_198 vdd gnd cell_6t
Xbit_r199_c211 bl_211 br_211 wl_199 vdd gnd cell_6t
Xbit_r200_c211 bl_211 br_211 wl_200 vdd gnd cell_6t
Xbit_r201_c211 bl_211 br_211 wl_201 vdd gnd cell_6t
Xbit_r202_c211 bl_211 br_211 wl_202 vdd gnd cell_6t
Xbit_r203_c211 bl_211 br_211 wl_203 vdd gnd cell_6t
Xbit_r204_c211 bl_211 br_211 wl_204 vdd gnd cell_6t
Xbit_r205_c211 bl_211 br_211 wl_205 vdd gnd cell_6t
Xbit_r206_c211 bl_211 br_211 wl_206 vdd gnd cell_6t
Xbit_r207_c211 bl_211 br_211 wl_207 vdd gnd cell_6t
Xbit_r208_c211 bl_211 br_211 wl_208 vdd gnd cell_6t
Xbit_r209_c211 bl_211 br_211 wl_209 vdd gnd cell_6t
Xbit_r210_c211 bl_211 br_211 wl_210 vdd gnd cell_6t
Xbit_r211_c211 bl_211 br_211 wl_211 vdd gnd cell_6t
Xbit_r212_c211 bl_211 br_211 wl_212 vdd gnd cell_6t
Xbit_r213_c211 bl_211 br_211 wl_213 vdd gnd cell_6t
Xbit_r214_c211 bl_211 br_211 wl_214 vdd gnd cell_6t
Xbit_r215_c211 bl_211 br_211 wl_215 vdd gnd cell_6t
Xbit_r216_c211 bl_211 br_211 wl_216 vdd gnd cell_6t
Xbit_r217_c211 bl_211 br_211 wl_217 vdd gnd cell_6t
Xbit_r218_c211 bl_211 br_211 wl_218 vdd gnd cell_6t
Xbit_r219_c211 bl_211 br_211 wl_219 vdd gnd cell_6t
Xbit_r220_c211 bl_211 br_211 wl_220 vdd gnd cell_6t
Xbit_r221_c211 bl_211 br_211 wl_221 vdd gnd cell_6t
Xbit_r222_c211 bl_211 br_211 wl_222 vdd gnd cell_6t
Xbit_r223_c211 bl_211 br_211 wl_223 vdd gnd cell_6t
Xbit_r224_c211 bl_211 br_211 wl_224 vdd gnd cell_6t
Xbit_r225_c211 bl_211 br_211 wl_225 vdd gnd cell_6t
Xbit_r226_c211 bl_211 br_211 wl_226 vdd gnd cell_6t
Xbit_r227_c211 bl_211 br_211 wl_227 vdd gnd cell_6t
Xbit_r228_c211 bl_211 br_211 wl_228 vdd gnd cell_6t
Xbit_r229_c211 bl_211 br_211 wl_229 vdd gnd cell_6t
Xbit_r230_c211 bl_211 br_211 wl_230 vdd gnd cell_6t
Xbit_r231_c211 bl_211 br_211 wl_231 vdd gnd cell_6t
Xbit_r232_c211 bl_211 br_211 wl_232 vdd gnd cell_6t
Xbit_r233_c211 bl_211 br_211 wl_233 vdd gnd cell_6t
Xbit_r234_c211 bl_211 br_211 wl_234 vdd gnd cell_6t
Xbit_r235_c211 bl_211 br_211 wl_235 vdd gnd cell_6t
Xbit_r236_c211 bl_211 br_211 wl_236 vdd gnd cell_6t
Xbit_r237_c211 bl_211 br_211 wl_237 vdd gnd cell_6t
Xbit_r238_c211 bl_211 br_211 wl_238 vdd gnd cell_6t
Xbit_r239_c211 bl_211 br_211 wl_239 vdd gnd cell_6t
Xbit_r240_c211 bl_211 br_211 wl_240 vdd gnd cell_6t
Xbit_r241_c211 bl_211 br_211 wl_241 vdd gnd cell_6t
Xbit_r242_c211 bl_211 br_211 wl_242 vdd gnd cell_6t
Xbit_r243_c211 bl_211 br_211 wl_243 vdd gnd cell_6t
Xbit_r244_c211 bl_211 br_211 wl_244 vdd gnd cell_6t
Xbit_r245_c211 bl_211 br_211 wl_245 vdd gnd cell_6t
Xbit_r246_c211 bl_211 br_211 wl_246 vdd gnd cell_6t
Xbit_r247_c211 bl_211 br_211 wl_247 vdd gnd cell_6t
Xbit_r248_c211 bl_211 br_211 wl_248 vdd gnd cell_6t
Xbit_r249_c211 bl_211 br_211 wl_249 vdd gnd cell_6t
Xbit_r250_c211 bl_211 br_211 wl_250 vdd gnd cell_6t
Xbit_r251_c211 bl_211 br_211 wl_251 vdd gnd cell_6t
Xbit_r252_c211 bl_211 br_211 wl_252 vdd gnd cell_6t
Xbit_r253_c211 bl_211 br_211 wl_253 vdd gnd cell_6t
Xbit_r254_c211 bl_211 br_211 wl_254 vdd gnd cell_6t
Xbit_r255_c211 bl_211 br_211 wl_255 vdd gnd cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd cell_6t
Xbit_r1_c212 bl_212 br_212 wl_1 vdd gnd cell_6t
Xbit_r2_c212 bl_212 br_212 wl_2 vdd gnd cell_6t
Xbit_r3_c212 bl_212 br_212 wl_3 vdd gnd cell_6t
Xbit_r4_c212 bl_212 br_212 wl_4 vdd gnd cell_6t
Xbit_r5_c212 bl_212 br_212 wl_5 vdd gnd cell_6t
Xbit_r6_c212 bl_212 br_212 wl_6 vdd gnd cell_6t
Xbit_r7_c212 bl_212 br_212 wl_7 vdd gnd cell_6t
Xbit_r8_c212 bl_212 br_212 wl_8 vdd gnd cell_6t
Xbit_r9_c212 bl_212 br_212 wl_9 vdd gnd cell_6t
Xbit_r10_c212 bl_212 br_212 wl_10 vdd gnd cell_6t
Xbit_r11_c212 bl_212 br_212 wl_11 vdd gnd cell_6t
Xbit_r12_c212 bl_212 br_212 wl_12 vdd gnd cell_6t
Xbit_r13_c212 bl_212 br_212 wl_13 vdd gnd cell_6t
Xbit_r14_c212 bl_212 br_212 wl_14 vdd gnd cell_6t
Xbit_r15_c212 bl_212 br_212 wl_15 vdd gnd cell_6t
Xbit_r16_c212 bl_212 br_212 wl_16 vdd gnd cell_6t
Xbit_r17_c212 bl_212 br_212 wl_17 vdd gnd cell_6t
Xbit_r18_c212 bl_212 br_212 wl_18 vdd gnd cell_6t
Xbit_r19_c212 bl_212 br_212 wl_19 vdd gnd cell_6t
Xbit_r20_c212 bl_212 br_212 wl_20 vdd gnd cell_6t
Xbit_r21_c212 bl_212 br_212 wl_21 vdd gnd cell_6t
Xbit_r22_c212 bl_212 br_212 wl_22 vdd gnd cell_6t
Xbit_r23_c212 bl_212 br_212 wl_23 vdd gnd cell_6t
Xbit_r24_c212 bl_212 br_212 wl_24 vdd gnd cell_6t
Xbit_r25_c212 bl_212 br_212 wl_25 vdd gnd cell_6t
Xbit_r26_c212 bl_212 br_212 wl_26 vdd gnd cell_6t
Xbit_r27_c212 bl_212 br_212 wl_27 vdd gnd cell_6t
Xbit_r28_c212 bl_212 br_212 wl_28 vdd gnd cell_6t
Xbit_r29_c212 bl_212 br_212 wl_29 vdd gnd cell_6t
Xbit_r30_c212 bl_212 br_212 wl_30 vdd gnd cell_6t
Xbit_r31_c212 bl_212 br_212 wl_31 vdd gnd cell_6t
Xbit_r32_c212 bl_212 br_212 wl_32 vdd gnd cell_6t
Xbit_r33_c212 bl_212 br_212 wl_33 vdd gnd cell_6t
Xbit_r34_c212 bl_212 br_212 wl_34 vdd gnd cell_6t
Xbit_r35_c212 bl_212 br_212 wl_35 vdd gnd cell_6t
Xbit_r36_c212 bl_212 br_212 wl_36 vdd gnd cell_6t
Xbit_r37_c212 bl_212 br_212 wl_37 vdd gnd cell_6t
Xbit_r38_c212 bl_212 br_212 wl_38 vdd gnd cell_6t
Xbit_r39_c212 bl_212 br_212 wl_39 vdd gnd cell_6t
Xbit_r40_c212 bl_212 br_212 wl_40 vdd gnd cell_6t
Xbit_r41_c212 bl_212 br_212 wl_41 vdd gnd cell_6t
Xbit_r42_c212 bl_212 br_212 wl_42 vdd gnd cell_6t
Xbit_r43_c212 bl_212 br_212 wl_43 vdd gnd cell_6t
Xbit_r44_c212 bl_212 br_212 wl_44 vdd gnd cell_6t
Xbit_r45_c212 bl_212 br_212 wl_45 vdd gnd cell_6t
Xbit_r46_c212 bl_212 br_212 wl_46 vdd gnd cell_6t
Xbit_r47_c212 bl_212 br_212 wl_47 vdd gnd cell_6t
Xbit_r48_c212 bl_212 br_212 wl_48 vdd gnd cell_6t
Xbit_r49_c212 bl_212 br_212 wl_49 vdd gnd cell_6t
Xbit_r50_c212 bl_212 br_212 wl_50 vdd gnd cell_6t
Xbit_r51_c212 bl_212 br_212 wl_51 vdd gnd cell_6t
Xbit_r52_c212 bl_212 br_212 wl_52 vdd gnd cell_6t
Xbit_r53_c212 bl_212 br_212 wl_53 vdd gnd cell_6t
Xbit_r54_c212 bl_212 br_212 wl_54 vdd gnd cell_6t
Xbit_r55_c212 bl_212 br_212 wl_55 vdd gnd cell_6t
Xbit_r56_c212 bl_212 br_212 wl_56 vdd gnd cell_6t
Xbit_r57_c212 bl_212 br_212 wl_57 vdd gnd cell_6t
Xbit_r58_c212 bl_212 br_212 wl_58 vdd gnd cell_6t
Xbit_r59_c212 bl_212 br_212 wl_59 vdd gnd cell_6t
Xbit_r60_c212 bl_212 br_212 wl_60 vdd gnd cell_6t
Xbit_r61_c212 bl_212 br_212 wl_61 vdd gnd cell_6t
Xbit_r62_c212 bl_212 br_212 wl_62 vdd gnd cell_6t
Xbit_r63_c212 bl_212 br_212 wl_63 vdd gnd cell_6t
Xbit_r64_c212 bl_212 br_212 wl_64 vdd gnd cell_6t
Xbit_r65_c212 bl_212 br_212 wl_65 vdd gnd cell_6t
Xbit_r66_c212 bl_212 br_212 wl_66 vdd gnd cell_6t
Xbit_r67_c212 bl_212 br_212 wl_67 vdd gnd cell_6t
Xbit_r68_c212 bl_212 br_212 wl_68 vdd gnd cell_6t
Xbit_r69_c212 bl_212 br_212 wl_69 vdd gnd cell_6t
Xbit_r70_c212 bl_212 br_212 wl_70 vdd gnd cell_6t
Xbit_r71_c212 bl_212 br_212 wl_71 vdd gnd cell_6t
Xbit_r72_c212 bl_212 br_212 wl_72 vdd gnd cell_6t
Xbit_r73_c212 bl_212 br_212 wl_73 vdd gnd cell_6t
Xbit_r74_c212 bl_212 br_212 wl_74 vdd gnd cell_6t
Xbit_r75_c212 bl_212 br_212 wl_75 vdd gnd cell_6t
Xbit_r76_c212 bl_212 br_212 wl_76 vdd gnd cell_6t
Xbit_r77_c212 bl_212 br_212 wl_77 vdd gnd cell_6t
Xbit_r78_c212 bl_212 br_212 wl_78 vdd gnd cell_6t
Xbit_r79_c212 bl_212 br_212 wl_79 vdd gnd cell_6t
Xbit_r80_c212 bl_212 br_212 wl_80 vdd gnd cell_6t
Xbit_r81_c212 bl_212 br_212 wl_81 vdd gnd cell_6t
Xbit_r82_c212 bl_212 br_212 wl_82 vdd gnd cell_6t
Xbit_r83_c212 bl_212 br_212 wl_83 vdd gnd cell_6t
Xbit_r84_c212 bl_212 br_212 wl_84 vdd gnd cell_6t
Xbit_r85_c212 bl_212 br_212 wl_85 vdd gnd cell_6t
Xbit_r86_c212 bl_212 br_212 wl_86 vdd gnd cell_6t
Xbit_r87_c212 bl_212 br_212 wl_87 vdd gnd cell_6t
Xbit_r88_c212 bl_212 br_212 wl_88 vdd gnd cell_6t
Xbit_r89_c212 bl_212 br_212 wl_89 vdd gnd cell_6t
Xbit_r90_c212 bl_212 br_212 wl_90 vdd gnd cell_6t
Xbit_r91_c212 bl_212 br_212 wl_91 vdd gnd cell_6t
Xbit_r92_c212 bl_212 br_212 wl_92 vdd gnd cell_6t
Xbit_r93_c212 bl_212 br_212 wl_93 vdd gnd cell_6t
Xbit_r94_c212 bl_212 br_212 wl_94 vdd gnd cell_6t
Xbit_r95_c212 bl_212 br_212 wl_95 vdd gnd cell_6t
Xbit_r96_c212 bl_212 br_212 wl_96 vdd gnd cell_6t
Xbit_r97_c212 bl_212 br_212 wl_97 vdd gnd cell_6t
Xbit_r98_c212 bl_212 br_212 wl_98 vdd gnd cell_6t
Xbit_r99_c212 bl_212 br_212 wl_99 vdd gnd cell_6t
Xbit_r100_c212 bl_212 br_212 wl_100 vdd gnd cell_6t
Xbit_r101_c212 bl_212 br_212 wl_101 vdd gnd cell_6t
Xbit_r102_c212 bl_212 br_212 wl_102 vdd gnd cell_6t
Xbit_r103_c212 bl_212 br_212 wl_103 vdd gnd cell_6t
Xbit_r104_c212 bl_212 br_212 wl_104 vdd gnd cell_6t
Xbit_r105_c212 bl_212 br_212 wl_105 vdd gnd cell_6t
Xbit_r106_c212 bl_212 br_212 wl_106 vdd gnd cell_6t
Xbit_r107_c212 bl_212 br_212 wl_107 vdd gnd cell_6t
Xbit_r108_c212 bl_212 br_212 wl_108 vdd gnd cell_6t
Xbit_r109_c212 bl_212 br_212 wl_109 vdd gnd cell_6t
Xbit_r110_c212 bl_212 br_212 wl_110 vdd gnd cell_6t
Xbit_r111_c212 bl_212 br_212 wl_111 vdd gnd cell_6t
Xbit_r112_c212 bl_212 br_212 wl_112 vdd gnd cell_6t
Xbit_r113_c212 bl_212 br_212 wl_113 vdd gnd cell_6t
Xbit_r114_c212 bl_212 br_212 wl_114 vdd gnd cell_6t
Xbit_r115_c212 bl_212 br_212 wl_115 vdd gnd cell_6t
Xbit_r116_c212 bl_212 br_212 wl_116 vdd gnd cell_6t
Xbit_r117_c212 bl_212 br_212 wl_117 vdd gnd cell_6t
Xbit_r118_c212 bl_212 br_212 wl_118 vdd gnd cell_6t
Xbit_r119_c212 bl_212 br_212 wl_119 vdd gnd cell_6t
Xbit_r120_c212 bl_212 br_212 wl_120 vdd gnd cell_6t
Xbit_r121_c212 bl_212 br_212 wl_121 vdd gnd cell_6t
Xbit_r122_c212 bl_212 br_212 wl_122 vdd gnd cell_6t
Xbit_r123_c212 bl_212 br_212 wl_123 vdd gnd cell_6t
Xbit_r124_c212 bl_212 br_212 wl_124 vdd gnd cell_6t
Xbit_r125_c212 bl_212 br_212 wl_125 vdd gnd cell_6t
Xbit_r126_c212 bl_212 br_212 wl_126 vdd gnd cell_6t
Xbit_r127_c212 bl_212 br_212 wl_127 vdd gnd cell_6t
Xbit_r128_c212 bl_212 br_212 wl_128 vdd gnd cell_6t
Xbit_r129_c212 bl_212 br_212 wl_129 vdd gnd cell_6t
Xbit_r130_c212 bl_212 br_212 wl_130 vdd gnd cell_6t
Xbit_r131_c212 bl_212 br_212 wl_131 vdd gnd cell_6t
Xbit_r132_c212 bl_212 br_212 wl_132 vdd gnd cell_6t
Xbit_r133_c212 bl_212 br_212 wl_133 vdd gnd cell_6t
Xbit_r134_c212 bl_212 br_212 wl_134 vdd gnd cell_6t
Xbit_r135_c212 bl_212 br_212 wl_135 vdd gnd cell_6t
Xbit_r136_c212 bl_212 br_212 wl_136 vdd gnd cell_6t
Xbit_r137_c212 bl_212 br_212 wl_137 vdd gnd cell_6t
Xbit_r138_c212 bl_212 br_212 wl_138 vdd gnd cell_6t
Xbit_r139_c212 bl_212 br_212 wl_139 vdd gnd cell_6t
Xbit_r140_c212 bl_212 br_212 wl_140 vdd gnd cell_6t
Xbit_r141_c212 bl_212 br_212 wl_141 vdd gnd cell_6t
Xbit_r142_c212 bl_212 br_212 wl_142 vdd gnd cell_6t
Xbit_r143_c212 bl_212 br_212 wl_143 vdd gnd cell_6t
Xbit_r144_c212 bl_212 br_212 wl_144 vdd gnd cell_6t
Xbit_r145_c212 bl_212 br_212 wl_145 vdd gnd cell_6t
Xbit_r146_c212 bl_212 br_212 wl_146 vdd gnd cell_6t
Xbit_r147_c212 bl_212 br_212 wl_147 vdd gnd cell_6t
Xbit_r148_c212 bl_212 br_212 wl_148 vdd gnd cell_6t
Xbit_r149_c212 bl_212 br_212 wl_149 vdd gnd cell_6t
Xbit_r150_c212 bl_212 br_212 wl_150 vdd gnd cell_6t
Xbit_r151_c212 bl_212 br_212 wl_151 vdd gnd cell_6t
Xbit_r152_c212 bl_212 br_212 wl_152 vdd gnd cell_6t
Xbit_r153_c212 bl_212 br_212 wl_153 vdd gnd cell_6t
Xbit_r154_c212 bl_212 br_212 wl_154 vdd gnd cell_6t
Xbit_r155_c212 bl_212 br_212 wl_155 vdd gnd cell_6t
Xbit_r156_c212 bl_212 br_212 wl_156 vdd gnd cell_6t
Xbit_r157_c212 bl_212 br_212 wl_157 vdd gnd cell_6t
Xbit_r158_c212 bl_212 br_212 wl_158 vdd gnd cell_6t
Xbit_r159_c212 bl_212 br_212 wl_159 vdd gnd cell_6t
Xbit_r160_c212 bl_212 br_212 wl_160 vdd gnd cell_6t
Xbit_r161_c212 bl_212 br_212 wl_161 vdd gnd cell_6t
Xbit_r162_c212 bl_212 br_212 wl_162 vdd gnd cell_6t
Xbit_r163_c212 bl_212 br_212 wl_163 vdd gnd cell_6t
Xbit_r164_c212 bl_212 br_212 wl_164 vdd gnd cell_6t
Xbit_r165_c212 bl_212 br_212 wl_165 vdd gnd cell_6t
Xbit_r166_c212 bl_212 br_212 wl_166 vdd gnd cell_6t
Xbit_r167_c212 bl_212 br_212 wl_167 vdd gnd cell_6t
Xbit_r168_c212 bl_212 br_212 wl_168 vdd gnd cell_6t
Xbit_r169_c212 bl_212 br_212 wl_169 vdd gnd cell_6t
Xbit_r170_c212 bl_212 br_212 wl_170 vdd gnd cell_6t
Xbit_r171_c212 bl_212 br_212 wl_171 vdd gnd cell_6t
Xbit_r172_c212 bl_212 br_212 wl_172 vdd gnd cell_6t
Xbit_r173_c212 bl_212 br_212 wl_173 vdd gnd cell_6t
Xbit_r174_c212 bl_212 br_212 wl_174 vdd gnd cell_6t
Xbit_r175_c212 bl_212 br_212 wl_175 vdd gnd cell_6t
Xbit_r176_c212 bl_212 br_212 wl_176 vdd gnd cell_6t
Xbit_r177_c212 bl_212 br_212 wl_177 vdd gnd cell_6t
Xbit_r178_c212 bl_212 br_212 wl_178 vdd gnd cell_6t
Xbit_r179_c212 bl_212 br_212 wl_179 vdd gnd cell_6t
Xbit_r180_c212 bl_212 br_212 wl_180 vdd gnd cell_6t
Xbit_r181_c212 bl_212 br_212 wl_181 vdd gnd cell_6t
Xbit_r182_c212 bl_212 br_212 wl_182 vdd gnd cell_6t
Xbit_r183_c212 bl_212 br_212 wl_183 vdd gnd cell_6t
Xbit_r184_c212 bl_212 br_212 wl_184 vdd gnd cell_6t
Xbit_r185_c212 bl_212 br_212 wl_185 vdd gnd cell_6t
Xbit_r186_c212 bl_212 br_212 wl_186 vdd gnd cell_6t
Xbit_r187_c212 bl_212 br_212 wl_187 vdd gnd cell_6t
Xbit_r188_c212 bl_212 br_212 wl_188 vdd gnd cell_6t
Xbit_r189_c212 bl_212 br_212 wl_189 vdd gnd cell_6t
Xbit_r190_c212 bl_212 br_212 wl_190 vdd gnd cell_6t
Xbit_r191_c212 bl_212 br_212 wl_191 vdd gnd cell_6t
Xbit_r192_c212 bl_212 br_212 wl_192 vdd gnd cell_6t
Xbit_r193_c212 bl_212 br_212 wl_193 vdd gnd cell_6t
Xbit_r194_c212 bl_212 br_212 wl_194 vdd gnd cell_6t
Xbit_r195_c212 bl_212 br_212 wl_195 vdd gnd cell_6t
Xbit_r196_c212 bl_212 br_212 wl_196 vdd gnd cell_6t
Xbit_r197_c212 bl_212 br_212 wl_197 vdd gnd cell_6t
Xbit_r198_c212 bl_212 br_212 wl_198 vdd gnd cell_6t
Xbit_r199_c212 bl_212 br_212 wl_199 vdd gnd cell_6t
Xbit_r200_c212 bl_212 br_212 wl_200 vdd gnd cell_6t
Xbit_r201_c212 bl_212 br_212 wl_201 vdd gnd cell_6t
Xbit_r202_c212 bl_212 br_212 wl_202 vdd gnd cell_6t
Xbit_r203_c212 bl_212 br_212 wl_203 vdd gnd cell_6t
Xbit_r204_c212 bl_212 br_212 wl_204 vdd gnd cell_6t
Xbit_r205_c212 bl_212 br_212 wl_205 vdd gnd cell_6t
Xbit_r206_c212 bl_212 br_212 wl_206 vdd gnd cell_6t
Xbit_r207_c212 bl_212 br_212 wl_207 vdd gnd cell_6t
Xbit_r208_c212 bl_212 br_212 wl_208 vdd gnd cell_6t
Xbit_r209_c212 bl_212 br_212 wl_209 vdd gnd cell_6t
Xbit_r210_c212 bl_212 br_212 wl_210 vdd gnd cell_6t
Xbit_r211_c212 bl_212 br_212 wl_211 vdd gnd cell_6t
Xbit_r212_c212 bl_212 br_212 wl_212 vdd gnd cell_6t
Xbit_r213_c212 bl_212 br_212 wl_213 vdd gnd cell_6t
Xbit_r214_c212 bl_212 br_212 wl_214 vdd gnd cell_6t
Xbit_r215_c212 bl_212 br_212 wl_215 vdd gnd cell_6t
Xbit_r216_c212 bl_212 br_212 wl_216 vdd gnd cell_6t
Xbit_r217_c212 bl_212 br_212 wl_217 vdd gnd cell_6t
Xbit_r218_c212 bl_212 br_212 wl_218 vdd gnd cell_6t
Xbit_r219_c212 bl_212 br_212 wl_219 vdd gnd cell_6t
Xbit_r220_c212 bl_212 br_212 wl_220 vdd gnd cell_6t
Xbit_r221_c212 bl_212 br_212 wl_221 vdd gnd cell_6t
Xbit_r222_c212 bl_212 br_212 wl_222 vdd gnd cell_6t
Xbit_r223_c212 bl_212 br_212 wl_223 vdd gnd cell_6t
Xbit_r224_c212 bl_212 br_212 wl_224 vdd gnd cell_6t
Xbit_r225_c212 bl_212 br_212 wl_225 vdd gnd cell_6t
Xbit_r226_c212 bl_212 br_212 wl_226 vdd gnd cell_6t
Xbit_r227_c212 bl_212 br_212 wl_227 vdd gnd cell_6t
Xbit_r228_c212 bl_212 br_212 wl_228 vdd gnd cell_6t
Xbit_r229_c212 bl_212 br_212 wl_229 vdd gnd cell_6t
Xbit_r230_c212 bl_212 br_212 wl_230 vdd gnd cell_6t
Xbit_r231_c212 bl_212 br_212 wl_231 vdd gnd cell_6t
Xbit_r232_c212 bl_212 br_212 wl_232 vdd gnd cell_6t
Xbit_r233_c212 bl_212 br_212 wl_233 vdd gnd cell_6t
Xbit_r234_c212 bl_212 br_212 wl_234 vdd gnd cell_6t
Xbit_r235_c212 bl_212 br_212 wl_235 vdd gnd cell_6t
Xbit_r236_c212 bl_212 br_212 wl_236 vdd gnd cell_6t
Xbit_r237_c212 bl_212 br_212 wl_237 vdd gnd cell_6t
Xbit_r238_c212 bl_212 br_212 wl_238 vdd gnd cell_6t
Xbit_r239_c212 bl_212 br_212 wl_239 vdd gnd cell_6t
Xbit_r240_c212 bl_212 br_212 wl_240 vdd gnd cell_6t
Xbit_r241_c212 bl_212 br_212 wl_241 vdd gnd cell_6t
Xbit_r242_c212 bl_212 br_212 wl_242 vdd gnd cell_6t
Xbit_r243_c212 bl_212 br_212 wl_243 vdd gnd cell_6t
Xbit_r244_c212 bl_212 br_212 wl_244 vdd gnd cell_6t
Xbit_r245_c212 bl_212 br_212 wl_245 vdd gnd cell_6t
Xbit_r246_c212 bl_212 br_212 wl_246 vdd gnd cell_6t
Xbit_r247_c212 bl_212 br_212 wl_247 vdd gnd cell_6t
Xbit_r248_c212 bl_212 br_212 wl_248 vdd gnd cell_6t
Xbit_r249_c212 bl_212 br_212 wl_249 vdd gnd cell_6t
Xbit_r250_c212 bl_212 br_212 wl_250 vdd gnd cell_6t
Xbit_r251_c212 bl_212 br_212 wl_251 vdd gnd cell_6t
Xbit_r252_c212 bl_212 br_212 wl_252 vdd gnd cell_6t
Xbit_r253_c212 bl_212 br_212 wl_253 vdd gnd cell_6t
Xbit_r254_c212 bl_212 br_212 wl_254 vdd gnd cell_6t
Xbit_r255_c212 bl_212 br_212 wl_255 vdd gnd cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd cell_6t
Xbit_r1_c213 bl_213 br_213 wl_1 vdd gnd cell_6t
Xbit_r2_c213 bl_213 br_213 wl_2 vdd gnd cell_6t
Xbit_r3_c213 bl_213 br_213 wl_3 vdd gnd cell_6t
Xbit_r4_c213 bl_213 br_213 wl_4 vdd gnd cell_6t
Xbit_r5_c213 bl_213 br_213 wl_5 vdd gnd cell_6t
Xbit_r6_c213 bl_213 br_213 wl_6 vdd gnd cell_6t
Xbit_r7_c213 bl_213 br_213 wl_7 vdd gnd cell_6t
Xbit_r8_c213 bl_213 br_213 wl_8 vdd gnd cell_6t
Xbit_r9_c213 bl_213 br_213 wl_9 vdd gnd cell_6t
Xbit_r10_c213 bl_213 br_213 wl_10 vdd gnd cell_6t
Xbit_r11_c213 bl_213 br_213 wl_11 vdd gnd cell_6t
Xbit_r12_c213 bl_213 br_213 wl_12 vdd gnd cell_6t
Xbit_r13_c213 bl_213 br_213 wl_13 vdd gnd cell_6t
Xbit_r14_c213 bl_213 br_213 wl_14 vdd gnd cell_6t
Xbit_r15_c213 bl_213 br_213 wl_15 vdd gnd cell_6t
Xbit_r16_c213 bl_213 br_213 wl_16 vdd gnd cell_6t
Xbit_r17_c213 bl_213 br_213 wl_17 vdd gnd cell_6t
Xbit_r18_c213 bl_213 br_213 wl_18 vdd gnd cell_6t
Xbit_r19_c213 bl_213 br_213 wl_19 vdd gnd cell_6t
Xbit_r20_c213 bl_213 br_213 wl_20 vdd gnd cell_6t
Xbit_r21_c213 bl_213 br_213 wl_21 vdd gnd cell_6t
Xbit_r22_c213 bl_213 br_213 wl_22 vdd gnd cell_6t
Xbit_r23_c213 bl_213 br_213 wl_23 vdd gnd cell_6t
Xbit_r24_c213 bl_213 br_213 wl_24 vdd gnd cell_6t
Xbit_r25_c213 bl_213 br_213 wl_25 vdd gnd cell_6t
Xbit_r26_c213 bl_213 br_213 wl_26 vdd gnd cell_6t
Xbit_r27_c213 bl_213 br_213 wl_27 vdd gnd cell_6t
Xbit_r28_c213 bl_213 br_213 wl_28 vdd gnd cell_6t
Xbit_r29_c213 bl_213 br_213 wl_29 vdd gnd cell_6t
Xbit_r30_c213 bl_213 br_213 wl_30 vdd gnd cell_6t
Xbit_r31_c213 bl_213 br_213 wl_31 vdd gnd cell_6t
Xbit_r32_c213 bl_213 br_213 wl_32 vdd gnd cell_6t
Xbit_r33_c213 bl_213 br_213 wl_33 vdd gnd cell_6t
Xbit_r34_c213 bl_213 br_213 wl_34 vdd gnd cell_6t
Xbit_r35_c213 bl_213 br_213 wl_35 vdd gnd cell_6t
Xbit_r36_c213 bl_213 br_213 wl_36 vdd gnd cell_6t
Xbit_r37_c213 bl_213 br_213 wl_37 vdd gnd cell_6t
Xbit_r38_c213 bl_213 br_213 wl_38 vdd gnd cell_6t
Xbit_r39_c213 bl_213 br_213 wl_39 vdd gnd cell_6t
Xbit_r40_c213 bl_213 br_213 wl_40 vdd gnd cell_6t
Xbit_r41_c213 bl_213 br_213 wl_41 vdd gnd cell_6t
Xbit_r42_c213 bl_213 br_213 wl_42 vdd gnd cell_6t
Xbit_r43_c213 bl_213 br_213 wl_43 vdd gnd cell_6t
Xbit_r44_c213 bl_213 br_213 wl_44 vdd gnd cell_6t
Xbit_r45_c213 bl_213 br_213 wl_45 vdd gnd cell_6t
Xbit_r46_c213 bl_213 br_213 wl_46 vdd gnd cell_6t
Xbit_r47_c213 bl_213 br_213 wl_47 vdd gnd cell_6t
Xbit_r48_c213 bl_213 br_213 wl_48 vdd gnd cell_6t
Xbit_r49_c213 bl_213 br_213 wl_49 vdd gnd cell_6t
Xbit_r50_c213 bl_213 br_213 wl_50 vdd gnd cell_6t
Xbit_r51_c213 bl_213 br_213 wl_51 vdd gnd cell_6t
Xbit_r52_c213 bl_213 br_213 wl_52 vdd gnd cell_6t
Xbit_r53_c213 bl_213 br_213 wl_53 vdd gnd cell_6t
Xbit_r54_c213 bl_213 br_213 wl_54 vdd gnd cell_6t
Xbit_r55_c213 bl_213 br_213 wl_55 vdd gnd cell_6t
Xbit_r56_c213 bl_213 br_213 wl_56 vdd gnd cell_6t
Xbit_r57_c213 bl_213 br_213 wl_57 vdd gnd cell_6t
Xbit_r58_c213 bl_213 br_213 wl_58 vdd gnd cell_6t
Xbit_r59_c213 bl_213 br_213 wl_59 vdd gnd cell_6t
Xbit_r60_c213 bl_213 br_213 wl_60 vdd gnd cell_6t
Xbit_r61_c213 bl_213 br_213 wl_61 vdd gnd cell_6t
Xbit_r62_c213 bl_213 br_213 wl_62 vdd gnd cell_6t
Xbit_r63_c213 bl_213 br_213 wl_63 vdd gnd cell_6t
Xbit_r64_c213 bl_213 br_213 wl_64 vdd gnd cell_6t
Xbit_r65_c213 bl_213 br_213 wl_65 vdd gnd cell_6t
Xbit_r66_c213 bl_213 br_213 wl_66 vdd gnd cell_6t
Xbit_r67_c213 bl_213 br_213 wl_67 vdd gnd cell_6t
Xbit_r68_c213 bl_213 br_213 wl_68 vdd gnd cell_6t
Xbit_r69_c213 bl_213 br_213 wl_69 vdd gnd cell_6t
Xbit_r70_c213 bl_213 br_213 wl_70 vdd gnd cell_6t
Xbit_r71_c213 bl_213 br_213 wl_71 vdd gnd cell_6t
Xbit_r72_c213 bl_213 br_213 wl_72 vdd gnd cell_6t
Xbit_r73_c213 bl_213 br_213 wl_73 vdd gnd cell_6t
Xbit_r74_c213 bl_213 br_213 wl_74 vdd gnd cell_6t
Xbit_r75_c213 bl_213 br_213 wl_75 vdd gnd cell_6t
Xbit_r76_c213 bl_213 br_213 wl_76 vdd gnd cell_6t
Xbit_r77_c213 bl_213 br_213 wl_77 vdd gnd cell_6t
Xbit_r78_c213 bl_213 br_213 wl_78 vdd gnd cell_6t
Xbit_r79_c213 bl_213 br_213 wl_79 vdd gnd cell_6t
Xbit_r80_c213 bl_213 br_213 wl_80 vdd gnd cell_6t
Xbit_r81_c213 bl_213 br_213 wl_81 vdd gnd cell_6t
Xbit_r82_c213 bl_213 br_213 wl_82 vdd gnd cell_6t
Xbit_r83_c213 bl_213 br_213 wl_83 vdd gnd cell_6t
Xbit_r84_c213 bl_213 br_213 wl_84 vdd gnd cell_6t
Xbit_r85_c213 bl_213 br_213 wl_85 vdd gnd cell_6t
Xbit_r86_c213 bl_213 br_213 wl_86 vdd gnd cell_6t
Xbit_r87_c213 bl_213 br_213 wl_87 vdd gnd cell_6t
Xbit_r88_c213 bl_213 br_213 wl_88 vdd gnd cell_6t
Xbit_r89_c213 bl_213 br_213 wl_89 vdd gnd cell_6t
Xbit_r90_c213 bl_213 br_213 wl_90 vdd gnd cell_6t
Xbit_r91_c213 bl_213 br_213 wl_91 vdd gnd cell_6t
Xbit_r92_c213 bl_213 br_213 wl_92 vdd gnd cell_6t
Xbit_r93_c213 bl_213 br_213 wl_93 vdd gnd cell_6t
Xbit_r94_c213 bl_213 br_213 wl_94 vdd gnd cell_6t
Xbit_r95_c213 bl_213 br_213 wl_95 vdd gnd cell_6t
Xbit_r96_c213 bl_213 br_213 wl_96 vdd gnd cell_6t
Xbit_r97_c213 bl_213 br_213 wl_97 vdd gnd cell_6t
Xbit_r98_c213 bl_213 br_213 wl_98 vdd gnd cell_6t
Xbit_r99_c213 bl_213 br_213 wl_99 vdd gnd cell_6t
Xbit_r100_c213 bl_213 br_213 wl_100 vdd gnd cell_6t
Xbit_r101_c213 bl_213 br_213 wl_101 vdd gnd cell_6t
Xbit_r102_c213 bl_213 br_213 wl_102 vdd gnd cell_6t
Xbit_r103_c213 bl_213 br_213 wl_103 vdd gnd cell_6t
Xbit_r104_c213 bl_213 br_213 wl_104 vdd gnd cell_6t
Xbit_r105_c213 bl_213 br_213 wl_105 vdd gnd cell_6t
Xbit_r106_c213 bl_213 br_213 wl_106 vdd gnd cell_6t
Xbit_r107_c213 bl_213 br_213 wl_107 vdd gnd cell_6t
Xbit_r108_c213 bl_213 br_213 wl_108 vdd gnd cell_6t
Xbit_r109_c213 bl_213 br_213 wl_109 vdd gnd cell_6t
Xbit_r110_c213 bl_213 br_213 wl_110 vdd gnd cell_6t
Xbit_r111_c213 bl_213 br_213 wl_111 vdd gnd cell_6t
Xbit_r112_c213 bl_213 br_213 wl_112 vdd gnd cell_6t
Xbit_r113_c213 bl_213 br_213 wl_113 vdd gnd cell_6t
Xbit_r114_c213 bl_213 br_213 wl_114 vdd gnd cell_6t
Xbit_r115_c213 bl_213 br_213 wl_115 vdd gnd cell_6t
Xbit_r116_c213 bl_213 br_213 wl_116 vdd gnd cell_6t
Xbit_r117_c213 bl_213 br_213 wl_117 vdd gnd cell_6t
Xbit_r118_c213 bl_213 br_213 wl_118 vdd gnd cell_6t
Xbit_r119_c213 bl_213 br_213 wl_119 vdd gnd cell_6t
Xbit_r120_c213 bl_213 br_213 wl_120 vdd gnd cell_6t
Xbit_r121_c213 bl_213 br_213 wl_121 vdd gnd cell_6t
Xbit_r122_c213 bl_213 br_213 wl_122 vdd gnd cell_6t
Xbit_r123_c213 bl_213 br_213 wl_123 vdd gnd cell_6t
Xbit_r124_c213 bl_213 br_213 wl_124 vdd gnd cell_6t
Xbit_r125_c213 bl_213 br_213 wl_125 vdd gnd cell_6t
Xbit_r126_c213 bl_213 br_213 wl_126 vdd gnd cell_6t
Xbit_r127_c213 bl_213 br_213 wl_127 vdd gnd cell_6t
Xbit_r128_c213 bl_213 br_213 wl_128 vdd gnd cell_6t
Xbit_r129_c213 bl_213 br_213 wl_129 vdd gnd cell_6t
Xbit_r130_c213 bl_213 br_213 wl_130 vdd gnd cell_6t
Xbit_r131_c213 bl_213 br_213 wl_131 vdd gnd cell_6t
Xbit_r132_c213 bl_213 br_213 wl_132 vdd gnd cell_6t
Xbit_r133_c213 bl_213 br_213 wl_133 vdd gnd cell_6t
Xbit_r134_c213 bl_213 br_213 wl_134 vdd gnd cell_6t
Xbit_r135_c213 bl_213 br_213 wl_135 vdd gnd cell_6t
Xbit_r136_c213 bl_213 br_213 wl_136 vdd gnd cell_6t
Xbit_r137_c213 bl_213 br_213 wl_137 vdd gnd cell_6t
Xbit_r138_c213 bl_213 br_213 wl_138 vdd gnd cell_6t
Xbit_r139_c213 bl_213 br_213 wl_139 vdd gnd cell_6t
Xbit_r140_c213 bl_213 br_213 wl_140 vdd gnd cell_6t
Xbit_r141_c213 bl_213 br_213 wl_141 vdd gnd cell_6t
Xbit_r142_c213 bl_213 br_213 wl_142 vdd gnd cell_6t
Xbit_r143_c213 bl_213 br_213 wl_143 vdd gnd cell_6t
Xbit_r144_c213 bl_213 br_213 wl_144 vdd gnd cell_6t
Xbit_r145_c213 bl_213 br_213 wl_145 vdd gnd cell_6t
Xbit_r146_c213 bl_213 br_213 wl_146 vdd gnd cell_6t
Xbit_r147_c213 bl_213 br_213 wl_147 vdd gnd cell_6t
Xbit_r148_c213 bl_213 br_213 wl_148 vdd gnd cell_6t
Xbit_r149_c213 bl_213 br_213 wl_149 vdd gnd cell_6t
Xbit_r150_c213 bl_213 br_213 wl_150 vdd gnd cell_6t
Xbit_r151_c213 bl_213 br_213 wl_151 vdd gnd cell_6t
Xbit_r152_c213 bl_213 br_213 wl_152 vdd gnd cell_6t
Xbit_r153_c213 bl_213 br_213 wl_153 vdd gnd cell_6t
Xbit_r154_c213 bl_213 br_213 wl_154 vdd gnd cell_6t
Xbit_r155_c213 bl_213 br_213 wl_155 vdd gnd cell_6t
Xbit_r156_c213 bl_213 br_213 wl_156 vdd gnd cell_6t
Xbit_r157_c213 bl_213 br_213 wl_157 vdd gnd cell_6t
Xbit_r158_c213 bl_213 br_213 wl_158 vdd gnd cell_6t
Xbit_r159_c213 bl_213 br_213 wl_159 vdd gnd cell_6t
Xbit_r160_c213 bl_213 br_213 wl_160 vdd gnd cell_6t
Xbit_r161_c213 bl_213 br_213 wl_161 vdd gnd cell_6t
Xbit_r162_c213 bl_213 br_213 wl_162 vdd gnd cell_6t
Xbit_r163_c213 bl_213 br_213 wl_163 vdd gnd cell_6t
Xbit_r164_c213 bl_213 br_213 wl_164 vdd gnd cell_6t
Xbit_r165_c213 bl_213 br_213 wl_165 vdd gnd cell_6t
Xbit_r166_c213 bl_213 br_213 wl_166 vdd gnd cell_6t
Xbit_r167_c213 bl_213 br_213 wl_167 vdd gnd cell_6t
Xbit_r168_c213 bl_213 br_213 wl_168 vdd gnd cell_6t
Xbit_r169_c213 bl_213 br_213 wl_169 vdd gnd cell_6t
Xbit_r170_c213 bl_213 br_213 wl_170 vdd gnd cell_6t
Xbit_r171_c213 bl_213 br_213 wl_171 vdd gnd cell_6t
Xbit_r172_c213 bl_213 br_213 wl_172 vdd gnd cell_6t
Xbit_r173_c213 bl_213 br_213 wl_173 vdd gnd cell_6t
Xbit_r174_c213 bl_213 br_213 wl_174 vdd gnd cell_6t
Xbit_r175_c213 bl_213 br_213 wl_175 vdd gnd cell_6t
Xbit_r176_c213 bl_213 br_213 wl_176 vdd gnd cell_6t
Xbit_r177_c213 bl_213 br_213 wl_177 vdd gnd cell_6t
Xbit_r178_c213 bl_213 br_213 wl_178 vdd gnd cell_6t
Xbit_r179_c213 bl_213 br_213 wl_179 vdd gnd cell_6t
Xbit_r180_c213 bl_213 br_213 wl_180 vdd gnd cell_6t
Xbit_r181_c213 bl_213 br_213 wl_181 vdd gnd cell_6t
Xbit_r182_c213 bl_213 br_213 wl_182 vdd gnd cell_6t
Xbit_r183_c213 bl_213 br_213 wl_183 vdd gnd cell_6t
Xbit_r184_c213 bl_213 br_213 wl_184 vdd gnd cell_6t
Xbit_r185_c213 bl_213 br_213 wl_185 vdd gnd cell_6t
Xbit_r186_c213 bl_213 br_213 wl_186 vdd gnd cell_6t
Xbit_r187_c213 bl_213 br_213 wl_187 vdd gnd cell_6t
Xbit_r188_c213 bl_213 br_213 wl_188 vdd gnd cell_6t
Xbit_r189_c213 bl_213 br_213 wl_189 vdd gnd cell_6t
Xbit_r190_c213 bl_213 br_213 wl_190 vdd gnd cell_6t
Xbit_r191_c213 bl_213 br_213 wl_191 vdd gnd cell_6t
Xbit_r192_c213 bl_213 br_213 wl_192 vdd gnd cell_6t
Xbit_r193_c213 bl_213 br_213 wl_193 vdd gnd cell_6t
Xbit_r194_c213 bl_213 br_213 wl_194 vdd gnd cell_6t
Xbit_r195_c213 bl_213 br_213 wl_195 vdd gnd cell_6t
Xbit_r196_c213 bl_213 br_213 wl_196 vdd gnd cell_6t
Xbit_r197_c213 bl_213 br_213 wl_197 vdd gnd cell_6t
Xbit_r198_c213 bl_213 br_213 wl_198 vdd gnd cell_6t
Xbit_r199_c213 bl_213 br_213 wl_199 vdd gnd cell_6t
Xbit_r200_c213 bl_213 br_213 wl_200 vdd gnd cell_6t
Xbit_r201_c213 bl_213 br_213 wl_201 vdd gnd cell_6t
Xbit_r202_c213 bl_213 br_213 wl_202 vdd gnd cell_6t
Xbit_r203_c213 bl_213 br_213 wl_203 vdd gnd cell_6t
Xbit_r204_c213 bl_213 br_213 wl_204 vdd gnd cell_6t
Xbit_r205_c213 bl_213 br_213 wl_205 vdd gnd cell_6t
Xbit_r206_c213 bl_213 br_213 wl_206 vdd gnd cell_6t
Xbit_r207_c213 bl_213 br_213 wl_207 vdd gnd cell_6t
Xbit_r208_c213 bl_213 br_213 wl_208 vdd gnd cell_6t
Xbit_r209_c213 bl_213 br_213 wl_209 vdd gnd cell_6t
Xbit_r210_c213 bl_213 br_213 wl_210 vdd gnd cell_6t
Xbit_r211_c213 bl_213 br_213 wl_211 vdd gnd cell_6t
Xbit_r212_c213 bl_213 br_213 wl_212 vdd gnd cell_6t
Xbit_r213_c213 bl_213 br_213 wl_213 vdd gnd cell_6t
Xbit_r214_c213 bl_213 br_213 wl_214 vdd gnd cell_6t
Xbit_r215_c213 bl_213 br_213 wl_215 vdd gnd cell_6t
Xbit_r216_c213 bl_213 br_213 wl_216 vdd gnd cell_6t
Xbit_r217_c213 bl_213 br_213 wl_217 vdd gnd cell_6t
Xbit_r218_c213 bl_213 br_213 wl_218 vdd gnd cell_6t
Xbit_r219_c213 bl_213 br_213 wl_219 vdd gnd cell_6t
Xbit_r220_c213 bl_213 br_213 wl_220 vdd gnd cell_6t
Xbit_r221_c213 bl_213 br_213 wl_221 vdd gnd cell_6t
Xbit_r222_c213 bl_213 br_213 wl_222 vdd gnd cell_6t
Xbit_r223_c213 bl_213 br_213 wl_223 vdd gnd cell_6t
Xbit_r224_c213 bl_213 br_213 wl_224 vdd gnd cell_6t
Xbit_r225_c213 bl_213 br_213 wl_225 vdd gnd cell_6t
Xbit_r226_c213 bl_213 br_213 wl_226 vdd gnd cell_6t
Xbit_r227_c213 bl_213 br_213 wl_227 vdd gnd cell_6t
Xbit_r228_c213 bl_213 br_213 wl_228 vdd gnd cell_6t
Xbit_r229_c213 bl_213 br_213 wl_229 vdd gnd cell_6t
Xbit_r230_c213 bl_213 br_213 wl_230 vdd gnd cell_6t
Xbit_r231_c213 bl_213 br_213 wl_231 vdd gnd cell_6t
Xbit_r232_c213 bl_213 br_213 wl_232 vdd gnd cell_6t
Xbit_r233_c213 bl_213 br_213 wl_233 vdd gnd cell_6t
Xbit_r234_c213 bl_213 br_213 wl_234 vdd gnd cell_6t
Xbit_r235_c213 bl_213 br_213 wl_235 vdd gnd cell_6t
Xbit_r236_c213 bl_213 br_213 wl_236 vdd gnd cell_6t
Xbit_r237_c213 bl_213 br_213 wl_237 vdd gnd cell_6t
Xbit_r238_c213 bl_213 br_213 wl_238 vdd gnd cell_6t
Xbit_r239_c213 bl_213 br_213 wl_239 vdd gnd cell_6t
Xbit_r240_c213 bl_213 br_213 wl_240 vdd gnd cell_6t
Xbit_r241_c213 bl_213 br_213 wl_241 vdd gnd cell_6t
Xbit_r242_c213 bl_213 br_213 wl_242 vdd gnd cell_6t
Xbit_r243_c213 bl_213 br_213 wl_243 vdd gnd cell_6t
Xbit_r244_c213 bl_213 br_213 wl_244 vdd gnd cell_6t
Xbit_r245_c213 bl_213 br_213 wl_245 vdd gnd cell_6t
Xbit_r246_c213 bl_213 br_213 wl_246 vdd gnd cell_6t
Xbit_r247_c213 bl_213 br_213 wl_247 vdd gnd cell_6t
Xbit_r248_c213 bl_213 br_213 wl_248 vdd gnd cell_6t
Xbit_r249_c213 bl_213 br_213 wl_249 vdd gnd cell_6t
Xbit_r250_c213 bl_213 br_213 wl_250 vdd gnd cell_6t
Xbit_r251_c213 bl_213 br_213 wl_251 vdd gnd cell_6t
Xbit_r252_c213 bl_213 br_213 wl_252 vdd gnd cell_6t
Xbit_r253_c213 bl_213 br_213 wl_253 vdd gnd cell_6t
Xbit_r254_c213 bl_213 br_213 wl_254 vdd gnd cell_6t
Xbit_r255_c213 bl_213 br_213 wl_255 vdd gnd cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd cell_6t
Xbit_r1_c214 bl_214 br_214 wl_1 vdd gnd cell_6t
Xbit_r2_c214 bl_214 br_214 wl_2 vdd gnd cell_6t
Xbit_r3_c214 bl_214 br_214 wl_3 vdd gnd cell_6t
Xbit_r4_c214 bl_214 br_214 wl_4 vdd gnd cell_6t
Xbit_r5_c214 bl_214 br_214 wl_5 vdd gnd cell_6t
Xbit_r6_c214 bl_214 br_214 wl_6 vdd gnd cell_6t
Xbit_r7_c214 bl_214 br_214 wl_7 vdd gnd cell_6t
Xbit_r8_c214 bl_214 br_214 wl_8 vdd gnd cell_6t
Xbit_r9_c214 bl_214 br_214 wl_9 vdd gnd cell_6t
Xbit_r10_c214 bl_214 br_214 wl_10 vdd gnd cell_6t
Xbit_r11_c214 bl_214 br_214 wl_11 vdd gnd cell_6t
Xbit_r12_c214 bl_214 br_214 wl_12 vdd gnd cell_6t
Xbit_r13_c214 bl_214 br_214 wl_13 vdd gnd cell_6t
Xbit_r14_c214 bl_214 br_214 wl_14 vdd gnd cell_6t
Xbit_r15_c214 bl_214 br_214 wl_15 vdd gnd cell_6t
Xbit_r16_c214 bl_214 br_214 wl_16 vdd gnd cell_6t
Xbit_r17_c214 bl_214 br_214 wl_17 vdd gnd cell_6t
Xbit_r18_c214 bl_214 br_214 wl_18 vdd gnd cell_6t
Xbit_r19_c214 bl_214 br_214 wl_19 vdd gnd cell_6t
Xbit_r20_c214 bl_214 br_214 wl_20 vdd gnd cell_6t
Xbit_r21_c214 bl_214 br_214 wl_21 vdd gnd cell_6t
Xbit_r22_c214 bl_214 br_214 wl_22 vdd gnd cell_6t
Xbit_r23_c214 bl_214 br_214 wl_23 vdd gnd cell_6t
Xbit_r24_c214 bl_214 br_214 wl_24 vdd gnd cell_6t
Xbit_r25_c214 bl_214 br_214 wl_25 vdd gnd cell_6t
Xbit_r26_c214 bl_214 br_214 wl_26 vdd gnd cell_6t
Xbit_r27_c214 bl_214 br_214 wl_27 vdd gnd cell_6t
Xbit_r28_c214 bl_214 br_214 wl_28 vdd gnd cell_6t
Xbit_r29_c214 bl_214 br_214 wl_29 vdd gnd cell_6t
Xbit_r30_c214 bl_214 br_214 wl_30 vdd gnd cell_6t
Xbit_r31_c214 bl_214 br_214 wl_31 vdd gnd cell_6t
Xbit_r32_c214 bl_214 br_214 wl_32 vdd gnd cell_6t
Xbit_r33_c214 bl_214 br_214 wl_33 vdd gnd cell_6t
Xbit_r34_c214 bl_214 br_214 wl_34 vdd gnd cell_6t
Xbit_r35_c214 bl_214 br_214 wl_35 vdd gnd cell_6t
Xbit_r36_c214 bl_214 br_214 wl_36 vdd gnd cell_6t
Xbit_r37_c214 bl_214 br_214 wl_37 vdd gnd cell_6t
Xbit_r38_c214 bl_214 br_214 wl_38 vdd gnd cell_6t
Xbit_r39_c214 bl_214 br_214 wl_39 vdd gnd cell_6t
Xbit_r40_c214 bl_214 br_214 wl_40 vdd gnd cell_6t
Xbit_r41_c214 bl_214 br_214 wl_41 vdd gnd cell_6t
Xbit_r42_c214 bl_214 br_214 wl_42 vdd gnd cell_6t
Xbit_r43_c214 bl_214 br_214 wl_43 vdd gnd cell_6t
Xbit_r44_c214 bl_214 br_214 wl_44 vdd gnd cell_6t
Xbit_r45_c214 bl_214 br_214 wl_45 vdd gnd cell_6t
Xbit_r46_c214 bl_214 br_214 wl_46 vdd gnd cell_6t
Xbit_r47_c214 bl_214 br_214 wl_47 vdd gnd cell_6t
Xbit_r48_c214 bl_214 br_214 wl_48 vdd gnd cell_6t
Xbit_r49_c214 bl_214 br_214 wl_49 vdd gnd cell_6t
Xbit_r50_c214 bl_214 br_214 wl_50 vdd gnd cell_6t
Xbit_r51_c214 bl_214 br_214 wl_51 vdd gnd cell_6t
Xbit_r52_c214 bl_214 br_214 wl_52 vdd gnd cell_6t
Xbit_r53_c214 bl_214 br_214 wl_53 vdd gnd cell_6t
Xbit_r54_c214 bl_214 br_214 wl_54 vdd gnd cell_6t
Xbit_r55_c214 bl_214 br_214 wl_55 vdd gnd cell_6t
Xbit_r56_c214 bl_214 br_214 wl_56 vdd gnd cell_6t
Xbit_r57_c214 bl_214 br_214 wl_57 vdd gnd cell_6t
Xbit_r58_c214 bl_214 br_214 wl_58 vdd gnd cell_6t
Xbit_r59_c214 bl_214 br_214 wl_59 vdd gnd cell_6t
Xbit_r60_c214 bl_214 br_214 wl_60 vdd gnd cell_6t
Xbit_r61_c214 bl_214 br_214 wl_61 vdd gnd cell_6t
Xbit_r62_c214 bl_214 br_214 wl_62 vdd gnd cell_6t
Xbit_r63_c214 bl_214 br_214 wl_63 vdd gnd cell_6t
Xbit_r64_c214 bl_214 br_214 wl_64 vdd gnd cell_6t
Xbit_r65_c214 bl_214 br_214 wl_65 vdd gnd cell_6t
Xbit_r66_c214 bl_214 br_214 wl_66 vdd gnd cell_6t
Xbit_r67_c214 bl_214 br_214 wl_67 vdd gnd cell_6t
Xbit_r68_c214 bl_214 br_214 wl_68 vdd gnd cell_6t
Xbit_r69_c214 bl_214 br_214 wl_69 vdd gnd cell_6t
Xbit_r70_c214 bl_214 br_214 wl_70 vdd gnd cell_6t
Xbit_r71_c214 bl_214 br_214 wl_71 vdd gnd cell_6t
Xbit_r72_c214 bl_214 br_214 wl_72 vdd gnd cell_6t
Xbit_r73_c214 bl_214 br_214 wl_73 vdd gnd cell_6t
Xbit_r74_c214 bl_214 br_214 wl_74 vdd gnd cell_6t
Xbit_r75_c214 bl_214 br_214 wl_75 vdd gnd cell_6t
Xbit_r76_c214 bl_214 br_214 wl_76 vdd gnd cell_6t
Xbit_r77_c214 bl_214 br_214 wl_77 vdd gnd cell_6t
Xbit_r78_c214 bl_214 br_214 wl_78 vdd gnd cell_6t
Xbit_r79_c214 bl_214 br_214 wl_79 vdd gnd cell_6t
Xbit_r80_c214 bl_214 br_214 wl_80 vdd gnd cell_6t
Xbit_r81_c214 bl_214 br_214 wl_81 vdd gnd cell_6t
Xbit_r82_c214 bl_214 br_214 wl_82 vdd gnd cell_6t
Xbit_r83_c214 bl_214 br_214 wl_83 vdd gnd cell_6t
Xbit_r84_c214 bl_214 br_214 wl_84 vdd gnd cell_6t
Xbit_r85_c214 bl_214 br_214 wl_85 vdd gnd cell_6t
Xbit_r86_c214 bl_214 br_214 wl_86 vdd gnd cell_6t
Xbit_r87_c214 bl_214 br_214 wl_87 vdd gnd cell_6t
Xbit_r88_c214 bl_214 br_214 wl_88 vdd gnd cell_6t
Xbit_r89_c214 bl_214 br_214 wl_89 vdd gnd cell_6t
Xbit_r90_c214 bl_214 br_214 wl_90 vdd gnd cell_6t
Xbit_r91_c214 bl_214 br_214 wl_91 vdd gnd cell_6t
Xbit_r92_c214 bl_214 br_214 wl_92 vdd gnd cell_6t
Xbit_r93_c214 bl_214 br_214 wl_93 vdd gnd cell_6t
Xbit_r94_c214 bl_214 br_214 wl_94 vdd gnd cell_6t
Xbit_r95_c214 bl_214 br_214 wl_95 vdd gnd cell_6t
Xbit_r96_c214 bl_214 br_214 wl_96 vdd gnd cell_6t
Xbit_r97_c214 bl_214 br_214 wl_97 vdd gnd cell_6t
Xbit_r98_c214 bl_214 br_214 wl_98 vdd gnd cell_6t
Xbit_r99_c214 bl_214 br_214 wl_99 vdd gnd cell_6t
Xbit_r100_c214 bl_214 br_214 wl_100 vdd gnd cell_6t
Xbit_r101_c214 bl_214 br_214 wl_101 vdd gnd cell_6t
Xbit_r102_c214 bl_214 br_214 wl_102 vdd gnd cell_6t
Xbit_r103_c214 bl_214 br_214 wl_103 vdd gnd cell_6t
Xbit_r104_c214 bl_214 br_214 wl_104 vdd gnd cell_6t
Xbit_r105_c214 bl_214 br_214 wl_105 vdd gnd cell_6t
Xbit_r106_c214 bl_214 br_214 wl_106 vdd gnd cell_6t
Xbit_r107_c214 bl_214 br_214 wl_107 vdd gnd cell_6t
Xbit_r108_c214 bl_214 br_214 wl_108 vdd gnd cell_6t
Xbit_r109_c214 bl_214 br_214 wl_109 vdd gnd cell_6t
Xbit_r110_c214 bl_214 br_214 wl_110 vdd gnd cell_6t
Xbit_r111_c214 bl_214 br_214 wl_111 vdd gnd cell_6t
Xbit_r112_c214 bl_214 br_214 wl_112 vdd gnd cell_6t
Xbit_r113_c214 bl_214 br_214 wl_113 vdd gnd cell_6t
Xbit_r114_c214 bl_214 br_214 wl_114 vdd gnd cell_6t
Xbit_r115_c214 bl_214 br_214 wl_115 vdd gnd cell_6t
Xbit_r116_c214 bl_214 br_214 wl_116 vdd gnd cell_6t
Xbit_r117_c214 bl_214 br_214 wl_117 vdd gnd cell_6t
Xbit_r118_c214 bl_214 br_214 wl_118 vdd gnd cell_6t
Xbit_r119_c214 bl_214 br_214 wl_119 vdd gnd cell_6t
Xbit_r120_c214 bl_214 br_214 wl_120 vdd gnd cell_6t
Xbit_r121_c214 bl_214 br_214 wl_121 vdd gnd cell_6t
Xbit_r122_c214 bl_214 br_214 wl_122 vdd gnd cell_6t
Xbit_r123_c214 bl_214 br_214 wl_123 vdd gnd cell_6t
Xbit_r124_c214 bl_214 br_214 wl_124 vdd gnd cell_6t
Xbit_r125_c214 bl_214 br_214 wl_125 vdd gnd cell_6t
Xbit_r126_c214 bl_214 br_214 wl_126 vdd gnd cell_6t
Xbit_r127_c214 bl_214 br_214 wl_127 vdd gnd cell_6t
Xbit_r128_c214 bl_214 br_214 wl_128 vdd gnd cell_6t
Xbit_r129_c214 bl_214 br_214 wl_129 vdd gnd cell_6t
Xbit_r130_c214 bl_214 br_214 wl_130 vdd gnd cell_6t
Xbit_r131_c214 bl_214 br_214 wl_131 vdd gnd cell_6t
Xbit_r132_c214 bl_214 br_214 wl_132 vdd gnd cell_6t
Xbit_r133_c214 bl_214 br_214 wl_133 vdd gnd cell_6t
Xbit_r134_c214 bl_214 br_214 wl_134 vdd gnd cell_6t
Xbit_r135_c214 bl_214 br_214 wl_135 vdd gnd cell_6t
Xbit_r136_c214 bl_214 br_214 wl_136 vdd gnd cell_6t
Xbit_r137_c214 bl_214 br_214 wl_137 vdd gnd cell_6t
Xbit_r138_c214 bl_214 br_214 wl_138 vdd gnd cell_6t
Xbit_r139_c214 bl_214 br_214 wl_139 vdd gnd cell_6t
Xbit_r140_c214 bl_214 br_214 wl_140 vdd gnd cell_6t
Xbit_r141_c214 bl_214 br_214 wl_141 vdd gnd cell_6t
Xbit_r142_c214 bl_214 br_214 wl_142 vdd gnd cell_6t
Xbit_r143_c214 bl_214 br_214 wl_143 vdd gnd cell_6t
Xbit_r144_c214 bl_214 br_214 wl_144 vdd gnd cell_6t
Xbit_r145_c214 bl_214 br_214 wl_145 vdd gnd cell_6t
Xbit_r146_c214 bl_214 br_214 wl_146 vdd gnd cell_6t
Xbit_r147_c214 bl_214 br_214 wl_147 vdd gnd cell_6t
Xbit_r148_c214 bl_214 br_214 wl_148 vdd gnd cell_6t
Xbit_r149_c214 bl_214 br_214 wl_149 vdd gnd cell_6t
Xbit_r150_c214 bl_214 br_214 wl_150 vdd gnd cell_6t
Xbit_r151_c214 bl_214 br_214 wl_151 vdd gnd cell_6t
Xbit_r152_c214 bl_214 br_214 wl_152 vdd gnd cell_6t
Xbit_r153_c214 bl_214 br_214 wl_153 vdd gnd cell_6t
Xbit_r154_c214 bl_214 br_214 wl_154 vdd gnd cell_6t
Xbit_r155_c214 bl_214 br_214 wl_155 vdd gnd cell_6t
Xbit_r156_c214 bl_214 br_214 wl_156 vdd gnd cell_6t
Xbit_r157_c214 bl_214 br_214 wl_157 vdd gnd cell_6t
Xbit_r158_c214 bl_214 br_214 wl_158 vdd gnd cell_6t
Xbit_r159_c214 bl_214 br_214 wl_159 vdd gnd cell_6t
Xbit_r160_c214 bl_214 br_214 wl_160 vdd gnd cell_6t
Xbit_r161_c214 bl_214 br_214 wl_161 vdd gnd cell_6t
Xbit_r162_c214 bl_214 br_214 wl_162 vdd gnd cell_6t
Xbit_r163_c214 bl_214 br_214 wl_163 vdd gnd cell_6t
Xbit_r164_c214 bl_214 br_214 wl_164 vdd gnd cell_6t
Xbit_r165_c214 bl_214 br_214 wl_165 vdd gnd cell_6t
Xbit_r166_c214 bl_214 br_214 wl_166 vdd gnd cell_6t
Xbit_r167_c214 bl_214 br_214 wl_167 vdd gnd cell_6t
Xbit_r168_c214 bl_214 br_214 wl_168 vdd gnd cell_6t
Xbit_r169_c214 bl_214 br_214 wl_169 vdd gnd cell_6t
Xbit_r170_c214 bl_214 br_214 wl_170 vdd gnd cell_6t
Xbit_r171_c214 bl_214 br_214 wl_171 vdd gnd cell_6t
Xbit_r172_c214 bl_214 br_214 wl_172 vdd gnd cell_6t
Xbit_r173_c214 bl_214 br_214 wl_173 vdd gnd cell_6t
Xbit_r174_c214 bl_214 br_214 wl_174 vdd gnd cell_6t
Xbit_r175_c214 bl_214 br_214 wl_175 vdd gnd cell_6t
Xbit_r176_c214 bl_214 br_214 wl_176 vdd gnd cell_6t
Xbit_r177_c214 bl_214 br_214 wl_177 vdd gnd cell_6t
Xbit_r178_c214 bl_214 br_214 wl_178 vdd gnd cell_6t
Xbit_r179_c214 bl_214 br_214 wl_179 vdd gnd cell_6t
Xbit_r180_c214 bl_214 br_214 wl_180 vdd gnd cell_6t
Xbit_r181_c214 bl_214 br_214 wl_181 vdd gnd cell_6t
Xbit_r182_c214 bl_214 br_214 wl_182 vdd gnd cell_6t
Xbit_r183_c214 bl_214 br_214 wl_183 vdd gnd cell_6t
Xbit_r184_c214 bl_214 br_214 wl_184 vdd gnd cell_6t
Xbit_r185_c214 bl_214 br_214 wl_185 vdd gnd cell_6t
Xbit_r186_c214 bl_214 br_214 wl_186 vdd gnd cell_6t
Xbit_r187_c214 bl_214 br_214 wl_187 vdd gnd cell_6t
Xbit_r188_c214 bl_214 br_214 wl_188 vdd gnd cell_6t
Xbit_r189_c214 bl_214 br_214 wl_189 vdd gnd cell_6t
Xbit_r190_c214 bl_214 br_214 wl_190 vdd gnd cell_6t
Xbit_r191_c214 bl_214 br_214 wl_191 vdd gnd cell_6t
Xbit_r192_c214 bl_214 br_214 wl_192 vdd gnd cell_6t
Xbit_r193_c214 bl_214 br_214 wl_193 vdd gnd cell_6t
Xbit_r194_c214 bl_214 br_214 wl_194 vdd gnd cell_6t
Xbit_r195_c214 bl_214 br_214 wl_195 vdd gnd cell_6t
Xbit_r196_c214 bl_214 br_214 wl_196 vdd gnd cell_6t
Xbit_r197_c214 bl_214 br_214 wl_197 vdd gnd cell_6t
Xbit_r198_c214 bl_214 br_214 wl_198 vdd gnd cell_6t
Xbit_r199_c214 bl_214 br_214 wl_199 vdd gnd cell_6t
Xbit_r200_c214 bl_214 br_214 wl_200 vdd gnd cell_6t
Xbit_r201_c214 bl_214 br_214 wl_201 vdd gnd cell_6t
Xbit_r202_c214 bl_214 br_214 wl_202 vdd gnd cell_6t
Xbit_r203_c214 bl_214 br_214 wl_203 vdd gnd cell_6t
Xbit_r204_c214 bl_214 br_214 wl_204 vdd gnd cell_6t
Xbit_r205_c214 bl_214 br_214 wl_205 vdd gnd cell_6t
Xbit_r206_c214 bl_214 br_214 wl_206 vdd gnd cell_6t
Xbit_r207_c214 bl_214 br_214 wl_207 vdd gnd cell_6t
Xbit_r208_c214 bl_214 br_214 wl_208 vdd gnd cell_6t
Xbit_r209_c214 bl_214 br_214 wl_209 vdd gnd cell_6t
Xbit_r210_c214 bl_214 br_214 wl_210 vdd gnd cell_6t
Xbit_r211_c214 bl_214 br_214 wl_211 vdd gnd cell_6t
Xbit_r212_c214 bl_214 br_214 wl_212 vdd gnd cell_6t
Xbit_r213_c214 bl_214 br_214 wl_213 vdd gnd cell_6t
Xbit_r214_c214 bl_214 br_214 wl_214 vdd gnd cell_6t
Xbit_r215_c214 bl_214 br_214 wl_215 vdd gnd cell_6t
Xbit_r216_c214 bl_214 br_214 wl_216 vdd gnd cell_6t
Xbit_r217_c214 bl_214 br_214 wl_217 vdd gnd cell_6t
Xbit_r218_c214 bl_214 br_214 wl_218 vdd gnd cell_6t
Xbit_r219_c214 bl_214 br_214 wl_219 vdd gnd cell_6t
Xbit_r220_c214 bl_214 br_214 wl_220 vdd gnd cell_6t
Xbit_r221_c214 bl_214 br_214 wl_221 vdd gnd cell_6t
Xbit_r222_c214 bl_214 br_214 wl_222 vdd gnd cell_6t
Xbit_r223_c214 bl_214 br_214 wl_223 vdd gnd cell_6t
Xbit_r224_c214 bl_214 br_214 wl_224 vdd gnd cell_6t
Xbit_r225_c214 bl_214 br_214 wl_225 vdd gnd cell_6t
Xbit_r226_c214 bl_214 br_214 wl_226 vdd gnd cell_6t
Xbit_r227_c214 bl_214 br_214 wl_227 vdd gnd cell_6t
Xbit_r228_c214 bl_214 br_214 wl_228 vdd gnd cell_6t
Xbit_r229_c214 bl_214 br_214 wl_229 vdd gnd cell_6t
Xbit_r230_c214 bl_214 br_214 wl_230 vdd gnd cell_6t
Xbit_r231_c214 bl_214 br_214 wl_231 vdd gnd cell_6t
Xbit_r232_c214 bl_214 br_214 wl_232 vdd gnd cell_6t
Xbit_r233_c214 bl_214 br_214 wl_233 vdd gnd cell_6t
Xbit_r234_c214 bl_214 br_214 wl_234 vdd gnd cell_6t
Xbit_r235_c214 bl_214 br_214 wl_235 vdd gnd cell_6t
Xbit_r236_c214 bl_214 br_214 wl_236 vdd gnd cell_6t
Xbit_r237_c214 bl_214 br_214 wl_237 vdd gnd cell_6t
Xbit_r238_c214 bl_214 br_214 wl_238 vdd gnd cell_6t
Xbit_r239_c214 bl_214 br_214 wl_239 vdd gnd cell_6t
Xbit_r240_c214 bl_214 br_214 wl_240 vdd gnd cell_6t
Xbit_r241_c214 bl_214 br_214 wl_241 vdd gnd cell_6t
Xbit_r242_c214 bl_214 br_214 wl_242 vdd gnd cell_6t
Xbit_r243_c214 bl_214 br_214 wl_243 vdd gnd cell_6t
Xbit_r244_c214 bl_214 br_214 wl_244 vdd gnd cell_6t
Xbit_r245_c214 bl_214 br_214 wl_245 vdd gnd cell_6t
Xbit_r246_c214 bl_214 br_214 wl_246 vdd gnd cell_6t
Xbit_r247_c214 bl_214 br_214 wl_247 vdd gnd cell_6t
Xbit_r248_c214 bl_214 br_214 wl_248 vdd gnd cell_6t
Xbit_r249_c214 bl_214 br_214 wl_249 vdd gnd cell_6t
Xbit_r250_c214 bl_214 br_214 wl_250 vdd gnd cell_6t
Xbit_r251_c214 bl_214 br_214 wl_251 vdd gnd cell_6t
Xbit_r252_c214 bl_214 br_214 wl_252 vdd gnd cell_6t
Xbit_r253_c214 bl_214 br_214 wl_253 vdd gnd cell_6t
Xbit_r254_c214 bl_214 br_214 wl_254 vdd gnd cell_6t
Xbit_r255_c214 bl_214 br_214 wl_255 vdd gnd cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd cell_6t
Xbit_r1_c215 bl_215 br_215 wl_1 vdd gnd cell_6t
Xbit_r2_c215 bl_215 br_215 wl_2 vdd gnd cell_6t
Xbit_r3_c215 bl_215 br_215 wl_3 vdd gnd cell_6t
Xbit_r4_c215 bl_215 br_215 wl_4 vdd gnd cell_6t
Xbit_r5_c215 bl_215 br_215 wl_5 vdd gnd cell_6t
Xbit_r6_c215 bl_215 br_215 wl_6 vdd gnd cell_6t
Xbit_r7_c215 bl_215 br_215 wl_7 vdd gnd cell_6t
Xbit_r8_c215 bl_215 br_215 wl_8 vdd gnd cell_6t
Xbit_r9_c215 bl_215 br_215 wl_9 vdd gnd cell_6t
Xbit_r10_c215 bl_215 br_215 wl_10 vdd gnd cell_6t
Xbit_r11_c215 bl_215 br_215 wl_11 vdd gnd cell_6t
Xbit_r12_c215 bl_215 br_215 wl_12 vdd gnd cell_6t
Xbit_r13_c215 bl_215 br_215 wl_13 vdd gnd cell_6t
Xbit_r14_c215 bl_215 br_215 wl_14 vdd gnd cell_6t
Xbit_r15_c215 bl_215 br_215 wl_15 vdd gnd cell_6t
Xbit_r16_c215 bl_215 br_215 wl_16 vdd gnd cell_6t
Xbit_r17_c215 bl_215 br_215 wl_17 vdd gnd cell_6t
Xbit_r18_c215 bl_215 br_215 wl_18 vdd gnd cell_6t
Xbit_r19_c215 bl_215 br_215 wl_19 vdd gnd cell_6t
Xbit_r20_c215 bl_215 br_215 wl_20 vdd gnd cell_6t
Xbit_r21_c215 bl_215 br_215 wl_21 vdd gnd cell_6t
Xbit_r22_c215 bl_215 br_215 wl_22 vdd gnd cell_6t
Xbit_r23_c215 bl_215 br_215 wl_23 vdd gnd cell_6t
Xbit_r24_c215 bl_215 br_215 wl_24 vdd gnd cell_6t
Xbit_r25_c215 bl_215 br_215 wl_25 vdd gnd cell_6t
Xbit_r26_c215 bl_215 br_215 wl_26 vdd gnd cell_6t
Xbit_r27_c215 bl_215 br_215 wl_27 vdd gnd cell_6t
Xbit_r28_c215 bl_215 br_215 wl_28 vdd gnd cell_6t
Xbit_r29_c215 bl_215 br_215 wl_29 vdd gnd cell_6t
Xbit_r30_c215 bl_215 br_215 wl_30 vdd gnd cell_6t
Xbit_r31_c215 bl_215 br_215 wl_31 vdd gnd cell_6t
Xbit_r32_c215 bl_215 br_215 wl_32 vdd gnd cell_6t
Xbit_r33_c215 bl_215 br_215 wl_33 vdd gnd cell_6t
Xbit_r34_c215 bl_215 br_215 wl_34 vdd gnd cell_6t
Xbit_r35_c215 bl_215 br_215 wl_35 vdd gnd cell_6t
Xbit_r36_c215 bl_215 br_215 wl_36 vdd gnd cell_6t
Xbit_r37_c215 bl_215 br_215 wl_37 vdd gnd cell_6t
Xbit_r38_c215 bl_215 br_215 wl_38 vdd gnd cell_6t
Xbit_r39_c215 bl_215 br_215 wl_39 vdd gnd cell_6t
Xbit_r40_c215 bl_215 br_215 wl_40 vdd gnd cell_6t
Xbit_r41_c215 bl_215 br_215 wl_41 vdd gnd cell_6t
Xbit_r42_c215 bl_215 br_215 wl_42 vdd gnd cell_6t
Xbit_r43_c215 bl_215 br_215 wl_43 vdd gnd cell_6t
Xbit_r44_c215 bl_215 br_215 wl_44 vdd gnd cell_6t
Xbit_r45_c215 bl_215 br_215 wl_45 vdd gnd cell_6t
Xbit_r46_c215 bl_215 br_215 wl_46 vdd gnd cell_6t
Xbit_r47_c215 bl_215 br_215 wl_47 vdd gnd cell_6t
Xbit_r48_c215 bl_215 br_215 wl_48 vdd gnd cell_6t
Xbit_r49_c215 bl_215 br_215 wl_49 vdd gnd cell_6t
Xbit_r50_c215 bl_215 br_215 wl_50 vdd gnd cell_6t
Xbit_r51_c215 bl_215 br_215 wl_51 vdd gnd cell_6t
Xbit_r52_c215 bl_215 br_215 wl_52 vdd gnd cell_6t
Xbit_r53_c215 bl_215 br_215 wl_53 vdd gnd cell_6t
Xbit_r54_c215 bl_215 br_215 wl_54 vdd gnd cell_6t
Xbit_r55_c215 bl_215 br_215 wl_55 vdd gnd cell_6t
Xbit_r56_c215 bl_215 br_215 wl_56 vdd gnd cell_6t
Xbit_r57_c215 bl_215 br_215 wl_57 vdd gnd cell_6t
Xbit_r58_c215 bl_215 br_215 wl_58 vdd gnd cell_6t
Xbit_r59_c215 bl_215 br_215 wl_59 vdd gnd cell_6t
Xbit_r60_c215 bl_215 br_215 wl_60 vdd gnd cell_6t
Xbit_r61_c215 bl_215 br_215 wl_61 vdd gnd cell_6t
Xbit_r62_c215 bl_215 br_215 wl_62 vdd gnd cell_6t
Xbit_r63_c215 bl_215 br_215 wl_63 vdd gnd cell_6t
Xbit_r64_c215 bl_215 br_215 wl_64 vdd gnd cell_6t
Xbit_r65_c215 bl_215 br_215 wl_65 vdd gnd cell_6t
Xbit_r66_c215 bl_215 br_215 wl_66 vdd gnd cell_6t
Xbit_r67_c215 bl_215 br_215 wl_67 vdd gnd cell_6t
Xbit_r68_c215 bl_215 br_215 wl_68 vdd gnd cell_6t
Xbit_r69_c215 bl_215 br_215 wl_69 vdd gnd cell_6t
Xbit_r70_c215 bl_215 br_215 wl_70 vdd gnd cell_6t
Xbit_r71_c215 bl_215 br_215 wl_71 vdd gnd cell_6t
Xbit_r72_c215 bl_215 br_215 wl_72 vdd gnd cell_6t
Xbit_r73_c215 bl_215 br_215 wl_73 vdd gnd cell_6t
Xbit_r74_c215 bl_215 br_215 wl_74 vdd gnd cell_6t
Xbit_r75_c215 bl_215 br_215 wl_75 vdd gnd cell_6t
Xbit_r76_c215 bl_215 br_215 wl_76 vdd gnd cell_6t
Xbit_r77_c215 bl_215 br_215 wl_77 vdd gnd cell_6t
Xbit_r78_c215 bl_215 br_215 wl_78 vdd gnd cell_6t
Xbit_r79_c215 bl_215 br_215 wl_79 vdd gnd cell_6t
Xbit_r80_c215 bl_215 br_215 wl_80 vdd gnd cell_6t
Xbit_r81_c215 bl_215 br_215 wl_81 vdd gnd cell_6t
Xbit_r82_c215 bl_215 br_215 wl_82 vdd gnd cell_6t
Xbit_r83_c215 bl_215 br_215 wl_83 vdd gnd cell_6t
Xbit_r84_c215 bl_215 br_215 wl_84 vdd gnd cell_6t
Xbit_r85_c215 bl_215 br_215 wl_85 vdd gnd cell_6t
Xbit_r86_c215 bl_215 br_215 wl_86 vdd gnd cell_6t
Xbit_r87_c215 bl_215 br_215 wl_87 vdd gnd cell_6t
Xbit_r88_c215 bl_215 br_215 wl_88 vdd gnd cell_6t
Xbit_r89_c215 bl_215 br_215 wl_89 vdd gnd cell_6t
Xbit_r90_c215 bl_215 br_215 wl_90 vdd gnd cell_6t
Xbit_r91_c215 bl_215 br_215 wl_91 vdd gnd cell_6t
Xbit_r92_c215 bl_215 br_215 wl_92 vdd gnd cell_6t
Xbit_r93_c215 bl_215 br_215 wl_93 vdd gnd cell_6t
Xbit_r94_c215 bl_215 br_215 wl_94 vdd gnd cell_6t
Xbit_r95_c215 bl_215 br_215 wl_95 vdd gnd cell_6t
Xbit_r96_c215 bl_215 br_215 wl_96 vdd gnd cell_6t
Xbit_r97_c215 bl_215 br_215 wl_97 vdd gnd cell_6t
Xbit_r98_c215 bl_215 br_215 wl_98 vdd gnd cell_6t
Xbit_r99_c215 bl_215 br_215 wl_99 vdd gnd cell_6t
Xbit_r100_c215 bl_215 br_215 wl_100 vdd gnd cell_6t
Xbit_r101_c215 bl_215 br_215 wl_101 vdd gnd cell_6t
Xbit_r102_c215 bl_215 br_215 wl_102 vdd gnd cell_6t
Xbit_r103_c215 bl_215 br_215 wl_103 vdd gnd cell_6t
Xbit_r104_c215 bl_215 br_215 wl_104 vdd gnd cell_6t
Xbit_r105_c215 bl_215 br_215 wl_105 vdd gnd cell_6t
Xbit_r106_c215 bl_215 br_215 wl_106 vdd gnd cell_6t
Xbit_r107_c215 bl_215 br_215 wl_107 vdd gnd cell_6t
Xbit_r108_c215 bl_215 br_215 wl_108 vdd gnd cell_6t
Xbit_r109_c215 bl_215 br_215 wl_109 vdd gnd cell_6t
Xbit_r110_c215 bl_215 br_215 wl_110 vdd gnd cell_6t
Xbit_r111_c215 bl_215 br_215 wl_111 vdd gnd cell_6t
Xbit_r112_c215 bl_215 br_215 wl_112 vdd gnd cell_6t
Xbit_r113_c215 bl_215 br_215 wl_113 vdd gnd cell_6t
Xbit_r114_c215 bl_215 br_215 wl_114 vdd gnd cell_6t
Xbit_r115_c215 bl_215 br_215 wl_115 vdd gnd cell_6t
Xbit_r116_c215 bl_215 br_215 wl_116 vdd gnd cell_6t
Xbit_r117_c215 bl_215 br_215 wl_117 vdd gnd cell_6t
Xbit_r118_c215 bl_215 br_215 wl_118 vdd gnd cell_6t
Xbit_r119_c215 bl_215 br_215 wl_119 vdd gnd cell_6t
Xbit_r120_c215 bl_215 br_215 wl_120 vdd gnd cell_6t
Xbit_r121_c215 bl_215 br_215 wl_121 vdd gnd cell_6t
Xbit_r122_c215 bl_215 br_215 wl_122 vdd gnd cell_6t
Xbit_r123_c215 bl_215 br_215 wl_123 vdd gnd cell_6t
Xbit_r124_c215 bl_215 br_215 wl_124 vdd gnd cell_6t
Xbit_r125_c215 bl_215 br_215 wl_125 vdd gnd cell_6t
Xbit_r126_c215 bl_215 br_215 wl_126 vdd gnd cell_6t
Xbit_r127_c215 bl_215 br_215 wl_127 vdd gnd cell_6t
Xbit_r128_c215 bl_215 br_215 wl_128 vdd gnd cell_6t
Xbit_r129_c215 bl_215 br_215 wl_129 vdd gnd cell_6t
Xbit_r130_c215 bl_215 br_215 wl_130 vdd gnd cell_6t
Xbit_r131_c215 bl_215 br_215 wl_131 vdd gnd cell_6t
Xbit_r132_c215 bl_215 br_215 wl_132 vdd gnd cell_6t
Xbit_r133_c215 bl_215 br_215 wl_133 vdd gnd cell_6t
Xbit_r134_c215 bl_215 br_215 wl_134 vdd gnd cell_6t
Xbit_r135_c215 bl_215 br_215 wl_135 vdd gnd cell_6t
Xbit_r136_c215 bl_215 br_215 wl_136 vdd gnd cell_6t
Xbit_r137_c215 bl_215 br_215 wl_137 vdd gnd cell_6t
Xbit_r138_c215 bl_215 br_215 wl_138 vdd gnd cell_6t
Xbit_r139_c215 bl_215 br_215 wl_139 vdd gnd cell_6t
Xbit_r140_c215 bl_215 br_215 wl_140 vdd gnd cell_6t
Xbit_r141_c215 bl_215 br_215 wl_141 vdd gnd cell_6t
Xbit_r142_c215 bl_215 br_215 wl_142 vdd gnd cell_6t
Xbit_r143_c215 bl_215 br_215 wl_143 vdd gnd cell_6t
Xbit_r144_c215 bl_215 br_215 wl_144 vdd gnd cell_6t
Xbit_r145_c215 bl_215 br_215 wl_145 vdd gnd cell_6t
Xbit_r146_c215 bl_215 br_215 wl_146 vdd gnd cell_6t
Xbit_r147_c215 bl_215 br_215 wl_147 vdd gnd cell_6t
Xbit_r148_c215 bl_215 br_215 wl_148 vdd gnd cell_6t
Xbit_r149_c215 bl_215 br_215 wl_149 vdd gnd cell_6t
Xbit_r150_c215 bl_215 br_215 wl_150 vdd gnd cell_6t
Xbit_r151_c215 bl_215 br_215 wl_151 vdd gnd cell_6t
Xbit_r152_c215 bl_215 br_215 wl_152 vdd gnd cell_6t
Xbit_r153_c215 bl_215 br_215 wl_153 vdd gnd cell_6t
Xbit_r154_c215 bl_215 br_215 wl_154 vdd gnd cell_6t
Xbit_r155_c215 bl_215 br_215 wl_155 vdd gnd cell_6t
Xbit_r156_c215 bl_215 br_215 wl_156 vdd gnd cell_6t
Xbit_r157_c215 bl_215 br_215 wl_157 vdd gnd cell_6t
Xbit_r158_c215 bl_215 br_215 wl_158 vdd gnd cell_6t
Xbit_r159_c215 bl_215 br_215 wl_159 vdd gnd cell_6t
Xbit_r160_c215 bl_215 br_215 wl_160 vdd gnd cell_6t
Xbit_r161_c215 bl_215 br_215 wl_161 vdd gnd cell_6t
Xbit_r162_c215 bl_215 br_215 wl_162 vdd gnd cell_6t
Xbit_r163_c215 bl_215 br_215 wl_163 vdd gnd cell_6t
Xbit_r164_c215 bl_215 br_215 wl_164 vdd gnd cell_6t
Xbit_r165_c215 bl_215 br_215 wl_165 vdd gnd cell_6t
Xbit_r166_c215 bl_215 br_215 wl_166 vdd gnd cell_6t
Xbit_r167_c215 bl_215 br_215 wl_167 vdd gnd cell_6t
Xbit_r168_c215 bl_215 br_215 wl_168 vdd gnd cell_6t
Xbit_r169_c215 bl_215 br_215 wl_169 vdd gnd cell_6t
Xbit_r170_c215 bl_215 br_215 wl_170 vdd gnd cell_6t
Xbit_r171_c215 bl_215 br_215 wl_171 vdd gnd cell_6t
Xbit_r172_c215 bl_215 br_215 wl_172 vdd gnd cell_6t
Xbit_r173_c215 bl_215 br_215 wl_173 vdd gnd cell_6t
Xbit_r174_c215 bl_215 br_215 wl_174 vdd gnd cell_6t
Xbit_r175_c215 bl_215 br_215 wl_175 vdd gnd cell_6t
Xbit_r176_c215 bl_215 br_215 wl_176 vdd gnd cell_6t
Xbit_r177_c215 bl_215 br_215 wl_177 vdd gnd cell_6t
Xbit_r178_c215 bl_215 br_215 wl_178 vdd gnd cell_6t
Xbit_r179_c215 bl_215 br_215 wl_179 vdd gnd cell_6t
Xbit_r180_c215 bl_215 br_215 wl_180 vdd gnd cell_6t
Xbit_r181_c215 bl_215 br_215 wl_181 vdd gnd cell_6t
Xbit_r182_c215 bl_215 br_215 wl_182 vdd gnd cell_6t
Xbit_r183_c215 bl_215 br_215 wl_183 vdd gnd cell_6t
Xbit_r184_c215 bl_215 br_215 wl_184 vdd gnd cell_6t
Xbit_r185_c215 bl_215 br_215 wl_185 vdd gnd cell_6t
Xbit_r186_c215 bl_215 br_215 wl_186 vdd gnd cell_6t
Xbit_r187_c215 bl_215 br_215 wl_187 vdd gnd cell_6t
Xbit_r188_c215 bl_215 br_215 wl_188 vdd gnd cell_6t
Xbit_r189_c215 bl_215 br_215 wl_189 vdd gnd cell_6t
Xbit_r190_c215 bl_215 br_215 wl_190 vdd gnd cell_6t
Xbit_r191_c215 bl_215 br_215 wl_191 vdd gnd cell_6t
Xbit_r192_c215 bl_215 br_215 wl_192 vdd gnd cell_6t
Xbit_r193_c215 bl_215 br_215 wl_193 vdd gnd cell_6t
Xbit_r194_c215 bl_215 br_215 wl_194 vdd gnd cell_6t
Xbit_r195_c215 bl_215 br_215 wl_195 vdd gnd cell_6t
Xbit_r196_c215 bl_215 br_215 wl_196 vdd gnd cell_6t
Xbit_r197_c215 bl_215 br_215 wl_197 vdd gnd cell_6t
Xbit_r198_c215 bl_215 br_215 wl_198 vdd gnd cell_6t
Xbit_r199_c215 bl_215 br_215 wl_199 vdd gnd cell_6t
Xbit_r200_c215 bl_215 br_215 wl_200 vdd gnd cell_6t
Xbit_r201_c215 bl_215 br_215 wl_201 vdd gnd cell_6t
Xbit_r202_c215 bl_215 br_215 wl_202 vdd gnd cell_6t
Xbit_r203_c215 bl_215 br_215 wl_203 vdd gnd cell_6t
Xbit_r204_c215 bl_215 br_215 wl_204 vdd gnd cell_6t
Xbit_r205_c215 bl_215 br_215 wl_205 vdd gnd cell_6t
Xbit_r206_c215 bl_215 br_215 wl_206 vdd gnd cell_6t
Xbit_r207_c215 bl_215 br_215 wl_207 vdd gnd cell_6t
Xbit_r208_c215 bl_215 br_215 wl_208 vdd gnd cell_6t
Xbit_r209_c215 bl_215 br_215 wl_209 vdd gnd cell_6t
Xbit_r210_c215 bl_215 br_215 wl_210 vdd gnd cell_6t
Xbit_r211_c215 bl_215 br_215 wl_211 vdd gnd cell_6t
Xbit_r212_c215 bl_215 br_215 wl_212 vdd gnd cell_6t
Xbit_r213_c215 bl_215 br_215 wl_213 vdd gnd cell_6t
Xbit_r214_c215 bl_215 br_215 wl_214 vdd gnd cell_6t
Xbit_r215_c215 bl_215 br_215 wl_215 vdd gnd cell_6t
Xbit_r216_c215 bl_215 br_215 wl_216 vdd gnd cell_6t
Xbit_r217_c215 bl_215 br_215 wl_217 vdd gnd cell_6t
Xbit_r218_c215 bl_215 br_215 wl_218 vdd gnd cell_6t
Xbit_r219_c215 bl_215 br_215 wl_219 vdd gnd cell_6t
Xbit_r220_c215 bl_215 br_215 wl_220 vdd gnd cell_6t
Xbit_r221_c215 bl_215 br_215 wl_221 vdd gnd cell_6t
Xbit_r222_c215 bl_215 br_215 wl_222 vdd gnd cell_6t
Xbit_r223_c215 bl_215 br_215 wl_223 vdd gnd cell_6t
Xbit_r224_c215 bl_215 br_215 wl_224 vdd gnd cell_6t
Xbit_r225_c215 bl_215 br_215 wl_225 vdd gnd cell_6t
Xbit_r226_c215 bl_215 br_215 wl_226 vdd gnd cell_6t
Xbit_r227_c215 bl_215 br_215 wl_227 vdd gnd cell_6t
Xbit_r228_c215 bl_215 br_215 wl_228 vdd gnd cell_6t
Xbit_r229_c215 bl_215 br_215 wl_229 vdd gnd cell_6t
Xbit_r230_c215 bl_215 br_215 wl_230 vdd gnd cell_6t
Xbit_r231_c215 bl_215 br_215 wl_231 vdd gnd cell_6t
Xbit_r232_c215 bl_215 br_215 wl_232 vdd gnd cell_6t
Xbit_r233_c215 bl_215 br_215 wl_233 vdd gnd cell_6t
Xbit_r234_c215 bl_215 br_215 wl_234 vdd gnd cell_6t
Xbit_r235_c215 bl_215 br_215 wl_235 vdd gnd cell_6t
Xbit_r236_c215 bl_215 br_215 wl_236 vdd gnd cell_6t
Xbit_r237_c215 bl_215 br_215 wl_237 vdd gnd cell_6t
Xbit_r238_c215 bl_215 br_215 wl_238 vdd gnd cell_6t
Xbit_r239_c215 bl_215 br_215 wl_239 vdd gnd cell_6t
Xbit_r240_c215 bl_215 br_215 wl_240 vdd gnd cell_6t
Xbit_r241_c215 bl_215 br_215 wl_241 vdd gnd cell_6t
Xbit_r242_c215 bl_215 br_215 wl_242 vdd gnd cell_6t
Xbit_r243_c215 bl_215 br_215 wl_243 vdd gnd cell_6t
Xbit_r244_c215 bl_215 br_215 wl_244 vdd gnd cell_6t
Xbit_r245_c215 bl_215 br_215 wl_245 vdd gnd cell_6t
Xbit_r246_c215 bl_215 br_215 wl_246 vdd gnd cell_6t
Xbit_r247_c215 bl_215 br_215 wl_247 vdd gnd cell_6t
Xbit_r248_c215 bl_215 br_215 wl_248 vdd gnd cell_6t
Xbit_r249_c215 bl_215 br_215 wl_249 vdd gnd cell_6t
Xbit_r250_c215 bl_215 br_215 wl_250 vdd gnd cell_6t
Xbit_r251_c215 bl_215 br_215 wl_251 vdd gnd cell_6t
Xbit_r252_c215 bl_215 br_215 wl_252 vdd gnd cell_6t
Xbit_r253_c215 bl_215 br_215 wl_253 vdd gnd cell_6t
Xbit_r254_c215 bl_215 br_215 wl_254 vdd gnd cell_6t
Xbit_r255_c215 bl_215 br_215 wl_255 vdd gnd cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd cell_6t
Xbit_r1_c216 bl_216 br_216 wl_1 vdd gnd cell_6t
Xbit_r2_c216 bl_216 br_216 wl_2 vdd gnd cell_6t
Xbit_r3_c216 bl_216 br_216 wl_3 vdd gnd cell_6t
Xbit_r4_c216 bl_216 br_216 wl_4 vdd gnd cell_6t
Xbit_r5_c216 bl_216 br_216 wl_5 vdd gnd cell_6t
Xbit_r6_c216 bl_216 br_216 wl_6 vdd gnd cell_6t
Xbit_r7_c216 bl_216 br_216 wl_7 vdd gnd cell_6t
Xbit_r8_c216 bl_216 br_216 wl_8 vdd gnd cell_6t
Xbit_r9_c216 bl_216 br_216 wl_9 vdd gnd cell_6t
Xbit_r10_c216 bl_216 br_216 wl_10 vdd gnd cell_6t
Xbit_r11_c216 bl_216 br_216 wl_11 vdd gnd cell_6t
Xbit_r12_c216 bl_216 br_216 wl_12 vdd gnd cell_6t
Xbit_r13_c216 bl_216 br_216 wl_13 vdd gnd cell_6t
Xbit_r14_c216 bl_216 br_216 wl_14 vdd gnd cell_6t
Xbit_r15_c216 bl_216 br_216 wl_15 vdd gnd cell_6t
Xbit_r16_c216 bl_216 br_216 wl_16 vdd gnd cell_6t
Xbit_r17_c216 bl_216 br_216 wl_17 vdd gnd cell_6t
Xbit_r18_c216 bl_216 br_216 wl_18 vdd gnd cell_6t
Xbit_r19_c216 bl_216 br_216 wl_19 vdd gnd cell_6t
Xbit_r20_c216 bl_216 br_216 wl_20 vdd gnd cell_6t
Xbit_r21_c216 bl_216 br_216 wl_21 vdd gnd cell_6t
Xbit_r22_c216 bl_216 br_216 wl_22 vdd gnd cell_6t
Xbit_r23_c216 bl_216 br_216 wl_23 vdd gnd cell_6t
Xbit_r24_c216 bl_216 br_216 wl_24 vdd gnd cell_6t
Xbit_r25_c216 bl_216 br_216 wl_25 vdd gnd cell_6t
Xbit_r26_c216 bl_216 br_216 wl_26 vdd gnd cell_6t
Xbit_r27_c216 bl_216 br_216 wl_27 vdd gnd cell_6t
Xbit_r28_c216 bl_216 br_216 wl_28 vdd gnd cell_6t
Xbit_r29_c216 bl_216 br_216 wl_29 vdd gnd cell_6t
Xbit_r30_c216 bl_216 br_216 wl_30 vdd gnd cell_6t
Xbit_r31_c216 bl_216 br_216 wl_31 vdd gnd cell_6t
Xbit_r32_c216 bl_216 br_216 wl_32 vdd gnd cell_6t
Xbit_r33_c216 bl_216 br_216 wl_33 vdd gnd cell_6t
Xbit_r34_c216 bl_216 br_216 wl_34 vdd gnd cell_6t
Xbit_r35_c216 bl_216 br_216 wl_35 vdd gnd cell_6t
Xbit_r36_c216 bl_216 br_216 wl_36 vdd gnd cell_6t
Xbit_r37_c216 bl_216 br_216 wl_37 vdd gnd cell_6t
Xbit_r38_c216 bl_216 br_216 wl_38 vdd gnd cell_6t
Xbit_r39_c216 bl_216 br_216 wl_39 vdd gnd cell_6t
Xbit_r40_c216 bl_216 br_216 wl_40 vdd gnd cell_6t
Xbit_r41_c216 bl_216 br_216 wl_41 vdd gnd cell_6t
Xbit_r42_c216 bl_216 br_216 wl_42 vdd gnd cell_6t
Xbit_r43_c216 bl_216 br_216 wl_43 vdd gnd cell_6t
Xbit_r44_c216 bl_216 br_216 wl_44 vdd gnd cell_6t
Xbit_r45_c216 bl_216 br_216 wl_45 vdd gnd cell_6t
Xbit_r46_c216 bl_216 br_216 wl_46 vdd gnd cell_6t
Xbit_r47_c216 bl_216 br_216 wl_47 vdd gnd cell_6t
Xbit_r48_c216 bl_216 br_216 wl_48 vdd gnd cell_6t
Xbit_r49_c216 bl_216 br_216 wl_49 vdd gnd cell_6t
Xbit_r50_c216 bl_216 br_216 wl_50 vdd gnd cell_6t
Xbit_r51_c216 bl_216 br_216 wl_51 vdd gnd cell_6t
Xbit_r52_c216 bl_216 br_216 wl_52 vdd gnd cell_6t
Xbit_r53_c216 bl_216 br_216 wl_53 vdd gnd cell_6t
Xbit_r54_c216 bl_216 br_216 wl_54 vdd gnd cell_6t
Xbit_r55_c216 bl_216 br_216 wl_55 vdd gnd cell_6t
Xbit_r56_c216 bl_216 br_216 wl_56 vdd gnd cell_6t
Xbit_r57_c216 bl_216 br_216 wl_57 vdd gnd cell_6t
Xbit_r58_c216 bl_216 br_216 wl_58 vdd gnd cell_6t
Xbit_r59_c216 bl_216 br_216 wl_59 vdd gnd cell_6t
Xbit_r60_c216 bl_216 br_216 wl_60 vdd gnd cell_6t
Xbit_r61_c216 bl_216 br_216 wl_61 vdd gnd cell_6t
Xbit_r62_c216 bl_216 br_216 wl_62 vdd gnd cell_6t
Xbit_r63_c216 bl_216 br_216 wl_63 vdd gnd cell_6t
Xbit_r64_c216 bl_216 br_216 wl_64 vdd gnd cell_6t
Xbit_r65_c216 bl_216 br_216 wl_65 vdd gnd cell_6t
Xbit_r66_c216 bl_216 br_216 wl_66 vdd gnd cell_6t
Xbit_r67_c216 bl_216 br_216 wl_67 vdd gnd cell_6t
Xbit_r68_c216 bl_216 br_216 wl_68 vdd gnd cell_6t
Xbit_r69_c216 bl_216 br_216 wl_69 vdd gnd cell_6t
Xbit_r70_c216 bl_216 br_216 wl_70 vdd gnd cell_6t
Xbit_r71_c216 bl_216 br_216 wl_71 vdd gnd cell_6t
Xbit_r72_c216 bl_216 br_216 wl_72 vdd gnd cell_6t
Xbit_r73_c216 bl_216 br_216 wl_73 vdd gnd cell_6t
Xbit_r74_c216 bl_216 br_216 wl_74 vdd gnd cell_6t
Xbit_r75_c216 bl_216 br_216 wl_75 vdd gnd cell_6t
Xbit_r76_c216 bl_216 br_216 wl_76 vdd gnd cell_6t
Xbit_r77_c216 bl_216 br_216 wl_77 vdd gnd cell_6t
Xbit_r78_c216 bl_216 br_216 wl_78 vdd gnd cell_6t
Xbit_r79_c216 bl_216 br_216 wl_79 vdd gnd cell_6t
Xbit_r80_c216 bl_216 br_216 wl_80 vdd gnd cell_6t
Xbit_r81_c216 bl_216 br_216 wl_81 vdd gnd cell_6t
Xbit_r82_c216 bl_216 br_216 wl_82 vdd gnd cell_6t
Xbit_r83_c216 bl_216 br_216 wl_83 vdd gnd cell_6t
Xbit_r84_c216 bl_216 br_216 wl_84 vdd gnd cell_6t
Xbit_r85_c216 bl_216 br_216 wl_85 vdd gnd cell_6t
Xbit_r86_c216 bl_216 br_216 wl_86 vdd gnd cell_6t
Xbit_r87_c216 bl_216 br_216 wl_87 vdd gnd cell_6t
Xbit_r88_c216 bl_216 br_216 wl_88 vdd gnd cell_6t
Xbit_r89_c216 bl_216 br_216 wl_89 vdd gnd cell_6t
Xbit_r90_c216 bl_216 br_216 wl_90 vdd gnd cell_6t
Xbit_r91_c216 bl_216 br_216 wl_91 vdd gnd cell_6t
Xbit_r92_c216 bl_216 br_216 wl_92 vdd gnd cell_6t
Xbit_r93_c216 bl_216 br_216 wl_93 vdd gnd cell_6t
Xbit_r94_c216 bl_216 br_216 wl_94 vdd gnd cell_6t
Xbit_r95_c216 bl_216 br_216 wl_95 vdd gnd cell_6t
Xbit_r96_c216 bl_216 br_216 wl_96 vdd gnd cell_6t
Xbit_r97_c216 bl_216 br_216 wl_97 vdd gnd cell_6t
Xbit_r98_c216 bl_216 br_216 wl_98 vdd gnd cell_6t
Xbit_r99_c216 bl_216 br_216 wl_99 vdd gnd cell_6t
Xbit_r100_c216 bl_216 br_216 wl_100 vdd gnd cell_6t
Xbit_r101_c216 bl_216 br_216 wl_101 vdd gnd cell_6t
Xbit_r102_c216 bl_216 br_216 wl_102 vdd gnd cell_6t
Xbit_r103_c216 bl_216 br_216 wl_103 vdd gnd cell_6t
Xbit_r104_c216 bl_216 br_216 wl_104 vdd gnd cell_6t
Xbit_r105_c216 bl_216 br_216 wl_105 vdd gnd cell_6t
Xbit_r106_c216 bl_216 br_216 wl_106 vdd gnd cell_6t
Xbit_r107_c216 bl_216 br_216 wl_107 vdd gnd cell_6t
Xbit_r108_c216 bl_216 br_216 wl_108 vdd gnd cell_6t
Xbit_r109_c216 bl_216 br_216 wl_109 vdd gnd cell_6t
Xbit_r110_c216 bl_216 br_216 wl_110 vdd gnd cell_6t
Xbit_r111_c216 bl_216 br_216 wl_111 vdd gnd cell_6t
Xbit_r112_c216 bl_216 br_216 wl_112 vdd gnd cell_6t
Xbit_r113_c216 bl_216 br_216 wl_113 vdd gnd cell_6t
Xbit_r114_c216 bl_216 br_216 wl_114 vdd gnd cell_6t
Xbit_r115_c216 bl_216 br_216 wl_115 vdd gnd cell_6t
Xbit_r116_c216 bl_216 br_216 wl_116 vdd gnd cell_6t
Xbit_r117_c216 bl_216 br_216 wl_117 vdd gnd cell_6t
Xbit_r118_c216 bl_216 br_216 wl_118 vdd gnd cell_6t
Xbit_r119_c216 bl_216 br_216 wl_119 vdd gnd cell_6t
Xbit_r120_c216 bl_216 br_216 wl_120 vdd gnd cell_6t
Xbit_r121_c216 bl_216 br_216 wl_121 vdd gnd cell_6t
Xbit_r122_c216 bl_216 br_216 wl_122 vdd gnd cell_6t
Xbit_r123_c216 bl_216 br_216 wl_123 vdd gnd cell_6t
Xbit_r124_c216 bl_216 br_216 wl_124 vdd gnd cell_6t
Xbit_r125_c216 bl_216 br_216 wl_125 vdd gnd cell_6t
Xbit_r126_c216 bl_216 br_216 wl_126 vdd gnd cell_6t
Xbit_r127_c216 bl_216 br_216 wl_127 vdd gnd cell_6t
Xbit_r128_c216 bl_216 br_216 wl_128 vdd gnd cell_6t
Xbit_r129_c216 bl_216 br_216 wl_129 vdd gnd cell_6t
Xbit_r130_c216 bl_216 br_216 wl_130 vdd gnd cell_6t
Xbit_r131_c216 bl_216 br_216 wl_131 vdd gnd cell_6t
Xbit_r132_c216 bl_216 br_216 wl_132 vdd gnd cell_6t
Xbit_r133_c216 bl_216 br_216 wl_133 vdd gnd cell_6t
Xbit_r134_c216 bl_216 br_216 wl_134 vdd gnd cell_6t
Xbit_r135_c216 bl_216 br_216 wl_135 vdd gnd cell_6t
Xbit_r136_c216 bl_216 br_216 wl_136 vdd gnd cell_6t
Xbit_r137_c216 bl_216 br_216 wl_137 vdd gnd cell_6t
Xbit_r138_c216 bl_216 br_216 wl_138 vdd gnd cell_6t
Xbit_r139_c216 bl_216 br_216 wl_139 vdd gnd cell_6t
Xbit_r140_c216 bl_216 br_216 wl_140 vdd gnd cell_6t
Xbit_r141_c216 bl_216 br_216 wl_141 vdd gnd cell_6t
Xbit_r142_c216 bl_216 br_216 wl_142 vdd gnd cell_6t
Xbit_r143_c216 bl_216 br_216 wl_143 vdd gnd cell_6t
Xbit_r144_c216 bl_216 br_216 wl_144 vdd gnd cell_6t
Xbit_r145_c216 bl_216 br_216 wl_145 vdd gnd cell_6t
Xbit_r146_c216 bl_216 br_216 wl_146 vdd gnd cell_6t
Xbit_r147_c216 bl_216 br_216 wl_147 vdd gnd cell_6t
Xbit_r148_c216 bl_216 br_216 wl_148 vdd gnd cell_6t
Xbit_r149_c216 bl_216 br_216 wl_149 vdd gnd cell_6t
Xbit_r150_c216 bl_216 br_216 wl_150 vdd gnd cell_6t
Xbit_r151_c216 bl_216 br_216 wl_151 vdd gnd cell_6t
Xbit_r152_c216 bl_216 br_216 wl_152 vdd gnd cell_6t
Xbit_r153_c216 bl_216 br_216 wl_153 vdd gnd cell_6t
Xbit_r154_c216 bl_216 br_216 wl_154 vdd gnd cell_6t
Xbit_r155_c216 bl_216 br_216 wl_155 vdd gnd cell_6t
Xbit_r156_c216 bl_216 br_216 wl_156 vdd gnd cell_6t
Xbit_r157_c216 bl_216 br_216 wl_157 vdd gnd cell_6t
Xbit_r158_c216 bl_216 br_216 wl_158 vdd gnd cell_6t
Xbit_r159_c216 bl_216 br_216 wl_159 vdd gnd cell_6t
Xbit_r160_c216 bl_216 br_216 wl_160 vdd gnd cell_6t
Xbit_r161_c216 bl_216 br_216 wl_161 vdd gnd cell_6t
Xbit_r162_c216 bl_216 br_216 wl_162 vdd gnd cell_6t
Xbit_r163_c216 bl_216 br_216 wl_163 vdd gnd cell_6t
Xbit_r164_c216 bl_216 br_216 wl_164 vdd gnd cell_6t
Xbit_r165_c216 bl_216 br_216 wl_165 vdd gnd cell_6t
Xbit_r166_c216 bl_216 br_216 wl_166 vdd gnd cell_6t
Xbit_r167_c216 bl_216 br_216 wl_167 vdd gnd cell_6t
Xbit_r168_c216 bl_216 br_216 wl_168 vdd gnd cell_6t
Xbit_r169_c216 bl_216 br_216 wl_169 vdd gnd cell_6t
Xbit_r170_c216 bl_216 br_216 wl_170 vdd gnd cell_6t
Xbit_r171_c216 bl_216 br_216 wl_171 vdd gnd cell_6t
Xbit_r172_c216 bl_216 br_216 wl_172 vdd gnd cell_6t
Xbit_r173_c216 bl_216 br_216 wl_173 vdd gnd cell_6t
Xbit_r174_c216 bl_216 br_216 wl_174 vdd gnd cell_6t
Xbit_r175_c216 bl_216 br_216 wl_175 vdd gnd cell_6t
Xbit_r176_c216 bl_216 br_216 wl_176 vdd gnd cell_6t
Xbit_r177_c216 bl_216 br_216 wl_177 vdd gnd cell_6t
Xbit_r178_c216 bl_216 br_216 wl_178 vdd gnd cell_6t
Xbit_r179_c216 bl_216 br_216 wl_179 vdd gnd cell_6t
Xbit_r180_c216 bl_216 br_216 wl_180 vdd gnd cell_6t
Xbit_r181_c216 bl_216 br_216 wl_181 vdd gnd cell_6t
Xbit_r182_c216 bl_216 br_216 wl_182 vdd gnd cell_6t
Xbit_r183_c216 bl_216 br_216 wl_183 vdd gnd cell_6t
Xbit_r184_c216 bl_216 br_216 wl_184 vdd gnd cell_6t
Xbit_r185_c216 bl_216 br_216 wl_185 vdd gnd cell_6t
Xbit_r186_c216 bl_216 br_216 wl_186 vdd gnd cell_6t
Xbit_r187_c216 bl_216 br_216 wl_187 vdd gnd cell_6t
Xbit_r188_c216 bl_216 br_216 wl_188 vdd gnd cell_6t
Xbit_r189_c216 bl_216 br_216 wl_189 vdd gnd cell_6t
Xbit_r190_c216 bl_216 br_216 wl_190 vdd gnd cell_6t
Xbit_r191_c216 bl_216 br_216 wl_191 vdd gnd cell_6t
Xbit_r192_c216 bl_216 br_216 wl_192 vdd gnd cell_6t
Xbit_r193_c216 bl_216 br_216 wl_193 vdd gnd cell_6t
Xbit_r194_c216 bl_216 br_216 wl_194 vdd gnd cell_6t
Xbit_r195_c216 bl_216 br_216 wl_195 vdd gnd cell_6t
Xbit_r196_c216 bl_216 br_216 wl_196 vdd gnd cell_6t
Xbit_r197_c216 bl_216 br_216 wl_197 vdd gnd cell_6t
Xbit_r198_c216 bl_216 br_216 wl_198 vdd gnd cell_6t
Xbit_r199_c216 bl_216 br_216 wl_199 vdd gnd cell_6t
Xbit_r200_c216 bl_216 br_216 wl_200 vdd gnd cell_6t
Xbit_r201_c216 bl_216 br_216 wl_201 vdd gnd cell_6t
Xbit_r202_c216 bl_216 br_216 wl_202 vdd gnd cell_6t
Xbit_r203_c216 bl_216 br_216 wl_203 vdd gnd cell_6t
Xbit_r204_c216 bl_216 br_216 wl_204 vdd gnd cell_6t
Xbit_r205_c216 bl_216 br_216 wl_205 vdd gnd cell_6t
Xbit_r206_c216 bl_216 br_216 wl_206 vdd gnd cell_6t
Xbit_r207_c216 bl_216 br_216 wl_207 vdd gnd cell_6t
Xbit_r208_c216 bl_216 br_216 wl_208 vdd gnd cell_6t
Xbit_r209_c216 bl_216 br_216 wl_209 vdd gnd cell_6t
Xbit_r210_c216 bl_216 br_216 wl_210 vdd gnd cell_6t
Xbit_r211_c216 bl_216 br_216 wl_211 vdd gnd cell_6t
Xbit_r212_c216 bl_216 br_216 wl_212 vdd gnd cell_6t
Xbit_r213_c216 bl_216 br_216 wl_213 vdd gnd cell_6t
Xbit_r214_c216 bl_216 br_216 wl_214 vdd gnd cell_6t
Xbit_r215_c216 bl_216 br_216 wl_215 vdd gnd cell_6t
Xbit_r216_c216 bl_216 br_216 wl_216 vdd gnd cell_6t
Xbit_r217_c216 bl_216 br_216 wl_217 vdd gnd cell_6t
Xbit_r218_c216 bl_216 br_216 wl_218 vdd gnd cell_6t
Xbit_r219_c216 bl_216 br_216 wl_219 vdd gnd cell_6t
Xbit_r220_c216 bl_216 br_216 wl_220 vdd gnd cell_6t
Xbit_r221_c216 bl_216 br_216 wl_221 vdd gnd cell_6t
Xbit_r222_c216 bl_216 br_216 wl_222 vdd gnd cell_6t
Xbit_r223_c216 bl_216 br_216 wl_223 vdd gnd cell_6t
Xbit_r224_c216 bl_216 br_216 wl_224 vdd gnd cell_6t
Xbit_r225_c216 bl_216 br_216 wl_225 vdd gnd cell_6t
Xbit_r226_c216 bl_216 br_216 wl_226 vdd gnd cell_6t
Xbit_r227_c216 bl_216 br_216 wl_227 vdd gnd cell_6t
Xbit_r228_c216 bl_216 br_216 wl_228 vdd gnd cell_6t
Xbit_r229_c216 bl_216 br_216 wl_229 vdd gnd cell_6t
Xbit_r230_c216 bl_216 br_216 wl_230 vdd gnd cell_6t
Xbit_r231_c216 bl_216 br_216 wl_231 vdd gnd cell_6t
Xbit_r232_c216 bl_216 br_216 wl_232 vdd gnd cell_6t
Xbit_r233_c216 bl_216 br_216 wl_233 vdd gnd cell_6t
Xbit_r234_c216 bl_216 br_216 wl_234 vdd gnd cell_6t
Xbit_r235_c216 bl_216 br_216 wl_235 vdd gnd cell_6t
Xbit_r236_c216 bl_216 br_216 wl_236 vdd gnd cell_6t
Xbit_r237_c216 bl_216 br_216 wl_237 vdd gnd cell_6t
Xbit_r238_c216 bl_216 br_216 wl_238 vdd gnd cell_6t
Xbit_r239_c216 bl_216 br_216 wl_239 vdd gnd cell_6t
Xbit_r240_c216 bl_216 br_216 wl_240 vdd gnd cell_6t
Xbit_r241_c216 bl_216 br_216 wl_241 vdd gnd cell_6t
Xbit_r242_c216 bl_216 br_216 wl_242 vdd gnd cell_6t
Xbit_r243_c216 bl_216 br_216 wl_243 vdd gnd cell_6t
Xbit_r244_c216 bl_216 br_216 wl_244 vdd gnd cell_6t
Xbit_r245_c216 bl_216 br_216 wl_245 vdd gnd cell_6t
Xbit_r246_c216 bl_216 br_216 wl_246 vdd gnd cell_6t
Xbit_r247_c216 bl_216 br_216 wl_247 vdd gnd cell_6t
Xbit_r248_c216 bl_216 br_216 wl_248 vdd gnd cell_6t
Xbit_r249_c216 bl_216 br_216 wl_249 vdd gnd cell_6t
Xbit_r250_c216 bl_216 br_216 wl_250 vdd gnd cell_6t
Xbit_r251_c216 bl_216 br_216 wl_251 vdd gnd cell_6t
Xbit_r252_c216 bl_216 br_216 wl_252 vdd gnd cell_6t
Xbit_r253_c216 bl_216 br_216 wl_253 vdd gnd cell_6t
Xbit_r254_c216 bl_216 br_216 wl_254 vdd gnd cell_6t
Xbit_r255_c216 bl_216 br_216 wl_255 vdd gnd cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd cell_6t
Xbit_r1_c217 bl_217 br_217 wl_1 vdd gnd cell_6t
Xbit_r2_c217 bl_217 br_217 wl_2 vdd gnd cell_6t
Xbit_r3_c217 bl_217 br_217 wl_3 vdd gnd cell_6t
Xbit_r4_c217 bl_217 br_217 wl_4 vdd gnd cell_6t
Xbit_r5_c217 bl_217 br_217 wl_5 vdd gnd cell_6t
Xbit_r6_c217 bl_217 br_217 wl_6 vdd gnd cell_6t
Xbit_r7_c217 bl_217 br_217 wl_7 vdd gnd cell_6t
Xbit_r8_c217 bl_217 br_217 wl_8 vdd gnd cell_6t
Xbit_r9_c217 bl_217 br_217 wl_9 vdd gnd cell_6t
Xbit_r10_c217 bl_217 br_217 wl_10 vdd gnd cell_6t
Xbit_r11_c217 bl_217 br_217 wl_11 vdd gnd cell_6t
Xbit_r12_c217 bl_217 br_217 wl_12 vdd gnd cell_6t
Xbit_r13_c217 bl_217 br_217 wl_13 vdd gnd cell_6t
Xbit_r14_c217 bl_217 br_217 wl_14 vdd gnd cell_6t
Xbit_r15_c217 bl_217 br_217 wl_15 vdd gnd cell_6t
Xbit_r16_c217 bl_217 br_217 wl_16 vdd gnd cell_6t
Xbit_r17_c217 bl_217 br_217 wl_17 vdd gnd cell_6t
Xbit_r18_c217 bl_217 br_217 wl_18 vdd gnd cell_6t
Xbit_r19_c217 bl_217 br_217 wl_19 vdd gnd cell_6t
Xbit_r20_c217 bl_217 br_217 wl_20 vdd gnd cell_6t
Xbit_r21_c217 bl_217 br_217 wl_21 vdd gnd cell_6t
Xbit_r22_c217 bl_217 br_217 wl_22 vdd gnd cell_6t
Xbit_r23_c217 bl_217 br_217 wl_23 vdd gnd cell_6t
Xbit_r24_c217 bl_217 br_217 wl_24 vdd gnd cell_6t
Xbit_r25_c217 bl_217 br_217 wl_25 vdd gnd cell_6t
Xbit_r26_c217 bl_217 br_217 wl_26 vdd gnd cell_6t
Xbit_r27_c217 bl_217 br_217 wl_27 vdd gnd cell_6t
Xbit_r28_c217 bl_217 br_217 wl_28 vdd gnd cell_6t
Xbit_r29_c217 bl_217 br_217 wl_29 vdd gnd cell_6t
Xbit_r30_c217 bl_217 br_217 wl_30 vdd gnd cell_6t
Xbit_r31_c217 bl_217 br_217 wl_31 vdd gnd cell_6t
Xbit_r32_c217 bl_217 br_217 wl_32 vdd gnd cell_6t
Xbit_r33_c217 bl_217 br_217 wl_33 vdd gnd cell_6t
Xbit_r34_c217 bl_217 br_217 wl_34 vdd gnd cell_6t
Xbit_r35_c217 bl_217 br_217 wl_35 vdd gnd cell_6t
Xbit_r36_c217 bl_217 br_217 wl_36 vdd gnd cell_6t
Xbit_r37_c217 bl_217 br_217 wl_37 vdd gnd cell_6t
Xbit_r38_c217 bl_217 br_217 wl_38 vdd gnd cell_6t
Xbit_r39_c217 bl_217 br_217 wl_39 vdd gnd cell_6t
Xbit_r40_c217 bl_217 br_217 wl_40 vdd gnd cell_6t
Xbit_r41_c217 bl_217 br_217 wl_41 vdd gnd cell_6t
Xbit_r42_c217 bl_217 br_217 wl_42 vdd gnd cell_6t
Xbit_r43_c217 bl_217 br_217 wl_43 vdd gnd cell_6t
Xbit_r44_c217 bl_217 br_217 wl_44 vdd gnd cell_6t
Xbit_r45_c217 bl_217 br_217 wl_45 vdd gnd cell_6t
Xbit_r46_c217 bl_217 br_217 wl_46 vdd gnd cell_6t
Xbit_r47_c217 bl_217 br_217 wl_47 vdd gnd cell_6t
Xbit_r48_c217 bl_217 br_217 wl_48 vdd gnd cell_6t
Xbit_r49_c217 bl_217 br_217 wl_49 vdd gnd cell_6t
Xbit_r50_c217 bl_217 br_217 wl_50 vdd gnd cell_6t
Xbit_r51_c217 bl_217 br_217 wl_51 vdd gnd cell_6t
Xbit_r52_c217 bl_217 br_217 wl_52 vdd gnd cell_6t
Xbit_r53_c217 bl_217 br_217 wl_53 vdd gnd cell_6t
Xbit_r54_c217 bl_217 br_217 wl_54 vdd gnd cell_6t
Xbit_r55_c217 bl_217 br_217 wl_55 vdd gnd cell_6t
Xbit_r56_c217 bl_217 br_217 wl_56 vdd gnd cell_6t
Xbit_r57_c217 bl_217 br_217 wl_57 vdd gnd cell_6t
Xbit_r58_c217 bl_217 br_217 wl_58 vdd gnd cell_6t
Xbit_r59_c217 bl_217 br_217 wl_59 vdd gnd cell_6t
Xbit_r60_c217 bl_217 br_217 wl_60 vdd gnd cell_6t
Xbit_r61_c217 bl_217 br_217 wl_61 vdd gnd cell_6t
Xbit_r62_c217 bl_217 br_217 wl_62 vdd gnd cell_6t
Xbit_r63_c217 bl_217 br_217 wl_63 vdd gnd cell_6t
Xbit_r64_c217 bl_217 br_217 wl_64 vdd gnd cell_6t
Xbit_r65_c217 bl_217 br_217 wl_65 vdd gnd cell_6t
Xbit_r66_c217 bl_217 br_217 wl_66 vdd gnd cell_6t
Xbit_r67_c217 bl_217 br_217 wl_67 vdd gnd cell_6t
Xbit_r68_c217 bl_217 br_217 wl_68 vdd gnd cell_6t
Xbit_r69_c217 bl_217 br_217 wl_69 vdd gnd cell_6t
Xbit_r70_c217 bl_217 br_217 wl_70 vdd gnd cell_6t
Xbit_r71_c217 bl_217 br_217 wl_71 vdd gnd cell_6t
Xbit_r72_c217 bl_217 br_217 wl_72 vdd gnd cell_6t
Xbit_r73_c217 bl_217 br_217 wl_73 vdd gnd cell_6t
Xbit_r74_c217 bl_217 br_217 wl_74 vdd gnd cell_6t
Xbit_r75_c217 bl_217 br_217 wl_75 vdd gnd cell_6t
Xbit_r76_c217 bl_217 br_217 wl_76 vdd gnd cell_6t
Xbit_r77_c217 bl_217 br_217 wl_77 vdd gnd cell_6t
Xbit_r78_c217 bl_217 br_217 wl_78 vdd gnd cell_6t
Xbit_r79_c217 bl_217 br_217 wl_79 vdd gnd cell_6t
Xbit_r80_c217 bl_217 br_217 wl_80 vdd gnd cell_6t
Xbit_r81_c217 bl_217 br_217 wl_81 vdd gnd cell_6t
Xbit_r82_c217 bl_217 br_217 wl_82 vdd gnd cell_6t
Xbit_r83_c217 bl_217 br_217 wl_83 vdd gnd cell_6t
Xbit_r84_c217 bl_217 br_217 wl_84 vdd gnd cell_6t
Xbit_r85_c217 bl_217 br_217 wl_85 vdd gnd cell_6t
Xbit_r86_c217 bl_217 br_217 wl_86 vdd gnd cell_6t
Xbit_r87_c217 bl_217 br_217 wl_87 vdd gnd cell_6t
Xbit_r88_c217 bl_217 br_217 wl_88 vdd gnd cell_6t
Xbit_r89_c217 bl_217 br_217 wl_89 vdd gnd cell_6t
Xbit_r90_c217 bl_217 br_217 wl_90 vdd gnd cell_6t
Xbit_r91_c217 bl_217 br_217 wl_91 vdd gnd cell_6t
Xbit_r92_c217 bl_217 br_217 wl_92 vdd gnd cell_6t
Xbit_r93_c217 bl_217 br_217 wl_93 vdd gnd cell_6t
Xbit_r94_c217 bl_217 br_217 wl_94 vdd gnd cell_6t
Xbit_r95_c217 bl_217 br_217 wl_95 vdd gnd cell_6t
Xbit_r96_c217 bl_217 br_217 wl_96 vdd gnd cell_6t
Xbit_r97_c217 bl_217 br_217 wl_97 vdd gnd cell_6t
Xbit_r98_c217 bl_217 br_217 wl_98 vdd gnd cell_6t
Xbit_r99_c217 bl_217 br_217 wl_99 vdd gnd cell_6t
Xbit_r100_c217 bl_217 br_217 wl_100 vdd gnd cell_6t
Xbit_r101_c217 bl_217 br_217 wl_101 vdd gnd cell_6t
Xbit_r102_c217 bl_217 br_217 wl_102 vdd gnd cell_6t
Xbit_r103_c217 bl_217 br_217 wl_103 vdd gnd cell_6t
Xbit_r104_c217 bl_217 br_217 wl_104 vdd gnd cell_6t
Xbit_r105_c217 bl_217 br_217 wl_105 vdd gnd cell_6t
Xbit_r106_c217 bl_217 br_217 wl_106 vdd gnd cell_6t
Xbit_r107_c217 bl_217 br_217 wl_107 vdd gnd cell_6t
Xbit_r108_c217 bl_217 br_217 wl_108 vdd gnd cell_6t
Xbit_r109_c217 bl_217 br_217 wl_109 vdd gnd cell_6t
Xbit_r110_c217 bl_217 br_217 wl_110 vdd gnd cell_6t
Xbit_r111_c217 bl_217 br_217 wl_111 vdd gnd cell_6t
Xbit_r112_c217 bl_217 br_217 wl_112 vdd gnd cell_6t
Xbit_r113_c217 bl_217 br_217 wl_113 vdd gnd cell_6t
Xbit_r114_c217 bl_217 br_217 wl_114 vdd gnd cell_6t
Xbit_r115_c217 bl_217 br_217 wl_115 vdd gnd cell_6t
Xbit_r116_c217 bl_217 br_217 wl_116 vdd gnd cell_6t
Xbit_r117_c217 bl_217 br_217 wl_117 vdd gnd cell_6t
Xbit_r118_c217 bl_217 br_217 wl_118 vdd gnd cell_6t
Xbit_r119_c217 bl_217 br_217 wl_119 vdd gnd cell_6t
Xbit_r120_c217 bl_217 br_217 wl_120 vdd gnd cell_6t
Xbit_r121_c217 bl_217 br_217 wl_121 vdd gnd cell_6t
Xbit_r122_c217 bl_217 br_217 wl_122 vdd gnd cell_6t
Xbit_r123_c217 bl_217 br_217 wl_123 vdd gnd cell_6t
Xbit_r124_c217 bl_217 br_217 wl_124 vdd gnd cell_6t
Xbit_r125_c217 bl_217 br_217 wl_125 vdd gnd cell_6t
Xbit_r126_c217 bl_217 br_217 wl_126 vdd gnd cell_6t
Xbit_r127_c217 bl_217 br_217 wl_127 vdd gnd cell_6t
Xbit_r128_c217 bl_217 br_217 wl_128 vdd gnd cell_6t
Xbit_r129_c217 bl_217 br_217 wl_129 vdd gnd cell_6t
Xbit_r130_c217 bl_217 br_217 wl_130 vdd gnd cell_6t
Xbit_r131_c217 bl_217 br_217 wl_131 vdd gnd cell_6t
Xbit_r132_c217 bl_217 br_217 wl_132 vdd gnd cell_6t
Xbit_r133_c217 bl_217 br_217 wl_133 vdd gnd cell_6t
Xbit_r134_c217 bl_217 br_217 wl_134 vdd gnd cell_6t
Xbit_r135_c217 bl_217 br_217 wl_135 vdd gnd cell_6t
Xbit_r136_c217 bl_217 br_217 wl_136 vdd gnd cell_6t
Xbit_r137_c217 bl_217 br_217 wl_137 vdd gnd cell_6t
Xbit_r138_c217 bl_217 br_217 wl_138 vdd gnd cell_6t
Xbit_r139_c217 bl_217 br_217 wl_139 vdd gnd cell_6t
Xbit_r140_c217 bl_217 br_217 wl_140 vdd gnd cell_6t
Xbit_r141_c217 bl_217 br_217 wl_141 vdd gnd cell_6t
Xbit_r142_c217 bl_217 br_217 wl_142 vdd gnd cell_6t
Xbit_r143_c217 bl_217 br_217 wl_143 vdd gnd cell_6t
Xbit_r144_c217 bl_217 br_217 wl_144 vdd gnd cell_6t
Xbit_r145_c217 bl_217 br_217 wl_145 vdd gnd cell_6t
Xbit_r146_c217 bl_217 br_217 wl_146 vdd gnd cell_6t
Xbit_r147_c217 bl_217 br_217 wl_147 vdd gnd cell_6t
Xbit_r148_c217 bl_217 br_217 wl_148 vdd gnd cell_6t
Xbit_r149_c217 bl_217 br_217 wl_149 vdd gnd cell_6t
Xbit_r150_c217 bl_217 br_217 wl_150 vdd gnd cell_6t
Xbit_r151_c217 bl_217 br_217 wl_151 vdd gnd cell_6t
Xbit_r152_c217 bl_217 br_217 wl_152 vdd gnd cell_6t
Xbit_r153_c217 bl_217 br_217 wl_153 vdd gnd cell_6t
Xbit_r154_c217 bl_217 br_217 wl_154 vdd gnd cell_6t
Xbit_r155_c217 bl_217 br_217 wl_155 vdd gnd cell_6t
Xbit_r156_c217 bl_217 br_217 wl_156 vdd gnd cell_6t
Xbit_r157_c217 bl_217 br_217 wl_157 vdd gnd cell_6t
Xbit_r158_c217 bl_217 br_217 wl_158 vdd gnd cell_6t
Xbit_r159_c217 bl_217 br_217 wl_159 vdd gnd cell_6t
Xbit_r160_c217 bl_217 br_217 wl_160 vdd gnd cell_6t
Xbit_r161_c217 bl_217 br_217 wl_161 vdd gnd cell_6t
Xbit_r162_c217 bl_217 br_217 wl_162 vdd gnd cell_6t
Xbit_r163_c217 bl_217 br_217 wl_163 vdd gnd cell_6t
Xbit_r164_c217 bl_217 br_217 wl_164 vdd gnd cell_6t
Xbit_r165_c217 bl_217 br_217 wl_165 vdd gnd cell_6t
Xbit_r166_c217 bl_217 br_217 wl_166 vdd gnd cell_6t
Xbit_r167_c217 bl_217 br_217 wl_167 vdd gnd cell_6t
Xbit_r168_c217 bl_217 br_217 wl_168 vdd gnd cell_6t
Xbit_r169_c217 bl_217 br_217 wl_169 vdd gnd cell_6t
Xbit_r170_c217 bl_217 br_217 wl_170 vdd gnd cell_6t
Xbit_r171_c217 bl_217 br_217 wl_171 vdd gnd cell_6t
Xbit_r172_c217 bl_217 br_217 wl_172 vdd gnd cell_6t
Xbit_r173_c217 bl_217 br_217 wl_173 vdd gnd cell_6t
Xbit_r174_c217 bl_217 br_217 wl_174 vdd gnd cell_6t
Xbit_r175_c217 bl_217 br_217 wl_175 vdd gnd cell_6t
Xbit_r176_c217 bl_217 br_217 wl_176 vdd gnd cell_6t
Xbit_r177_c217 bl_217 br_217 wl_177 vdd gnd cell_6t
Xbit_r178_c217 bl_217 br_217 wl_178 vdd gnd cell_6t
Xbit_r179_c217 bl_217 br_217 wl_179 vdd gnd cell_6t
Xbit_r180_c217 bl_217 br_217 wl_180 vdd gnd cell_6t
Xbit_r181_c217 bl_217 br_217 wl_181 vdd gnd cell_6t
Xbit_r182_c217 bl_217 br_217 wl_182 vdd gnd cell_6t
Xbit_r183_c217 bl_217 br_217 wl_183 vdd gnd cell_6t
Xbit_r184_c217 bl_217 br_217 wl_184 vdd gnd cell_6t
Xbit_r185_c217 bl_217 br_217 wl_185 vdd gnd cell_6t
Xbit_r186_c217 bl_217 br_217 wl_186 vdd gnd cell_6t
Xbit_r187_c217 bl_217 br_217 wl_187 vdd gnd cell_6t
Xbit_r188_c217 bl_217 br_217 wl_188 vdd gnd cell_6t
Xbit_r189_c217 bl_217 br_217 wl_189 vdd gnd cell_6t
Xbit_r190_c217 bl_217 br_217 wl_190 vdd gnd cell_6t
Xbit_r191_c217 bl_217 br_217 wl_191 vdd gnd cell_6t
Xbit_r192_c217 bl_217 br_217 wl_192 vdd gnd cell_6t
Xbit_r193_c217 bl_217 br_217 wl_193 vdd gnd cell_6t
Xbit_r194_c217 bl_217 br_217 wl_194 vdd gnd cell_6t
Xbit_r195_c217 bl_217 br_217 wl_195 vdd gnd cell_6t
Xbit_r196_c217 bl_217 br_217 wl_196 vdd gnd cell_6t
Xbit_r197_c217 bl_217 br_217 wl_197 vdd gnd cell_6t
Xbit_r198_c217 bl_217 br_217 wl_198 vdd gnd cell_6t
Xbit_r199_c217 bl_217 br_217 wl_199 vdd gnd cell_6t
Xbit_r200_c217 bl_217 br_217 wl_200 vdd gnd cell_6t
Xbit_r201_c217 bl_217 br_217 wl_201 vdd gnd cell_6t
Xbit_r202_c217 bl_217 br_217 wl_202 vdd gnd cell_6t
Xbit_r203_c217 bl_217 br_217 wl_203 vdd gnd cell_6t
Xbit_r204_c217 bl_217 br_217 wl_204 vdd gnd cell_6t
Xbit_r205_c217 bl_217 br_217 wl_205 vdd gnd cell_6t
Xbit_r206_c217 bl_217 br_217 wl_206 vdd gnd cell_6t
Xbit_r207_c217 bl_217 br_217 wl_207 vdd gnd cell_6t
Xbit_r208_c217 bl_217 br_217 wl_208 vdd gnd cell_6t
Xbit_r209_c217 bl_217 br_217 wl_209 vdd gnd cell_6t
Xbit_r210_c217 bl_217 br_217 wl_210 vdd gnd cell_6t
Xbit_r211_c217 bl_217 br_217 wl_211 vdd gnd cell_6t
Xbit_r212_c217 bl_217 br_217 wl_212 vdd gnd cell_6t
Xbit_r213_c217 bl_217 br_217 wl_213 vdd gnd cell_6t
Xbit_r214_c217 bl_217 br_217 wl_214 vdd gnd cell_6t
Xbit_r215_c217 bl_217 br_217 wl_215 vdd gnd cell_6t
Xbit_r216_c217 bl_217 br_217 wl_216 vdd gnd cell_6t
Xbit_r217_c217 bl_217 br_217 wl_217 vdd gnd cell_6t
Xbit_r218_c217 bl_217 br_217 wl_218 vdd gnd cell_6t
Xbit_r219_c217 bl_217 br_217 wl_219 vdd gnd cell_6t
Xbit_r220_c217 bl_217 br_217 wl_220 vdd gnd cell_6t
Xbit_r221_c217 bl_217 br_217 wl_221 vdd gnd cell_6t
Xbit_r222_c217 bl_217 br_217 wl_222 vdd gnd cell_6t
Xbit_r223_c217 bl_217 br_217 wl_223 vdd gnd cell_6t
Xbit_r224_c217 bl_217 br_217 wl_224 vdd gnd cell_6t
Xbit_r225_c217 bl_217 br_217 wl_225 vdd gnd cell_6t
Xbit_r226_c217 bl_217 br_217 wl_226 vdd gnd cell_6t
Xbit_r227_c217 bl_217 br_217 wl_227 vdd gnd cell_6t
Xbit_r228_c217 bl_217 br_217 wl_228 vdd gnd cell_6t
Xbit_r229_c217 bl_217 br_217 wl_229 vdd gnd cell_6t
Xbit_r230_c217 bl_217 br_217 wl_230 vdd gnd cell_6t
Xbit_r231_c217 bl_217 br_217 wl_231 vdd gnd cell_6t
Xbit_r232_c217 bl_217 br_217 wl_232 vdd gnd cell_6t
Xbit_r233_c217 bl_217 br_217 wl_233 vdd gnd cell_6t
Xbit_r234_c217 bl_217 br_217 wl_234 vdd gnd cell_6t
Xbit_r235_c217 bl_217 br_217 wl_235 vdd gnd cell_6t
Xbit_r236_c217 bl_217 br_217 wl_236 vdd gnd cell_6t
Xbit_r237_c217 bl_217 br_217 wl_237 vdd gnd cell_6t
Xbit_r238_c217 bl_217 br_217 wl_238 vdd gnd cell_6t
Xbit_r239_c217 bl_217 br_217 wl_239 vdd gnd cell_6t
Xbit_r240_c217 bl_217 br_217 wl_240 vdd gnd cell_6t
Xbit_r241_c217 bl_217 br_217 wl_241 vdd gnd cell_6t
Xbit_r242_c217 bl_217 br_217 wl_242 vdd gnd cell_6t
Xbit_r243_c217 bl_217 br_217 wl_243 vdd gnd cell_6t
Xbit_r244_c217 bl_217 br_217 wl_244 vdd gnd cell_6t
Xbit_r245_c217 bl_217 br_217 wl_245 vdd gnd cell_6t
Xbit_r246_c217 bl_217 br_217 wl_246 vdd gnd cell_6t
Xbit_r247_c217 bl_217 br_217 wl_247 vdd gnd cell_6t
Xbit_r248_c217 bl_217 br_217 wl_248 vdd gnd cell_6t
Xbit_r249_c217 bl_217 br_217 wl_249 vdd gnd cell_6t
Xbit_r250_c217 bl_217 br_217 wl_250 vdd gnd cell_6t
Xbit_r251_c217 bl_217 br_217 wl_251 vdd gnd cell_6t
Xbit_r252_c217 bl_217 br_217 wl_252 vdd gnd cell_6t
Xbit_r253_c217 bl_217 br_217 wl_253 vdd gnd cell_6t
Xbit_r254_c217 bl_217 br_217 wl_254 vdd gnd cell_6t
Xbit_r255_c217 bl_217 br_217 wl_255 vdd gnd cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd cell_6t
Xbit_r1_c218 bl_218 br_218 wl_1 vdd gnd cell_6t
Xbit_r2_c218 bl_218 br_218 wl_2 vdd gnd cell_6t
Xbit_r3_c218 bl_218 br_218 wl_3 vdd gnd cell_6t
Xbit_r4_c218 bl_218 br_218 wl_4 vdd gnd cell_6t
Xbit_r5_c218 bl_218 br_218 wl_5 vdd gnd cell_6t
Xbit_r6_c218 bl_218 br_218 wl_6 vdd gnd cell_6t
Xbit_r7_c218 bl_218 br_218 wl_7 vdd gnd cell_6t
Xbit_r8_c218 bl_218 br_218 wl_8 vdd gnd cell_6t
Xbit_r9_c218 bl_218 br_218 wl_9 vdd gnd cell_6t
Xbit_r10_c218 bl_218 br_218 wl_10 vdd gnd cell_6t
Xbit_r11_c218 bl_218 br_218 wl_11 vdd gnd cell_6t
Xbit_r12_c218 bl_218 br_218 wl_12 vdd gnd cell_6t
Xbit_r13_c218 bl_218 br_218 wl_13 vdd gnd cell_6t
Xbit_r14_c218 bl_218 br_218 wl_14 vdd gnd cell_6t
Xbit_r15_c218 bl_218 br_218 wl_15 vdd gnd cell_6t
Xbit_r16_c218 bl_218 br_218 wl_16 vdd gnd cell_6t
Xbit_r17_c218 bl_218 br_218 wl_17 vdd gnd cell_6t
Xbit_r18_c218 bl_218 br_218 wl_18 vdd gnd cell_6t
Xbit_r19_c218 bl_218 br_218 wl_19 vdd gnd cell_6t
Xbit_r20_c218 bl_218 br_218 wl_20 vdd gnd cell_6t
Xbit_r21_c218 bl_218 br_218 wl_21 vdd gnd cell_6t
Xbit_r22_c218 bl_218 br_218 wl_22 vdd gnd cell_6t
Xbit_r23_c218 bl_218 br_218 wl_23 vdd gnd cell_6t
Xbit_r24_c218 bl_218 br_218 wl_24 vdd gnd cell_6t
Xbit_r25_c218 bl_218 br_218 wl_25 vdd gnd cell_6t
Xbit_r26_c218 bl_218 br_218 wl_26 vdd gnd cell_6t
Xbit_r27_c218 bl_218 br_218 wl_27 vdd gnd cell_6t
Xbit_r28_c218 bl_218 br_218 wl_28 vdd gnd cell_6t
Xbit_r29_c218 bl_218 br_218 wl_29 vdd gnd cell_6t
Xbit_r30_c218 bl_218 br_218 wl_30 vdd gnd cell_6t
Xbit_r31_c218 bl_218 br_218 wl_31 vdd gnd cell_6t
Xbit_r32_c218 bl_218 br_218 wl_32 vdd gnd cell_6t
Xbit_r33_c218 bl_218 br_218 wl_33 vdd gnd cell_6t
Xbit_r34_c218 bl_218 br_218 wl_34 vdd gnd cell_6t
Xbit_r35_c218 bl_218 br_218 wl_35 vdd gnd cell_6t
Xbit_r36_c218 bl_218 br_218 wl_36 vdd gnd cell_6t
Xbit_r37_c218 bl_218 br_218 wl_37 vdd gnd cell_6t
Xbit_r38_c218 bl_218 br_218 wl_38 vdd gnd cell_6t
Xbit_r39_c218 bl_218 br_218 wl_39 vdd gnd cell_6t
Xbit_r40_c218 bl_218 br_218 wl_40 vdd gnd cell_6t
Xbit_r41_c218 bl_218 br_218 wl_41 vdd gnd cell_6t
Xbit_r42_c218 bl_218 br_218 wl_42 vdd gnd cell_6t
Xbit_r43_c218 bl_218 br_218 wl_43 vdd gnd cell_6t
Xbit_r44_c218 bl_218 br_218 wl_44 vdd gnd cell_6t
Xbit_r45_c218 bl_218 br_218 wl_45 vdd gnd cell_6t
Xbit_r46_c218 bl_218 br_218 wl_46 vdd gnd cell_6t
Xbit_r47_c218 bl_218 br_218 wl_47 vdd gnd cell_6t
Xbit_r48_c218 bl_218 br_218 wl_48 vdd gnd cell_6t
Xbit_r49_c218 bl_218 br_218 wl_49 vdd gnd cell_6t
Xbit_r50_c218 bl_218 br_218 wl_50 vdd gnd cell_6t
Xbit_r51_c218 bl_218 br_218 wl_51 vdd gnd cell_6t
Xbit_r52_c218 bl_218 br_218 wl_52 vdd gnd cell_6t
Xbit_r53_c218 bl_218 br_218 wl_53 vdd gnd cell_6t
Xbit_r54_c218 bl_218 br_218 wl_54 vdd gnd cell_6t
Xbit_r55_c218 bl_218 br_218 wl_55 vdd gnd cell_6t
Xbit_r56_c218 bl_218 br_218 wl_56 vdd gnd cell_6t
Xbit_r57_c218 bl_218 br_218 wl_57 vdd gnd cell_6t
Xbit_r58_c218 bl_218 br_218 wl_58 vdd gnd cell_6t
Xbit_r59_c218 bl_218 br_218 wl_59 vdd gnd cell_6t
Xbit_r60_c218 bl_218 br_218 wl_60 vdd gnd cell_6t
Xbit_r61_c218 bl_218 br_218 wl_61 vdd gnd cell_6t
Xbit_r62_c218 bl_218 br_218 wl_62 vdd gnd cell_6t
Xbit_r63_c218 bl_218 br_218 wl_63 vdd gnd cell_6t
Xbit_r64_c218 bl_218 br_218 wl_64 vdd gnd cell_6t
Xbit_r65_c218 bl_218 br_218 wl_65 vdd gnd cell_6t
Xbit_r66_c218 bl_218 br_218 wl_66 vdd gnd cell_6t
Xbit_r67_c218 bl_218 br_218 wl_67 vdd gnd cell_6t
Xbit_r68_c218 bl_218 br_218 wl_68 vdd gnd cell_6t
Xbit_r69_c218 bl_218 br_218 wl_69 vdd gnd cell_6t
Xbit_r70_c218 bl_218 br_218 wl_70 vdd gnd cell_6t
Xbit_r71_c218 bl_218 br_218 wl_71 vdd gnd cell_6t
Xbit_r72_c218 bl_218 br_218 wl_72 vdd gnd cell_6t
Xbit_r73_c218 bl_218 br_218 wl_73 vdd gnd cell_6t
Xbit_r74_c218 bl_218 br_218 wl_74 vdd gnd cell_6t
Xbit_r75_c218 bl_218 br_218 wl_75 vdd gnd cell_6t
Xbit_r76_c218 bl_218 br_218 wl_76 vdd gnd cell_6t
Xbit_r77_c218 bl_218 br_218 wl_77 vdd gnd cell_6t
Xbit_r78_c218 bl_218 br_218 wl_78 vdd gnd cell_6t
Xbit_r79_c218 bl_218 br_218 wl_79 vdd gnd cell_6t
Xbit_r80_c218 bl_218 br_218 wl_80 vdd gnd cell_6t
Xbit_r81_c218 bl_218 br_218 wl_81 vdd gnd cell_6t
Xbit_r82_c218 bl_218 br_218 wl_82 vdd gnd cell_6t
Xbit_r83_c218 bl_218 br_218 wl_83 vdd gnd cell_6t
Xbit_r84_c218 bl_218 br_218 wl_84 vdd gnd cell_6t
Xbit_r85_c218 bl_218 br_218 wl_85 vdd gnd cell_6t
Xbit_r86_c218 bl_218 br_218 wl_86 vdd gnd cell_6t
Xbit_r87_c218 bl_218 br_218 wl_87 vdd gnd cell_6t
Xbit_r88_c218 bl_218 br_218 wl_88 vdd gnd cell_6t
Xbit_r89_c218 bl_218 br_218 wl_89 vdd gnd cell_6t
Xbit_r90_c218 bl_218 br_218 wl_90 vdd gnd cell_6t
Xbit_r91_c218 bl_218 br_218 wl_91 vdd gnd cell_6t
Xbit_r92_c218 bl_218 br_218 wl_92 vdd gnd cell_6t
Xbit_r93_c218 bl_218 br_218 wl_93 vdd gnd cell_6t
Xbit_r94_c218 bl_218 br_218 wl_94 vdd gnd cell_6t
Xbit_r95_c218 bl_218 br_218 wl_95 vdd gnd cell_6t
Xbit_r96_c218 bl_218 br_218 wl_96 vdd gnd cell_6t
Xbit_r97_c218 bl_218 br_218 wl_97 vdd gnd cell_6t
Xbit_r98_c218 bl_218 br_218 wl_98 vdd gnd cell_6t
Xbit_r99_c218 bl_218 br_218 wl_99 vdd gnd cell_6t
Xbit_r100_c218 bl_218 br_218 wl_100 vdd gnd cell_6t
Xbit_r101_c218 bl_218 br_218 wl_101 vdd gnd cell_6t
Xbit_r102_c218 bl_218 br_218 wl_102 vdd gnd cell_6t
Xbit_r103_c218 bl_218 br_218 wl_103 vdd gnd cell_6t
Xbit_r104_c218 bl_218 br_218 wl_104 vdd gnd cell_6t
Xbit_r105_c218 bl_218 br_218 wl_105 vdd gnd cell_6t
Xbit_r106_c218 bl_218 br_218 wl_106 vdd gnd cell_6t
Xbit_r107_c218 bl_218 br_218 wl_107 vdd gnd cell_6t
Xbit_r108_c218 bl_218 br_218 wl_108 vdd gnd cell_6t
Xbit_r109_c218 bl_218 br_218 wl_109 vdd gnd cell_6t
Xbit_r110_c218 bl_218 br_218 wl_110 vdd gnd cell_6t
Xbit_r111_c218 bl_218 br_218 wl_111 vdd gnd cell_6t
Xbit_r112_c218 bl_218 br_218 wl_112 vdd gnd cell_6t
Xbit_r113_c218 bl_218 br_218 wl_113 vdd gnd cell_6t
Xbit_r114_c218 bl_218 br_218 wl_114 vdd gnd cell_6t
Xbit_r115_c218 bl_218 br_218 wl_115 vdd gnd cell_6t
Xbit_r116_c218 bl_218 br_218 wl_116 vdd gnd cell_6t
Xbit_r117_c218 bl_218 br_218 wl_117 vdd gnd cell_6t
Xbit_r118_c218 bl_218 br_218 wl_118 vdd gnd cell_6t
Xbit_r119_c218 bl_218 br_218 wl_119 vdd gnd cell_6t
Xbit_r120_c218 bl_218 br_218 wl_120 vdd gnd cell_6t
Xbit_r121_c218 bl_218 br_218 wl_121 vdd gnd cell_6t
Xbit_r122_c218 bl_218 br_218 wl_122 vdd gnd cell_6t
Xbit_r123_c218 bl_218 br_218 wl_123 vdd gnd cell_6t
Xbit_r124_c218 bl_218 br_218 wl_124 vdd gnd cell_6t
Xbit_r125_c218 bl_218 br_218 wl_125 vdd gnd cell_6t
Xbit_r126_c218 bl_218 br_218 wl_126 vdd gnd cell_6t
Xbit_r127_c218 bl_218 br_218 wl_127 vdd gnd cell_6t
Xbit_r128_c218 bl_218 br_218 wl_128 vdd gnd cell_6t
Xbit_r129_c218 bl_218 br_218 wl_129 vdd gnd cell_6t
Xbit_r130_c218 bl_218 br_218 wl_130 vdd gnd cell_6t
Xbit_r131_c218 bl_218 br_218 wl_131 vdd gnd cell_6t
Xbit_r132_c218 bl_218 br_218 wl_132 vdd gnd cell_6t
Xbit_r133_c218 bl_218 br_218 wl_133 vdd gnd cell_6t
Xbit_r134_c218 bl_218 br_218 wl_134 vdd gnd cell_6t
Xbit_r135_c218 bl_218 br_218 wl_135 vdd gnd cell_6t
Xbit_r136_c218 bl_218 br_218 wl_136 vdd gnd cell_6t
Xbit_r137_c218 bl_218 br_218 wl_137 vdd gnd cell_6t
Xbit_r138_c218 bl_218 br_218 wl_138 vdd gnd cell_6t
Xbit_r139_c218 bl_218 br_218 wl_139 vdd gnd cell_6t
Xbit_r140_c218 bl_218 br_218 wl_140 vdd gnd cell_6t
Xbit_r141_c218 bl_218 br_218 wl_141 vdd gnd cell_6t
Xbit_r142_c218 bl_218 br_218 wl_142 vdd gnd cell_6t
Xbit_r143_c218 bl_218 br_218 wl_143 vdd gnd cell_6t
Xbit_r144_c218 bl_218 br_218 wl_144 vdd gnd cell_6t
Xbit_r145_c218 bl_218 br_218 wl_145 vdd gnd cell_6t
Xbit_r146_c218 bl_218 br_218 wl_146 vdd gnd cell_6t
Xbit_r147_c218 bl_218 br_218 wl_147 vdd gnd cell_6t
Xbit_r148_c218 bl_218 br_218 wl_148 vdd gnd cell_6t
Xbit_r149_c218 bl_218 br_218 wl_149 vdd gnd cell_6t
Xbit_r150_c218 bl_218 br_218 wl_150 vdd gnd cell_6t
Xbit_r151_c218 bl_218 br_218 wl_151 vdd gnd cell_6t
Xbit_r152_c218 bl_218 br_218 wl_152 vdd gnd cell_6t
Xbit_r153_c218 bl_218 br_218 wl_153 vdd gnd cell_6t
Xbit_r154_c218 bl_218 br_218 wl_154 vdd gnd cell_6t
Xbit_r155_c218 bl_218 br_218 wl_155 vdd gnd cell_6t
Xbit_r156_c218 bl_218 br_218 wl_156 vdd gnd cell_6t
Xbit_r157_c218 bl_218 br_218 wl_157 vdd gnd cell_6t
Xbit_r158_c218 bl_218 br_218 wl_158 vdd gnd cell_6t
Xbit_r159_c218 bl_218 br_218 wl_159 vdd gnd cell_6t
Xbit_r160_c218 bl_218 br_218 wl_160 vdd gnd cell_6t
Xbit_r161_c218 bl_218 br_218 wl_161 vdd gnd cell_6t
Xbit_r162_c218 bl_218 br_218 wl_162 vdd gnd cell_6t
Xbit_r163_c218 bl_218 br_218 wl_163 vdd gnd cell_6t
Xbit_r164_c218 bl_218 br_218 wl_164 vdd gnd cell_6t
Xbit_r165_c218 bl_218 br_218 wl_165 vdd gnd cell_6t
Xbit_r166_c218 bl_218 br_218 wl_166 vdd gnd cell_6t
Xbit_r167_c218 bl_218 br_218 wl_167 vdd gnd cell_6t
Xbit_r168_c218 bl_218 br_218 wl_168 vdd gnd cell_6t
Xbit_r169_c218 bl_218 br_218 wl_169 vdd gnd cell_6t
Xbit_r170_c218 bl_218 br_218 wl_170 vdd gnd cell_6t
Xbit_r171_c218 bl_218 br_218 wl_171 vdd gnd cell_6t
Xbit_r172_c218 bl_218 br_218 wl_172 vdd gnd cell_6t
Xbit_r173_c218 bl_218 br_218 wl_173 vdd gnd cell_6t
Xbit_r174_c218 bl_218 br_218 wl_174 vdd gnd cell_6t
Xbit_r175_c218 bl_218 br_218 wl_175 vdd gnd cell_6t
Xbit_r176_c218 bl_218 br_218 wl_176 vdd gnd cell_6t
Xbit_r177_c218 bl_218 br_218 wl_177 vdd gnd cell_6t
Xbit_r178_c218 bl_218 br_218 wl_178 vdd gnd cell_6t
Xbit_r179_c218 bl_218 br_218 wl_179 vdd gnd cell_6t
Xbit_r180_c218 bl_218 br_218 wl_180 vdd gnd cell_6t
Xbit_r181_c218 bl_218 br_218 wl_181 vdd gnd cell_6t
Xbit_r182_c218 bl_218 br_218 wl_182 vdd gnd cell_6t
Xbit_r183_c218 bl_218 br_218 wl_183 vdd gnd cell_6t
Xbit_r184_c218 bl_218 br_218 wl_184 vdd gnd cell_6t
Xbit_r185_c218 bl_218 br_218 wl_185 vdd gnd cell_6t
Xbit_r186_c218 bl_218 br_218 wl_186 vdd gnd cell_6t
Xbit_r187_c218 bl_218 br_218 wl_187 vdd gnd cell_6t
Xbit_r188_c218 bl_218 br_218 wl_188 vdd gnd cell_6t
Xbit_r189_c218 bl_218 br_218 wl_189 vdd gnd cell_6t
Xbit_r190_c218 bl_218 br_218 wl_190 vdd gnd cell_6t
Xbit_r191_c218 bl_218 br_218 wl_191 vdd gnd cell_6t
Xbit_r192_c218 bl_218 br_218 wl_192 vdd gnd cell_6t
Xbit_r193_c218 bl_218 br_218 wl_193 vdd gnd cell_6t
Xbit_r194_c218 bl_218 br_218 wl_194 vdd gnd cell_6t
Xbit_r195_c218 bl_218 br_218 wl_195 vdd gnd cell_6t
Xbit_r196_c218 bl_218 br_218 wl_196 vdd gnd cell_6t
Xbit_r197_c218 bl_218 br_218 wl_197 vdd gnd cell_6t
Xbit_r198_c218 bl_218 br_218 wl_198 vdd gnd cell_6t
Xbit_r199_c218 bl_218 br_218 wl_199 vdd gnd cell_6t
Xbit_r200_c218 bl_218 br_218 wl_200 vdd gnd cell_6t
Xbit_r201_c218 bl_218 br_218 wl_201 vdd gnd cell_6t
Xbit_r202_c218 bl_218 br_218 wl_202 vdd gnd cell_6t
Xbit_r203_c218 bl_218 br_218 wl_203 vdd gnd cell_6t
Xbit_r204_c218 bl_218 br_218 wl_204 vdd gnd cell_6t
Xbit_r205_c218 bl_218 br_218 wl_205 vdd gnd cell_6t
Xbit_r206_c218 bl_218 br_218 wl_206 vdd gnd cell_6t
Xbit_r207_c218 bl_218 br_218 wl_207 vdd gnd cell_6t
Xbit_r208_c218 bl_218 br_218 wl_208 vdd gnd cell_6t
Xbit_r209_c218 bl_218 br_218 wl_209 vdd gnd cell_6t
Xbit_r210_c218 bl_218 br_218 wl_210 vdd gnd cell_6t
Xbit_r211_c218 bl_218 br_218 wl_211 vdd gnd cell_6t
Xbit_r212_c218 bl_218 br_218 wl_212 vdd gnd cell_6t
Xbit_r213_c218 bl_218 br_218 wl_213 vdd gnd cell_6t
Xbit_r214_c218 bl_218 br_218 wl_214 vdd gnd cell_6t
Xbit_r215_c218 bl_218 br_218 wl_215 vdd gnd cell_6t
Xbit_r216_c218 bl_218 br_218 wl_216 vdd gnd cell_6t
Xbit_r217_c218 bl_218 br_218 wl_217 vdd gnd cell_6t
Xbit_r218_c218 bl_218 br_218 wl_218 vdd gnd cell_6t
Xbit_r219_c218 bl_218 br_218 wl_219 vdd gnd cell_6t
Xbit_r220_c218 bl_218 br_218 wl_220 vdd gnd cell_6t
Xbit_r221_c218 bl_218 br_218 wl_221 vdd gnd cell_6t
Xbit_r222_c218 bl_218 br_218 wl_222 vdd gnd cell_6t
Xbit_r223_c218 bl_218 br_218 wl_223 vdd gnd cell_6t
Xbit_r224_c218 bl_218 br_218 wl_224 vdd gnd cell_6t
Xbit_r225_c218 bl_218 br_218 wl_225 vdd gnd cell_6t
Xbit_r226_c218 bl_218 br_218 wl_226 vdd gnd cell_6t
Xbit_r227_c218 bl_218 br_218 wl_227 vdd gnd cell_6t
Xbit_r228_c218 bl_218 br_218 wl_228 vdd gnd cell_6t
Xbit_r229_c218 bl_218 br_218 wl_229 vdd gnd cell_6t
Xbit_r230_c218 bl_218 br_218 wl_230 vdd gnd cell_6t
Xbit_r231_c218 bl_218 br_218 wl_231 vdd gnd cell_6t
Xbit_r232_c218 bl_218 br_218 wl_232 vdd gnd cell_6t
Xbit_r233_c218 bl_218 br_218 wl_233 vdd gnd cell_6t
Xbit_r234_c218 bl_218 br_218 wl_234 vdd gnd cell_6t
Xbit_r235_c218 bl_218 br_218 wl_235 vdd gnd cell_6t
Xbit_r236_c218 bl_218 br_218 wl_236 vdd gnd cell_6t
Xbit_r237_c218 bl_218 br_218 wl_237 vdd gnd cell_6t
Xbit_r238_c218 bl_218 br_218 wl_238 vdd gnd cell_6t
Xbit_r239_c218 bl_218 br_218 wl_239 vdd gnd cell_6t
Xbit_r240_c218 bl_218 br_218 wl_240 vdd gnd cell_6t
Xbit_r241_c218 bl_218 br_218 wl_241 vdd gnd cell_6t
Xbit_r242_c218 bl_218 br_218 wl_242 vdd gnd cell_6t
Xbit_r243_c218 bl_218 br_218 wl_243 vdd gnd cell_6t
Xbit_r244_c218 bl_218 br_218 wl_244 vdd gnd cell_6t
Xbit_r245_c218 bl_218 br_218 wl_245 vdd gnd cell_6t
Xbit_r246_c218 bl_218 br_218 wl_246 vdd gnd cell_6t
Xbit_r247_c218 bl_218 br_218 wl_247 vdd gnd cell_6t
Xbit_r248_c218 bl_218 br_218 wl_248 vdd gnd cell_6t
Xbit_r249_c218 bl_218 br_218 wl_249 vdd gnd cell_6t
Xbit_r250_c218 bl_218 br_218 wl_250 vdd gnd cell_6t
Xbit_r251_c218 bl_218 br_218 wl_251 vdd gnd cell_6t
Xbit_r252_c218 bl_218 br_218 wl_252 vdd gnd cell_6t
Xbit_r253_c218 bl_218 br_218 wl_253 vdd gnd cell_6t
Xbit_r254_c218 bl_218 br_218 wl_254 vdd gnd cell_6t
Xbit_r255_c218 bl_218 br_218 wl_255 vdd gnd cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd cell_6t
Xbit_r1_c219 bl_219 br_219 wl_1 vdd gnd cell_6t
Xbit_r2_c219 bl_219 br_219 wl_2 vdd gnd cell_6t
Xbit_r3_c219 bl_219 br_219 wl_3 vdd gnd cell_6t
Xbit_r4_c219 bl_219 br_219 wl_4 vdd gnd cell_6t
Xbit_r5_c219 bl_219 br_219 wl_5 vdd gnd cell_6t
Xbit_r6_c219 bl_219 br_219 wl_6 vdd gnd cell_6t
Xbit_r7_c219 bl_219 br_219 wl_7 vdd gnd cell_6t
Xbit_r8_c219 bl_219 br_219 wl_8 vdd gnd cell_6t
Xbit_r9_c219 bl_219 br_219 wl_9 vdd gnd cell_6t
Xbit_r10_c219 bl_219 br_219 wl_10 vdd gnd cell_6t
Xbit_r11_c219 bl_219 br_219 wl_11 vdd gnd cell_6t
Xbit_r12_c219 bl_219 br_219 wl_12 vdd gnd cell_6t
Xbit_r13_c219 bl_219 br_219 wl_13 vdd gnd cell_6t
Xbit_r14_c219 bl_219 br_219 wl_14 vdd gnd cell_6t
Xbit_r15_c219 bl_219 br_219 wl_15 vdd gnd cell_6t
Xbit_r16_c219 bl_219 br_219 wl_16 vdd gnd cell_6t
Xbit_r17_c219 bl_219 br_219 wl_17 vdd gnd cell_6t
Xbit_r18_c219 bl_219 br_219 wl_18 vdd gnd cell_6t
Xbit_r19_c219 bl_219 br_219 wl_19 vdd gnd cell_6t
Xbit_r20_c219 bl_219 br_219 wl_20 vdd gnd cell_6t
Xbit_r21_c219 bl_219 br_219 wl_21 vdd gnd cell_6t
Xbit_r22_c219 bl_219 br_219 wl_22 vdd gnd cell_6t
Xbit_r23_c219 bl_219 br_219 wl_23 vdd gnd cell_6t
Xbit_r24_c219 bl_219 br_219 wl_24 vdd gnd cell_6t
Xbit_r25_c219 bl_219 br_219 wl_25 vdd gnd cell_6t
Xbit_r26_c219 bl_219 br_219 wl_26 vdd gnd cell_6t
Xbit_r27_c219 bl_219 br_219 wl_27 vdd gnd cell_6t
Xbit_r28_c219 bl_219 br_219 wl_28 vdd gnd cell_6t
Xbit_r29_c219 bl_219 br_219 wl_29 vdd gnd cell_6t
Xbit_r30_c219 bl_219 br_219 wl_30 vdd gnd cell_6t
Xbit_r31_c219 bl_219 br_219 wl_31 vdd gnd cell_6t
Xbit_r32_c219 bl_219 br_219 wl_32 vdd gnd cell_6t
Xbit_r33_c219 bl_219 br_219 wl_33 vdd gnd cell_6t
Xbit_r34_c219 bl_219 br_219 wl_34 vdd gnd cell_6t
Xbit_r35_c219 bl_219 br_219 wl_35 vdd gnd cell_6t
Xbit_r36_c219 bl_219 br_219 wl_36 vdd gnd cell_6t
Xbit_r37_c219 bl_219 br_219 wl_37 vdd gnd cell_6t
Xbit_r38_c219 bl_219 br_219 wl_38 vdd gnd cell_6t
Xbit_r39_c219 bl_219 br_219 wl_39 vdd gnd cell_6t
Xbit_r40_c219 bl_219 br_219 wl_40 vdd gnd cell_6t
Xbit_r41_c219 bl_219 br_219 wl_41 vdd gnd cell_6t
Xbit_r42_c219 bl_219 br_219 wl_42 vdd gnd cell_6t
Xbit_r43_c219 bl_219 br_219 wl_43 vdd gnd cell_6t
Xbit_r44_c219 bl_219 br_219 wl_44 vdd gnd cell_6t
Xbit_r45_c219 bl_219 br_219 wl_45 vdd gnd cell_6t
Xbit_r46_c219 bl_219 br_219 wl_46 vdd gnd cell_6t
Xbit_r47_c219 bl_219 br_219 wl_47 vdd gnd cell_6t
Xbit_r48_c219 bl_219 br_219 wl_48 vdd gnd cell_6t
Xbit_r49_c219 bl_219 br_219 wl_49 vdd gnd cell_6t
Xbit_r50_c219 bl_219 br_219 wl_50 vdd gnd cell_6t
Xbit_r51_c219 bl_219 br_219 wl_51 vdd gnd cell_6t
Xbit_r52_c219 bl_219 br_219 wl_52 vdd gnd cell_6t
Xbit_r53_c219 bl_219 br_219 wl_53 vdd gnd cell_6t
Xbit_r54_c219 bl_219 br_219 wl_54 vdd gnd cell_6t
Xbit_r55_c219 bl_219 br_219 wl_55 vdd gnd cell_6t
Xbit_r56_c219 bl_219 br_219 wl_56 vdd gnd cell_6t
Xbit_r57_c219 bl_219 br_219 wl_57 vdd gnd cell_6t
Xbit_r58_c219 bl_219 br_219 wl_58 vdd gnd cell_6t
Xbit_r59_c219 bl_219 br_219 wl_59 vdd gnd cell_6t
Xbit_r60_c219 bl_219 br_219 wl_60 vdd gnd cell_6t
Xbit_r61_c219 bl_219 br_219 wl_61 vdd gnd cell_6t
Xbit_r62_c219 bl_219 br_219 wl_62 vdd gnd cell_6t
Xbit_r63_c219 bl_219 br_219 wl_63 vdd gnd cell_6t
Xbit_r64_c219 bl_219 br_219 wl_64 vdd gnd cell_6t
Xbit_r65_c219 bl_219 br_219 wl_65 vdd gnd cell_6t
Xbit_r66_c219 bl_219 br_219 wl_66 vdd gnd cell_6t
Xbit_r67_c219 bl_219 br_219 wl_67 vdd gnd cell_6t
Xbit_r68_c219 bl_219 br_219 wl_68 vdd gnd cell_6t
Xbit_r69_c219 bl_219 br_219 wl_69 vdd gnd cell_6t
Xbit_r70_c219 bl_219 br_219 wl_70 vdd gnd cell_6t
Xbit_r71_c219 bl_219 br_219 wl_71 vdd gnd cell_6t
Xbit_r72_c219 bl_219 br_219 wl_72 vdd gnd cell_6t
Xbit_r73_c219 bl_219 br_219 wl_73 vdd gnd cell_6t
Xbit_r74_c219 bl_219 br_219 wl_74 vdd gnd cell_6t
Xbit_r75_c219 bl_219 br_219 wl_75 vdd gnd cell_6t
Xbit_r76_c219 bl_219 br_219 wl_76 vdd gnd cell_6t
Xbit_r77_c219 bl_219 br_219 wl_77 vdd gnd cell_6t
Xbit_r78_c219 bl_219 br_219 wl_78 vdd gnd cell_6t
Xbit_r79_c219 bl_219 br_219 wl_79 vdd gnd cell_6t
Xbit_r80_c219 bl_219 br_219 wl_80 vdd gnd cell_6t
Xbit_r81_c219 bl_219 br_219 wl_81 vdd gnd cell_6t
Xbit_r82_c219 bl_219 br_219 wl_82 vdd gnd cell_6t
Xbit_r83_c219 bl_219 br_219 wl_83 vdd gnd cell_6t
Xbit_r84_c219 bl_219 br_219 wl_84 vdd gnd cell_6t
Xbit_r85_c219 bl_219 br_219 wl_85 vdd gnd cell_6t
Xbit_r86_c219 bl_219 br_219 wl_86 vdd gnd cell_6t
Xbit_r87_c219 bl_219 br_219 wl_87 vdd gnd cell_6t
Xbit_r88_c219 bl_219 br_219 wl_88 vdd gnd cell_6t
Xbit_r89_c219 bl_219 br_219 wl_89 vdd gnd cell_6t
Xbit_r90_c219 bl_219 br_219 wl_90 vdd gnd cell_6t
Xbit_r91_c219 bl_219 br_219 wl_91 vdd gnd cell_6t
Xbit_r92_c219 bl_219 br_219 wl_92 vdd gnd cell_6t
Xbit_r93_c219 bl_219 br_219 wl_93 vdd gnd cell_6t
Xbit_r94_c219 bl_219 br_219 wl_94 vdd gnd cell_6t
Xbit_r95_c219 bl_219 br_219 wl_95 vdd gnd cell_6t
Xbit_r96_c219 bl_219 br_219 wl_96 vdd gnd cell_6t
Xbit_r97_c219 bl_219 br_219 wl_97 vdd gnd cell_6t
Xbit_r98_c219 bl_219 br_219 wl_98 vdd gnd cell_6t
Xbit_r99_c219 bl_219 br_219 wl_99 vdd gnd cell_6t
Xbit_r100_c219 bl_219 br_219 wl_100 vdd gnd cell_6t
Xbit_r101_c219 bl_219 br_219 wl_101 vdd gnd cell_6t
Xbit_r102_c219 bl_219 br_219 wl_102 vdd gnd cell_6t
Xbit_r103_c219 bl_219 br_219 wl_103 vdd gnd cell_6t
Xbit_r104_c219 bl_219 br_219 wl_104 vdd gnd cell_6t
Xbit_r105_c219 bl_219 br_219 wl_105 vdd gnd cell_6t
Xbit_r106_c219 bl_219 br_219 wl_106 vdd gnd cell_6t
Xbit_r107_c219 bl_219 br_219 wl_107 vdd gnd cell_6t
Xbit_r108_c219 bl_219 br_219 wl_108 vdd gnd cell_6t
Xbit_r109_c219 bl_219 br_219 wl_109 vdd gnd cell_6t
Xbit_r110_c219 bl_219 br_219 wl_110 vdd gnd cell_6t
Xbit_r111_c219 bl_219 br_219 wl_111 vdd gnd cell_6t
Xbit_r112_c219 bl_219 br_219 wl_112 vdd gnd cell_6t
Xbit_r113_c219 bl_219 br_219 wl_113 vdd gnd cell_6t
Xbit_r114_c219 bl_219 br_219 wl_114 vdd gnd cell_6t
Xbit_r115_c219 bl_219 br_219 wl_115 vdd gnd cell_6t
Xbit_r116_c219 bl_219 br_219 wl_116 vdd gnd cell_6t
Xbit_r117_c219 bl_219 br_219 wl_117 vdd gnd cell_6t
Xbit_r118_c219 bl_219 br_219 wl_118 vdd gnd cell_6t
Xbit_r119_c219 bl_219 br_219 wl_119 vdd gnd cell_6t
Xbit_r120_c219 bl_219 br_219 wl_120 vdd gnd cell_6t
Xbit_r121_c219 bl_219 br_219 wl_121 vdd gnd cell_6t
Xbit_r122_c219 bl_219 br_219 wl_122 vdd gnd cell_6t
Xbit_r123_c219 bl_219 br_219 wl_123 vdd gnd cell_6t
Xbit_r124_c219 bl_219 br_219 wl_124 vdd gnd cell_6t
Xbit_r125_c219 bl_219 br_219 wl_125 vdd gnd cell_6t
Xbit_r126_c219 bl_219 br_219 wl_126 vdd gnd cell_6t
Xbit_r127_c219 bl_219 br_219 wl_127 vdd gnd cell_6t
Xbit_r128_c219 bl_219 br_219 wl_128 vdd gnd cell_6t
Xbit_r129_c219 bl_219 br_219 wl_129 vdd gnd cell_6t
Xbit_r130_c219 bl_219 br_219 wl_130 vdd gnd cell_6t
Xbit_r131_c219 bl_219 br_219 wl_131 vdd gnd cell_6t
Xbit_r132_c219 bl_219 br_219 wl_132 vdd gnd cell_6t
Xbit_r133_c219 bl_219 br_219 wl_133 vdd gnd cell_6t
Xbit_r134_c219 bl_219 br_219 wl_134 vdd gnd cell_6t
Xbit_r135_c219 bl_219 br_219 wl_135 vdd gnd cell_6t
Xbit_r136_c219 bl_219 br_219 wl_136 vdd gnd cell_6t
Xbit_r137_c219 bl_219 br_219 wl_137 vdd gnd cell_6t
Xbit_r138_c219 bl_219 br_219 wl_138 vdd gnd cell_6t
Xbit_r139_c219 bl_219 br_219 wl_139 vdd gnd cell_6t
Xbit_r140_c219 bl_219 br_219 wl_140 vdd gnd cell_6t
Xbit_r141_c219 bl_219 br_219 wl_141 vdd gnd cell_6t
Xbit_r142_c219 bl_219 br_219 wl_142 vdd gnd cell_6t
Xbit_r143_c219 bl_219 br_219 wl_143 vdd gnd cell_6t
Xbit_r144_c219 bl_219 br_219 wl_144 vdd gnd cell_6t
Xbit_r145_c219 bl_219 br_219 wl_145 vdd gnd cell_6t
Xbit_r146_c219 bl_219 br_219 wl_146 vdd gnd cell_6t
Xbit_r147_c219 bl_219 br_219 wl_147 vdd gnd cell_6t
Xbit_r148_c219 bl_219 br_219 wl_148 vdd gnd cell_6t
Xbit_r149_c219 bl_219 br_219 wl_149 vdd gnd cell_6t
Xbit_r150_c219 bl_219 br_219 wl_150 vdd gnd cell_6t
Xbit_r151_c219 bl_219 br_219 wl_151 vdd gnd cell_6t
Xbit_r152_c219 bl_219 br_219 wl_152 vdd gnd cell_6t
Xbit_r153_c219 bl_219 br_219 wl_153 vdd gnd cell_6t
Xbit_r154_c219 bl_219 br_219 wl_154 vdd gnd cell_6t
Xbit_r155_c219 bl_219 br_219 wl_155 vdd gnd cell_6t
Xbit_r156_c219 bl_219 br_219 wl_156 vdd gnd cell_6t
Xbit_r157_c219 bl_219 br_219 wl_157 vdd gnd cell_6t
Xbit_r158_c219 bl_219 br_219 wl_158 vdd gnd cell_6t
Xbit_r159_c219 bl_219 br_219 wl_159 vdd gnd cell_6t
Xbit_r160_c219 bl_219 br_219 wl_160 vdd gnd cell_6t
Xbit_r161_c219 bl_219 br_219 wl_161 vdd gnd cell_6t
Xbit_r162_c219 bl_219 br_219 wl_162 vdd gnd cell_6t
Xbit_r163_c219 bl_219 br_219 wl_163 vdd gnd cell_6t
Xbit_r164_c219 bl_219 br_219 wl_164 vdd gnd cell_6t
Xbit_r165_c219 bl_219 br_219 wl_165 vdd gnd cell_6t
Xbit_r166_c219 bl_219 br_219 wl_166 vdd gnd cell_6t
Xbit_r167_c219 bl_219 br_219 wl_167 vdd gnd cell_6t
Xbit_r168_c219 bl_219 br_219 wl_168 vdd gnd cell_6t
Xbit_r169_c219 bl_219 br_219 wl_169 vdd gnd cell_6t
Xbit_r170_c219 bl_219 br_219 wl_170 vdd gnd cell_6t
Xbit_r171_c219 bl_219 br_219 wl_171 vdd gnd cell_6t
Xbit_r172_c219 bl_219 br_219 wl_172 vdd gnd cell_6t
Xbit_r173_c219 bl_219 br_219 wl_173 vdd gnd cell_6t
Xbit_r174_c219 bl_219 br_219 wl_174 vdd gnd cell_6t
Xbit_r175_c219 bl_219 br_219 wl_175 vdd gnd cell_6t
Xbit_r176_c219 bl_219 br_219 wl_176 vdd gnd cell_6t
Xbit_r177_c219 bl_219 br_219 wl_177 vdd gnd cell_6t
Xbit_r178_c219 bl_219 br_219 wl_178 vdd gnd cell_6t
Xbit_r179_c219 bl_219 br_219 wl_179 vdd gnd cell_6t
Xbit_r180_c219 bl_219 br_219 wl_180 vdd gnd cell_6t
Xbit_r181_c219 bl_219 br_219 wl_181 vdd gnd cell_6t
Xbit_r182_c219 bl_219 br_219 wl_182 vdd gnd cell_6t
Xbit_r183_c219 bl_219 br_219 wl_183 vdd gnd cell_6t
Xbit_r184_c219 bl_219 br_219 wl_184 vdd gnd cell_6t
Xbit_r185_c219 bl_219 br_219 wl_185 vdd gnd cell_6t
Xbit_r186_c219 bl_219 br_219 wl_186 vdd gnd cell_6t
Xbit_r187_c219 bl_219 br_219 wl_187 vdd gnd cell_6t
Xbit_r188_c219 bl_219 br_219 wl_188 vdd gnd cell_6t
Xbit_r189_c219 bl_219 br_219 wl_189 vdd gnd cell_6t
Xbit_r190_c219 bl_219 br_219 wl_190 vdd gnd cell_6t
Xbit_r191_c219 bl_219 br_219 wl_191 vdd gnd cell_6t
Xbit_r192_c219 bl_219 br_219 wl_192 vdd gnd cell_6t
Xbit_r193_c219 bl_219 br_219 wl_193 vdd gnd cell_6t
Xbit_r194_c219 bl_219 br_219 wl_194 vdd gnd cell_6t
Xbit_r195_c219 bl_219 br_219 wl_195 vdd gnd cell_6t
Xbit_r196_c219 bl_219 br_219 wl_196 vdd gnd cell_6t
Xbit_r197_c219 bl_219 br_219 wl_197 vdd gnd cell_6t
Xbit_r198_c219 bl_219 br_219 wl_198 vdd gnd cell_6t
Xbit_r199_c219 bl_219 br_219 wl_199 vdd gnd cell_6t
Xbit_r200_c219 bl_219 br_219 wl_200 vdd gnd cell_6t
Xbit_r201_c219 bl_219 br_219 wl_201 vdd gnd cell_6t
Xbit_r202_c219 bl_219 br_219 wl_202 vdd gnd cell_6t
Xbit_r203_c219 bl_219 br_219 wl_203 vdd gnd cell_6t
Xbit_r204_c219 bl_219 br_219 wl_204 vdd gnd cell_6t
Xbit_r205_c219 bl_219 br_219 wl_205 vdd gnd cell_6t
Xbit_r206_c219 bl_219 br_219 wl_206 vdd gnd cell_6t
Xbit_r207_c219 bl_219 br_219 wl_207 vdd gnd cell_6t
Xbit_r208_c219 bl_219 br_219 wl_208 vdd gnd cell_6t
Xbit_r209_c219 bl_219 br_219 wl_209 vdd gnd cell_6t
Xbit_r210_c219 bl_219 br_219 wl_210 vdd gnd cell_6t
Xbit_r211_c219 bl_219 br_219 wl_211 vdd gnd cell_6t
Xbit_r212_c219 bl_219 br_219 wl_212 vdd gnd cell_6t
Xbit_r213_c219 bl_219 br_219 wl_213 vdd gnd cell_6t
Xbit_r214_c219 bl_219 br_219 wl_214 vdd gnd cell_6t
Xbit_r215_c219 bl_219 br_219 wl_215 vdd gnd cell_6t
Xbit_r216_c219 bl_219 br_219 wl_216 vdd gnd cell_6t
Xbit_r217_c219 bl_219 br_219 wl_217 vdd gnd cell_6t
Xbit_r218_c219 bl_219 br_219 wl_218 vdd gnd cell_6t
Xbit_r219_c219 bl_219 br_219 wl_219 vdd gnd cell_6t
Xbit_r220_c219 bl_219 br_219 wl_220 vdd gnd cell_6t
Xbit_r221_c219 bl_219 br_219 wl_221 vdd gnd cell_6t
Xbit_r222_c219 bl_219 br_219 wl_222 vdd gnd cell_6t
Xbit_r223_c219 bl_219 br_219 wl_223 vdd gnd cell_6t
Xbit_r224_c219 bl_219 br_219 wl_224 vdd gnd cell_6t
Xbit_r225_c219 bl_219 br_219 wl_225 vdd gnd cell_6t
Xbit_r226_c219 bl_219 br_219 wl_226 vdd gnd cell_6t
Xbit_r227_c219 bl_219 br_219 wl_227 vdd gnd cell_6t
Xbit_r228_c219 bl_219 br_219 wl_228 vdd gnd cell_6t
Xbit_r229_c219 bl_219 br_219 wl_229 vdd gnd cell_6t
Xbit_r230_c219 bl_219 br_219 wl_230 vdd gnd cell_6t
Xbit_r231_c219 bl_219 br_219 wl_231 vdd gnd cell_6t
Xbit_r232_c219 bl_219 br_219 wl_232 vdd gnd cell_6t
Xbit_r233_c219 bl_219 br_219 wl_233 vdd gnd cell_6t
Xbit_r234_c219 bl_219 br_219 wl_234 vdd gnd cell_6t
Xbit_r235_c219 bl_219 br_219 wl_235 vdd gnd cell_6t
Xbit_r236_c219 bl_219 br_219 wl_236 vdd gnd cell_6t
Xbit_r237_c219 bl_219 br_219 wl_237 vdd gnd cell_6t
Xbit_r238_c219 bl_219 br_219 wl_238 vdd gnd cell_6t
Xbit_r239_c219 bl_219 br_219 wl_239 vdd gnd cell_6t
Xbit_r240_c219 bl_219 br_219 wl_240 vdd gnd cell_6t
Xbit_r241_c219 bl_219 br_219 wl_241 vdd gnd cell_6t
Xbit_r242_c219 bl_219 br_219 wl_242 vdd gnd cell_6t
Xbit_r243_c219 bl_219 br_219 wl_243 vdd gnd cell_6t
Xbit_r244_c219 bl_219 br_219 wl_244 vdd gnd cell_6t
Xbit_r245_c219 bl_219 br_219 wl_245 vdd gnd cell_6t
Xbit_r246_c219 bl_219 br_219 wl_246 vdd gnd cell_6t
Xbit_r247_c219 bl_219 br_219 wl_247 vdd gnd cell_6t
Xbit_r248_c219 bl_219 br_219 wl_248 vdd gnd cell_6t
Xbit_r249_c219 bl_219 br_219 wl_249 vdd gnd cell_6t
Xbit_r250_c219 bl_219 br_219 wl_250 vdd gnd cell_6t
Xbit_r251_c219 bl_219 br_219 wl_251 vdd gnd cell_6t
Xbit_r252_c219 bl_219 br_219 wl_252 vdd gnd cell_6t
Xbit_r253_c219 bl_219 br_219 wl_253 vdd gnd cell_6t
Xbit_r254_c219 bl_219 br_219 wl_254 vdd gnd cell_6t
Xbit_r255_c219 bl_219 br_219 wl_255 vdd gnd cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd cell_6t
Xbit_r1_c220 bl_220 br_220 wl_1 vdd gnd cell_6t
Xbit_r2_c220 bl_220 br_220 wl_2 vdd gnd cell_6t
Xbit_r3_c220 bl_220 br_220 wl_3 vdd gnd cell_6t
Xbit_r4_c220 bl_220 br_220 wl_4 vdd gnd cell_6t
Xbit_r5_c220 bl_220 br_220 wl_5 vdd gnd cell_6t
Xbit_r6_c220 bl_220 br_220 wl_6 vdd gnd cell_6t
Xbit_r7_c220 bl_220 br_220 wl_7 vdd gnd cell_6t
Xbit_r8_c220 bl_220 br_220 wl_8 vdd gnd cell_6t
Xbit_r9_c220 bl_220 br_220 wl_9 vdd gnd cell_6t
Xbit_r10_c220 bl_220 br_220 wl_10 vdd gnd cell_6t
Xbit_r11_c220 bl_220 br_220 wl_11 vdd gnd cell_6t
Xbit_r12_c220 bl_220 br_220 wl_12 vdd gnd cell_6t
Xbit_r13_c220 bl_220 br_220 wl_13 vdd gnd cell_6t
Xbit_r14_c220 bl_220 br_220 wl_14 vdd gnd cell_6t
Xbit_r15_c220 bl_220 br_220 wl_15 vdd gnd cell_6t
Xbit_r16_c220 bl_220 br_220 wl_16 vdd gnd cell_6t
Xbit_r17_c220 bl_220 br_220 wl_17 vdd gnd cell_6t
Xbit_r18_c220 bl_220 br_220 wl_18 vdd gnd cell_6t
Xbit_r19_c220 bl_220 br_220 wl_19 vdd gnd cell_6t
Xbit_r20_c220 bl_220 br_220 wl_20 vdd gnd cell_6t
Xbit_r21_c220 bl_220 br_220 wl_21 vdd gnd cell_6t
Xbit_r22_c220 bl_220 br_220 wl_22 vdd gnd cell_6t
Xbit_r23_c220 bl_220 br_220 wl_23 vdd gnd cell_6t
Xbit_r24_c220 bl_220 br_220 wl_24 vdd gnd cell_6t
Xbit_r25_c220 bl_220 br_220 wl_25 vdd gnd cell_6t
Xbit_r26_c220 bl_220 br_220 wl_26 vdd gnd cell_6t
Xbit_r27_c220 bl_220 br_220 wl_27 vdd gnd cell_6t
Xbit_r28_c220 bl_220 br_220 wl_28 vdd gnd cell_6t
Xbit_r29_c220 bl_220 br_220 wl_29 vdd gnd cell_6t
Xbit_r30_c220 bl_220 br_220 wl_30 vdd gnd cell_6t
Xbit_r31_c220 bl_220 br_220 wl_31 vdd gnd cell_6t
Xbit_r32_c220 bl_220 br_220 wl_32 vdd gnd cell_6t
Xbit_r33_c220 bl_220 br_220 wl_33 vdd gnd cell_6t
Xbit_r34_c220 bl_220 br_220 wl_34 vdd gnd cell_6t
Xbit_r35_c220 bl_220 br_220 wl_35 vdd gnd cell_6t
Xbit_r36_c220 bl_220 br_220 wl_36 vdd gnd cell_6t
Xbit_r37_c220 bl_220 br_220 wl_37 vdd gnd cell_6t
Xbit_r38_c220 bl_220 br_220 wl_38 vdd gnd cell_6t
Xbit_r39_c220 bl_220 br_220 wl_39 vdd gnd cell_6t
Xbit_r40_c220 bl_220 br_220 wl_40 vdd gnd cell_6t
Xbit_r41_c220 bl_220 br_220 wl_41 vdd gnd cell_6t
Xbit_r42_c220 bl_220 br_220 wl_42 vdd gnd cell_6t
Xbit_r43_c220 bl_220 br_220 wl_43 vdd gnd cell_6t
Xbit_r44_c220 bl_220 br_220 wl_44 vdd gnd cell_6t
Xbit_r45_c220 bl_220 br_220 wl_45 vdd gnd cell_6t
Xbit_r46_c220 bl_220 br_220 wl_46 vdd gnd cell_6t
Xbit_r47_c220 bl_220 br_220 wl_47 vdd gnd cell_6t
Xbit_r48_c220 bl_220 br_220 wl_48 vdd gnd cell_6t
Xbit_r49_c220 bl_220 br_220 wl_49 vdd gnd cell_6t
Xbit_r50_c220 bl_220 br_220 wl_50 vdd gnd cell_6t
Xbit_r51_c220 bl_220 br_220 wl_51 vdd gnd cell_6t
Xbit_r52_c220 bl_220 br_220 wl_52 vdd gnd cell_6t
Xbit_r53_c220 bl_220 br_220 wl_53 vdd gnd cell_6t
Xbit_r54_c220 bl_220 br_220 wl_54 vdd gnd cell_6t
Xbit_r55_c220 bl_220 br_220 wl_55 vdd gnd cell_6t
Xbit_r56_c220 bl_220 br_220 wl_56 vdd gnd cell_6t
Xbit_r57_c220 bl_220 br_220 wl_57 vdd gnd cell_6t
Xbit_r58_c220 bl_220 br_220 wl_58 vdd gnd cell_6t
Xbit_r59_c220 bl_220 br_220 wl_59 vdd gnd cell_6t
Xbit_r60_c220 bl_220 br_220 wl_60 vdd gnd cell_6t
Xbit_r61_c220 bl_220 br_220 wl_61 vdd gnd cell_6t
Xbit_r62_c220 bl_220 br_220 wl_62 vdd gnd cell_6t
Xbit_r63_c220 bl_220 br_220 wl_63 vdd gnd cell_6t
Xbit_r64_c220 bl_220 br_220 wl_64 vdd gnd cell_6t
Xbit_r65_c220 bl_220 br_220 wl_65 vdd gnd cell_6t
Xbit_r66_c220 bl_220 br_220 wl_66 vdd gnd cell_6t
Xbit_r67_c220 bl_220 br_220 wl_67 vdd gnd cell_6t
Xbit_r68_c220 bl_220 br_220 wl_68 vdd gnd cell_6t
Xbit_r69_c220 bl_220 br_220 wl_69 vdd gnd cell_6t
Xbit_r70_c220 bl_220 br_220 wl_70 vdd gnd cell_6t
Xbit_r71_c220 bl_220 br_220 wl_71 vdd gnd cell_6t
Xbit_r72_c220 bl_220 br_220 wl_72 vdd gnd cell_6t
Xbit_r73_c220 bl_220 br_220 wl_73 vdd gnd cell_6t
Xbit_r74_c220 bl_220 br_220 wl_74 vdd gnd cell_6t
Xbit_r75_c220 bl_220 br_220 wl_75 vdd gnd cell_6t
Xbit_r76_c220 bl_220 br_220 wl_76 vdd gnd cell_6t
Xbit_r77_c220 bl_220 br_220 wl_77 vdd gnd cell_6t
Xbit_r78_c220 bl_220 br_220 wl_78 vdd gnd cell_6t
Xbit_r79_c220 bl_220 br_220 wl_79 vdd gnd cell_6t
Xbit_r80_c220 bl_220 br_220 wl_80 vdd gnd cell_6t
Xbit_r81_c220 bl_220 br_220 wl_81 vdd gnd cell_6t
Xbit_r82_c220 bl_220 br_220 wl_82 vdd gnd cell_6t
Xbit_r83_c220 bl_220 br_220 wl_83 vdd gnd cell_6t
Xbit_r84_c220 bl_220 br_220 wl_84 vdd gnd cell_6t
Xbit_r85_c220 bl_220 br_220 wl_85 vdd gnd cell_6t
Xbit_r86_c220 bl_220 br_220 wl_86 vdd gnd cell_6t
Xbit_r87_c220 bl_220 br_220 wl_87 vdd gnd cell_6t
Xbit_r88_c220 bl_220 br_220 wl_88 vdd gnd cell_6t
Xbit_r89_c220 bl_220 br_220 wl_89 vdd gnd cell_6t
Xbit_r90_c220 bl_220 br_220 wl_90 vdd gnd cell_6t
Xbit_r91_c220 bl_220 br_220 wl_91 vdd gnd cell_6t
Xbit_r92_c220 bl_220 br_220 wl_92 vdd gnd cell_6t
Xbit_r93_c220 bl_220 br_220 wl_93 vdd gnd cell_6t
Xbit_r94_c220 bl_220 br_220 wl_94 vdd gnd cell_6t
Xbit_r95_c220 bl_220 br_220 wl_95 vdd gnd cell_6t
Xbit_r96_c220 bl_220 br_220 wl_96 vdd gnd cell_6t
Xbit_r97_c220 bl_220 br_220 wl_97 vdd gnd cell_6t
Xbit_r98_c220 bl_220 br_220 wl_98 vdd gnd cell_6t
Xbit_r99_c220 bl_220 br_220 wl_99 vdd gnd cell_6t
Xbit_r100_c220 bl_220 br_220 wl_100 vdd gnd cell_6t
Xbit_r101_c220 bl_220 br_220 wl_101 vdd gnd cell_6t
Xbit_r102_c220 bl_220 br_220 wl_102 vdd gnd cell_6t
Xbit_r103_c220 bl_220 br_220 wl_103 vdd gnd cell_6t
Xbit_r104_c220 bl_220 br_220 wl_104 vdd gnd cell_6t
Xbit_r105_c220 bl_220 br_220 wl_105 vdd gnd cell_6t
Xbit_r106_c220 bl_220 br_220 wl_106 vdd gnd cell_6t
Xbit_r107_c220 bl_220 br_220 wl_107 vdd gnd cell_6t
Xbit_r108_c220 bl_220 br_220 wl_108 vdd gnd cell_6t
Xbit_r109_c220 bl_220 br_220 wl_109 vdd gnd cell_6t
Xbit_r110_c220 bl_220 br_220 wl_110 vdd gnd cell_6t
Xbit_r111_c220 bl_220 br_220 wl_111 vdd gnd cell_6t
Xbit_r112_c220 bl_220 br_220 wl_112 vdd gnd cell_6t
Xbit_r113_c220 bl_220 br_220 wl_113 vdd gnd cell_6t
Xbit_r114_c220 bl_220 br_220 wl_114 vdd gnd cell_6t
Xbit_r115_c220 bl_220 br_220 wl_115 vdd gnd cell_6t
Xbit_r116_c220 bl_220 br_220 wl_116 vdd gnd cell_6t
Xbit_r117_c220 bl_220 br_220 wl_117 vdd gnd cell_6t
Xbit_r118_c220 bl_220 br_220 wl_118 vdd gnd cell_6t
Xbit_r119_c220 bl_220 br_220 wl_119 vdd gnd cell_6t
Xbit_r120_c220 bl_220 br_220 wl_120 vdd gnd cell_6t
Xbit_r121_c220 bl_220 br_220 wl_121 vdd gnd cell_6t
Xbit_r122_c220 bl_220 br_220 wl_122 vdd gnd cell_6t
Xbit_r123_c220 bl_220 br_220 wl_123 vdd gnd cell_6t
Xbit_r124_c220 bl_220 br_220 wl_124 vdd gnd cell_6t
Xbit_r125_c220 bl_220 br_220 wl_125 vdd gnd cell_6t
Xbit_r126_c220 bl_220 br_220 wl_126 vdd gnd cell_6t
Xbit_r127_c220 bl_220 br_220 wl_127 vdd gnd cell_6t
Xbit_r128_c220 bl_220 br_220 wl_128 vdd gnd cell_6t
Xbit_r129_c220 bl_220 br_220 wl_129 vdd gnd cell_6t
Xbit_r130_c220 bl_220 br_220 wl_130 vdd gnd cell_6t
Xbit_r131_c220 bl_220 br_220 wl_131 vdd gnd cell_6t
Xbit_r132_c220 bl_220 br_220 wl_132 vdd gnd cell_6t
Xbit_r133_c220 bl_220 br_220 wl_133 vdd gnd cell_6t
Xbit_r134_c220 bl_220 br_220 wl_134 vdd gnd cell_6t
Xbit_r135_c220 bl_220 br_220 wl_135 vdd gnd cell_6t
Xbit_r136_c220 bl_220 br_220 wl_136 vdd gnd cell_6t
Xbit_r137_c220 bl_220 br_220 wl_137 vdd gnd cell_6t
Xbit_r138_c220 bl_220 br_220 wl_138 vdd gnd cell_6t
Xbit_r139_c220 bl_220 br_220 wl_139 vdd gnd cell_6t
Xbit_r140_c220 bl_220 br_220 wl_140 vdd gnd cell_6t
Xbit_r141_c220 bl_220 br_220 wl_141 vdd gnd cell_6t
Xbit_r142_c220 bl_220 br_220 wl_142 vdd gnd cell_6t
Xbit_r143_c220 bl_220 br_220 wl_143 vdd gnd cell_6t
Xbit_r144_c220 bl_220 br_220 wl_144 vdd gnd cell_6t
Xbit_r145_c220 bl_220 br_220 wl_145 vdd gnd cell_6t
Xbit_r146_c220 bl_220 br_220 wl_146 vdd gnd cell_6t
Xbit_r147_c220 bl_220 br_220 wl_147 vdd gnd cell_6t
Xbit_r148_c220 bl_220 br_220 wl_148 vdd gnd cell_6t
Xbit_r149_c220 bl_220 br_220 wl_149 vdd gnd cell_6t
Xbit_r150_c220 bl_220 br_220 wl_150 vdd gnd cell_6t
Xbit_r151_c220 bl_220 br_220 wl_151 vdd gnd cell_6t
Xbit_r152_c220 bl_220 br_220 wl_152 vdd gnd cell_6t
Xbit_r153_c220 bl_220 br_220 wl_153 vdd gnd cell_6t
Xbit_r154_c220 bl_220 br_220 wl_154 vdd gnd cell_6t
Xbit_r155_c220 bl_220 br_220 wl_155 vdd gnd cell_6t
Xbit_r156_c220 bl_220 br_220 wl_156 vdd gnd cell_6t
Xbit_r157_c220 bl_220 br_220 wl_157 vdd gnd cell_6t
Xbit_r158_c220 bl_220 br_220 wl_158 vdd gnd cell_6t
Xbit_r159_c220 bl_220 br_220 wl_159 vdd gnd cell_6t
Xbit_r160_c220 bl_220 br_220 wl_160 vdd gnd cell_6t
Xbit_r161_c220 bl_220 br_220 wl_161 vdd gnd cell_6t
Xbit_r162_c220 bl_220 br_220 wl_162 vdd gnd cell_6t
Xbit_r163_c220 bl_220 br_220 wl_163 vdd gnd cell_6t
Xbit_r164_c220 bl_220 br_220 wl_164 vdd gnd cell_6t
Xbit_r165_c220 bl_220 br_220 wl_165 vdd gnd cell_6t
Xbit_r166_c220 bl_220 br_220 wl_166 vdd gnd cell_6t
Xbit_r167_c220 bl_220 br_220 wl_167 vdd gnd cell_6t
Xbit_r168_c220 bl_220 br_220 wl_168 vdd gnd cell_6t
Xbit_r169_c220 bl_220 br_220 wl_169 vdd gnd cell_6t
Xbit_r170_c220 bl_220 br_220 wl_170 vdd gnd cell_6t
Xbit_r171_c220 bl_220 br_220 wl_171 vdd gnd cell_6t
Xbit_r172_c220 bl_220 br_220 wl_172 vdd gnd cell_6t
Xbit_r173_c220 bl_220 br_220 wl_173 vdd gnd cell_6t
Xbit_r174_c220 bl_220 br_220 wl_174 vdd gnd cell_6t
Xbit_r175_c220 bl_220 br_220 wl_175 vdd gnd cell_6t
Xbit_r176_c220 bl_220 br_220 wl_176 vdd gnd cell_6t
Xbit_r177_c220 bl_220 br_220 wl_177 vdd gnd cell_6t
Xbit_r178_c220 bl_220 br_220 wl_178 vdd gnd cell_6t
Xbit_r179_c220 bl_220 br_220 wl_179 vdd gnd cell_6t
Xbit_r180_c220 bl_220 br_220 wl_180 vdd gnd cell_6t
Xbit_r181_c220 bl_220 br_220 wl_181 vdd gnd cell_6t
Xbit_r182_c220 bl_220 br_220 wl_182 vdd gnd cell_6t
Xbit_r183_c220 bl_220 br_220 wl_183 vdd gnd cell_6t
Xbit_r184_c220 bl_220 br_220 wl_184 vdd gnd cell_6t
Xbit_r185_c220 bl_220 br_220 wl_185 vdd gnd cell_6t
Xbit_r186_c220 bl_220 br_220 wl_186 vdd gnd cell_6t
Xbit_r187_c220 bl_220 br_220 wl_187 vdd gnd cell_6t
Xbit_r188_c220 bl_220 br_220 wl_188 vdd gnd cell_6t
Xbit_r189_c220 bl_220 br_220 wl_189 vdd gnd cell_6t
Xbit_r190_c220 bl_220 br_220 wl_190 vdd gnd cell_6t
Xbit_r191_c220 bl_220 br_220 wl_191 vdd gnd cell_6t
Xbit_r192_c220 bl_220 br_220 wl_192 vdd gnd cell_6t
Xbit_r193_c220 bl_220 br_220 wl_193 vdd gnd cell_6t
Xbit_r194_c220 bl_220 br_220 wl_194 vdd gnd cell_6t
Xbit_r195_c220 bl_220 br_220 wl_195 vdd gnd cell_6t
Xbit_r196_c220 bl_220 br_220 wl_196 vdd gnd cell_6t
Xbit_r197_c220 bl_220 br_220 wl_197 vdd gnd cell_6t
Xbit_r198_c220 bl_220 br_220 wl_198 vdd gnd cell_6t
Xbit_r199_c220 bl_220 br_220 wl_199 vdd gnd cell_6t
Xbit_r200_c220 bl_220 br_220 wl_200 vdd gnd cell_6t
Xbit_r201_c220 bl_220 br_220 wl_201 vdd gnd cell_6t
Xbit_r202_c220 bl_220 br_220 wl_202 vdd gnd cell_6t
Xbit_r203_c220 bl_220 br_220 wl_203 vdd gnd cell_6t
Xbit_r204_c220 bl_220 br_220 wl_204 vdd gnd cell_6t
Xbit_r205_c220 bl_220 br_220 wl_205 vdd gnd cell_6t
Xbit_r206_c220 bl_220 br_220 wl_206 vdd gnd cell_6t
Xbit_r207_c220 bl_220 br_220 wl_207 vdd gnd cell_6t
Xbit_r208_c220 bl_220 br_220 wl_208 vdd gnd cell_6t
Xbit_r209_c220 bl_220 br_220 wl_209 vdd gnd cell_6t
Xbit_r210_c220 bl_220 br_220 wl_210 vdd gnd cell_6t
Xbit_r211_c220 bl_220 br_220 wl_211 vdd gnd cell_6t
Xbit_r212_c220 bl_220 br_220 wl_212 vdd gnd cell_6t
Xbit_r213_c220 bl_220 br_220 wl_213 vdd gnd cell_6t
Xbit_r214_c220 bl_220 br_220 wl_214 vdd gnd cell_6t
Xbit_r215_c220 bl_220 br_220 wl_215 vdd gnd cell_6t
Xbit_r216_c220 bl_220 br_220 wl_216 vdd gnd cell_6t
Xbit_r217_c220 bl_220 br_220 wl_217 vdd gnd cell_6t
Xbit_r218_c220 bl_220 br_220 wl_218 vdd gnd cell_6t
Xbit_r219_c220 bl_220 br_220 wl_219 vdd gnd cell_6t
Xbit_r220_c220 bl_220 br_220 wl_220 vdd gnd cell_6t
Xbit_r221_c220 bl_220 br_220 wl_221 vdd gnd cell_6t
Xbit_r222_c220 bl_220 br_220 wl_222 vdd gnd cell_6t
Xbit_r223_c220 bl_220 br_220 wl_223 vdd gnd cell_6t
Xbit_r224_c220 bl_220 br_220 wl_224 vdd gnd cell_6t
Xbit_r225_c220 bl_220 br_220 wl_225 vdd gnd cell_6t
Xbit_r226_c220 bl_220 br_220 wl_226 vdd gnd cell_6t
Xbit_r227_c220 bl_220 br_220 wl_227 vdd gnd cell_6t
Xbit_r228_c220 bl_220 br_220 wl_228 vdd gnd cell_6t
Xbit_r229_c220 bl_220 br_220 wl_229 vdd gnd cell_6t
Xbit_r230_c220 bl_220 br_220 wl_230 vdd gnd cell_6t
Xbit_r231_c220 bl_220 br_220 wl_231 vdd gnd cell_6t
Xbit_r232_c220 bl_220 br_220 wl_232 vdd gnd cell_6t
Xbit_r233_c220 bl_220 br_220 wl_233 vdd gnd cell_6t
Xbit_r234_c220 bl_220 br_220 wl_234 vdd gnd cell_6t
Xbit_r235_c220 bl_220 br_220 wl_235 vdd gnd cell_6t
Xbit_r236_c220 bl_220 br_220 wl_236 vdd gnd cell_6t
Xbit_r237_c220 bl_220 br_220 wl_237 vdd gnd cell_6t
Xbit_r238_c220 bl_220 br_220 wl_238 vdd gnd cell_6t
Xbit_r239_c220 bl_220 br_220 wl_239 vdd gnd cell_6t
Xbit_r240_c220 bl_220 br_220 wl_240 vdd gnd cell_6t
Xbit_r241_c220 bl_220 br_220 wl_241 vdd gnd cell_6t
Xbit_r242_c220 bl_220 br_220 wl_242 vdd gnd cell_6t
Xbit_r243_c220 bl_220 br_220 wl_243 vdd gnd cell_6t
Xbit_r244_c220 bl_220 br_220 wl_244 vdd gnd cell_6t
Xbit_r245_c220 bl_220 br_220 wl_245 vdd gnd cell_6t
Xbit_r246_c220 bl_220 br_220 wl_246 vdd gnd cell_6t
Xbit_r247_c220 bl_220 br_220 wl_247 vdd gnd cell_6t
Xbit_r248_c220 bl_220 br_220 wl_248 vdd gnd cell_6t
Xbit_r249_c220 bl_220 br_220 wl_249 vdd gnd cell_6t
Xbit_r250_c220 bl_220 br_220 wl_250 vdd gnd cell_6t
Xbit_r251_c220 bl_220 br_220 wl_251 vdd gnd cell_6t
Xbit_r252_c220 bl_220 br_220 wl_252 vdd gnd cell_6t
Xbit_r253_c220 bl_220 br_220 wl_253 vdd gnd cell_6t
Xbit_r254_c220 bl_220 br_220 wl_254 vdd gnd cell_6t
Xbit_r255_c220 bl_220 br_220 wl_255 vdd gnd cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd cell_6t
Xbit_r1_c221 bl_221 br_221 wl_1 vdd gnd cell_6t
Xbit_r2_c221 bl_221 br_221 wl_2 vdd gnd cell_6t
Xbit_r3_c221 bl_221 br_221 wl_3 vdd gnd cell_6t
Xbit_r4_c221 bl_221 br_221 wl_4 vdd gnd cell_6t
Xbit_r5_c221 bl_221 br_221 wl_5 vdd gnd cell_6t
Xbit_r6_c221 bl_221 br_221 wl_6 vdd gnd cell_6t
Xbit_r7_c221 bl_221 br_221 wl_7 vdd gnd cell_6t
Xbit_r8_c221 bl_221 br_221 wl_8 vdd gnd cell_6t
Xbit_r9_c221 bl_221 br_221 wl_9 vdd gnd cell_6t
Xbit_r10_c221 bl_221 br_221 wl_10 vdd gnd cell_6t
Xbit_r11_c221 bl_221 br_221 wl_11 vdd gnd cell_6t
Xbit_r12_c221 bl_221 br_221 wl_12 vdd gnd cell_6t
Xbit_r13_c221 bl_221 br_221 wl_13 vdd gnd cell_6t
Xbit_r14_c221 bl_221 br_221 wl_14 vdd gnd cell_6t
Xbit_r15_c221 bl_221 br_221 wl_15 vdd gnd cell_6t
Xbit_r16_c221 bl_221 br_221 wl_16 vdd gnd cell_6t
Xbit_r17_c221 bl_221 br_221 wl_17 vdd gnd cell_6t
Xbit_r18_c221 bl_221 br_221 wl_18 vdd gnd cell_6t
Xbit_r19_c221 bl_221 br_221 wl_19 vdd gnd cell_6t
Xbit_r20_c221 bl_221 br_221 wl_20 vdd gnd cell_6t
Xbit_r21_c221 bl_221 br_221 wl_21 vdd gnd cell_6t
Xbit_r22_c221 bl_221 br_221 wl_22 vdd gnd cell_6t
Xbit_r23_c221 bl_221 br_221 wl_23 vdd gnd cell_6t
Xbit_r24_c221 bl_221 br_221 wl_24 vdd gnd cell_6t
Xbit_r25_c221 bl_221 br_221 wl_25 vdd gnd cell_6t
Xbit_r26_c221 bl_221 br_221 wl_26 vdd gnd cell_6t
Xbit_r27_c221 bl_221 br_221 wl_27 vdd gnd cell_6t
Xbit_r28_c221 bl_221 br_221 wl_28 vdd gnd cell_6t
Xbit_r29_c221 bl_221 br_221 wl_29 vdd gnd cell_6t
Xbit_r30_c221 bl_221 br_221 wl_30 vdd gnd cell_6t
Xbit_r31_c221 bl_221 br_221 wl_31 vdd gnd cell_6t
Xbit_r32_c221 bl_221 br_221 wl_32 vdd gnd cell_6t
Xbit_r33_c221 bl_221 br_221 wl_33 vdd gnd cell_6t
Xbit_r34_c221 bl_221 br_221 wl_34 vdd gnd cell_6t
Xbit_r35_c221 bl_221 br_221 wl_35 vdd gnd cell_6t
Xbit_r36_c221 bl_221 br_221 wl_36 vdd gnd cell_6t
Xbit_r37_c221 bl_221 br_221 wl_37 vdd gnd cell_6t
Xbit_r38_c221 bl_221 br_221 wl_38 vdd gnd cell_6t
Xbit_r39_c221 bl_221 br_221 wl_39 vdd gnd cell_6t
Xbit_r40_c221 bl_221 br_221 wl_40 vdd gnd cell_6t
Xbit_r41_c221 bl_221 br_221 wl_41 vdd gnd cell_6t
Xbit_r42_c221 bl_221 br_221 wl_42 vdd gnd cell_6t
Xbit_r43_c221 bl_221 br_221 wl_43 vdd gnd cell_6t
Xbit_r44_c221 bl_221 br_221 wl_44 vdd gnd cell_6t
Xbit_r45_c221 bl_221 br_221 wl_45 vdd gnd cell_6t
Xbit_r46_c221 bl_221 br_221 wl_46 vdd gnd cell_6t
Xbit_r47_c221 bl_221 br_221 wl_47 vdd gnd cell_6t
Xbit_r48_c221 bl_221 br_221 wl_48 vdd gnd cell_6t
Xbit_r49_c221 bl_221 br_221 wl_49 vdd gnd cell_6t
Xbit_r50_c221 bl_221 br_221 wl_50 vdd gnd cell_6t
Xbit_r51_c221 bl_221 br_221 wl_51 vdd gnd cell_6t
Xbit_r52_c221 bl_221 br_221 wl_52 vdd gnd cell_6t
Xbit_r53_c221 bl_221 br_221 wl_53 vdd gnd cell_6t
Xbit_r54_c221 bl_221 br_221 wl_54 vdd gnd cell_6t
Xbit_r55_c221 bl_221 br_221 wl_55 vdd gnd cell_6t
Xbit_r56_c221 bl_221 br_221 wl_56 vdd gnd cell_6t
Xbit_r57_c221 bl_221 br_221 wl_57 vdd gnd cell_6t
Xbit_r58_c221 bl_221 br_221 wl_58 vdd gnd cell_6t
Xbit_r59_c221 bl_221 br_221 wl_59 vdd gnd cell_6t
Xbit_r60_c221 bl_221 br_221 wl_60 vdd gnd cell_6t
Xbit_r61_c221 bl_221 br_221 wl_61 vdd gnd cell_6t
Xbit_r62_c221 bl_221 br_221 wl_62 vdd gnd cell_6t
Xbit_r63_c221 bl_221 br_221 wl_63 vdd gnd cell_6t
Xbit_r64_c221 bl_221 br_221 wl_64 vdd gnd cell_6t
Xbit_r65_c221 bl_221 br_221 wl_65 vdd gnd cell_6t
Xbit_r66_c221 bl_221 br_221 wl_66 vdd gnd cell_6t
Xbit_r67_c221 bl_221 br_221 wl_67 vdd gnd cell_6t
Xbit_r68_c221 bl_221 br_221 wl_68 vdd gnd cell_6t
Xbit_r69_c221 bl_221 br_221 wl_69 vdd gnd cell_6t
Xbit_r70_c221 bl_221 br_221 wl_70 vdd gnd cell_6t
Xbit_r71_c221 bl_221 br_221 wl_71 vdd gnd cell_6t
Xbit_r72_c221 bl_221 br_221 wl_72 vdd gnd cell_6t
Xbit_r73_c221 bl_221 br_221 wl_73 vdd gnd cell_6t
Xbit_r74_c221 bl_221 br_221 wl_74 vdd gnd cell_6t
Xbit_r75_c221 bl_221 br_221 wl_75 vdd gnd cell_6t
Xbit_r76_c221 bl_221 br_221 wl_76 vdd gnd cell_6t
Xbit_r77_c221 bl_221 br_221 wl_77 vdd gnd cell_6t
Xbit_r78_c221 bl_221 br_221 wl_78 vdd gnd cell_6t
Xbit_r79_c221 bl_221 br_221 wl_79 vdd gnd cell_6t
Xbit_r80_c221 bl_221 br_221 wl_80 vdd gnd cell_6t
Xbit_r81_c221 bl_221 br_221 wl_81 vdd gnd cell_6t
Xbit_r82_c221 bl_221 br_221 wl_82 vdd gnd cell_6t
Xbit_r83_c221 bl_221 br_221 wl_83 vdd gnd cell_6t
Xbit_r84_c221 bl_221 br_221 wl_84 vdd gnd cell_6t
Xbit_r85_c221 bl_221 br_221 wl_85 vdd gnd cell_6t
Xbit_r86_c221 bl_221 br_221 wl_86 vdd gnd cell_6t
Xbit_r87_c221 bl_221 br_221 wl_87 vdd gnd cell_6t
Xbit_r88_c221 bl_221 br_221 wl_88 vdd gnd cell_6t
Xbit_r89_c221 bl_221 br_221 wl_89 vdd gnd cell_6t
Xbit_r90_c221 bl_221 br_221 wl_90 vdd gnd cell_6t
Xbit_r91_c221 bl_221 br_221 wl_91 vdd gnd cell_6t
Xbit_r92_c221 bl_221 br_221 wl_92 vdd gnd cell_6t
Xbit_r93_c221 bl_221 br_221 wl_93 vdd gnd cell_6t
Xbit_r94_c221 bl_221 br_221 wl_94 vdd gnd cell_6t
Xbit_r95_c221 bl_221 br_221 wl_95 vdd gnd cell_6t
Xbit_r96_c221 bl_221 br_221 wl_96 vdd gnd cell_6t
Xbit_r97_c221 bl_221 br_221 wl_97 vdd gnd cell_6t
Xbit_r98_c221 bl_221 br_221 wl_98 vdd gnd cell_6t
Xbit_r99_c221 bl_221 br_221 wl_99 vdd gnd cell_6t
Xbit_r100_c221 bl_221 br_221 wl_100 vdd gnd cell_6t
Xbit_r101_c221 bl_221 br_221 wl_101 vdd gnd cell_6t
Xbit_r102_c221 bl_221 br_221 wl_102 vdd gnd cell_6t
Xbit_r103_c221 bl_221 br_221 wl_103 vdd gnd cell_6t
Xbit_r104_c221 bl_221 br_221 wl_104 vdd gnd cell_6t
Xbit_r105_c221 bl_221 br_221 wl_105 vdd gnd cell_6t
Xbit_r106_c221 bl_221 br_221 wl_106 vdd gnd cell_6t
Xbit_r107_c221 bl_221 br_221 wl_107 vdd gnd cell_6t
Xbit_r108_c221 bl_221 br_221 wl_108 vdd gnd cell_6t
Xbit_r109_c221 bl_221 br_221 wl_109 vdd gnd cell_6t
Xbit_r110_c221 bl_221 br_221 wl_110 vdd gnd cell_6t
Xbit_r111_c221 bl_221 br_221 wl_111 vdd gnd cell_6t
Xbit_r112_c221 bl_221 br_221 wl_112 vdd gnd cell_6t
Xbit_r113_c221 bl_221 br_221 wl_113 vdd gnd cell_6t
Xbit_r114_c221 bl_221 br_221 wl_114 vdd gnd cell_6t
Xbit_r115_c221 bl_221 br_221 wl_115 vdd gnd cell_6t
Xbit_r116_c221 bl_221 br_221 wl_116 vdd gnd cell_6t
Xbit_r117_c221 bl_221 br_221 wl_117 vdd gnd cell_6t
Xbit_r118_c221 bl_221 br_221 wl_118 vdd gnd cell_6t
Xbit_r119_c221 bl_221 br_221 wl_119 vdd gnd cell_6t
Xbit_r120_c221 bl_221 br_221 wl_120 vdd gnd cell_6t
Xbit_r121_c221 bl_221 br_221 wl_121 vdd gnd cell_6t
Xbit_r122_c221 bl_221 br_221 wl_122 vdd gnd cell_6t
Xbit_r123_c221 bl_221 br_221 wl_123 vdd gnd cell_6t
Xbit_r124_c221 bl_221 br_221 wl_124 vdd gnd cell_6t
Xbit_r125_c221 bl_221 br_221 wl_125 vdd gnd cell_6t
Xbit_r126_c221 bl_221 br_221 wl_126 vdd gnd cell_6t
Xbit_r127_c221 bl_221 br_221 wl_127 vdd gnd cell_6t
Xbit_r128_c221 bl_221 br_221 wl_128 vdd gnd cell_6t
Xbit_r129_c221 bl_221 br_221 wl_129 vdd gnd cell_6t
Xbit_r130_c221 bl_221 br_221 wl_130 vdd gnd cell_6t
Xbit_r131_c221 bl_221 br_221 wl_131 vdd gnd cell_6t
Xbit_r132_c221 bl_221 br_221 wl_132 vdd gnd cell_6t
Xbit_r133_c221 bl_221 br_221 wl_133 vdd gnd cell_6t
Xbit_r134_c221 bl_221 br_221 wl_134 vdd gnd cell_6t
Xbit_r135_c221 bl_221 br_221 wl_135 vdd gnd cell_6t
Xbit_r136_c221 bl_221 br_221 wl_136 vdd gnd cell_6t
Xbit_r137_c221 bl_221 br_221 wl_137 vdd gnd cell_6t
Xbit_r138_c221 bl_221 br_221 wl_138 vdd gnd cell_6t
Xbit_r139_c221 bl_221 br_221 wl_139 vdd gnd cell_6t
Xbit_r140_c221 bl_221 br_221 wl_140 vdd gnd cell_6t
Xbit_r141_c221 bl_221 br_221 wl_141 vdd gnd cell_6t
Xbit_r142_c221 bl_221 br_221 wl_142 vdd gnd cell_6t
Xbit_r143_c221 bl_221 br_221 wl_143 vdd gnd cell_6t
Xbit_r144_c221 bl_221 br_221 wl_144 vdd gnd cell_6t
Xbit_r145_c221 bl_221 br_221 wl_145 vdd gnd cell_6t
Xbit_r146_c221 bl_221 br_221 wl_146 vdd gnd cell_6t
Xbit_r147_c221 bl_221 br_221 wl_147 vdd gnd cell_6t
Xbit_r148_c221 bl_221 br_221 wl_148 vdd gnd cell_6t
Xbit_r149_c221 bl_221 br_221 wl_149 vdd gnd cell_6t
Xbit_r150_c221 bl_221 br_221 wl_150 vdd gnd cell_6t
Xbit_r151_c221 bl_221 br_221 wl_151 vdd gnd cell_6t
Xbit_r152_c221 bl_221 br_221 wl_152 vdd gnd cell_6t
Xbit_r153_c221 bl_221 br_221 wl_153 vdd gnd cell_6t
Xbit_r154_c221 bl_221 br_221 wl_154 vdd gnd cell_6t
Xbit_r155_c221 bl_221 br_221 wl_155 vdd gnd cell_6t
Xbit_r156_c221 bl_221 br_221 wl_156 vdd gnd cell_6t
Xbit_r157_c221 bl_221 br_221 wl_157 vdd gnd cell_6t
Xbit_r158_c221 bl_221 br_221 wl_158 vdd gnd cell_6t
Xbit_r159_c221 bl_221 br_221 wl_159 vdd gnd cell_6t
Xbit_r160_c221 bl_221 br_221 wl_160 vdd gnd cell_6t
Xbit_r161_c221 bl_221 br_221 wl_161 vdd gnd cell_6t
Xbit_r162_c221 bl_221 br_221 wl_162 vdd gnd cell_6t
Xbit_r163_c221 bl_221 br_221 wl_163 vdd gnd cell_6t
Xbit_r164_c221 bl_221 br_221 wl_164 vdd gnd cell_6t
Xbit_r165_c221 bl_221 br_221 wl_165 vdd gnd cell_6t
Xbit_r166_c221 bl_221 br_221 wl_166 vdd gnd cell_6t
Xbit_r167_c221 bl_221 br_221 wl_167 vdd gnd cell_6t
Xbit_r168_c221 bl_221 br_221 wl_168 vdd gnd cell_6t
Xbit_r169_c221 bl_221 br_221 wl_169 vdd gnd cell_6t
Xbit_r170_c221 bl_221 br_221 wl_170 vdd gnd cell_6t
Xbit_r171_c221 bl_221 br_221 wl_171 vdd gnd cell_6t
Xbit_r172_c221 bl_221 br_221 wl_172 vdd gnd cell_6t
Xbit_r173_c221 bl_221 br_221 wl_173 vdd gnd cell_6t
Xbit_r174_c221 bl_221 br_221 wl_174 vdd gnd cell_6t
Xbit_r175_c221 bl_221 br_221 wl_175 vdd gnd cell_6t
Xbit_r176_c221 bl_221 br_221 wl_176 vdd gnd cell_6t
Xbit_r177_c221 bl_221 br_221 wl_177 vdd gnd cell_6t
Xbit_r178_c221 bl_221 br_221 wl_178 vdd gnd cell_6t
Xbit_r179_c221 bl_221 br_221 wl_179 vdd gnd cell_6t
Xbit_r180_c221 bl_221 br_221 wl_180 vdd gnd cell_6t
Xbit_r181_c221 bl_221 br_221 wl_181 vdd gnd cell_6t
Xbit_r182_c221 bl_221 br_221 wl_182 vdd gnd cell_6t
Xbit_r183_c221 bl_221 br_221 wl_183 vdd gnd cell_6t
Xbit_r184_c221 bl_221 br_221 wl_184 vdd gnd cell_6t
Xbit_r185_c221 bl_221 br_221 wl_185 vdd gnd cell_6t
Xbit_r186_c221 bl_221 br_221 wl_186 vdd gnd cell_6t
Xbit_r187_c221 bl_221 br_221 wl_187 vdd gnd cell_6t
Xbit_r188_c221 bl_221 br_221 wl_188 vdd gnd cell_6t
Xbit_r189_c221 bl_221 br_221 wl_189 vdd gnd cell_6t
Xbit_r190_c221 bl_221 br_221 wl_190 vdd gnd cell_6t
Xbit_r191_c221 bl_221 br_221 wl_191 vdd gnd cell_6t
Xbit_r192_c221 bl_221 br_221 wl_192 vdd gnd cell_6t
Xbit_r193_c221 bl_221 br_221 wl_193 vdd gnd cell_6t
Xbit_r194_c221 bl_221 br_221 wl_194 vdd gnd cell_6t
Xbit_r195_c221 bl_221 br_221 wl_195 vdd gnd cell_6t
Xbit_r196_c221 bl_221 br_221 wl_196 vdd gnd cell_6t
Xbit_r197_c221 bl_221 br_221 wl_197 vdd gnd cell_6t
Xbit_r198_c221 bl_221 br_221 wl_198 vdd gnd cell_6t
Xbit_r199_c221 bl_221 br_221 wl_199 vdd gnd cell_6t
Xbit_r200_c221 bl_221 br_221 wl_200 vdd gnd cell_6t
Xbit_r201_c221 bl_221 br_221 wl_201 vdd gnd cell_6t
Xbit_r202_c221 bl_221 br_221 wl_202 vdd gnd cell_6t
Xbit_r203_c221 bl_221 br_221 wl_203 vdd gnd cell_6t
Xbit_r204_c221 bl_221 br_221 wl_204 vdd gnd cell_6t
Xbit_r205_c221 bl_221 br_221 wl_205 vdd gnd cell_6t
Xbit_r206_c221 bl_221 br_221 wl_206 vdd gnd cell_6t
Xbit_r207_c221 bl_221 br_221 wl_207 vdd gnd cell_6t
Xbit_r208_c221 bl_221 br_221 wl_208 vdd gnd cell_6t
Xbit_r209_c221 bl_221 br_221 wl_209 vdd gnd cell_6t
Xbit_r210_c221 bl_221 br_221 wl_210 vdd gnd cell_6t
Xbit_r211_c221 bl_221 br_221 wl_211 vdd gnd cell_6t
Xbit_r212_c221 bl_221 br_221 wl_212 vdd gnd cell_6t
Xbit_r213_c221 bl_221 br_221 wl_213 vdd gnd cell_6t
Xbit_r214_c221 bl_221 br_221 wl_214 vdd gnd cell_6t
Xbit_r215_c221 bl_221 br_221 wl_215 vdd gnd cell_6t
Xbit_r216_c221 bl_221 br_221 wl_216 vdd gnd cell_6t
Xbit_r217_c221 bl_221 br_221 wl_217 vdd gnd cell_6t
Xbit_r218_c221 bl_221 br_221 wl_218 vdd gnd cell_6t
Xbit_r219_c221 bl_221 br_221 wl_219 vdd gnd cell_6t
Xbit_r220_c221 bl_221 br_221 wl_220 vdd gnd cell_6t
Xbit_r221_c221 bl_221 br_221 wl_221 vdd gnd cell_6t
Xbit_r222_c221 bl_221 br_221 wl_222 vdd gnd cell_6t
Xbit_r223_c221 bl_221 br_221 wl_223 vdd gnd cell_6t
Xbit_r224_c221 bl_221 br_221 wl_224 vdd gnd cell_6t
Xbit_r225_c221 bl_221 br_221 wl_225 vdd gnd cell_6t
Xbit_r226_c221 bl_221 br_221 wl_226 vdd gnd cell_6t
Xbit_r227_c221 bl_221 br_221 wl_227 vdd gnd cell_6t
Xbit_r228_c221 bl_221 br_221 wl_228 vdd gnd cell_6t
Xbit_r229_c221 bl_221 br_221 wl_229 vdd gnd cell_6t
Xbit_r230_c221 bl_221 br_221 wl_230 vdd gnd cell_6t
Xbit_r231_c221 bl_221 br_221 wl_231 vdd gnd cell_6t
Xbit_r232_c221 bl_221 br_221 wl_232 vdd gnd cell_6t
Xbit_r233_c221 bl_221 br_221 wl_233 vdd gnd cell_6t
Xbit_r234_c221 bl_221 br_221 wl_234 vdd gnd cell_6t
Xbit_r235_c221 bl_221 br_221 wl_235 vdd gnd cell_6t
Xbit_r236_c221 bl_221 br_221 wl_236 vdd gnd cell_6t
Xbit_r237_c221 bl_221 br_221 wl_237 vdd gnd cell_6t
Xbit_r238_c221 bl_221 br_221 wl_238 vdd gnd cell_6t
Xbit_r239_c221 bl_221 br_221 wl_239 vdd gnd cell_6t
Xbit_r240_c221 bl_221 br_221 wl_240 vdd gnd cell_6t
Xbit_r241_c221 bl_221 br_221 wl_241 vdd gnd cell_6t
Xbit_r242_c221 bl_221 br_221 wl_242 vdd gnd cell_6t
Xbit_r243_c221 bl_221 br_221 wl_243 vdd gnd cell_6t
Xbit_r244_c221 bl_221 br_221 wl_244 vdd gnd cell_6t
Xbit_r245_c221 bl_221 br_221 wl_245 vdd gnd cell_6t
Xbit_r246_c221 bl_221 br_221 wl_246 vdd gnd cell_6t
Xbit_r247_c221 bl_221 br_221 wl_247 vdd gnd cell_6t
Xbit_r248_c221 bl_221 br_221 wl_248 vdd gnd cell_6t
Xbit_r249_c221 bl_221 br_221 wl_249 vdd gnd cell_6t
Xbit_r250_c221 bl_221 br_221 wl_250 vdd gnd cell_6t
Xbit_r251_c221 bl_221 br_221 wl_251 vdd gnd cell_6t
Xbit_r252_c221 bl_221 br_221 wl_252 vdd gnd cell_6t
Xbit_r253_c221 bl_221 br_221 wl_253 vdd gnd cell_6t
Xbit_r254_c221 bl_221 br_221 wl_254 vdd gnd cell_6t
Xbit_r255_c221 bl_221 br_221 wl_255 vdd gnd cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd cell_6t
Xbit_r1_c222 bl_222 br_222 wl_1 vdd gnd cell_6t
Xbit_r2_c222 bl_222 br_222 wl_2 vdd gnd cell_6t
Xbit_r3_c222 bl_222 br_222 wl_3 vdd gnd cell_6t
Xbit_r4_c222 bl_222 br_222 wl_4 vdd gnd cell_6t
Xbit_r5_c222 bl_222 br_222 wl_5 vdd gnd cell_6t
Xbit_r6_c222 bl_222 br_222 wl_6 vdd gnd cell_6t
Xbit_r7_c222 bl_222 br_222 wl_7 vdd gnd cell_6t
Xbit_r8_c222 bl_222 br_222 wl_8 vdd gnd cell_6t
Xbit_r9_c222 bl_222 br_222 wl_9 vdd gnd cell_6t
Xbit_r10_c222 bl_222 br_222 wl_10 vdd gnd cell_6t
Xbit_r11_c222 bl_222 br_222 wl_11 vdd gnd cell_6t
Xbit_r12_c222 bl_222 br_222 wl_12 vdd gnd cell_6t
Xbit_r13_c222 bl_222 br_222 wl_13 vdd gnd cell_6t
Xbit_r14_c222 bl_222 br_222 wl_14 vdd gnd cell_6t
Xbit_r15_c222 bl_222 br_222 wl_15 vdd gnd cell_6t
Xbit_r16_c222 bl_222 br_222 wl_16 vdd gnd cell_6t
Xbit_r17_c222 bl_222 br_222 wl_17 vdd gnd cell_6t
Xbit_r18_c222 bl_222 br_222 wl_18 vdd gnd cell_6t
Xbit_r19_c222 bl_222 br_222 wl_19 vdd gnd cell_6t
Xbit_r20_c222 bl_222 br_222 wl_20 vdd gnd cell_6t
Xbit_r21_c222 bl_222 br_222 wl_21 vdd gnd cell_6t
Xbit_r22_c222 bl_222 br_222 wl_22 vdd gnd cell_6t
Xbit_r23_c222 bl_222 br_222 wl_23 vdd gnd cell_6t
Xbit_r24_c222 bl_222 br_222 wl_24 vdd gnd cell_6t
Xbit_r25_c222 bl_222 br_222 wl_25 vdd gnd cell_6t
Xbit_r26_c222 bl_222 br_222 wl_26 vdd gnd cell_6t
Xbit_r27_c222 bl_222 br_222 wl_27 vdd gnd cell_6t
Xbit_r28_c222 bl_222 br_222 wl_28 vdd gnd cell_6t
Xbit_r29_c222 bl_222 br_222 wl_29 vdd gnd cell_6t
Xbit_r30_c222 bl_222 br_222 wl_30 vdd gnd cell_6t
Xbit_r31_c222 bl_222 br_222 wl_31 vdd gnd cell_6t
Xbit_r32_c222 bl_222 br_222 wl_32 vdd gnd cell_6t
Xbit_r33_c222 bl_222 br_222 wl_33 vdd gnd cell_6t
Xbit_r34_c222 bl_222 br_222 wl_34 vdd gnd cell_6t
Xbit_r35_c222 bl_222 br_222 wl_35 vdd gnd cell_6t
Xbit_r36_c222 bl_222 br_222 wl_36 vdd gnd cell_6t
Xbit_r37_c222 bl_222 br_222 wl_37 vdd gnd cell_6t
Xbit_r38_c222 bl_222 br_222 wl_38 vdd gnd cell_6t
Xbit_r39_c222 bl_222 br_222 wl_39 vdd gnd cell_6t
Xbit_r40_c222 bl_222 br_222 wl_40 vdd gnd cell_6t
Xbit_r41_c222 bl_222 br_222 wl_41 vdd gnd cell_6t
Xbit_r42_c222 bl_222 br_222 wl_42 vdd gnd cell_6t
Xbit_r43_c222 bl_222 br_222 wl_43 vdd gnd cell_6t
Xbit_r44_c222 bl_222 br_222 wl_44 vdd gnd cell_6t
Xbit_r45_c222 bl_222 br_222 wl_45 vdd gnd cell_6t
Xbit_r46_c222 bl_222 br_222 wl_46 vdd gnd cell_6t
Xbit_r47_c222 bl_222 br_222 wl_47 vdd gnd cell_6t
Xbit_r48_c222 bl_222 br_222 wl_48 vdd gnd cell_6t
Xbit_r49_c222 bl_222 br_222 wl_49 vdd gnd cell_6t
Xbit_r50_c222 bl_222 br_222 wl_50 vdd gnd cell_6t
Xbit_r51_c222 bl_222 br_222 wl_51 vdd gnd cell_6t
Xbit_r52_c222 bl_222 br_222 wl_52 vdd gnd cell_6t
Xbit_r53_c222 bl_222 br_222 wl_53 vdd gnd cell_6t
Xbit_r54_c222 bl_222 br_222 wl_54 vdd gnd cell_6t
Xbit_r55_c222 bl_222 br_222 wl_55 vdd gnd cell_6t
Xbit_r56_c222 bl_222 br_222 wl_56 vdd gnd cell_6t
Xbit_r57_c222 bl_222 br_222 wl_57 vdd gnd cell_6t
Xbit_r58_c222 bl_222 br_222 wl_58 vdd gnd cell_6t
Xbit_r59_c222 bl_222 br_222 wl_59 vdd gnd cell_6t
Xbit_r60_c222 bl_222 br_222 wl_60 vdd gnd cell_6t
Xbit_r61_c222 bl_222 br_222 wl_61 vdd gnd cell_6t
Xbit_r62_c222 bl_222 br_222 wl_62 vdd gnd cell_6t
Xbit_r63_c222 bl_222 br_222 wl_63 vdd gnd cell_6t
Xbit_r64_c222 bl_222 br_222 wl_64 vdd gnd cell_6t
Xbit_r65_c222 bl_222 br_222 wl_65 vdd gnd cell_6t
Xbit_r66_c222 bl_222 br_222 wl_66 vdd gnd cell_6t
Xbit_r67_c222 bl_222 br_222 wl_67 vdd gnd cell_6t
Xbit_r68_c222 bl_222 br_222 wl_68 vdd gnd cell_6t
Xbit_r69_c222 bl_222 br_222 wl_69 vdd gnd cell_6t
Xbit_r70_c222 bl_222 br_222 wl_70 vdd gnd cell_6t
Xbit_r71_c222 bl_222 br_222 wl_71 vdd gnd cell_6t
Xbit_r72_c222 bl_222 br_222 wl_72 vdd gnd cell_6t
Xbit_r73_c222 bl_222 br_222 wl_73 vdd gnd cell_6t
Xbit_r74_c222 bl_222 br_222 wl_74 vdd gnd cell_6t
Xbit_r75_c222 bl_222 br_222 wl_75 vdd gnd cell_6t
Xbit_r76_c222 bl_222 br_222 wl_76 vdd gnd cell_6t
Xbit_r77_c222 bl_222 br_222 wl_77 vdd gnd cell_6t
Xbit_r78_c222 bl_222 br_222 wl_78 vdd gnd cell_6t
Xbit_r79_c222 bl_222 br_222 wl_79 vdd gnd cell_6t
Xbit_r80_c222 bl_222 br_222 wl_80 vdd gnd cell_6t
Xbit_r81_c222 bl_222 br_222 wl_81 vdd gnd cell_6t
Xbit_r82_c222 bl_222 br_222 wl_82 vdd gnd cell_6t
Xbit_r83_c222 bl_222 br_222 wl_83 vdd gnd cell_6t
Xbit_r84_c222 bl_222 br_222 wl_84 vdd gnd cell_6t
Xbit_r85_c222 bl_222 br_222 wl_85 vdd gnd cell_6t
Xbit_r86_c222 bl_222 br_222 wl_86 vdd gnd cell_6t
Xbit_r87_c222 bl_222 br_222 wl_87 vdd gnd cell_6t
Xbit_r88_c222 bl_222 br_222 wl_88 vdd gnd cell_6t
Xbit_r89_c222 bl_222 br_222 wl_89 vdd gnd cell_6t
Xbit_r90_c222 bl_222 br_222 wl_90 vdd gnd cell_6t
Xbit_r91_c222 bl_222 br_222 wl_91 vdd gnd cell_6t
Xbit_r92_c222 bl_222 br_222 wl_92 vdd gnd cell_6t
Xbit_r93_c222 bl_222 br_222 wl_93 vdd gnd cell_6t
Xbit_r94_c222 bl_222 br_222 wl_94 vdd gnd cell_6t
Xbit_r95_c222 bl_222 br_222 wl_95 vdd gnd cell_6t
Xbit_r96_c222 bl_222 br_222 wl_96 vdd gnd cell_6t
Xbit_r97_c222 bl_222 br_222 wl_97 vdd gnd cell_6t
Xbit_r98_c222 bl_222 br_222 wl_98 vdd gnd cell_6t
Xbit_r99_c222 bl_222 br_222 wl_99 vdd gnd cell_6t
Xbit_r100_c222 bl_222 br_222 wl_100 vdd gnd cell_6t
Xbit_r101_c222 bl_222 br_222 wl_101 vdd gnd cell_6t
Xbit_r102_c222 bl_222 br_222 wl_102 vdd gnd cell_6t
Xbit_r103_c222 bl_222 br_222 wl_103 vdd gnd cell_6t
Xbit_r104_c222 bl_222 br_222 wl_104 vdd gnd cell_6t
Xbit_r105_c222 bl_222 br_222 wl_105 vdd gnd cell_6t
Xbit_r106_c222 bl_222 br_222 wl_106 vdd gnd cell_6t
Xbit_r107_c222 bl_222 br_222 wl_107 vdd gnd cell_6t
Xbit_r108_c222 bl_222 br_222 wl_108 vdd gnd cell_6t
Xbit_r109_c222 bl_222 br_222 wl_109 vdd gnd cell_6t
Xbit_r110_c222 bl_222 br_222 wl_110 vdd gnd cell_6t
Xbit_r111_c222 bl_222 br_222 wl_111 vdd gnd cell_6t
Xbit_r112_c222 bl_222 br_222 wl_112 vdd gnd cell_6t
Xbit_r113_c222 bl_222 br_222 wl_113 vdd gnd cell_6t
Xbit_r114_c222 bl_222 br_222 wl_114 vdd gnd cell_6t
Xbit_r115_c222 bl_222 br_222 wl_115 vdd gnd cell_6t
Xbit_r116_c222 bl_222 br_222 wl_116 vdd gnd cell_6t
Xbit_r117_c222 bl_222 br_222 wl_117 vdd gnd cell_6t
Xbit_r118_c222 bl_222 br_222 wl_118 vdd gnd cell_6t
Xbit_r119_c222 bl_222 br_222 wl_119 vdd gnd cell_6t
Xbit_r120_c222 bl_222 br_222 wl_120 vdd gnd cell_6t
Xbit_r121_c222 bl_222 br_222 wl_121 vdd gnd cell_6t
Xbit_r122_c222 bl_222 br_222 wl_122 vdd gnd cell_6t
Xbit_r123_c222 bl_222 br_222 wl_123 vdd gnd cell_6t
Xbit_r124_c222 bl_222 br_222 wl_124 vdd gnd cell_6t
Xbit_r125_c222 bl_222 br_222 wl_125 vdd gnd cell_6t
Xbit_r126_c222 bl_222 br_222 wl_126 vdd gnd cell_6t
Xbit_r127_c222 bl_222 br_222 wl_127 vdd gnd cell_6t
Xbit_r128_c222 bl_222 br_222 wl_128 vdd gnd cell_6t
Xbit_r129_c222 bl_222 br_222 wl_129 vdd gnd cell_6t
Xbit_r130_c222 bl_222 br_222 wl_130 vdd gnd cell_6t
Xbit_r131_c222 bl_222 br_222 wl_131 vdd gnd cell_6t
Xbit_r132_c222 bl_222 br_222 wl_132 vdd gnd cell_6t
Xbit_r133_c222 bl_222 br_222 wl_133 vdd gnd cell_6t
Xbit_r134_c222 bl_222 br_222 wl_134 vdd gnd cell_6t
Xbit_r135_c222 bl_222 br_222 wl_135 vdd gnd cell_6t
Xbit_r136_c222 bl_222 br_222 wl_136 vdd gnd cell_6t
Xbit_r137_c222 bl_222 br_222 wl_137 vdd gnd cell_6t
Xbit_r138_c222 bl_222 br_222 wl_138 vdd gnd cell_6t
Xbit_r139_c222 bl_222 br_222 wl_139 vdd gnd cell_6t
Xbit_r140_c222 bl_222 br_222 wl_140 vdd gnd cell_6t
Xbit_r141_c222 bl_222 br_222 wl_141 vdd gnd cell_6t
Xbit_r142_c222 bl_222 br_222 wl_142 vdd gnd cell_6t
Xbit_r143_c222 bl_222 br_222 wl_143 vdd gnd cell_6t
Xbit_r144_c222 bl_222 br_222 wl_144 vdd gnd cell_6t
Xbit_r145_c222 bl_222 br_222 wl_145 vdd gnd cell_6t
Xbit_r146_c222 bl_222 br_222 wl_146 vdd gnd cell_6t
Xbit_r147_c222 bl_222 br_222 wl_147 vdd gnd cell_6t
Xbit_r148_c222 bl_222 br_222 wl_148 vdd gnd cell_6t
Xbit_r149_c222 bl_222 br_222 wl_149 vdd gnd cell_6t
Xbit_r150_c222 bl_222 br_222 wl_150 vdd gnd cell_6t
Xbit_r151_c222 bl_222 br_222 wl_151 vdd gnd cell_6t
Xbit_r152_c222 bl_222 br_222 wl_152 vdd gnd cell_6t
Xbit_r153_c222 bl_222 br_222 wl_153 vdd gnd cell_6t
Xbit_r154_c222 bl_222 br_222 wl_154 vdd gnd cell_6t
Xbit_r155_c222 bl_222 br_222 wl_155 vdd gnd cell_6t
Xbit_r156_c222 bl_222 br_222 wl_156 vdd gnd cell_6t
Xbit_r157_c222 bl_222 br_222 wl_157 vdd gnd cell_6t
Xbit_r158_c222 bl_222 br_222 wl_158 vdd gnd cell_6t
Xbit_r159_c222 bl_222 br_222 wl_159 vdd gnd cell_6t
Xbit_r160_c222 bl_222 br_222 wl_160 vdd gnd cell_6t
Xbit_r161_c222 bl_222 br_222 wl_161 vdd gnd cell_6t
Xbit_r162_c222 bl_222 br_222 wl_162 vdd gnd cell_6t
Xbit_r163_c222 bl_222 br_222 wl_163 vdd gnd cell_6t
Xbit_r164_c222 bl_222 br_222 wl_164 vdd gnd cell_6t
Xbit_r165_c222 bl_222 br_222 wl_165 vdd gnd cell_6t
Xbit_r166_c222 bl_222 br_222 wl_166 vdd gnd cell_6t
Xbit_r167_c222 bl_222 br_222 wl_167 vdd gnd cell_6t
Xbit_r168_c222 bl_222 br_222 wl_168 vdd gnd cell_6t
Xbit_r169_c222 bl_222 br_222 wl_169 vdd gnd cell_6t
Xbit_r170_c222 bl_222 br_222 wl_170 vdd gnd cell_6t
Xbit_r171_c222 bl_222 br_222 wl_171 vdd gnd cell_6t
Xbit_r172_c222 bl_222 br_222 wl_172 vdd gnd cell_6t
Xbit_r173_c222 bl_222 br_222 wl_173 vdd gnd cell_6t
Xbit_r174_c222 bl_222 br_222 wl_174 vdd gnd cell_6t
Xbit_r175_c222 bl_222 br_222 wl_175 vdd gnd cell_6t
Xbit_r176_c222 bl_222 br_222 wl_176 vdd gnd cell_6t
Xbit_r177_c222 bl_222 br_222 wl_177 vdd gnd cell_6t
Xbit_r178_c222 bl_222 br_222 wl_178 vdd gnd cell_6t
Xbit_r179_c222 bl_222 br_222 wl_179 vdd gnd cell_6t
Xbit_r180_c222 bl_222 br_222 wl_180 vdd gnd cell_6t
Xbit_r181_c222 bl_222 br_222 wl_181 vdd gnd cell_6t
Xbit_r182_c222 bl_222 br_222 wl_182 vdd gnd cell_6t
Xbit_r183_c222 bl_222 br_222 wl_183 vdd gnd cell_6t
Xbit_r184_c222 bl_222 br_222 wl_184 vdd gnd cell_6t
Xbit_r185_c222 bl_222 br_222 wl_185 vdd gnd cell_6t
Xbit_r186_c222 bl_222 br_222 wl_186 vdd gnd cell_6t
Xbit_r187_c222 bl_222 br_222 wl_187 vdd gnd cell_6t
Xbit_r188_c222 bl_222 br_222 wl_188 vdd gnd cell_6t
Xbit_r189_c222 bl_222 br_222 wl_189 vdd gnd cell_6t
Xbit_r190_c222 bl_222 br_222 wl_190 vdd gnd cell_6t
Xbit_r191_c222 bl_222 br_222 wl_191 vdd gnd cell_6t
Xbit_r192_c222 bl_222 br_222 wl_192 vdd gnd cell_6t
Xbit_r193_c222 bl_222 br_222 wl_193 vdd gnd cell_6t
Xbit_r194_c222 bl_222 br_222 wl_194 vdd gnd cell_6t
Xbit_r195_c222 bl_222 br_222 wl_195 vdd gnd cell_6t
Xbit_r196_c222 bl_222 br_222 wl_196 vdd gnd cell_6t
Xbit_r197_c222 bl_222 br_222 wl_197 vdd gnd cell_6t
Xbit_r198_c222 bl_222 br_222 wl_198 vdd gnd cell_6t
Xbit_r199_c222 bl_222 br_222 wl_199 vdd gnd cell_6t
Xbit_r200_c222 bl_222 br_222 wl_200 vdd gnd cell_6t
Xbit_r201_c222 bl_222 br_222 wl_201 vdd gnd cell_6t
Xbit_r202_c222 bl_222 br_222 wl_202 vdd gnd cell_6t
Xbit_r203_c222 bl_222 br_222 wl_203 vdd gnd cell_6t
Xbit_r204_c222 bl_222 br_222 wl_204 vdd gnd cell_6t
Xbit_r205_c222 bl_222 br_222 wl_205 vdd gnd cell_6t
Xbit_r206_c222 bl_222 br_222 wl_206 vdd gnd cell_6t
Xbit_r207_c222 bl_222 br_222 wl_207 vdd gnd cell_6t
Xbit_r208_c222 bl_222 br_222 wl_208 vdd gnd cell_6t
Xbit_r209_c222 bl_222 br_222 wl_209 vdd gnd cell_6t
Xbit_r210_c222 bl_222 br_222 wl_210 vdd gnd cell_6t
Xbit_r211_c222 bl_222 br_222 wl_211 vdd gnd cell_6t
Xbit_r212_c222 bl_222 br_222 wl_212 vdd gnd cell_6t
Xbit_r213_c222 bl_222 br_222 wl_213 vdd gnd cell_6t
Xbit_r214_c222 bl_222 br_222 wl_214 vdd gnd cell_6t
Xbit_r215_c222 bl_222 br_222 wl_215 vdd gnd cell_6t
Xbit_r216_c222 bl_222 br_222 wl_216 vdd gnd cell_6t
Xbit_r217_c222 bl_222 br_222 wl_217 vdd gnd cell_6t
Xbit_r218_c222 bl_222 br_222 wl_218 vdd gnd cell_6t
Xbit_r219_c222 bl_222 br_222 wl_219 vdd gnd cell_6t
Xbit_r220_c222 bl_222 br_222 wl_220 vdd gnd cell_6t
Xbit_r221_c222 bl_222 br_222 wl_221 vdd gnd cell_6t
Xbit_r222_c222 bl_222 br_222 wl_222 vdd gnd cell_6t
Xbit_r223_c222 bl_222 br_222 wl_223 vdd gnd cell_6t
Xbit_r224_c222 bl_222 br_222 wl_224 vdd gnd cell_6t
Xbit_r225_c222 bl_222 br_222 wl_225 vdd gnd cell_6t
Xbit_r226_c222 bl_222 br_222 wl_226 vdd gnd cell_6t
Xbit_r227_c222 bl_222 br_222 wl_227 vdd gnd cell_6t
Xbit_r228_c222 bl_222 br_222 wl_228 vdd gnd cell_6t
Xbit_r229_c222 bl_222 br_222 wl_229 vdd gnd cell_6t
Xbit_r230_c222 bl_222 br_222 wl_230 vdd gnd cell_6t
Xbit_r231_c222 bl_222 br_222 wl_231 vdd gnd cell_6t
Xbit_r232_c222 bl_222 br_222 wl_232 vdd gnd cell_6t
Xbit_r233_c222 bl_222 br_222 wl_233 vdd gnd cell_6t
Xbit_r234_c222 bl_222 br_222 wl_234 vdd gnd cell_6t
Xbit_r235_c222 bl_222 br_222 wl_235 vdd gnd cell_6t
Xbit_r236_c222 bl_222 br_222 wl_236 vdd gnd cell_6t
Xbit_r237_c222 bl_222 br_222 wl_237 vdd gnd cell_6t
Xbit_r238_c222 bl_222 br_222 wl_238 vdd gnd cell_6t
Xbit_r239_c222 bl_222 br_222 wl_239 vdd gnd cell_6t
Xbit_r240_c222 bl_222 br_222 wl_240 vdd gnd cell_6t
Xbit_r241_c222 bl_222 br_222 wl_241 vdd gnd cell_6t
Xbit_r242_c222 bl_222 br_222 wl_242 vdd gnd cell_6t
Xbit_r243_c222 bl_222 br_222 wl_243 vdd gnd cell_6t
Xbit_r244_c222 bl_222 br_222 wl_244 vdd gnd cell_6t
Xbit_r245_c222 bl_222 br_222 wl_245 vdd gnd cell_6t
Xbit_r246_c222 bl_222 br_222 wl_246 vdd gnd cell_6t
Xbit_r247_c222 bl_222 br_222 wl_247 vdd gnd cell_6t
Xbit_r248_c222 bl_222 br_222 wl_248 vdd gnd cell_6t
Xbit_r249_c222 bl_222 br_222 wl_249 vdd gnd cell_6t
Xbit_r250_c222 bl_222 br_222 wl_250 vdd gnd cell_6t
Xbit_r251_c222 bl_222 br_222 wl_251 vdd gnd cell_6t
Xbit_r252_c222 bl_222 br_222 wl_252 vdd gnd cell_6t
Xbit_r253_c222 bl_222 br_222 wl_253 vdd gnd cell_6t
Xbit_r254_c222 bl_222 br_222 wl_254 vdd gnd cell_6t
Xbit_r255_c222 bl_222 br_222 wl_255 vdd gnd cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd cell_6t
Xbit_r1_c223 bl_223 br_223 wl_1 vdd gnd cell_6t
Xbit_r2_c223 bl_223 br_223 wl_2 vdd gnd cell_6t
Xbit_r3_c223 bl_223 br_223 wl_3 vdd gnd cell_6t
Xbit_r4_c223 bl_223 br_223 wl_4 vdd gnd cell_6t
Xbit_r5_c223 bl_223 br_223 wl_5 vdd gnd cell_6t
Xbit_r6_c223 bl_223 br_223 wl_6 vdd gnd cell_6t
Xbit_r7_c223 bl_223 br_223 wl_7 vdd gnd cell_6t
Xbit_r8_c223 bl_223 br_223 wl_8 vdd gnd cell_6t
Xbit_r9_c223 bl_223 br_223 wl_9 vdd gnd cell_6t
Xbit_r10_c223 bl_223 br_223 wl_10 vdd gnd cell_6t
Xbit_r11_c223 bl_223 br_223 wl_11 vdd gnd cell_6t
Xbit_r12_c223 bl_223 br_223 wl_12 vdd gnd cell_6t
Xbit_r13_c223 bl_223 br_223 wl_13 vdd gnd cell_6t
Xbit_r14_c223 bl_223 br_223 wl_14 vdd gnd cell_6t
Xbit_r15_c223 bl_223 br_223 wl_15 vdd gnd cell_6t
Xbit_r16_c223 bl_223 br_223 wl_16 vdd gnd cell_6t
Xbit_r17_c223 bl_223 br_223 wl_17 vdd gnd cell_6t
Xbit_r18_c223 bl_223 br_223 wl_18 vdd gnd cell_6t
Xbit_r19_c223 bl_223 br_223 wl_19 vdd gnd cell_6t
Xbit_r20_c223 bl_223 br_223 wl_20 vdd gnd cell_6t
Xbit_r21_c223 bl_223 br_223 wl_21 vdd gnd cell_6t
Xbit_r22_c223 bl_223 br_223 wl_22 vdd gnd cell_6t
Xbit_r23_c223 bl_223 br_223 wl_23 vdd gnd cell_6t
Xbit_r24_c223 bl_223 br_223 wl_24 vdd gnd cell_6t
Xbit_r25_c223 bl_223 br_223 wl_25 vdd gnd cell_6t
Xbit_r26_c223 bl_223 br_223 wl_26 vdd gnd cell_6t
Xbit_r27_c223 bl_223 br_223 wl_27 vdd gnd cell_6t
Xbit_r28_c223 bl_223 br_223 wl_28 vdd gnd cell_6t
Xbit_r29_c223 bl_223 br_223 wl_29 vdd gnd cell_6t
Xbit_r30_c223 bl_223 br_223 wl_30 vdd gnd cell_6t
Xbit_r31_c223 bl_223 br_223 wl_31 vdd gnd cell_6t
Xbit_r32_c223 bl_223 br_223 wl_32 vdd gnd cell_6t
Xbit_r33_c223 bl_223 br_223 wl_33 vdd gnd cell_6t
Xbit_r34_c223 bl_223 br_223 wl_34 vdd gnd cell_6t
Xbit_r35_c223 bl_223 br_223 wl_35 vdd gnd cell_6t
Xbit_r36_c223 bl_223 br_223 wl_36 vdd gnd cell_6t
Xbit_r37_c223 bl_223 br_223 wl_37 vdd gnd cell_6t
Xbit_r38_c223 bl_223 br_223 wl_38 vdd gnd cell_6t
Xbit_r39_c223 bl_223 br_223 wl_39 vdd gnd cell_6t
Xbit_r40_c223 bl_223 br_223 wl_40 vdd gnd cell_6t
Xbit_r41_c223 bl_223 br_223 wl_41 vdd gnd cell_6t
Xbit_r42_c223 bl_223 br_223 wl_42 vdd gnd cell_6t
Xbit_r43_c223 bl_223 br_223 wl_43 vdd gnd cell_6t
Xbit_r44_c223 bl_223 br_223 wl_44 vdd gnd cell_6t
Xbit_r45_c223 bl_223 br_223 wl_45 vdd gnd cell_6t
Xbit_r46_c223 bl_223 br_223 wl_46 vdd gnd cell_6t
Xbit_r47_c223 bl_223 br_223 wl_47 vdd gnd cell_6t
Xbit_r48_c223 bl_223 br_223 wl_48 vdd gnd cell_6t
Xbit_r49_c223 bl_223 br_223 wl_49 vdd gnd cell_6t
Xbit_r50_c223 bl_223 br_223 wl_50 vdd gnd cell_6t
Xbit_r51_c223 bl_223 br_223 wl_51 vdd gnd cell_6t
Xbit_r52_c223 bl_223 br_223 wl_52 vdd gnd cell_6t
Xbit_r53_c223 bl_223 br_223 wl_53 vdd gnd cell_6t
Xbit_r54_c223 bl_223 br_223 wl_54 vdd gnd cell_6t
Xbit_r55_c223 bl_223 br_223 wl_55 vdd gnd cell_6t
Xbit_r56_c223 bl_223 br_223 wl_56 vdd gnd cell_6t
Xbit_r57_c223 bl_223 br_223 wl_57 vdd gnd cell_6t
Xbit_r58_c223 bl_223 br_223 wl_58 vdd gnd cell_6t
Xbit_r59_c223 bl_223 br_223 wl_59 vdd gnd cell_6t
Xbit_r60_c223 bl_223 br_223 wl_60 vdd gnd cell_6t
Xbit_r61_c223 bl_223 br_223 wl_61 vdd gnd cell_6t
Xbit_r62_c223 bl_223 br_223 wl_62 vdd gnd cell_6t
Xbit_r63_c223 bl_223 br_223 wl_63 vdd gnd cell_6t
Xbit_r64_c223 bl_223 br_223 wl_64 vdd gnd cell_6t
Xbit_r65_c223 bl_223 br_223 wl_65 vdd gnd cell_6t
Xbit_r66_c223 bl_223 br_223 wl_66 vdd gnd cell_6t
Xbit_r67_c223 bl_223 br_223 wl_67 vdd gnd cell_6t
Xbit_r68_c223 bl_223 br_223 wl_68 vdd gnd cell_6t
Xbit_r69_c223 bl_223 br_223 wl_69 vdd gnd cell_6t
Xbit_r70_c223 bl_223 br_223 wl_70 vdd gnd cell_6t
Xbit_r71_c223 bl_223 br_223 wl_71 vdd gnd cell_6t
Xbit_r72_c223 bl_223 br_223 wl_72 vdd gnd cell_6t
Xbit_r73_c223 bl_223 br_223 wl_73 vdd gnd cell_6t
Xbit_r74_c223 bl_223 br_223 wl_74 vdd gnd cell_6t
Xbit_r75_c223 bl_223 br_223 wl_75 vdd gnd cell_6t
Xbit_r76_c223 bl_223 br_223 wl_76 vdd gnd cell_6t
Xbit_r77_c223 bl_223 br_223 wl_77 vdd gnd cell_6t
Xbit_r78_c223 bl_223 br_223 wl_78 vdd gnd cell_6t
Xbit_r79_c223 bl_223 br_223 wl_79 vdd gnd cell_6t
Xbit_r80_c223 bl_223 br_223 wl_80 vdd gnd cell_6t
Xbit_r81_c223 bl_223 br_223 wl_81 vdd gnd cell_6t
Xbit_r82_c223 bl_223 br_223 wl_82 vdd gnd cell_6t
Xbit_r83_c223 bl_223 br_223 wl_83 vdd gnd cell_6t
Xbit_r84_c223 bl_223 br_223 wl_84 vdd gnd cell_6t
Xbit_r85_c223 bl_223 br_223 wl_85 vdd gnd cell_6t
Xbit_r86_c223 bl_223 br_223 wl_86 vdd gnd cell_6t
Xbit_r87_c223 bl_223 br_223 wl_87 vdd gnd cell_6t
Xbit_r88_c223 bl_223 br_223 wl_88 vdd gnd cell_6t
Xbit_r89_c223 bl_223 br_223 wl_89 vdd gnd cell_6t
Xbit_r90_c223 bl_223 br_223 wl_90 vdd gnd cell_6t
Xbit_r91_c223 bl_223 br_223 wl_91 vdd gnd cell_6t
Xbit_r92_c223 bl_223 br_223 wl_92 vdd gnd cell_6t
Xbit_r93_c223 bl_223 br_223 wl_93 vdd gnd cell_6t
Xbit_r94_c223 bl_223 br_223 wl_94 vdd gnd cell_6t
Xbit_r95_c223 bl_223 br_223 wl_95 vdd gnd cell_6t
Xbit_r96_c223 bl_223 br_223 wl_96 vdd gnd cell_6t
Xbit_r97_c223 bl_223 br_223 wl_97 vdd gnd cell_6t
Xbit_r98_c223 bl_223 br_223 wl_98 vdd gnd cell_6t
Xbit_r99_c223 bl_223 br_223 wl_99 vdd gnd cell_6t
Xbit_r100_c223 bl_223 br_223 wl_100 vdd gnd cell_6t
Xbit_r101_c223 bl_223 br_223 wl_101 vdd gnd cell_6t
Xbit_r102_c223 bl_223 br_223 wl_102 vdd gnd cell_6t
Xbit_r103_c223 bl_223 br_223 wl_103 vdd gnd cell_6t
Xbit_r104_c223 bl_223 br_223 wl_104 vdd gnd cell_6t
Xbit_r105_c223 bl_223 br_223 wl_105 vdd gnd cell_6t
Xbit_r106_c223 bl_223 br_223 wl_106 vdd gnd cell_6t
Xbit_r107_c223 bl_223 br_223 wl_107 vdd gnd cell_6t
Xbit_r108_c223 bl_223 br_223 wl_108 vdd gnd cell_6t
Xbit_r109_c223 bl_223 br_223 wl_109 vdd gnd cell_6t
Xbit_r110_c223 bl_223 br_223 wl_110 vdd gnd cell_6t
Xbit_r111_c223 bl_223 br_223 wl_111 vdd gnd cell_6t
Xbit_r112_c223 bl_223 br_223 wl_112 vdd gnd cell_6t
Xbit_r113_c223 bl_223 br_223 wl_113 vdd gnd cell_6t
Xbit_r114_c223 bl_223 br_223 wl_114 vdd gnd cell_6t
Xbit_r115_c223 bl_223 br_223 wl_115 vdd gnd cell_6t
Xbit_r116_c223 bl_223 br_223 wl_116 vdd gnd cell_6t
Xbit_r117_c223 bl_223 br_223 wl_117 vdd gnd cell_6t
Xbit_r118_c223 bl_223 br_223 wl_118 vdd gnd cell_6t
Xbit_r119_c223 bl_223 br_223 wl_119 vdd gnd cell_6t
Xbit_r120_c223 bl_223 br_223 wl_120 vdd gnd cell_6t
Xbit_r121_c223 bl_223 br_223 wl_121 vdd gnd cell_6t
Xbit_r122_c223 bl_223 br_223 wl_122 vdd gnd cell_6t
Xbit_r123_c223 bl_223 br_223 wl_123 vdd gnd cell_6t
Xbit_r124_c223 bl_223 br_223 wl_124 vdd gnd cell_6t
Xbit_r125_c223 bl_223 br_223 wl_125 vdd gnd cell_6t
Xbit_r126_c223 bl_223 br_223 wl_126 vdd gnd cell_6t
Xbit_r127_c223 bl_223 br_223 wl_127 vdd gnd cell_6t
Xbit_r128_c223 bl_223 br_223 wl_128 vdd gnd cell_6t
Xbit_r129_c223 bl_223 br_223 wl_129 vdd gnd cell_6t
Xbit_r130_c223 bl_223 br_223 wl_130 vdd gnd cell_6t
Xbit_r131_c223 bl_223 br_223 wl_131 vdd gnd cell_6t
Xbit_r132_c223 bl_223 br_223 wl_132 vdd gnd cell_6t
Xbit_r133_c223 bl_223 br_223 wl_133 vdd gnd cell_6t
Xbit_r134_c223 bl_223 br_223 wl_134 vdd gnd cell_6t
Xbit_r135_c223 bl_223 br_223 wl_135 vdd gnd cell_6t
Xbit_r136_c223 bl_223 br_223 wl_136 vdd gnd cell_6t
Xbit_r137_c223 bl_223 br_223 wl_137 vdd gnd cell_6t
Xbit_r138_c223 bl_223 br_223 wl_138 vdd gnd cell_6t
Xbit_r139_c223 bl_223 br_223 wl_139 vdd gnd cell_6t
Xbit_r140_c223 bl_223 br_223 wl_140 vdd gnd cell_6t
Xbit_r141_c223 bl_223 br_223 wl_141 vdd gnd cell_6t
Xbit_r142_c223 bl_223 br_223 wl_142 vdd gnd cell_6t
Xbit_r143_c223 bl_223 br_223 wl_143 vdd gnd cell_6t
Xbit_r144_c223 bl_223 br_223 wl_144 vdd gnd cell_6t
Xbit_r145_c223 bl_223 br_223 wl_145 vdd gnd cell_6t
Xbit_r146_c223 bl_223 br_223 wl_146 vdd gnd cell_6t
Xbit_r147_c223 bl_223 br_223 wl_147 vdd gnd cell_6t
Xbit_r148_c223 bl_223 br_223 wl_148 vdd gnd cell_6t
Xbit_r149_c223 bl_223 br_223 wl_149 vdd gnd cell_6t
Xbit_r150_c223 bl_223 br_223 wl_150 vdd gnd cell_6t
Xbit_r151_c223 bl_223 br_223 wl_151 vdd gnd cell_6t
Xbit_r152_c223 bl_223 br_223 wl_152 vdd gnd cell_6t
Xbit_r153_c223 bl_223 br_223 wl_153 vdd gnd cell_6t
Xbit_r154_c223 bl_223 br_223 wl_154 vdd gnd cell_6t
Xbit_r155_c223 bl_223 br_223 wl_155 vdd gnd cell_6t
Xbit_r156_c223 bl_223 br_223 wl_156 vdd gnd cell_6t
Xbit_r157_c223 bl_223 br_223 wl_157 vdd gnd cell_6t
Xbit_r158_c223 bl_223 br_223 wl_158 vdd gnd cell_6t
Xbit_r159_c223 bl_223 br_223 wl_159 vdd gnd cell_6t
Xbit_r160_c223 bl_223 br_223 wl_160 vdd gnd cell_6t
Xbit_r161_c223 bl_223 br_223 wl_161 vdd gnd cell_6t
Xbit_r162_c223 bl_223 br_223 wl_162 vdd gnd cell_6t
Xbit_r163_c223 bl_223 br_223 wl_163 vdd gnd cell_6t
Xbit_r164_c223 bl_223 br_223 wl_164 vdd gnd cell_6t
Xbit_r165_c223 bl_223 br_223 wl_165 vdd gnd cell_6t
Xbit_r166_c223 bl_223 br_223 wl_166 vdd gnd cell_6t
Xbit_r167_c223 bl_223 br_223 wl_167 vdd gnd cell_6t
Xbit_r168_c223 bl_223 br_223 wl_168 vdd gnd cell_6t
Xbit_r169_c223 bl_223 br_223 wl_169 vdd gnd cell_6t
Xbit_r170_c223 bl_223 br_223 wl_170 vdd gnd cell_6t
Xbit_r171_c223 bl_223 br_223 wl_171 vdd gnd cell_6t
Xbit_r172_c223 bl_223 br_223 wl_172 vdd gnd cell_6t
Xbit_r173_c223 bl_223 br_223 wl_173 vdd gnd cell_6t
Xbit_r174_c223 bl_223 br_223 wl_174 vdd gnd cell_6t
Xbit_r175_c223 bl_223 br_223 wl_175 vdd gnd cell_6t
Xbit_r176_c223 bl_223 br_223 wl_176 vdd gnd cell_6t
Xbit_r177_c223 bl_223 br_223 wl_177 vdd gnd cell_6t
Xbit_r178_c223 bl_223 br_223 wl_178 vdd gnd cell_6t
Xbit_r179_c223 bl_223 br_223 wl_179 vdd gnd cell_6t
Xbit_r180_c223 bl_223 br_223 wl_180 vdd gnd cell_6t
Xbit_r181_c223 bl_223 br_223 wl_181 vdd gnd cell_6t
Xbit_r182_c223 bl_223 br_223 wl_182 vdd gnd cell_6t
Xbit_r183_c223 bl_223 br_223 wl_183 vdd gnd cell_6t
Xbit_r184_c223 bl_223 br_223 wl_184 vdd gnd cell_6t
Xbit_r185_c223 bl_223 br_223 wl_185 vdd gnd cell_6t
Xbit_r186_c223 bl_223 br_223 wl_186 vdd gnd cell_6t
Xbit_r187_c223 bl_223 br_223 wl_187 vdd gnd cell_6t
Xbit_r188_c223 bl_223 br_223 wl_188 vdd gnd cell_6t
Xbit_r189_c223 bl_223 br_223 wl_189 vdd gnd cell_6t
Xbit_r190_c223 bl_223 br_223 wl_190 vdd gnd cell_6t
Xbit_r191_c223 bl_223 br_223 wl_191 vdd gnd cell_6t
Xbit_r192_c223 bl_223 br_223 wl_192 vdd gnd cell_6t
Xbit_r193_c223 bl_223 br_223 wl_193 vdd gnd cell_6t
Xbit_r194_c223 bl_223 br_223 wl_194 vdd gnd cell_6t
Xbit_r195_c223 bl_223 br_223 wl_195 vdd gnd cell_6t
Xbit_r196_c223 bl_223 br_223 wl_196 vdd gnd cell_6t
Xbit_r197_c223 bl_223 br_223 wl_197 vdd gnd cell_6t
Xbit_r198_c223 bl_223 br_223 wl_198 vdd gnd cell_6t
Xbit_r199_c223 bl_223 br_223 wl_199 vdd gnd cell_6t
Xbit_r200_c223 bl_223 br_223 wl_200 vdd gnd cell_6t
Xbit_r201_c223 bl_223 br_223 wl_201 vdd gnd cell_6t
Xbit_r202_c223 bl_223 br_223 wl_202 vdd gnd cell_6t
Xbit_r203_c223 bl_223 br_223 wl_203 vdd gnd cell_6t
Xbit_r204_c223 bl_223 br_223 wl_204 vdd gnd cell_6t
Xbit_r205_c223 bl_223 br_223 wl_205 vdd gnd cell_6t
Xbit_r206_c223 bl_223 br_223 wl_206 vdd gnd cell_6t
Xbit_r207_c223 bl_223 br_223 wl_207 vdd gnd cell_6t
Xbit_r208_c223 bl_223 br_223 wl_208 vdd gnd cell_6t
Xbit_r209_c223 bl_223 br_223 wl_209 vdd gnd cell_6t
Xbit_r210_c223 bl_223 br_223 wl_210 vdd gnd cell_6t
Xbit_r211_c223 bl_223 br_223 wl_211 vdd gnd cell_6t
Xbit_r212_c223 bl_223 br_223 wl_212 vdd gnd cell_6t
Xbit_r213_c223 bl_223 br_223 wl_213 vdd gnd cell_6t
Xbit_r214_c223 bl_223 br_223 wl_214 vdd gnd cell_6t
Xbit_r215_c223 bl_223 br_223 wl_215 vdd gnd cell_6t
Xbit_r216_c223 bl_223 br_223 wl_216 vdd gnd cell_6t
Xbit_r217_c223 bl_223 br_223 wl_217 vdd gnd cell_6t
Xbit_r218_c223 bl_223 br_223 wl_218 vdd gnd cell_6t
Xbit_r219_c223 bl_223 br_223 wl_219 vdd gnd cell_6t
Xbit_r220_c223 bl_223 br_223 wl_220 vdd gnd cell_6t
Xbit_r221_c223 bl_223 br_223 wl_221 vdd gnd cell_6t
Xbit_r222_c223 bl_223 br_223 wl_222 vdd gnd cell_6t
Xbit_r223_c223 bl_223 br_223 wl_223 vdd gnd cell_6t
Xbit_r224_c223 bl_223 br_223 wl_224 vdd gnd cell_6t
Xbit_r225_c223 bl_223 br_223 wl_225 vdd gnd cell_6t
Xbit_r226_c223 bl_223 br_223 wl_226 vdd gnd cell_6t
Xbit_r227_c223 bl_223 br_223 wl_227 vdd gnd cell_6t
Xbit_r228_c223 bl_223 br_223 wl_228 vdd gnd cell_6t
Xbit_r229_c223 bl_223 br_223 wl_229 vdd gnd cell_6t
Xbit_r230_c223 bl_223 br_223 wl_230 vdd gnd cell_6t
Xbit_r231_c223 bl_223 br_223 wl_231 vdd gnd cell_6t
Xbit_r232_c223 bl_223 br_223 wl_232 vdd gnd cell_6t
Xbit_r233_c223 bl_223 br_223 wl_233 vdd gnd cell_6t
Xbit_r234_c223 bl_223 br_223 wl_234 vdd gnd cell_6t
Xbit_r235_c223 bl_223 br_223 wl_235 vdd gnd cell_6t
Xbit_r236_c223 bl_223 br_223 wl_236 vdd gnd cell_6t
Xbit_r237_c223 bl_223 br_223 wl_237 vdd gnd cell_6t
Xbit_r238_c223 bl_223 br_223 wl_238 vdd gnd cell_6t
Xbit_r239_c223 bl_223 br_223 wl_239 vdd gnd cell_6t
Xbit_r240_c223 bl_223 br_223 wl_240 vdd gnd cell_6t
Xbit_r241_c223 bl_223 br_223 wl_241 vdd gnd cell_6t
Xbit_r242_c223 bl_223 br_223 wl_242 vdd gnd cell_6t
Xbit_r243_c223 bl_223 br_223 wl_243 vdd gnd cell_6t
Xbit_r244_c223 bl_223 br_223 wl_244 vdd gnd cell_6t
Xbit_r245_c223 bl_223 br_223 wl_245 vdd gnd cell_6t
Xbit_r246_c223 bl_223 br_223 wl_246 vdd gnd cell_6t
Xbit_r247_c223 bl_223 br_223 wl_247 vdd gnd cell_6t
Xbit_r248_c223 bl_223 br_223 wl_248 vdd gnd cell_6t
Xbit_r249_c223 bl_223 br_223 wl_249 vdd gnd cell_6t
Xbit_r250_c223 bl_223 br_223 wl_250 vdd gnd cell_6t
Xbit_r251_c223 bl_223 br_223 wl_251 vdd gnd cell_6t
Xbit_r252_c223 bl_223 br_223 wl_252 vdd gnd cell_6t
Xbit_r253_c223 bl_223 br_223 wl_253 vdd gnd cell_6t
Xbit_r254_c223 bl_223 br_223 wl_254 vdd gnd cell_6t
Xbit_r255_c223 bl_223 br_223 wl_255 vdd gnd cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd cell_6t
Xbit_r1_c224 bl_224 br_224 wl_1 vdd gnd cell_6t
Xbit_r2_c224 bl_224 br_224 wl_2 vdd gnd cell_6t
Xbit_r3_c224 bl_224 br_224 wl_3 vdd gnd cell_6t
Xbit_r4_c224 bl_224 br_224 wl_4 vdd gnd cell_6t
Xbit_r5_c224 bl_224 br_224 wl_5 vdd gnd cell_6t
Xbit_r6_c224 bl_224 br_224 wl_6 vdd gnd cell_6t
Xbit_r7_c224 bl_224 br_224 wl_7 vdd gnd cell_6t
Xbit_r8_c224 bl_224 br_224 wl_8 vdd gnd cell_6t
Xbit_r9_c224 bl_224 br_224 wl_9 vdd gnd cell_6t
Xbit_r10_c224 bl_224 br_224 wl_10 vdd gnd cell_6t
Xbit_r11_c224 bl_224 br_224 wl_11 vdd gnd cell_6t
Xbit_r12_c224 bl_224 br_224 wl_12 vdd gnd cell_6t
Xbit_r13_c224 bl_224 br_224 wl_13 vdd gnd cell_6t
Xbit_r14_c224 bl_224 br_224 wl_14 vdd gnd cell_6t
Xbit_r15_c224 bl_224 br_224 wl_15 vdd gnd cell_6t
Xbit_r16_c224 bl_224 br_224 wl_16 vdd gnd cell_6t
Xbit_r17_c224 bl_224 br_224 wl_17 vdd gnd cell_6t
Xbit_r18_c224 bl_224 br_224 wl_18 vdd gnd cell_6t
Xbit_r19_c224 bl_224 br_224 wl_19 vdd gnd cell_6t
Xbit_r20_c224 bl_224 br_224 wl_20 vdd gnd cell_6t
Xbit_r21_c224 bl_224 br_224 wl_21 vdd gnd cell_6t
Xbit_r22_c224 bl_224 br_224 wl_22 vdd gnd cell_6t
Xbit_r23_c224 bl_224 br_224 wl_23 vdd gnd cell_6t
Xbit_r24_c224 bl_224 br_224 wl_24 vdd gnd cell_6t
Xbit_r25_c224 bl_224 br_224 wl_25 vdd gnd cell_6t
Xbit_r26_c224 bl_224 br_224 wl_26 vdd gnd cell_6t
Xbit_r27_c224 bl_224 br_224 wl_27 vdd gnd cell_6t
Xbit_r28_c224 bl_224 br_224 wl_28 vdd gnd cell_6t
Xbit_r29_c224 bl_224 br_224 wl_29 vdd gnd cell_6t
Xbit_r30_c224 bl_224 br_224 wl_30 vdd gnd cell_6t
Xbit_r31_c224 bl_224 br_224 wl_31 vdd gnd cell_6t
Xbit_r32_c224 bl_224 br_224 wl_32 vdd gnd cell_6t
Xbit_r33_c224 bl_224 br_224 wl_33 vdd gnd cell_6t
Xbit_r34_c224 bl_224 br_224 wl_34 vdd gnd cell_6t
Xbit_r35_c224 bl_224 br_224 wl_35 vdd gnd cell_6t
Xbit_r36_c224 bl_224 br_224 wl_36 vdd gnd cell_6t
Xbit_r37_c224 bl_224 br_224 wl_37 vdd gnd cell_6t
Xbit_r38_c224 bl_224 br_224 wl_38 vdd gnd cell_6t
Xbit_r39_c224 bl_224 br_224 wl_39 vdd gnd cell_6t
Xbit_r40_c224 bl_224 br_224 wl_40 vdd gnd cell_6t
Xbit_r41_c224 bl_224 br_224 wl_41 vdd gnd cell_6t
Xbit_r42_c224 bl_224 br_224 wl_42 vdd gnd cell_6t
Xbit_r43_c224 bl_224 br_224 wl_43 vdd gnd cell_6t
Xbit_r44_c224 bl_224 br_224 wl_44 vdd gnd cell_6t
Xbit_r45_c224 bl_224 br_224 wl_45 vdd gnd cell_6t
Xbit_r46_c224 bl_224 br_224 wl_46 vdd gnd cell_6t
Xbit_r47_c224 bl_224 br_224 wl_47 vdd gnd cell_6t
Xbit_r48_c224 bl_224 br_224 wl_48 vdd gnd cell_6t
Xbit_r49_c224 bl_224 br_224 wl_49 vdd gnd cell_6t
Xbit_r50_c224 bl_224 br_224 wl_50 vdd gnd cell_6t
Xbit_r51_c224 bl_224 br_224 wl_51 vdd gnd cell_6t
Xbit_r52_c224 bl_224 br_224 wl_52 vdd gnd cell_6t
Xbit_r53_c224 bl_224 br_224 wl_53 vdd gnd cell_6t
Xbit_r54_c224 bl_224 br_224 wl_54 vdd gnd cell_6t
Xbit_r55_c224 bl_224 br_224 wl_55 vdd gnd cell_6t
Xbit_r56_c224 bl_224 br_224 wl_56 vdd gnd cell_6t
Xbit_r57_c224 bl_224 br_224 wl_57 vdd gnd cell_6t
Xbit_r58_c224 bl_224 br_224 wl_58 vdd gnd cell_6t
Xbit_r59_c224 bl_224 br_224 wl_59 vdd gnd cell_6t
Xbit_r60_c224 bl_224 br_224 wl_60 vdd gnd cell_6t
Xbit_r61_c224 bl_224 br_224 wl_61 vdd gnd cell_6t
Xbit_r62_c224 bl_224 br_224 wl_62 vdd gnd cell_6t
Xbit_r63_c224 bl_224 br_224 wl_63 vdd gnd cell_6t
Xbit_r64_c224 bl_224 br_224 wl_64 vdd gnd cell_6t
Xbit_r65_c224 bl_224 br_224 wl_65 vdd gnd cell_6t
Xbit_r66_c224 bl_224 br_224 wl_66 vdd gnd cell_6t
Xbit_r67_c224 bl_224 br_224 wl_67 vdd gnd cell_6t
Xbit_r68_c224 bl_224 br_224 wl_68 vdd gnd cell_6t
Xbit_r69_c224 bl_224 br_224 wl_69 vdd gnd cell_6t
Xbit_r70_c224 bl_224 br_224 wl_70 vdd gnd cell_6t
Xbit_r71_c224 bl_224 br_224 wl_71 vdd gnd cell_6t
Xbit_r72_c224 bl_224 br_224 wl_72 vdd gnd cell_6t
Xbit_r73_c224 bl_224 br_224 wl_73 vdd gnd cell_6t
Xbit_r74_c224 bl_224 br_224 wl_74 vdd gnd cell_6t
Xbit_r75_c224 bl_224 br_224 wl_75 vdd gnd cell_6t
Xbit_r76_c224 bl_224 br_224 wl_76 vdd gnd cell_6t
Xbit_r77_c224 bl_224 br_224 wl_77 vdd gnd cell_6t
Xbit_r78_c224 bl_224 br_224 wl_78 vdd gnd cell_6t
Xbit_r79_c224 bl_224 br_224 wl_79 vdd gnd cell_6t
Xbit_r80_c224 bl_224 br_224 wl_80 vdd gnd cell_6t
Xbit_r81_c224 bl_224 br_224 wl_81 vdd gnd cell_6t
Xbit_r82_c224 bl_224 br_224 wl_82 vdd gnd cell_6t
Xbit_r83_c224 bl_224 br_224 wl_83 vdd gnd cell_6t
Xbit_r84_c224 bl_224 br_224 wl_84 vdd gnd cell_6t
Xbit_r85_c224 bl_224 br_224 wl_85 vdd gnd cell_6t
Xbit_r86_c224 bl_224 br_224 wl_86 vdd gnd cell_6t
Xbit_r87_c224 bl_224 br_224 wl_87 vdd gnd cell_6t
Xbit_r88_c224 bl_224 br_224 wl_88 vdd gnd cell_6t
Xbit_r89_c224 bl_224 br_224 wl_89 vdd gnd cell_6t
Xbit_r90_c224 bl_224 br_224 wl_90 vdd gnd cell_6t
Xbit_r91_c224 bl_224 br_224 wl_91 vdd gnd cell_6t
Xbit_r92_c224 bl_224 br_224 wl_92 vdd gnd cell_6t
Xbit_r93_c224 bl_224 br_224 wl_93 vdd gnd cell_6t
Xbit_r94_c224 bl_224 br_224 wl_94 vdd gnd cell_6t
Xbit_r95_c224 bl_224 br_224 wl_95 vdd gnd cell_6t
Xbit_r96_c224 bl_224 br_224 wl_96 vdd gnd cell_6t
Xbit_r97_c224 bl_224 br_224 wl_97 vdd gnd cell_6t
Xbit_r98_c224 bl_224 br_224 wl_98 vdd gnd cell_6t
Xbit_r99_c224 bl_224 br_224 wl_99 vdd gnd cell_6t
Xbit_r100_c224 bl_224 br_224 wl_100 vdd gnd cell_6t
Xbit_r101_c224 bl_224 br_224 wl_101 vdd gnd cell_6t
Xbit_r102_c224 bl_224 br_224 wl_102 vdd gnd cell_6t
Xbit_r103_c224 bl_224 br_224 wl_103 vdd gnd cell_6t
Xbit_r104_c224 bl_224 br_224 wl_104 vdd gnd cell_6t
Xbit_r105_c224 bl_224 br_224 wl_105 vdd gnd cell_6t
Xbit_r106_c224 bl_224 br_224 wl_106 vdd gnd cell_6t
Xbit_r107_c224 bl_224 br_224 wl_107 vdd gnd cell_6t
Xbit_r108_c224 bl_224 br_224 wl_108 vdd gnd cell_6t
Xbit_r109_c224 bl_224 br_224 wl_109 vdd gnd cell_6t
Xbit_r110_c224 bl_224 br_224 wl_110 vdd gnd cell_6t
Xbit_r111_c224 bl_224 br_224 wl_111 vdd gnd cell_6t
Xbit_r112_c224 bl_224 br_224 wl_112 vdd gnd cell_6t
Xbit_r113_c224 bl_224 br_224 wl_113 vdd gnd cell_6t
Xbit_r114_c224 bl_224 br_224 wl_114 vdd gnd cell_6t
Xbit_r115_c224 bl_224 br_224 wl_115 vdd gnd cell_6t
Xbit_r116_c224 bl_224 br_224 wl_116 vdd gnd cell_6t
Xbit_r117_c224 bl_224 br_224 wl_117 vdd gnd cell_6t
Xbit_r118_c224 bl_224 br_224 wl_118 vdd gnd cell_6t
Xbit_r119_c224 bl_224 br_224 wl_119 vdd gnd cell_6t
Xbit_r120_c224 bl_224 br_224 wl_120 vdd gnd cell_6t
Xbit_r121_c224 bl_224 br_224 wl_121 vdd gnd cell_6t
Xbit_r122_c224 bl_224 br_224 wl_122 vdd gnd cell_6t
Xbit_r123_c224 bl_224 br_224 wl_123 vdd gnd cell_6t
Xbit_r124_c224 bl_224 br_224 wl_124 vdd gnd cell_6t
Xbit_r125_c224 bl_224 br_224 wl_125 vdd gnd cell_6t
Xbit_r126_c224 bl_224 br_224 wl_126 vdd gnd cell_6t
Xbit_r127_c224 bl_224 br_224 wl_127 vdd gnd cell_6t
Xbit_r128_c224 bl_224 br_224 wl_128 vdd gnd cell_6t
Xbit_r129_c224 bl_224 br_224 wl_129 vdd gnd cell_6t
Xbit_r130_c224 bl_224 br_224 wl_130 vdd gnd cell_6t
Xbit_r131_c224 bl_224 br_224 wl_131 vdd gnd cell_6t
Xbit_r132_c224 bl_224 br_224 wl_132 vdd gnd cell_6t
Xbit_r133_c224 bl_224 br_224 wl_133 vdd gnd cell_6t
Xbit_r134_c224 bl_224 br_224 wl_134 vdd gnd cell_6t
Xbit_r135_c224 bl_224 br_224 wl_135 vdd gnd cell_6t
Xbit_r136_c224 bl_224 br_224 wl_136 vdd gnd cell_6t
Xbit_r137_c224 bl_224 br_224 wl_137 vdd gnd cell_6t
Xbit_r138_c224 bl_224 br_224 wl_138 vdd gnd cell_6t
Xbit_r139_c224 bl_224 br_224 wl_139 vdd gnd cell_6t
Xbit_r140_c224 bl_224 br_224 wl_140 vdd gnd cell_6t
Xbit_r141_c224 bl_224 br_224 wl_141 vdd gnd cell_6t
Xbit_r142_c224 bl_224 br_224 wl_142 vdd gnd cell_6t
Xbit_r143_c224 bl_224 br_224 wl_143 vdd gnd cell_6t
Xbit_r144_c224 bl_224 br_224 wl_144 vdd gnd cell_6t
Xbit_r145_c224 bl_224 br_224 wl_145 vdd gnd cell_6t
Xbit_r146_c224 bl_224 br_224 wl_146 vdd gnd cell_6t
Xbit_r147_c224 bl_224 br_224 wl_147 vdd gnd cell_6t
Xbit_r148_c224 bl_224 br_224 wl_148 vdd gnd cell_6t
Xbit_r149_c224 bl_224 br_224 wl_149 vdd gnd cell_6t
Xbit_r150_c224 bl_224 br_224 wl_150 vdd gnd cell_6t
Xbit_r151_c224 bl_224 br_224 wl_151 vdd gnd cell_6t
Xbit_r152_c224 bl_224 br_224 wl_152 vdd gnd cell_6t
Xbit_r153_c224 bl_224 br_224 wl_153 vdd gnd cell_6t
Xbit_r154_c224 bl_224 br_224 wl_154 vdd gnd cell_6t
Xbit_r155_c224 bl_224 br_224 wl_155 vdd gnd cell_6t
Xbit_r156_c224 bl_224 br_224 wl_156 vdd gnd cell_6t
Xbit_r157_c224 bl_224 br_224 wl_157 vdd gnd cell_6t
Xbit_r158_c224 bl_224 br_224 wl_158 vdd gnd cell_6t
Xbit_r159_c224 bl_224 br_224 wl_159 vdd gnd cell_6t
Xbit_r160_c224 bl_224 br_224 wl_160 vdd gnd cell_6t
Xbit_r161_c224 bl_224 br_224 wl_161 vdd gnd cell_6t
Xbit_r162_c224 bl_224 br_224 wl_162 vdd gnd cell_6t
Xbit_r163_c224 bl_224 br_224 wl_163 vdd gnd cell_6t
Xbit_r164_c224 bl_224 br_224 wl_164 vdd gnd cell_6t
Xbit_r165_c224 bl_224 br_224 wl_165 vdd gnd cell_6t
Xbit_r166_c224 bl_224 br_224 wl_166 vdd gnd cell_6t
Xbit_r167_c224 bl_224 br_224 wl_167 vdd gnd cell_6t
Xbit_r168_c224 bl_224 br_224 wl_168 vdd gnd cell_6t
Xbit_r169_c224 bl_224 br_224 wl_169 vdd gnd cell_6t
Xbit_r170_c224 bl_224 br_224 wl_170 vdd gnd cell_6t
Xbit_r171_c224 bl_224 br_224 wl_171 vdd gnd cell_6t
Xbit_r172_c224 bl_224 br_224 wl_172 vdd gnd cell_6t
Xbit_r173_c224 bl_224 br_224 wl_173 vdd gnd cell_6t
Xbit_r174_c224 bl_224 br_224 wl_174 vdd gnd cell_6t
Xbit_r175_c224 bl_224 br_224 wl_175 vdd gnd cell_6t
Xbit_r176_c224 bl_224 br_224 wl_176 vdd gnd cell_6t
Xbit_r177_c224 bl_224 br_224 wl_177 vdd gnd cell_6t
Xbit_r178_c224 bl_224 br_224 wl_178 vdd gnd cell_6t
Xbit_r179_c224 bl_224 br_224 wl_179 vdd gnd cell_6t
Xbit_r180_c224 bl_224 br_224 wl_180 vdd gnd cell_6t
Xbit_r181_c224 bl_224 br_224 wl_181 vdd gnd cell_6t
Xbit_r182_c224 bl_224 br_224 wl_182 vdd gnd cell_6t
Xbit_r183_c224 bl_224 br_224 wl_183 vdd gnd cell_6t
Xbit_r184_c224 bl_224 br_224 wl_184 vdd gnd cell_6t
Xbit_r185_c224 bl_224 br_224 wl_185 vdd gnd cell_6t
Xbit_r186_c224 bl_224 br_224 wl_186 vdd gnd cell_6t
Xbit_r187_c224 bl_224 br_224 wl_187 vdd gnd cell_6t
Xbit_r188_c224 bl_224 br_224 wl_188 vdd gnd cell_6t
Xbit_r189_c224 bl_224 br_224 wl_189 vdd gnd cell_6t
Xbit_r190_c224 bl_224 br_224 wl_190 vdd gnd cell_6t
Xbit_r191_c224 bl_224 br_224 wl_191 vdd gnd cell_6t
Xbit_r192_c224 bl_224 br_224 wl_192 vdd gnd cell_6t
Xbit_r193_c224 bl_224 br_224 wl_193 vdd gnd cell_6t
Xbit_r194_c224 bl_224 br_224 wl_194 vdd gnd cell_6t
Xbit_r195_c224 bl_224 br_224 wl_195 vdd gnd cell_6t
Xbit_r196_c224 bl_224 br_224 wl_196 vdd gnd cell_6t
Xbit_r197_c224 bl_224 br_224 wl_197 vdd gnd cell_6t
Xbit_r198_c224 bl_224 br_224 wl_198 vdd gnd cell_6t
Xbit_r199_c224 bl_224 br_224 wl_199 vdd gnd cell_6t
Xbit_r200_c224 bl_224 br_224 wl_200 vdd gnd cell_6t
Xbit_r201_c224 bl_224 br_224 wl_201 vdd gnd cell_6t
Xbit_r202_c224 bl_224 br_224 wl_202 vdd gnd cell_6t
Xbit_r203_c224 bl_224 br_224 wl_203 vdd gnd cell_6t
Xbit_r204_c224 bl_224 br_224 wl_204 vdd gnd cell_6t
Xbit_r205_c224 bl_224 br_224 wl_205 vdd gnd cell_6t
Xbit_r206_c224 bl_224 br_224 wl_206 vdd gnd cell_6t
Xbit_r207_c224 bl_224 br_224 wl_207 vdd gnd cell_6t
Xbit_r208_c224 bl_224 br_224 wl_208 vdd gnd cell_6t
Xbit_r209_c224 bl_224 br_224 wl_209 vdd gnd cell_6t
Xbit_r210_c224 bl_224 br_224 wl_210 vdd gnd cell_6t
Xbit_r211_c224 bl_224 br_224 wl_211 vdd gnd cell_6t
Xbit_r212_c224 bl_224 br_224 wl_212 vdd gnd cell_6t
Xbit_r213_c224 bl_224 br_224 wl_213 vdd gnd cell_6t
Xbit_r214_c224 bl_224 br_224 wl_214 vdd gnd cell_6t
Xbit_r215_c224 bl_224 br_224 wl_215 vdd gnd cell_6t
Xbit_r216_c224 bl_224 br_224 wl_216 vdd gnd cell_6t
Xbit_r217_c224 bl_224 br_224 wl_217 vdd gnd cell_6t
Xbit_r218_c224 bl_224 br_224 wl_218 vdd gnd cell_6t
Xbit_r219_c224 bl_224 br_224 wl_219 vdd gnd cell_6t
Xbit_r220_c224 bl_224 br_224 wl_220 vdd gnd cell_6t
Xbit_r221_c224 bl_224 br_224 wl_221 vdd gnd cell_6t
Xbit_r222_c224 bl_224 br_224 wl_222 vdd gnd cell_6t
Xbit_r223_c224 bl_224 br_224 wl_223 vdd gnd cell_6t
Xbit_r224_c224 bl_224 br_224 wl_224 vdd gnd cell_6t
Xbit_r225_c224 bl_224 br_224 wl_225 vdd gnd cell_6t
Xbit_r226_c224 bl_224 br_224 wl_226 vdd gnd cell_6t
Xbit_r227_c224 bl_224 br_224 wl_227 vdd gnd cell_6t
Xbit_r228_c224 bl_224 br_224 wl_228 vdd gnd cell_6t
Xbit_r229_c224 bl_224 br_224 wl_229 vdd gnd cell_6t
Xbit_r230_c224 bl_224 br_224 wl_230 vdd gnd cell_6t
Xbit_r231_c224 bl_224 br_224 wl_231 vdd gnd cell_6t
Xbit_r232_c224 bl_224 br_224 wl_232 vdd gnd cell_6t
Xbit_r233_c224 bl_224 br_224 wl_233 vdd gnd cell_6t
Xbit_r234_c224 bl_224 br_224 wl_234 vdd gnd cell_6t
Xbit_r235_c224 bl_224 br_224 wl_235 vdd gnd cell_6t
Xbit_r236_c224 bl_224 br_224 wl_236 vdd gnd cell_6t
Xbit_r237_c224 bl_224 br_224 wl_237 vdd gnd cell_6t
Xbit_r238_c224 bl_224 br_224 wl_238 vdd gnd cell_6t
Xbit_r239_c224 bl_224 br_224 wl_239 vdd gnd cell_6t
Xbit_r240_c224 bl_224 br_224 wl_240 vdd gnd cell_6t
Xbit_r241_c224 bl_224 br_224 wl_241 vdd gnd cell_6t
Xbit_r242_c224 bl_224 br_224 wl_242 vdd gnd cell_6t
Xbit_r243_c224 bl_224 br_224 wl_243 vdd gnd cell_6t
Xbit_r244_c224 bl_224 br_224 wl_244 vdd gnd cell_6t
Xbit_r245_c224 bl_224 br_224 wl_245 vdd gnd cell_6t
Xbit_r246_c224 bl_224 br_224 wl_246 vdd gnd cell_6t
Xbit_r247_c224 bl_224 br_224 wl_247 vdd gnd cell_6t
Xbit_r248_c224 bl_224 br_224 wl_248 vdd gnd cell_6t
Xbit_r249_c224 bl_224 br_224 wl_249 vdd gnd cell_6t
Xbit_r250_c224 bl_224 br_224 wl_250 vdd gnd cell_6t
Xbit_r251_c224 bl_224 br_224 wl_251 vdd gnd cell_6t
Xbit_r252_c224 bl_224 br_224 wl_252 vdd gnd cell_6t
Xbit_r253_c224 bl_224 br_224 wl_253 vdd gnd cell_6t
Xbit_r254_c224 bl_224 br_224 wl_254 vdd gnd cell_6t
Xbit_r255_c224 bl_224 br_224 wl_255 vdd gnd cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd cell_6t
Xbit_r1_c225 bl_225 br_225 wl_1 vdd gnd cell_6t
Xbit_r2_c225 bl_225 br_225 wl_2 vdd gnd cell_6t
Xbit_r3_c225 bl_225 br_225 wl_3 vdd gnd cell_6t
Xbit_r4_c225 bl_225 br_225 wl_4 vdd gnd cell_6t
Xbit_r5_c225 bl_225 br_225 wl_5 vdd gnd cell_6t
Xbit_r6_c225 bl_225 br_225 wl_6 vdd gnd cell_6t
Xbit_r7_c225 bl_225 br_225 wl_7 vdd gnd cell_6t
Xbit_r8_c225 bl_225 br_225 wl_8 vdd gnd cell_6t
Xbit_r9_c225 bl_225 br_225 wl_9 vdd gnd cell_6t
Xbit_r10_c225 bl_225 br_225 wl_10 vdd gnd cell_6t
Xbit_r11_c225 bl_225 br_225 wl_11 vdd gnd cell_6t
Xbit_r12_c225 bl_225 br_225 wl_12 vdd gnd cell_6t
Xbit_r13_c225 bl_225 br_225 wl_13 vdd gnd cell_6t
Xbit_r14_c225 bl_225 br_225 wl_14 vdd gnd cell_6t
Xbit_r15_c225 bl_225 br_225 wl_15 vdd gnd cell_6t
Xbit_r16_c225 bl_225 br_225 wl_16 vdd gnd cell_6t
Xbit_r17_c225 bl_225 br_225 wl_17 vdd gnd cell_6t
Xbit_r18_c225 bl_225 br_225 wl_18 vdd gnd cell_6t
Xbit_r19_c225 bl_225 br_225 wl_19 vdd gnd cell_6t
Xbit_r20_c225 bl_225 br_225 wl_20 vdd gnd cell_6t
Xbit_r21_c225 bl_225 br_225 wl_21 vdd gnd cell_6t
Xbit_r22_c225 bl_225 br_225 wl_22 vdd gnd cell_6t
Xbit_r23_c225 bl_225 br_225 wl_23 vdd gnd cell_6t
Xbit_r24_c225 bl_225 br_225 wl_24 vdd gnd cell_6t
Xbit_r25_c225 bl_225 br_225 wl_25 vdd gnd cell_6t
Xbit_r26_c225 bl_225 br_225 wl_26 vdd gnd cell_6t
Xbit_r27_c225 bl_225 br_225 wl_27 vdd gnd cell_6t
Xbit_r28_c225 bl_225 br_225 wl_28 vdd gnd cell_6t
Xbit_r29_c225 bl_225 br_225 wl_29 vdd gnd cell_6t
Xbit_r30_c225 bl_225 br_225 wl_30 vdd gnd cell_6t
Xbit_r31_c225 bl_225 br_225 wl_31 vdd gnd cell_6t
Xbit_r32_c225 bl_225 br_225 wl_32 vdd gnd cell_6t
Xbit_r33_c225 bl_225 br_225 wl_33 vdd gnd cell_6t
Xbit_r34_c225 bl_225 br_225 wl_34 vdd gnd cell_6t
Xbit_r35_c225 bl_225 br_225 wl_35 vdd gnd cell_6t
Xbit_r36_c225 bl_225 br_225 wl_36 vdd gnd cell_6t
Xbit_r37_c225 bl_225 br_225 wl_37 vdd gnd cell_6t
Xbit_r38_c225 bl_225 br_225 wl_38 vdd gnd cell_6t
Xbit_r39_c225 bl_225 br_225 wl_39 vdd gnd cell_6t
Xbit_r40_c225 bl_225 br_225 wl_40 vdd gnd cell_6t
Xbit_r41_c225 bl_225 br_225 wl_41 vdd gnd cell_6t
Xbit_r42_c225 bl_225 br_225 wl_42 vdd gnd cell_6t
Xbit_r43_c225 bl_225 br_225 wl_43 vdd gnd cell_6t
Xbit_r44_c225 bl_225 br_225 wl_44 vdd gnd cell_6t
Xbit_r45_c225 bl_225 br_225 wl_45 vdd gnd cell_6t
Xbit_r46_c225 bl_225 br_225 wl_46 vdd gnd cell_6t
Xbit_r47_c225 bl_225 br_225 wl_47 vdd gnd cell_6t
Xbit_r48_c225 bl_225 br_225 wl_48 vdd gnd cell_6t
Xbit_r49_c225 bl_225 br_225 wl_49 vdd gnd cell_6t
Xbit_r50_c225 bl_225 br_225 wl_50 vdd gnd cell_6t
Xbit_r51_c225 bl_225 br_225 wl_51 vdd gnd cell_6t
Xbit_r52_c225 bl_225 br_225 wl_52 vdd gnd cell_6t
Xbit_r53_c225 bl_225 br_225 wl_53 vdd gnd cell_6t
Xbit_r54_c225 bl_225 br_225 wl_54 vdd gnd cell_6t
Xbit_r55_c225 bl_225 br_225 wl_55 vdd gnd cell_6t
Xbit_r56_c225 bl_225 br_225 wl_56 vdd gnd cell_6t
Xbit_r57_c225 bl_225 br_225 wl_57 vdd gnd cell_6t
Xbit_r58_c225 bl_225 br_225 wl_58 vdd gnd cell_6t
Xbit_r59_c225 bl_225 br_225 wl_59 vdd gnd cell_6t
Xbit_r60_c225 bl_225 br_225 wl_60 vdd gnd cell_6t
Xbit_r61_c225 bl_225 br_225 wl_61 vdd gnd cell_6t
Xbit_r62_c225 bl_225 br_225 wl_62 vdd gnd cell_6t
Xbit_r63_c225 bl_225 br_225 wl_63 vdd gnd cell_6t
Xbit_r64_c225 bl_225 br_225 wl_64 vdd gnd cell_6t
Xbit_r65_c225 bl_225 br_225 wl_65 vdd gnd cell_6t
Xbit_r66_c225 bl_225 br_225 wl_66 vdd gnd cell_6t
Xbit_r67_c225 bl_225 br_225 wl_67 vdd gnd cell_6t
Xbit_r68_c225 bl_225 br_225 wl_68 vdd gnd cell_6t
Xbit_r69_c225 bl_225 br_225 wl_69 vdd gnd cell_6t
Xbit_r70_c225 bl_225 br_225 wl_70 vdd gnd cell_6t
Xbit_r71_c225 bl_225 br_225 wl_71 vdd gnd cell_6t
Xbit_r72_c225 bl_225 br_225 wl_72 vdd gnd cell_6t
Xbit_r73_c225 bl_225 br_225 wl_73 vdd gnd cell_6t
Xbit_r74_c225 bl_225 br_225 wl_74 vdd gnd cell_6t
Xbit_r75_c225 bl_225 br_225 wl_75 vdd gnd cell_6t
Xbit_r76_c225 bl_225 br_225 wl_76 vdd gnd cell_6t
Xbit_r77_c225 bl_225 br_225 wl_77 vdd gnd cell_6t
Xbit_r78_c225 bl_225 br_225 wl_78 vdd gnd cell_6t
Xbit_r79_c225 bl_225 br_225 wl_79 vdd gnd cell_6t
Xbit_r80_c225 bl_225 br_225 wl_80 vdd gnd cell_6t
Xbit_r81_c225 bl_225 br_225 wl_81 vdd gnd cell_6t
Xbit_r82_c225 bl_225 br_225 wl_82 vdd gnd cell_6t
Xbit_r83_c225 bl_225 br_225 wl_83 vdd gnd cell_6t
Xbit_r84_c225 bl_225 br_225 wl_84 vdd gnd cell_6t
Xbit_r85_c225 bl_225 br_225 wl_85 vdd gnd cell_6t
Xbit_r86_c225 bl_225 br_225 wl_86 vdd gnd cell_6t
Xbit_r87_c225 bl_225 br_225 wl_87 vdd gnd cell_6t
Xbit_r88_c225 bl_225 br_225 wl_88 vdd gnd cell_6t
Xbit_r89_c225 bl_225 br_225 wl_89 vdd gnd cell_6t
Xbit_r90_c225 bl_225 br_225 wl_90 vdd gnd cell_6t
Xbit_r91_c225 bl_225 br_225 wl_91 vdd gnd cell_6t
Xbit_r92_c225 bl_225 br_225 wl_92 vdd gnd cell_6t
Xbit_r93_c225 bl_225 br_225 wl_93 vdd gnd cell_6t
Xbit_r94_c225 bl_225 br_225 wl_94 vdd gnd cell_6t
Xbit_r95_c225 bl_225 br_225 wl_95 vdd gnd cell_6t
Xbit_r96_c225 bl_225 br_225 wl_96 vdd gnd cell_6t
Xbit_r97_c225 bl_225 br_225 wl_97 vdd gnd cell_6t
Xbit_r98_c225 bl_225 br_225 wl_98 vdd gnd cell_6t
Xbit_r99_c225 bl_225 br_225 wl_99 vdd gnd cell_6t
Xbit_r100_c225 bl_225 br_225 wl_100 vdd gnd cell_6t
Xbit_r101_c225 bl_225 br_225 wl_101 vdd gnd cell_6t
Xbit_r102_c225 bl_225 br_225 wl_102 vdd gnd cell_6t
Xbit_r103_c225 bl_225 br_225 wl_103 vdd gnd cell_6t
Xbit_r104_c225 bl_225 br_225 wl_104 vdd gnd cell_6t
Xbit_r105_c225 bl_225 br_225 wl_105 vdd gnd cell_6t
Xbit_r106_c225 bl_225 br_225 wl_106 vdd gnd cell_6t
Xbit_r107_c225 bl_225 br_225 wl_107 vdd gnd cell_6t
Xbit_r108_c225 bl_225 br_225 wl_108 vdd gnd cell_6t
Xbit_r109_c225 bl_225 br_225 wl_109 vdd gnd cell_6t
Xbit_r110_c225 bl_225 br_225 wl_110 vdd gnd cell_6t
Xbit_r111_c225 bl_225 br_225 wl_111 vdd gnd cell_6t
Xbit_r112_c225 bl_225 br_225 wl_112 vdd gnd cell_6t
Xbit_r113_c225 bl_225 br_225 wl_113 vdd gnd cell_6t
Xbit_r114_c225 bl_225 br_225 wl_114 vdd gnd cell_6t
Xbit_r115_c225 bl_225 br_225 wl_115 vdd gnd cell_6t
Xbit_r116_c225 bl_225 br_225 wl_116 vdd gnd cell_6t
Xbit_r117_c225 bl_225 br_225 wl_117 vdd gnd cell_6t
Xbit_r118_c225 bl_225 br_225 wl_118 vdd gnd cell_6t
Xbit_r119_c225 bl_225 br_225 wl_119 vdd gnd cell_6t
Xbit_r120_c225 bl_225 br_225 wl_120 vdd gnd cell_6t
Xbit_r121_c225 bl_225 br_225 wl_121 vdd gnd cell_6t
Xbit_r122_c225 bl_225 br_225 wl_122 vdd gnd cell_6t
Xbit_r123_c225 bl_225 br_225 wl_123 vdd gnd cell_6t
Xbit_r124_c225 bl_225 br_225 wl_124 vdd gnd cell_6t
Xbit_r125_c225 bl_225 br_225 wl_125 vdd gnd cell_6t
Xbit_r126_c225 bl_225 br_225 wl_126 vdd gnd cell_6t
Xbit_r127_c225 bl_225 br_225 wl_127 vdd gnd cell_6t
Xbit_r128_c225 bl_225 br_225 wl_128 vdd gnd cell_6t
Xbit_r129_c225 bl_225 br_225 wl_129 vdd gnd cell_6t
Xbit_r130_c225 bl_225 br_225 wl_130 vdd gnd cell_6t
Xbit_r131_c225 bl_225 br_225 wl_131 vdd gnd cell_6t
Xbit_r132_c225 bl_225 br_225 wl_132 vdd gnd cell_6t
Xbit_r133_c225 bl_225 br_225 wl_133 vdd gnd cell_6t
Xbit_r134_c225 bl_225 br_225 wl_134 vdd gnd cell_6t
Xbit_r135_c225 bl_225 br_225 wl_135 vdd gnd cell_6t
Xbit_r136_c225 bl_225 br_225 wl_136 vdd gnd cell_6t
Xbit_r137_c225 bl_225 br_225 wl_137 vdd gnd cell_6t
Xbit_r138_c225 bl_225 br_225 wl_138 vdd gnd cell_6t
Xbit_r139_c225 bl_225 br_225 wl_139 vdd gnd cell_6t
Xbit_r140_c225 bl_225 br_225 wl_140 vdd gnd cell_6t
Xbit_r141_c225 bl_225 br_225 wl_141 vdd gnd cell_6t
Xbit_r142_c225 bl_225 br_225 wl_142 vdd gnd cell_6t
Xbit_r143_c225 bl_225 br_225 wl_143 vdd gnd cell_6t
Xbit_r144_c225 bl_225 br_225 wl_144 vdd gnd cell_6t
Xbit_r145_c225 bl_225 br_225 wl_145 vdd gnd cell_6t
Xbit_r146_c225 bl_225 br_225 wl_146 vdd gnd cell_6t
Xbit_r147_c225 bl_225 br_225 wl_147 vdd gnd cell_6t
Xbit_r148_c225 bl_225 br_225 wl_148 vdd gnd cell_6t
Xbit_r149_c225 bl_225 br_225 wl_149 vdd gnd cell_6t
Xbit_r150_c225 bl_225 br_225 wl_150 vdd gnd cell_6t
Xbit_r151_c225 bl_225 br_225 wl_151 vdd gnd cell_6t
Xbit_r152_c225 bl_225 br_225 wl_152 vdd gnd cell_6t
Xbit_r153_c225 bl_225 br_225 wl_153 vdd gnd cell_6t
Xbit_r154_c225 bl_225 br_225 wl_154 vdd gnd cell_6t
Xbit_r155_c225 bl_225 br_225 wl_155 vdd gnd cell_6t
Xbit_r156_c225 bl_225 br_225 wl_156 vdd gnd cell_6t
Xbit_r157_c225 bl_225 br_225 wl_157 vdd gnd cell_6t
Xbit_r158_c225 bl_225 br_225 wl_158 vdd gnd cell_6t
Xbit_r159_c225 bl_225 br_225 wl_159 vdd gnd cell_6t
Xbit_r160_c225 bl_225 br_225 wl_160 vdd gnd cell_6t
Xbit_r161_c225 bl_225 br_225 wl_161 vdd gnd cell_6t
Xbit_r162_c225 bl_225 br_225 wl_162 vdd gnd cell_6t
Xbit_r163_c225 bl_225 br_225 wl_163 vdd gnd cell_6t
Xbit_r164_c225 bl_225 br_225 wl_164 vdd gnd cell_6t
Xbit_r165_c225 bl_225 br_225 wl_165 vdd gnd cell_6t
Xbit_r166_c225 bl_225 br_225 wl_166 vdd gnd cell_6t
Xbit_r167_c225 bl_225 br_225 wl_167 vdd gnd cell_6t
Xbit_r168_c225 bl_225 br_225 wl_168 vdd gnd cell_6t
Xbit_r169_c225 bl_225 br_225 wl_169 vdd gnd cell_6t
Xbit_r170_c225 bl_225 br_225 wl_170 vdd gnd cell_6t
Xbit_r171_c225 bl_225 br_225 wl_171 vdd gnd cell_6t
Xbit_r172_c225 bl_225 br_225 wl_172 vdd gnd cell_6t
Xbit_r173_c225 bl_225 br_225 wl_173 vdd gnd cell_6t
Xbit_r174_c225 bl_225 br_225 wl_174 vdd gnd cell_6t
Xbit_r175_c225 bl_225 br_225 wl_175 vdd gnd cell_6t
Xbit_r176_c225 bl_225 br_225 wl_176 vdd gnd cell_6t
Xbit_r177_c225 bl_225 br_225 wl_177 vdd gnd cell_6t
Xbit_r178_c225 bl_225 br_225 wl_178 vdd gnd cell_6t
Xbit_r179_c225 bl_225 br_225 wl_179 vdd gnd cell_6t
Xbit_r180_c225 bl_225 br_225 wl_180 vdd gnd cell_6t
Xbit_r181_c225 bl_225 br_225 wl_181 vdd gnd cell_6t
Xbit_r182_c225 bl_225 br_225 wl_182 vdd gnd cell_6t
Xbit_r183_c225 bl_225 br_225 wl_183 vdd gnd cell_6t
Xbit_r184_c225 bl_225 br_225 wl_184 vdd gnd cell_6t
Xbit_r185_c225 bl_225 br_225 wl_185 vdd gnd cell_6t
Xbit_r186_c225 bl_225 br_225 wl_186 vdd gnd cell_6t
Xbit_r187_c225 bl_225 br_225 wl_187 vdd gnd cell_6t
Xbit_r188_c225 bl_225 br_225 wl_188 vdd gnd cell_6t
Xbit_r189_c225 bl_225 br_225 wl_189 vdd gnd cell_6t
Xbit_r190_c225 bl_225 br_225 wl_190 vdd gnd cell_6t
Xbit_r191_c225 bl_225 br_225 wl_191 vdd gnd cell_6t
Xbit_r192_c225 bl_225 br_225 wl_192 vdd gnd cell_6t
Xbit_r193_c225 bl_225 br_225 wl_193 vdd gnd cell_6t
Xbit_r194_c225 bl_225 br_225 wl_194 vdd gnd cell_6t
Xbit_r195_c225 bl_225 br_225 wl_195 vdd gnd cell_6t
Xbit_r196_c225 bl_225 br_225 wl_196 vdd gnd cell_6t
Xbit_r197_c225 bl_225 br_225 wl_197 vdd gnd cell_6t
Xbit_r198_c225 bl_225 br_225 wl_198 vdd gnd cell_6t
Xbit_r199_c225 bl_225 br_225 wl_199 vdd gnd cell_6t
Xbit_r200_c225 bl_225 br_225 wl_200 vdd gnd cell_6t
Xbit_r201_c225 bl_225 br_225 wl_201 vdd gnd cell_6t
Xbit_r202_c225 bl_225 br_225 wl_202 vdd gnd cell_6t
Xbit_r203_c225 bl_225 br_225 wl_203 vdd gnd cell_6t
Xbit_r204_c225 bl_225 br_225 wl_204 vdd gnd cell_6t
Xbit_r205_c225 bl_225 br_225 wl_205 vdd gnd cell_6t
Xbit_r206_c225 bl_225 br_225 wl_206 vdd gnd cell_6t
Xbit_r207_c225 bl_225 br_225 wl_207 vdd gnd cell_6t
Xbit_r208_c225 bl_225 br_225 wl_208 vdd gnd cell_6t
Xbit_r209_c225 bl_225 br_225 wl_209 vdd gnd cell_6t
Xbit_r210_c225 bl_225 br_225 wl_210 vdd gnd cell_6t
Xbit_r211_c225 bl_225 br_225 wl_211 vdd gnd cell_6t
Xbit_r212_c225 bl_225 br_225 wl_212 vdd gnd cell_6t
Xbit_r213_c225 bl_225 br_225 wl_213 vdd gnd cell_6t
Xbit_r214_c225 bl_225 br_225 wl_214 vdd gnd cell_6t
Xbit_r215_c225 bl_225 br_225 wl_215 vdd gnd cell_6t
Xbit_r216_c225 bl_225 br_225 wl_216 vdd gnd cell_6t
Xbit_r217_c225 bl_225 br_225 wl_217 vdd gnd cell_6t
Xbit_r218_c225 bl_225 br_225 wl_218 vdd gnd cell_6t
Xbit_r219_c225 bl_225 br_225 wl_219 vdd gnd cell_6t
Xbit_r220_c225 bl_225 br_225 wl_220 vdd gnd cell_6t
Xbit_r221_c225 bl_225 br_225 wl_221 vdd gnd cell_6t
Xbit_r222_c225 bl_225 br_225 wl_222 vdd gnd cell_6t
Xbit_r223_c225 bl_225 br_225 wl_223 vdd gnd cell_6t
Xbit_r224_c225 bl_225 br_225 wl_224 vdd gnd cell_6t
Xbit_r225_c225 bl_225 br_225 wl_225 vdd gnd cell_6t
Xbit_r226_c225 bl_225 br_225 wl_226 vdd gnd cell_6t
Xbit_r227_c225 bl_225 br_225 wl_227 vdd gnd cell_6t
Xbit_r228_c225 bl_225 br_225 wl_228 vdd gnd cell_6t
Xbit_r229_c225 bl_225 br_225 wl_229 vdd gnd cell_6t
Xbit_r230_c225 bl_225 br_225 wl_230 vdd gnd cell_6t
Xbit_r231_c225 bl_225 br_225 wl_231 vdd gnd cell_6t
Xbit_r232_c225 bl_225 br_225 wl_232 vdd gnd cell_6t
Xbit_r233_c225 bl_225 br_225 wl_233 vdd gnd cell_6t
Xbit_r234_c225 bl_225 br_225 wl_234 vdd gnd cell_6t
Xbit_r235_c225 bl_225 br_225 wl_235 vdd gnd cell_6t
Xbit_r236_c225 bl_225 br_225 wl_236 vdd gnd cell_6t
Xbit_r237_c225 bl_225 br_225 wl_237 vdd gnd cell_6t
Xbit_r238_c225 bl_225 br_225 wl_238 vdd gnd cell_6t
Xbit_r239_c225 bl_225 br_225 wl_239 vdd gnd cell_6t
Xbit_r240_c225 bl_225 br_225 wl_240 vdd gnd cell_6t
Xbit_r241_c225 bl_225 br_225 wl_241 vdd gnd cell_6t
Xbit_r242_c225 bl_225 br_225 wl_242 vdd gnd cell_6t
Xbit_r243_c225 bl_225 br_225 wl_243 vdd gnd cell_6t
Xbit_r244_c225 bl_225 br_225 wl_244 vdd gnd cell_6t
Xbit_r245_c225 bl_225 br_225 wl_245 vdd gnd cell_6t
Xbit_r246_c225 bl_225 br_225 wl_246 vdd gnd cell_6t
Xbit_r247_c225 bl_225 br_225 wl_247 vdd gnd cell_6t
Xbit_r248_c225 bl_225 br_225 wl_248 vdd gnd cell_6t
Xbit_r249_c225 bl_225 br_225 wl_249 vdd gnd cell_6t
Xbit_r250_c225 bl_225 br_225 wl_250 vdd gnd cell_6t
Xbit_r251_c225 bl_225 br_225 wl_251 vdd gnd cell_6t
Xbit_r252_c225 bl_225 br_225 wl_252 vdd gnd cell_6t
Xbit_r253_c225 bl_225 br_225 wl_253 vdd gnd cell_6t
Xbit_r254_c225 bl_225 br_225 wl_254 vdd gnd cell_6t
Xbit_r255_c225 bl_225 br_225 wl_255 vdd gnd cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd cell_6t
Xbit_r1_c226 bl_226 br_226 wl_1 vdd gnd cell_6t
Xbit_r2_c226 bl_226 br_226 wl_2 vdd gnd cell_6t
Xbit_r3_c226 bl_226 br_226 wl_3 vdd gnd cell_6t
Xbit_r4_c226 bl_226 br_226 wl_4 vdd gnd cell_6t
Xbit_r5_c226 bl_226 br_226 wl_5 vdd gnd cell_6t
Xbit_r6_c226 bl_226 br_226 wl_6 vdd gnd cell_6t
Xbit_r7_c226 bl_226 br_226 wl_7 vdd gnd cell_6t
Xbit_r8_c226 bl_226 br_226 wl_8 vdd gnd cell_6t
Xbit_r9_c226 bl_226 br_226 wl_9 vdd gnd cell_6t
Xbit_r10_c226 bl_226 br_226 wl_10 vdd gnd cell_6t
Xbit_r11_c226 bl_226 br_226 wl_11 vdd gnd cell_6t
Xbit_r12_c226 bl_226 br_226 wl_12 vdd gnd cell_6t
Xbit_r13_c226 bl_226 br_226 wl_13 vdd gnd cell_6t
Xbit_r14_c226 bl_226 br_226 wl_14 vdd gnd cell_6t
Xbit_r15_c226 bl_226 br_226 wl_15 vdd gnd cell_6t
Xbit_r16_c226 bl_226 br_226 wl_16 vdd gnd cell_6t
Xbit_r17_c226 bl_226 br_226 wl_17 vdd gnd cell_6t
Xbit_r18_c226 bl_226 br_226 wl_18 vdd gnd cell_6t
Xbit_r19_c226 bl_226 br_226 wl_19 vdd gnd cell_6t
Xbit_r20_c226 bl_226 br_226 wl_20 vdd gnd cell_6t
Xbit_r21_c226 bl_226 br_226 wl_21 vdd gnd cell_6t
Xbit_r22_c226 bl_226 br_226 wl_22 vdd gnd cell_6t
Xbit_r23_c226 bl_226 br_226 wl_23 vdd gnd cell_6t
Xbit_r24_c226 bl_226 br_226 wl_24 vdd gnd cell_6t
Xbit_r25_c226 bl_226 br_226 wl_25 vdd gnd cell_6t
Xbit_r26_c226 bl_226 br_226 wl_26 vdd gnd cell_6t
Xbit_r27_c226 bl_226 br_226 wl_27 vdd gnd cell_6t
Xbit_r28_c226 bl_226 br_226 wl_28 vdd gnd cell_6t
Xbit_r29_c226 bl_226 br_226 wl_29 vdd gnd cell_6t
Xbit_r30_c226 bl_226 br_226 wl_30 vdd gnd cell_6t
Xbit_r31_c226 bl_226 br_226 wl_31 vdd gnd cell_6t
Xbit_r32_c226 bl_226 br_226 wl_32 vdd gnd cell_6t
Xbit_r33_c226 bl_226 br_226 wl_33 vdd gnd cell_6t
Xbit_r34_c226 bl_226 br_226 wl_34 vdd gnd cell_6t
Xbit_r35_c226 bl_226 br_226 wl_35 vdd gnd cell_6t
Xbit_r36_c226 bl_226 br_226 wl_36 vdd gnd cell_6t
Xbit_r37_c226 bl_226 br_226 wl_37 vdd gnd cell_6t
Xbit_r38_c226 bl_226 br_226 wl_38 vdd gnd cell_6t
Xbit_r39_c226 bl_226 br_226 wl_39 vdd gnd cell_6t
Xbit_r40_c226 bl_226 br_226 wl_40 vdd gnd cell_6t
Xbit_r41_c226 bl_226 br_226 wl_41 vdd gnd cell_6t
Xbit_r42_c226 bl_226 br_226 wl_42 vdd gnd cell_6t
Xbit_r43_c226 bl_226 br_226 wl_43 vdd gnd cell_6t
Xbit_r44_c226 bl_226 br_226 wl_44 vdd gnd cell_6t
Xbit_r45_c226 bl_226 br_226 wl_45 vdd gnd cell_6t
Xbit_r46_c226 bl_226 br_226 wl_46 vdd gnd cell_6t
Xbit_r47_c226 bl_226 br_226 wl_47 vdd gnd cell_6t
Xbit_r48_c226 bl_226 br_226 wl_48 vdd gnd cell_6t
Xbit_r49_c226 bl_226 br_226 wl_49 vdd gnd cell_6t
Xbit_r50_c226 bl_226 br_226 wl_50 vdd gnd cell_6t
Xbit_r51_c226 bl_226 br_226 wl_51 vdd gnd cell_6t
Xbit_r52_c226 bl_226 br_226 wl_52 vdd gnd cell_6t
Xbit_r53_c226 bl_226 br_226 wl_53 vdd gnd cell_6t
Xbit_r54_c226 bl_226 br_226 wl_54 vdd gnd cell_6t
Xbit_r55_c226 bl_226 br_226 wl_55 vdd gnd cell_6t
Xbit_r56_c226 bl_226 br_226 wl_56 vdd gnd cell_6t
Xbit_r57_c226 bl_226 br_226 wl_57 vdd gnd cell_6t
Xbit_r58_c226 bl_226 br_226 wl_58 vdd gnd cell_6t
Xbit_r59_c226 bl_226 br_226 wl_59 vdd gnd cell_6t
Xbit_r60_c226 bl_226 br_226 wl_60 vdd gnd cell_6t
Xbit_r61_c226 bl_226 br_226 wl_61 vdd gnd cell_6t
Xbit_r62_c226 bl_226 br_226 wl_62 vdd gnd cell_6t
Xbit_r63_c226 bl_226 br_226 wl_63 vdd gnd cell_6t
Xbit_r64_c226 bl_226 br_226 wl_64 vdd gnd cell_6t
Xbit_r65_c226 bl_226 br_226 wl_65 vdd gnd cell_6t
Xbit_r66_c226 bl_226 br_226 wl_66 vdd gnd cell_6t
Xbit_r67_c226 bl_226 br_226 wl_67 vdd gnd cell_6t
Xbit_r68_c226 bl_226 br_226 wl_68 vdd gnd cell_6t
Xbit_r69_c226 bl_226 br_226 wl_69 vdd gnd cell_6t
Xbit_r70_c226 bl_226 br_226 wl_70 vdd gnd cell_6t
Xbit_r71_c226 bl_226 br_226 wl_71 vdd gnd cell_6t
Xbit_r72_c226 bl_226 br_226 wl_72 vdd gnd cell_6t
Xbit_r73_c226 bl_226 br_226 wl_73 vdd gnd cell_6t
Xbit_r74_c226 bl_226 br_226 wl_74 vdd gnd cell_6t
Xbit_r75_c226 bl_226 br_226 wl_75 vdd gnd cell_6t
Xbit_r76_c226 bl_226 br_226 wl_76 vdd gnd cell_6t
Xbit_r77_c226 bl_226 br_226 wl_77 vdd gnd cell_6t
Xbit_r78_c226 bl_226 br_226 wl_78 vdd gnd cell_6t
Xbit_r79_c226 bl_226 br_226 wl_79 vdd gnd cell_6t
Xbit_r80_c226 bl_226 br_226 wl_80 vdd gnd cell_6t
Xbit_r81_c226 bl_226 br_226 wl_81 vdd gnd cell_6t
Xbit_r82_c226 bl_226 br_226 wl_82 vdd gnd cell_6t
Xbit_r83_c226 bl_226 br_226 wl_83 vdd gnd cell_6t
Xbit_r84_c226 bl_226 br_226 wl_84 vdd gnd cell_6t
Xbit_r85_c226 bl_226 br_226 wl_85 vdd gnd cell_6t
Xbit_r86_c226 bl_226 br_226 wl_86 vdd gnd cell_6t
Xbit_r87_c226 bl_226 br_226 wl_87 vdd gnd cell_6t
Xbit_r88_c226 bl_226 br_226 wl_88 vdd gnd cell_6t
Xbit_r89_c226 bl_226 br_226 wl_89 vdd gnd cell_6t
Xbit_r90_c226 bl_226 br_226 wl_90 vdd gnd cell_6t
Xbit_r91_c226 bl_226 br_226 wl_91 vdd gnd cell_6t
Xbit_r92_c226 bl_226 br_226 wl_92 vdd gnd cell_6t
Xbit_r93_c226 bl_226 br_226 wl_93 vdd gnd cell_6t
Xbit_r94_c226 bl_226 br_226 wl_94 vdd gnd cell_6t
Xbit_r95_c226 bl_226 br_226 wl_95 vdd gnd cell_6t
Xbit_r96_c226 bl_226 br_226 wl_96 vdd gnd cell_6t
Xbit_r97_c226 bl_226 br_226 wl_97 vdd gnd cell_6t
Xbit_r98_c226 bl_226 br_226 wl_98 vdd gnd cell_6t
Xbit_r99_c226 bl_226 br_226 wl_99 vdd gnd cell_6t
Xbit_r100_c226 bl_226 br_226 wl_100 vdd gnd cell_6t
Xbit_r101_c226 bl_226 br_226 wl_101 vdd gnd cell_6t
Xbit_r102_c226 bl_226 br_226 wl_102 vdd gnd cell_6t
Xbit_r103_c226 bl_226 br_226 wl_103 vdd gnd cell_6t
Xbit_r104_c226 bl_226 br_226 wl_104 vdd gnd cell_6t
Xbit_r105_c226 bl_226 br_226 wl_105 vdd gnd cell_6t
Xbit_r106_c226 bl_226 br_226 wl_106 vdd gnd cell_6t
Xbit_r107_c226 bl_226 br_226 wl_107 vdd gnd cell_6t
Xbit_r108_c226 bl_226 br_226 wl_108 vdd gnd cell_6t
Xbit_r109_c226 bl_226 br_226 wl_109 vdd gnd cell_6t
Xbit_r110_c226 bl_226 br_226 wl_110 vdd gnd cell_6t
Xbit_r111_c226 bl_226 br_226 wl_111 vdd gnd cell_6t
Xbit_r112_c226 bl_226 br_226 wl_112 vdd gnd cell_6t
Xbit_r113_c226 bl_226 br_226 wl_113 vdd gnd cell_6t
Xbit_r114_c226 bl_226 br_226 wl_114 vdd gnd cell_6t
Xbit_r115_c226 bl_226 br_226 wl_115 vdd gnd cell_6t
Xbit_r116_c226 bl_226 br_226 wl_116 vdd gnd cell_6t
Xbit_r117_c226 bl_226 br_226 wl_117 vdd gnd cell_6t
Xbit_r118_c226 bl_226 br_226 wl_118 vdd gnd cell_6t
Xbit_r119_c226 bl_226 br_226 wl_119 vdd gnd cell_6t
Xbit_r120_c226 bl_226 br_226 wl_120 vdd gnd cell_6t
Xbit_r121_c226 bl_226 br_226 wl_121 vdd gnd cell_6t
Xbit_r122_c226 bl_226 br_226 wl_122 vdd gnd cell_6t
Xbit_r123_c226 bl_226 br_226 wl_123 vdd gnd cell_6t
Xbit_r124_c226 bl_226 br_226 wl_124 vdd gnd cell_6t
Xbit_r125_c226 bl_226 br_226 wl_125 vdd gnd cell_6t
Xbit_r126_c226 bl_226 br_226 wl_126 vdd gnd cell_6t
Xbit_r127_c226 bl_226 br_226 wl_127 vdd gnd cell_6t
Xbit_r128_c226 bl_226 br_226 wl_128 vdd gnd cell_6t
Xbit_r129_c226 bl_226 br_226 wl_129 vdd gnd cell_6t
Xbit_r130_c226 bl_226 br_226 wl_130 vdd gnd cell_6t
Xbit_r131_c226 bl_226 br_226 wl_131 vdd gnd cell_6t
Xbit_r132_c226 bl_226 br_226 wl_132 vdd gnd cell_6t
Xbit_r133_c226 bl_226 br_226 wl_133 vdd gnd cell_6t
Xbit_r134_c226 bl_226 br_226 wl_134 vdd gnd cell_6t
Xbit_r135_c226 bl_226 br_226 wl_135 vdd gnd cell_6t
Xbit_r136_c226 bl_226 br_226 wl_136 vdd gnd cell_6t
Xbit_r137_c226 bl_226 br_226 wl_137 vdd gnd cell_6t
Xbit_r138_c226 bl_226 br_226 wl_138 vdd gnd cell_6t
Xbit_r139_c226 bl_226 br_226 wl_139 vdd gnd cell_6t
Xbit_r140_c226 bl_226 br_226 wl_140 vdd gnd cell_6t
Xbit_r141_c226 bl_226 br_226 wl_141 vdd gnd cell_6t
Xbit_r142_c226 bl_226 br_226 wl_142 vdd gnd cell_6t
Xbit_r143_c226 bl_226 br_226 wl_143 vdd gnd cell_6t
Xbit_r144_c226 bl_226 br_226 wl_144 vdd gnd cell_6t
Xbit_r145_c226 bl_226 br_226 wl_145 vdd gnd cell_6t
Xbit_r146_c226 bl_226 br_226 wl_146 vdd gnd cell_6t
Xbit_r147_c226 bl_226 br_226 wl_147 vdd gnd cell_6t
Xbit_r148_c226 bl_226 br_226 wl_148 vdd gnd cell_6t
Xbit_r149_c226 bl_226 br_226 wl_149 vdd gnd cell_6t
Xbit_r150_c226 bl_226 br_226 wl_150 vdd gnd cell_6t
Xbit_r151_c226 bl_226 br_226 wl_151 vdd gnd cell_6t
Xbit_r152_c226 bl_226 br_226 wl_152 vdd gnd cell_6t
Xbit_r153_c226 bl_226 br_226 wl_153 vdd gnd cell_6t
Xbit_r154_c226 bl_226 br_226 wl_154 vdd gnd cell_6t
Xbit_r155_c226 bl_226 br_226 wl_155 vdd gnd cell_6t
Xbit_r156_c226 bl_226 br_226 wl_156 vdd gnd cell_6t
Xbit_r157_c226 bl_226 br_226 wl_157 vdd gnd cell_6t
Xbit_r158_c226 bl_226 br_226 wl_158 vdd gnd cell_6t
Xbit_r159_c226 bl_226 br_226 wl_159 vdd gnd cell_6t
Xbit_r160_c226 bl_226 br_226 wl_160 vdd gnd cell_6t
Xbit_r161_c226 bl_226 br_226 wl_161 vdd gnd cell_6t
Xbit_r162_c226 bl_226 br_226 wl_162 vdd gnd cell_6t
Xbit_r163_c226 bl_226 br_226 wl_163 vdd gnd cell_6t
Xbit_r164_c226 bl_226 br_226 wl_164 vdd gnd cell_6t
Xbit_r165_c226 bl_226 br_226 wl_165 vdd gnd cell_6t
Xbit_r166_c226 bl_226 br_226 wl_166 vdd gnd cell_6t
Xbit_r167_c226 bl_226 br_226 wl_167 vdd gnd cell_6t
Xbit_r168_c226 bl_226 br_226 wl_168 vdd gnd cell_6t
Xbit_r169_c226 bl_226 br_226 wl_169 vdd gnd cell_6t
Xbit_r170_c226 bl_226 br_226 wl_170 vdd gnd cell_6t
Xbit_r171_c226 bl_226 br_226 wl_171 vdd gnd cell_6t
Xbit_r172_c226 bl_226 br_226 wl_172 vdd gnd cell_6t
Xbit_r173_c226 bl_226 br_226 wl_173 vdd gnd cell_6t
Xbit_r174_c226 bl_226 br_226 wl_174 vdd gnd cell_6t
Xbit_r175_c226 bl_226 br_226 wl_175 vdd gnd cell_6t
Xbit_r176_c226 bl_226 br_226 wl_176 vdd gnd cell_6t
Xbit_r177_c226 bl_226 br_226 wl_177 vdd gnd cell_6t
Xbit_r178_c226 bl_226 br_226 wl_178 vdd gnd cell_6t
Xbit_r179_c226 bl_226 br_226 wl_179 vdd gnd cell_6t
Xbit_r180_c226 bl_226 br_226 wl_180 vdd gnd cell_6t
Xbit_r181_c226 bl_226 br_226 wl_181 vdd gnd cell_6t
Xbit_r182_c226 bl_226 br_226 wl_182 vdd gnd cell_6t
Xbit_r183_c226 bl_226 br_226 wl_183 vdd gnd cell_6t
Xbit_r184_c226 bl_226 br_226 wl_184 vdd gnd cell_6t
Xbit_r185_c226 bl_226 br_226 wl_185 vdd gnd cell_6t
Xbit_r186_c226 bl_226 br_226 wl_186 vdd gnd cell_6t
Xbit_r187_c226 bl_226 br_226 wl_187 vdd gnd cell_6t
Xbit_r188_c226 bl_226 br_226 wl_188 vdd gnd cell_6t
Xbit_r189_c226 bl_226 br_226 wl_189 vdd gnd cell_6t
Xbit_r190_c226 bl_226 br_226 wl_190 vdd gnd cell_6t
Xbit_r191_c226 bl_226 br_226 wl_191 vdd gnd cell_6t
Xbit_r192_c226 bl_226 br_226 wl_192 vdd gnd cell_6t
Xbit_r193_c226 bl_226 br_226 wl_193 vdd gnd cell_6t
Xbit_r194_c226 bl_226 br_226 wl_194 vdd gnd cell_6t
Xbit_r195_c226 bl_226 br_226 wl_195 vdd gnd cell_6t
Xbit_r196_c226 bl_226 br_226 wl_196 vdd gnd cell_6t
Xbit_r197_c226 bl_226 br_226 wl_197 vdd gnd cell_6t
Xbit_r198_c226 bl_226 br_226 wl_198 vdd gnd cell_6t
Xbit_r199_c226 bl_226 br_226 wl_199 vdd gnd cell_6t
Xbit_r200_c226 bl_226 br_226 wl_200 vdd gnd cell_6t
Xbit_r201_c226 bl_226 br_226 wl_201 vdd gnd cell_6t
Xbit_r202_c226 bl_226 br_226 wl_202 vdd gnd cell_6t
Xbit_r203_c226 bl_226 br_226 wl_203 vdd gnd cell_6t
Xbit_r204_c226 bl_226 br_226 wl_204 vdd gnd cell_6t
Xbit_r205_c226 bl_226 br_226 wl_205 vdd gnd cell_6t
Xbit_r206_c226 bl_226 br_226 wl_206 vdd gnd cell_6t
Xbit_r207_c226 bl_226 br_226 wl_207 vdd gnd cell_6t
Xbit_r208_c226 bl_226 br_226 wl_208 vdd gnd cell_6t
Xbit_r209_c226 bl_226 br_226 wl_209 vdd gnd cell_6t
Xbit_r210_c226 bl_226 br_226 wl_210 vdd gnd cell_6t
Xbit_r211_c226 bl_226 br_226 wl_211 vdd gnd cell_6t
Xbit_r212_c226 bl_226 br_226 wl_212 vdd gnd cell_6t
Xbit_r213_c226 bl_226 br_226 wl_213 vdd gnd cell_6t
Xbit_r214_c226 bl_226 br_226 wl_214 vdd gnd cell_6t
Xbit_r215_c226 bl_226 br_226 wl_215 vdd gnd cell_6t
Xbit_r216_c226 bl_226 br_226 wl_216 vdd gnd cell_6t
Xbit_r217_c226 bl_226 br_226 wl_217 vdd gnd cell_6t
Xbit_r218_c226 bl_226 br_226 wl_218 vdd gnd cell_6t
Xbit_r219_c226 bl_226 br_226 wl_219 vdd gnd cell_6t
Xbit_r220_c226 bl_226 br_226 wl_220 vdd gnd cell_6t
Xbit_r221_c226 bl_226 br_226 wl_221 vdd gnd cell_6t
Xbit_r222_c226 bl_226 br_226 wl_222 vdd gnd cell_6t
Xbit_r223_c226 bl_226 br_226 wl_223 vdd gnd cell_6t
Xbit_r224_c226 bl_226 br_226 wl_224 vdd gnd cell_6t
Xbit_r225_c226 bl_226 br_226 wl_225 vdd gnd cell_6t
Xbit_r226_c226 bl_226 br_226 wl_226 vdd gnd cell_6t
Xbit_r227_c226 bl_226 br_226 wl_227 vdd gnd cell_6t
Xbit_r228_c226 bl_226 br_226 wl_228 vdd gnd cell_6t
Xbit_r229_c226 bl_226 br_226 wl_229 vdd gnd cell_6t
Xbit_r230_c226 bl_226 br_226 wl_230 vdd gnd cell_6t
Xbit_r231_c226 bl_226 br_226 wl_231 vdd gnd cell_6t
Xbit_r232_c226 bl_226 br_226 wl_232 vdd gnd cell_6t
Xbit_r233_c226 bl_226 br_226 wl_233 vdd gnd cell_6t
Xbit_r234_c226 bl_226 br_226 wl_234 vdd gnd cell_6t
Xbit_r235_c226 bl_226 br_226 wl_235 vdd gnd cell_6t
Xbit_r236_c226 bl_226 br_226 wl_236 vdd gnd cell_6t
Xbit_r237_c226 bl_226 br_226 wl_237 vdd gnd cell_6t
Xbit_r238_c226 bl_226 br_226 wl_238 vdd gnd cell_6t
Xbit_r239_c226 bl_226 br_226 wl_239 vdd gnd cell_6t
Xbit_r240_c226 bl_226 br_226 wl_240 vdd gnd cell_6t
Xbit_r241_c226 bl_226 br_226 wl_241 vdd gnd cell_6t
Xbit_r242_c226 bl_226 br_226 wl_242 vdd gnd cell_6t
Xbit_r243_c226 bl_226 br_226 wl_243 vdd gnd cell_6t
Xbit_r244_c226 bl_226 br_226 wl_244 vdd gnd cell_6t
Xbit_r245_c226 bl_226 br_226 wl_245 vdd gnd cell_6t
Xbit_r246_c226 bl_226 br_226 wl_246 vdd gnd cell_6t
Xbit_r247_c226 bl_226 br_226 wl_247 vdd gnd cell_6t
Xbit_r248_c226 bl_226 br_226 wl_248 vdd gnd cell_6t
Xbit_r249_c226 bl_226 br_226 wl_249 vdd gnd cell_6t
Xbit_r250_c226 bl_226 br_226 wl_250 vdd gnd cell_6t
Xbit_r251_c226 bl_226 br_226 wl_251 vdd gnd cell_6t
Xbit_r252_c226 bl_226 br_226 wl_252 vdd gnd cell_6t
Xbit_r253_c226 bl_226 br_226 wl_253 vdd gnd cell_6t
Xbit_r254_c226 bl_226 br_226 wl_254 vdd gnd cell_6t
Xbit_r255_c226 bl_226 br_226 wl_255 vdd gnd cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd cell_6t
Xbit_r1_c227 bl_227 br_227 wl_1 vdd gnd cell_6t
Xbit_r2_c227 bl_227 br_227 wl_2 vdd gnd cell_6t
Xbit_r3_c227 bl_227 br_227 wl_3 vdd gnd cell_6t
Xbit_r4_c227 bl_227 br_227 wl_4 vdd gnd cell_6t
Xbit_r5_c227 bl_227 br_227 wl_5 vdd gnd cell_6t
Xbit_r6_c227 bl_227 br_227 wl_6 vdd gnd cell_6t
Xbit_r7_c227 bl_227 br_227 wl_7 vdd gnd cell_6t
Xbit_r8_c227 bl_227 br_227 wl_8 vdd gnd cell_6t
Xbit_r9_c227 bl_227 br_227 wl_9 vdd gnd cell_6t
Xbit_r10_c227 bl_227 br_227 wl_10 vdd gnd cell_6t
Xbit_r11_c227 bl_227 br_227 wl_11 vdd gnd cell_6t
Xbit_r12_c227 bl_227 br_227 wl_12 vdd gnd cell_6t
Xbit_r13_c227 bl_227 br_227 wl_13 vdd gnd cell_6t
Xbit_r14_c227 bl_227 br_227 wl_14 vdd gnd cell_6t
Xbit_r15_c227 bl_227 br_227 wl_15 vdd gnd cell_6t
Xbit_r16_c227 bl_227 br_227 wl_16 vdd gnd cell_6t
Xbit_r17_c227 bl_227 br_227 wl_17 vdd gnd cell_6t
Xbit_r18_c227 bl_227 br_227 wl_18 vdd gnd cell_6t
Xbit_r19_c227 bl_227 br_227 wl_19 vdd gnd cell_6t
Xbit_r20_c227 bl_227 br_227 wl_20 vdd gnd cell_6t
Xbit_r21_c227 bl_227 br_227 wl_21 vdd gnd cell_6t
Xbit_r22_c227 bl_227 br_227 wl_22 vdd gnd cell_6t
Xbit_r23_c227 bl_227 br_227 wl_23 vdd gnd cell_6t
Xbit_r24_c227 bl_227 br_227 wl_24 vdd gnd cell_6t
Xbit_r25_c227 bl_227 br_227 wl_25 vdd gnd cell_6t
Xbit_r26_c227 bl_227 br_227 wl_26 vdd gnd cell_6t
Xbit_r27_c227 bl_227 br_227 wl_27 vdd gnd cell_6t
Xbit_r28_c227 bl_227 br_227 wl_28 vdd gnd cell_6t
Xbit_r29_c227 bl_227 br_227 wl_29 vdd gnd cell_6t
Xbit_r30_c227 bl_227 br_227 wl_30 vdd gnd cell_6t
Xbit_r31_c227 bl_227 br_227 wl_31 vdd gnd cell_6t
Xbit_r32_c227 bl_227 br_227 wl_32 vdd gnd cell_6t
Xbit_r33_c227 bl_227 br_227 wl_33 vdd gnd cell_6t
Xbit_r34_c227 bl_227 br_227 wl_34 vdd gnd cell_6t
Xbit_r35_c227 bl_227 br_227 wl_35 vdd gnd cell_6t
Xbit_r36_c227 bl_227 br_227 wl_36 vdd gnd cell_6t
Xbit_r37_c227 bl_227 br_227 wl_37 vdd gnd cell_6t
Xbit_r38_c227 bl_227 br_227 wl_38 vdd gnd cell_6t
Xbit_r39_c227 bl_227 br_227 wl_39 vdd gnd cell_6t
Xbit_r40_c227 bl_227 br_227 wl_40 vdd gnd cell_6t
Xbit_r41_c227 bl_227 br_227 wl_41 vdd gnd cell_6t
Xbit_r42_c227 bl_227 br_227 wl_42 vdd gnd cell_6t
Xbit_r43_c227 bl_227 br_227 wl_43 vdd gnd cell_6t
Xbit_r44_c227 bl_227 br_227 wl_44 vdd gnd cell_6t
Xbit_r45_c227 bl_227 br_227 wl_45 vdd gnd cell_6t
Xbit_r46_c227 bl_227 br_227 wl_46 vdd gnd cell_6t
Xbit_r47_c227 bl_227 br_227 wl_47 vdd gnd cell_6t
Xbit_r48_c227 bl_227 br_227 wl_48 vdd gnd cell_6t
Xbit_r49_c227 bl_227 br_227 wl_49 vdd gnd cell_6t
Xbit_r50_c227 bl_227 br_227 wl_50 vdd gnd cell_6t
Xbit_r51_c227 bl_227 br_227 wl_51 vdd gnd cell_6t
Xbit_r52_c227 bl_227 br_227 wl_52 vdd gnd cell_6t
Xbit_r53_c227 bl_227 br_227 wl_53 vdd gnd cell_6t
Xbit_r54_c227 bl_227 br_227 wl_54 vdd gnd cell_6t
Xbit_r55_c227 bl_227 br_227 wl_55 vdd gnd cell_6t
Xbit_r56_c227 bl_227 br_227 wl_56 vdd gnd cell_6t
Xbit_r57_c227 bl_227 br_227 wl_57 vdd gnd cell_6t
Xbit_r58_c227 bl_227 br_227 wl_58 vdd gnd cell_6t
Xbit_r59_c227 bl_227 br_227 wl_59 vdd gnd cell_6t
Xbit_r60_c227 bl_227 br_227 wl_60 vdd gnd cell_6t
Xbit_r61_c227 bl_227 br_227 wl_61 vdd gnd cell_6t
Xbit_r62_c227 bl_227 br_227 wl_62 vdd gnd cell_6t
Xbit_r63_c227 bl_227 br_227 wl_63 vdd gnd cell_6t
Xbit_r64_c227 bl_227 br_227 wl_64 vdd gnd cell_6t
Xbit_r65_c227 bl_227 br_227 wl_65 vdd gnd cell_6t
Xbit_r66_c227 bl_227 br_227 wl_66 vdd gnd cell_6t
Xbit_r67_c227 bl_227 br_227 wl_67 vdd gnd cell_6t
Xbit_r68_c227 bl_227 br_227 wl_68 vdd gnd cell_6t
Xbit_r69_c227 bl_227 br_227 wl_69 vdd gnd cell_6t
Xbit_r70_c227 bl_227 br_227 wl_70 vdd gnd cell_6t
Xbit_r71_c227 bl_227 br_227 wl_71 vdd gnd cell_6t
Xbit_r72_c227 bl_227 br_227 wl_72 vdd gnd cell_6t
Xbit_r73_c227 bl_227 br_227 wl_73 vdd gnd cell_6t
Xbit_r74_c227 bl_227 br_227 wl_74 vdd gnd cell_6t
Xbit_r75_c227 bl_227 br_227 wl_75 vdd gnd cell_6t
Xbit_r76_c227 bl_227 br_227 wl_76 vdd gnd cell_6t
Xbit_r77_c227 bl_227 br_227 wl_77 vdd gnd cell_6t
Xbit_r78_c227 bl_227 br_227 wl_78 vdd gnd cell_6t
Xbit_r79_c227 bl_227 br_227 wl_79 vdd gnd cell_6t
Xbit_r80_c227 bl_227 br_227 wl_80 vdd gnd cell_6t
Xbit_r81_c227 bl_227 br_227 wl_81 vdd gnd cell_6t
Xbit_r82_c227 bl_227 br_227 wl_82 vdd gnd cell_6t
Xbit_r83_c227 bl_227 br_227 wl_83 vdd gnd cell_6t
Xbit_r84_c227 bl_227 br_227 wl_84 vdd gnd cell_6t
Xbit_r85_c227 bl_227 br_227 wl_85 vdd gnd cell_6t
Xbit_r86_c227 bl_227 br_227 wl_86 vdd gnd cell_6t
Xbit_r87_c227 bl_227 br_227 wl_87 vdd gnd cell_6t
Xbit_r88_c227 bl_227 br_227 wl_88 vdd gnd cell_6t
Xbit_r89_c227 bl_227 br_227 wl_89 vdd gnd cell_6t
Xbit_r90_c227 bl_227 br_227 wl_90 vdd gnd cell_6t
Xbit_r91_c227 bl_227 br_227 wl_91 vdd gnd cell_6t
Xbit_r92_c227 bl_227 br_227 wl_92 vdd gnd cell_6t
Xbit_r93_c227 bl_227 br_227 wl_93 vdd gnd cell_6t
Xbit_r94_c227 bl_227 br_227 wl_94 vdd gnd cell_6t
Xbit_r95_c227 bl_227 br_227 wl_95 vdd gnd cell_6t
Xbit_r96_c227 bl_227 br_227 wl_96 vdd gnd cell_6t
Xbit_r97_c227 bl_227 br_227 wl_97 vdd gnd cell_6t
Xbit_r98_c227 bl_227 br_227 wl_98 vdd gnd cell_6t
Xbit_r99_c227 bl_227 br_227 wl_99 vdd gnd cell_6t
Xbit_r100_c227 bl_227 br_227 wl_100 vdd gnd cell_6t
Xbit_r101_c227 bl_227 br_227 wl_101 vdd gnd cell_6t
Xbit_r102_c227 bl_227 br_227 wl_102 vdd gnd cell_6t
Xbit_r103_c227 bl_227 br_227 wl_103 vdd gnd cell_6t
Xbit_r104_c227 bl_227 br_227 wl_104 vdd gnd cell_6t
Xbit_r105_c227 bl_227 br_227 wl_105 vdd gnd cell_6t
Xbit_r106_c227 bl_227 br_227 wl_106 vdd gnd cell_6t
Xbit_r107_c227 bl_227 br_227 wl_107 vdd gnd cell_6t
Xbit_r108_c227 bl_227 br_227 wl_108 vdd gnd cell_6t
Xbit_r109_c227 bl_227 br_227 wl_109 vdd gnd cell_6t
Xbit_r110_c227 bl_227 br_227 wl_110 vdd gnd cell_6t
Xbit_r111_c227 bl_227 br_227 wl_111 vdd gnd cell_6t
Xbit_r112_c227 bl_227 br_227 wl_112 vdd gnd cell_6t
Xbit_r113_c227 bl_227 br_227 wl_113 vdd gnd cell_6t
Xbit_r114_c227 bl_227 br_227 wl_114 vdd gnd cell_6t
Xbit_r115_c227 bl_227 br_227 wl_115 vdd gnd cell_6t
Xbit_r116_c227 bl_227 br_227 wl_116 vdd gnd cell_6t
Xbit_r117_c227 bl_227 br_227 wl_117 vdd gnd cell_6t
Xbit_r118_c227 bl_227 br_227 wl_118 vdd gnd cell_6t
Xbit_r119_c227 bl_227 br_227 wl_119 vdd gnd cell_6t
Xbit_r120_c227 bl_227 br_227 wl_120 vdd gnd cell_6t
Xbit_r121_c227 bl_227 br_227 wl_121 vdd gnd cell_6t
Xbit_r122_c227 bl_227 br_227 wl_122 vdd gnd cell_6t
Xbit_r123_c227 bl_227 br_227 wl_123 vdd gnd cell_6t
Xbit_r124_c227 bl_227 br_227 wl_124 vdd gnd cell_6t
Xbit_r125_c227 bl_227 br_227 wl_125 vdd gnd cell_6t
Xbit_r126_c227 bl_227 br_227 wl_126 vdd gnd cell_6t
Xbit_r127_c227 bl_227 br_227 wl_127 vdd gnd cell_6t
Xbit_r128_c227 bl_227 br_227 wl_128 vdd gnd cell_6t
Xbit_r129_c227 bl_227 br_227 wl_129 vdd gnd cell_6t
Xbit_r130_c227 bl_227 br_227 wl_130 vdd gnd cell_6t
Xbit_r131_c227 bl_227 br_227 wl_131 vdd gnd cell_6t
Xbit_r132_c227 bl_227 br_227 wl_132 vdd gnd cell_6t
Xbit_r133_c227 bl_227 br_227 wl_133 vdd gnd cell_6t
Xbit_r134_c227 bl_227 br_227 wl_134 vdd gnd cell_6t
Xbit_r135_c227 bl_227 br_227 wl_135 vdd gnd cell_6t
Xbit_r136_c227 bl_227 br_227 wl_136 vdd gnd cell_6t
Xbit_r137_c227 bl_227 br_227 wl_137 vdd gnd cell_6t
Xbit_r138_c227 bl_227 br_227 wl_138 vdd gnd cell_6t
Xbit_r139_c227 bl_227 br_227 wl_139 vdd gnd cell_6t
Xbit_r140_c227 bl_227 br_227 wl_140 vdd gnd cell_6t
Xbit_r141_c227 bl_227 br_227 wl_141 vdd gnd cell_6t
Xbit_r142_c227 bl_227 br_227 wl_142 vdd gnd cell_6t
Xbit_r143_c227 bl_227 br_227 wl_143 vdd gnd cell_6t
Xbit_r144_c227 bl_227 br_227 wl_144 vdd gnd cell_6t
Xbit_r145_c227 bl_227 br_227 wl_145 vdd gnd cell_6t
Xbit_r146_c227 bl_227 br_227 wl_146 vdd gnd cell_6t
Xbit_r147_c227 bl_227 br_227 wl_147 vdd gnd cell_6t
Xbit_r148_c227 bl_227 br_227 wl_148 vdd gnd cell_6t
Xbit_r149_c227 bl_227 br_227 wl_149 vdd gnd cell_6t
Xbit_r150_c227 bl_227 br_227 wl_150 vdd gnd cell_6t
Xbit_r151_c227 bl_227 br_227 wl_151 vdd gnd cell_6t
Xbit_r152_c227 bl_227 br_227 wl_152 vdd gnd cell_6t
Xbit_r153_c227 bl_227 br_227 wl_153 vdd gnd cell_6t
Xbit_r154_c227 bl_227 br_227 wl_154 vdd gnd cell_6t
Xbit_r155_c227 bl_227 br_227 wl_155 vdd gnd cell_6t
Xbit_r156_c227 bl_227 br_227 wl_156 vdd gnd cell_6t
Xbit_r157_c227 bl_227 br_227 wl_157 vdd gnd cell_6t
Xbit_r158_c227 bl_227 br_227 wl_158 vdd gnd cell_6t
Xbit_r159_c227 bl_227 br_227 wl_159 vdd gnd cell_6t
Xbit_r160_c227 bl_227 br_227 wl_160 vdd gnd cell_6t
Xbit_r161_c227 bl_227 br_227 wl_161 vdd gnd cell_6t
Xbit_r162_c227 bl_227 br_227 wl_162 vdd gnd cell_6t
Xbit_r163_c227 bl_227 br_227 wl_163 vdd gnd cell_6t
Xbit_r164_c227 bl_227 br_227 wl_164 vdd gnd cell_6t
Xbit_r165_c227 bl_227 br_227 wl_165 vdd gnd cell_6t
Xbit_r166_c227 bl_227 br_227 wl_166 vdd gnd cell_6t
Xbit_r167_c227 bl_227 br_227 wl_167 vdd gnd cell_6t
Xbit_r168_c227 bl_227 br_227 wl_168 vdd gnd cell_6t
Xbit_r169_c227 bl_227 br_227 wl_169 vdd gnd cell_6t
Xbit_r170_c227 bl_227 br_227 wl_170 vdd gnd cell_6t
Xbit_r171_c227 bl_227 br_227 wl_171 vdd gnd cell_6t
Xbit_r172_c227 bl_227 br_227 wl_172 vdd gnd cell_6t
Xbit_r173_c227 bl_227 br_227 wl_173 vdd gnd cell_6t
Xbit_r174_c227 bl_227 br_227 wl_174 vdd gnd cell_6t
Xbit_r175_c227 bl_227 br_227 wl_175 vdd gnd cell_6t
Xbit_r176_c227 bl_227 br_227 wl_176 vdd gnd cell_6t
Xbit_r177_c227 bl_227 br_227 wl_177 vdd gnd cell_6t
Xbit_r178_c227 bl_227 br_227 wl_178 vdd gnd cell_6t
Xbit_r179_c227 bl_227 br_227 wl_179 vdd gnd cell_6t
Xbit_r180_c227 bl_227 br_227 wl_180 vdd gnd cell_6t
Xbit_r181_c227 bl_227 br_227 wl_181 vdd gnd cell_6t
Xbit_r182_c227 bl_227 br_227 wl_182 vdd gnd cell_6t
Xbit_r183_c227 bl_227 br_227 wl_183 vdd gnd cell_6t
Xbit_r184_c227 bl_227 br_227 wl_184 vdd gnd cell_6t
Xbit_r185_c227 bl_227 br_227 wl_185 vdd gnd cell_6t
Xbit_r186_c227 bl_227 br_227 wl_186 vdd gnd cell_6t
Xbit_r187_c227 bl_227 br_227 wl_187 vdd gnd cell_6t
Xbit_r188_c227 bl_227 br_227 wl_188 vdd gnd cell_6t
Xbit_r189_c227 bl_227 br_227 wl_189 vdd gnd cell_6t
Xbit_r190_c227 bl_227 br_227 wl_190 vdd gnd cell_6t
Xbit_r191_c227 bl_227 br_227 wl_191 vdd gnd cell_6t
Xbit_r192_c227 bl_227 br_227 wl_192 vdd gnd cell_6t
Xbit_r193_c227 bl_227 br_227 wl_193 vdd gnd cell_6t
Xbit_r194_c227 bl_227 br_227 wl_194 vdd gnd cell_6t
Xbit_r195_c227 bl_227 br_227 wl_195 vdd gnd cell_6t
Xbit_r196_c227 bl_227 br_227 wl_196 vdd gnd cell_6t
Xbit_r197_c227 bl_227 br_227 wl_197 vdd gnd cell_6t
Xbit_r198_c227 bl_227 br_227 wl_198 vdd gnd cell_6t
Xbit_r199_c227 bl_227 br_227 wl_199 vdd gnd cell_6t
Xbit_r200_c227 bl_227 br_227 wl_200 vdd gnd cell_6t
Xbit_r201_c227 bl_227 br_227 wl_201 vdd gnd cell_6t
Xbit_r202_c227 bl_227 br_227 wl_202 vdd gnd cell_6t
Xbit_r203_c227 bl_227 br_227 wl_203 vdd gnd cell_6t
Xbit_r204_c227 bl_227 br_227 wl_204 vdd gnd cell_6t
Xbit_r205_c227 bl_227 br_227 wl_205 vdd gnd cell_6t
Xbit_r206_c227 bl_227 br_227 wl_206 vdd gnd cell_6t
Xbit_r207_c227 bl_227 br_227 wl_207 vdd gnd cell_6t
Xbit_r208_c227 bl_227 br_227 wl_208 vdd gnd cell_6t
Xbit_r209_c227 bl_227 br_227 wl_209 vdd gnd cell_6t
Xbit_r210_c227 bl_227 br_227 wl_210 vdd gnd cell_6t
Xbit_r211_c227 bl_227 br_227 wl_211 vdd gnd cell_6t
Xbit_r212_c227 bl_227 br_227 wl_212 vdd gnd cell_6t
Xbit_r213_c227 bl_227 br_227 wl_213 vdd gnd cell_6t
Xbit_r214_c227 bl_227 br_227 wl_214 vdd gnd cell_6t
Xbit_r215_c227 bl_227 br_227 wl_215 vdd gnd cell_6t
Xbit_r216_c227 bl_227 br_227 wl_216 vdd gnd cell_6t
Xbit_r217_c227 bl_227 br_227 wl_217 vdd gnd cell_6t
Xbit_r218_c227 bl_227 br_227 wl_218 vdd gnd cell_6t
Xbit_r219_c227 bl_227 br_227 wl_219 vdd gnd cell_6t
Xbit_r220_c227 bl_227 br_227 wl_220 vdd gnd cell_6t
Xbit_r221_c227 bl_227 br_227 wl_221 vdd gnd cell_6t
Xbit_r222_c227 bl_227 br_227 wl_222 vdd gnd cell_6t
Xbit_r223_c227 bl_227 br_227 wl_223 vdd gnd cell_6t
Xbit_r224_c227 bl_227 br_227 wl_224 vdd gnd cell_6t
Xbit_r225_c227 bl_227 br_227 wl_225 vdd gnd cell_6t
Xbit_r226_c227 bl_227 br_227 wl_226 vdd gnd cell_6t
Xbit_r227_c227 bl_227 br_227 wl_227 vdd gnd cell_6t
Xbit_r228_c227 bl_227 br_227 wl_228 vdd gnd cell_6t
Xbit_r229_c227 bl_227 br_227 wl_229 vdd gnd cell_6t
Xbit_r230_c227 bl_227 br_227 wl_230 vdd gnd cell_6t
Xbit_r231_c227 bl_227 br_227 wl_231 vdd gnd cell_6t
Xbit_r232_c227 bl_227 br_227 wl_232 vdd gnd cell_6t
Xbit_r233_c227 bl_227 br_227 wl_233 vdd gnd cell_6t
Xbit_r234_c227 bl_227 br_227 wl_234 vdd gnd cell_6t
Xbit_r235_c227 bl_227 br_227 wl_235 vdd gnd cell_6t
Xbit_r236_c227 bl_227 br_227 wl_236 vdd gnd cell_6t
Xbit_r237_c227 bl_227 br_227 wl_237 vdd gnd cell_6t
Xbit_r238_c227 bl_227 br_227 wl_238 vdd gnd cell_6t
Xbit_r239_c227 bl_227 br_227 wl_239 vdd gnd cell_6t
Xbit_r240_c227 bl_227 br_227 wl_240 vdd gnd cell_6t
Xbit_r241_c227 bl_227 br_227 wl_241 vdd gnd cell_6t
Xbit_r242_c227 bl_227 br_227 wl_242 vdd gnd cell_6t
Xbit_r243_c227 bl_227 br_227 wl_243 vdd gnd cell_6t
Xbit_r244_c227 bl_227 br_227 wl_244 vdd gnd cell_6t
Xbit_r245_c227 bl_227 br_227 wl_245 vdd gnd cell_6t
Xbit_r246_c227 bl_227 br_227 wl_246 vdd gnd cell_6t
Xbit_r247_c227 bl_227 br_227 wl_247 vdd gnd cell_6t
Xbit_r248_c227 bl_227 br_227 wl_248 vdd gnd cell_6t
Xbit_r249_c227 bl_227 br_227 wl_249 vdd gnd cell_6t
Xbit_r250_c227 bl_227 br_227 wl_250 vdd gnd cell_6t
Xbit_r251_c227 bl_227 br_227 wl_251 vdd gnd cell_6t
Xbit_r252_c227 bl_227 br_227 wl_252 vdd gnd cell_6t
Xbit_r253_c227 bl_227 br_227 wl_253 vdd gnd cell_6t
Xbit_r254_c227 bl_227 br_227 wl_254 vdd gnd cell_6t
Xbit_r255_c227 bl_227 br_227 wl_255 vdd gnd cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd cell_6t
Xbit_r1_c228 bl_228 br_228 wl_1 vdd gnd cell_6t
Xbit_r2_c228 bl_228 br_228 wl_2 vdd gnd cell_6t
Xbit_r3_c228 bl_228 br_228 wl_3 vdd gnd cell_6t
Xbit_r4_c228 bl_228 br_228 wl_4 vdd gnd cell_6t
Xbit_r5_c228 bl_228 br_228 wl_5 vdd gnd cell_6t
Xbit_r6_c228 bl_228 br_228 wl_6 vdd gnd cell_6t
Xbit_r7_c228 bl_228 br_228 wl_7 vdd gnd cell_6t
Xbit_r8_c228 bl_228 br_228 wl_8 vdd gnd cell_6t
Xbit_r9_c228 bl_228 br_228 wl_9 vdd gnd cell_6t
Xbit_r10_c228 bl_228 br_228 wl_10 vdd gnd cell_6t
Xbit_r11_c228 bl_228 br_228 wl_11 vdd gnd cell_6t
Xbit_r12_c228 bl_228 br_228 wl_12 vdd gnd cell_6t
Xbit_r13_c228 bl_228 br_228 wl_13 vdd gnd cell_6t
Xbit_r14_c228 bl_228 br_228 wl_14 vdd gnd cell_6t
Xbit_r15_c228 bl_228 br_228 wl_15 vdd gnd cell_6t
Xbit_r16_c228 bl_228 br_228 wl_16 vdd gnd cell_6t
Xbit_r17_c228 bl_228 br_228 wl_17 vdd gnd cell_6t
Xbit_r18_c228 bl_228 br_228 wl_18 vdd gnd cell_6t
Xbit_r19_c228 bl_228 br_228 wl_19 vdd gnd cell_6t
Xbit_r20_c228 bl_228 br_228 wl_20 vdd gnd cell_6t
Xbit_r21_c228 bl_228 br_228 wl_21 vdd gnd cell_6t
Xbit_r22_c228 bl_228 br_228 wl_22 vdd gnd cell_6t
Xbit_r23_c228 bl_228 br_228 wl_23 vdd gnd cell_6t
Xbit_r24_c228 bl_228 br_228 wl_24 vdd gnd cell_6t
Xbit_r25_c228 bl_228 br_228 wl_25 vdd gnd cell_6t
Xbit_r26_c228 bl_228 br_228 wl_26 vdd gnd cell_6t
Xbit_r27_c228 bl_228 br_228 wl_27 vdd gnd cell_6t
Xbit_r28_c228 bl_228 br_228 wl_28 vdd gnd cell_6t
Xbit_r29_c228 bl_228 br_228 wl_29 vdd gnd cell_6t
Xbit_r30_c228 bl_228 br_228 wl_30 vdd gnd cell_6t
Xbit_r31_c228 bl_228 br_228 wl_31 vdd gnd cell_6t
Xbit_r32_c228 bl_228 br_228 wl_32 vdd gnd cell_6t
Xbit_r33_c228 bl_228 br_228 wl_33 vdd gnd cell_6t
Xbit_r34_c228 bl_228 br_228 wl_34 vdd gnd cell_6t
Xbit_r35_c228 bl_228 br_228 wl_35 vdd gnd cell_6t
Xbit_r36_c228 bl_228 br_228 wl_36 vdd gnd cell_6t
Xbit_r37_c228 bl_228 br_228 wl_37 vdd gnd cell_6t
Xbit_r38_c228 bl_228 br_228 wl_38 vdd gnd cell_6t
Xbit_r39_c228 bl_228 br_228 wl_39 vdd gnd cell_6t
Xbit_r40_c228 bl_228 br_228 wl_40 vdd gnd cell_6t
Xbit_r41_c228 bl_228 br_228 wl_41 vdd gnd cell_6t
Xbit_r42_c228 bl_228 br_228 wl_42 vdd gnd cell_6t
Xbit_r43_c228 bl_228 br_228 wl_43 vdd gnd cell_6t
Xbit_r44_c228 bl_228 br_228 wl_44 vdd gnd cell_6t
Xbit_r45_c228 bl_228 br_228 wl_45 vdd gnd cell_6t
Xbit_r46_c228 bl_228 br_228 wl_46 vdd gnd cell_6t
Xbit_r47_c228 bl_228 br_228 wl_47 vdd gnd cell_6t
Xbit_r48_c228 bl_228 br_228 wl_48 vdd gnd cell_6t
Xbit_r49_c228 bl_228 br_228 wl_49 vdd gnd cell_6t
Xbit_r50_c228 bl_228 br_228 wl_50 vdd gnd cell_6t
Xbit_r51_c228 bl_228 br_228 wl_51 vdd gnd cell_6t
Xbit_r52_c228 bl_228 br_228 wl_52 vdd gnd cell_6t
Xbit_r53_c228 bl_228 br_228 wl_53 vdd gnd cell_6t
Xbit_r54_c228 bl_228 br_228 wl_54 vdd gnd cell_6t
Xbit_r55_c228 bl_228 br_228 wl_55 vdd gnd cell_6t
Xbit_r56_c228 bl_228 br_228 wl_56 vdd gnd cell_6t
Xbit_r57_c228 bl_228 br_228 wl_57 vdd gnd cell_6t
Xbit_r58_c228 bl_228 br_228 wl_58 vdd gnd cell_6t
Xbit_r59_c228 bl_228 br_228 wl_59 vdd gnd cell_6t
Xbit_r60_c228 bl_228 br_228 wl_60 vdd gnd cell_6t
Xbit_r61_c228 bl_228 br_228 wl_61 vdd gnd cell_6t
Xbit_r62_c228 bl_228 br_228 wl_62 vdd gnd cell_6t
Xbit_r63_c228 bl_228 br_228 wl_63 vdd gnd cell_6t
Xbit_r64_c228 bl_228 br_228 wl_64 vdd gnd cell_6t
Xbit_r65_c228 bl_228 br_228 wl_65 vdd gnd cell_6t
Xbit_r66_c228 bl_228 br_228 wl_66 vdd gnd cell_6t
Xbit_r67_c228 bl_228 br_228 wl_67 vdd gnd cell_6t
Xbit_r68_c228 bl_228 br_228 wl_68 vdd gnd cell_6t
Xbit_r69_c228 bl_228 br_228 wl_69 vdd gnd cell_6t
Xbit_r70_c228 bl_228 br_228 wl_70 vdd gnd cell_6t
Xbit_r71_c228 bl_228 br_228 wl_71 vdd gnd cell_6t
Xbit_r72_c228 bl_228 br_228 wl_72 vdd gnd cell_6t
Xbit_r73_c228 bl_228 br_228 wl_73 vdd gnd cell_6t
Xbit_r74_c228 bl_228 br_228 wl_74 vdd gnd cell_6t
Xbit_r75_c228 bl_228 br_228 wl_75 vdd gnd cell_6t
Xbit_r76_c228 bl_228 br_228 wl_76 vdd gnd cell_6t
Xbit_r77_c228 bl_228 br_228 wl_77 vdd gnd cell_6t
Xbit_r78_c228 bl_228 br_228 wl_78 vdd gnd cell_6t
Xbit_r79_c228 bl_228 br_228 wl_79 vdd gnd cell_6t
Xbit_r80_c228 bl_228 br_228 wl_80 vdd gnd cell_6t
Xbit_r81_c228 bl_228 br_228 wl_81 vdd gnd cell_6t
Xbit_r82_c228 bl_228 br_228 wl_82 vdd gnd cell_6t
Xbit_r83_c228 bl_228 br_228 wl_83 vdd gnd cell_6t
Xbit_r84_c228 bl_228 br_228 wl_84 vdd gnd cell_6t
Xbit_r85_c228 bl_228 br_228 wl_85 vdd gnd cell_6t
Xbit_r86_c228 bl_228 br_228 wl_86 vdd gnd cell_6t
Xbit_r87_c228 bl_228 br_228 wl_87 vdd gnd cell_6t
Xbit_r88_c228 bl_228 br_228 wl_88 vdd gnd cell_6t
Xbit_r89_c228 bl_228 br_228 wl_89 vdd gnd cell_6t
Xbit_r90_c228 bl_228 br_228 wl_90 vdd gnd cell_6t
Xbit_r91_c228 bl_228 br_228 wl_91 vdd gnd cell_6t
Xbit_r92_c228 bl_228 br_228 wl_92 vdd gnd cell_6t
Xbit_r93_c228 bl_228 br_228 wl_93 vdd gnd cell_6t
Xbit_r94_c228 bl_228 br_228 wl_94 vdd gnd cell_6t
Xbit_r95_c228 bl_228 br_228 wl_95 vdd gnd cell_6t
Xbit_r96_c228 bl_228 br_228 wl_96 vdd gnd cell_6t
Xbit_r97_c228 bl_228 br_228 wl_97 vdd gnd cell_6t
Xbit_r98_c228 bl_228 br_228 wl_98 vdd gnd cell_6t
Xbit_r99_c228 bl_228 br_228 wl_99 vdd gnd cell_6t
Xbit_r100_c228 bl_228 br_228 wl_100 vdd gnd cell_6t
Xbit_r101_c228 bl_228 br_228 wl_101 vdd gnd cell_6t
Xbit_r102_c228 bl_228 br_228 wl_102 vdd gnd cell_6t
Xbit_r103_c228 bl_228 br_228 wl_103 vdd gnd cell_6t
Xbit_r104_c228 bl_228 br_228 wl_104 vdd gnd cell_6t
Xbit_r105_c228 bl_228 br_228 wl_105 vdd gnd cell_6t
Xbit_r106_c228 bl_228 br_228 wl_106 vdd gnd cell_6t
Xbit_r107_c228 bl_228 br_228 wl_107 vdd gnd cell_6t
Xbit_r108_c228 bl_228 br_228 wl_108 vdd gnd cell_6t
Xbit_r109_c228 bl_228 br_228 wl_109 vdd gnd cell_6t
Xbit_r110_c228 bl_228 br_228 wl_110 vdd gnd cell_6t
Xbit_r111_c228 bl_228 br_228 wl_111 vdd gnd cell_6t
Xbit_r112_c228 bl_228 br_228 wl_112 vdd gnd cell_6t
Xbit_r113_c228 bl_228 br_228 wl_113 vdd gnd cell_6t
Xbit_r114_c228 bl_228 br_228 wl_114 vdd gnd cell_6t
Xbit_r115_c228 bl_228 br_228 wl_115 vdd gnd cell_6t
Xbit_r116_c228 bl_228 br_228 wl_116 vdd gnd cell_6t
Xbit_r117_c228 bl_228 br_228 wl_117 vdd gnd cell_6t
Xbit_r118_c228 bl_228 br_228 wl_118 vdd gnd cell_6t
Xbit_r119_c228 bl_228 br_228 wl_119 vdd gnd cell_6t
Xbit_r120_c228 bl_228 br_228 wl_120 vdd gnd cell_6t
Xbit_r121_c228 bl_228 br_228 wl_121 vdd gnd cell_6t
Xbit_r122_c228 bl_228 br_228 wl_122 vdd gnd cell_6t
Xbit_r123_c228 bl_228 br_228 wl_123 vdd gnd cell_6t
Xbit_r124_c228 bl_228 br_228 wl_124 vdd gnd cell_6t
Xbit_r125_c228 bl_228 br_228 wl_125 vdd gnd cell_6t
Xbit_r126_c228 bl_228 br_228 wl_126 vdd gnd cell_6t
Xbit_r127_c228 bl_228 br_228 wl_127 vdd gnd cell_6t
Xbit_r128_c228 bl_228 br_228 wl_128 vdd gnd cell_6t
Xbit_r129_c228 bl_228 br_228 wl_129 vdd gnd cell_6t
Xbit_r130_c228 bl_228 br_228 wl_130 vdd gnd cell_6t
Xbit_r131_c228 bl_228 br_228 wl_131 vdd gnd cell_6t
Xbit_r132_c228 bl_228 br_228 wl_132 vdd gnd cell_6t
Xbit_r133_c228 bl_228 br_228 wl_133 vdd gnd cell_6t
Xbit_r134_c228 bl_228 br_228 wl_134 vdd gnd cell_6t
Xbit_r135_c228 bl_228 br_228 wl_135 vdd gnd cell_6t
Xbit_r136_c228 bl_228 br_228 wl_136 vdd gnd cell_6t
Xbit_r137_c228 bl_228 br_228 wl_137 vdd gnd cell_6t
Xbit_r138_c228 bl_228 br_228 wl_138 vdd gnd cell_6t
Xbit_r139_c228 bl_228 br_228 wl_139 vdd gnd cell_6t
Xbit_r140_c228 bl_228 br_228 wl_140 vdd gnd cell_6t
Xbit_r141_c228 bl_228 br_228 wl_141 vdd gnd cell_6t
Xbit_r142_c228 bl_228 br_228 wl_142 vdd gnd cell_6t
Xbit_r143_c228 bl_228 br_228 wl_143 vdd gnd cell_6t
Xbit_r144_c228 bl_228 br_228 wl_144 vdd gnd cell_6t
Xbit_r145_c228 bl_228 br_228 wl_145 vdd gnd cell_6t
Xbit_r146_c228 bl_228 br_228 wl_146 vdd gnd cell_6t
Xbit_r147_c228 bl_228 br_228 wl_147 vdd gnd cell_6t
Xbit_r148_c228 bl_228 br_228 wl_148 vdd gnd cell_6t
Xbit_r149_c228 bl_228 br_228 wl_149 vdd gnd cell_6t
Xbit_r150_c228 bl_228 br_228 wl_150 vdd gnd cell_6t
Xbit_r151_c228 bl_228 br_228 wl_151 vdd gnd cell_6t
Xbit_r152_c228 bl_228 br_228 wl_152 vdd gnd cell_6t
Xbit_r153_c228 bl_228 br_228 wl_153 vdd gnd cell_6t
Xbit_r154_c228 bl_228 br_228 wl_154 vdd gnd cell_6t
Xbit_r155_c228 bl_228 br_228 wl_155 vdd gnd cell_6t
Xbit_r156_c228 bl_228 br_228 wl_156 vdd gnd cell_6t
Xbit_r157_c228 bl_228 br_228 wl_157 vdd gnd cell_6t
Xbit_r158_c228 bl_228 br_228 wl_158 vdd gnd cell_6t
Xbit_r159_c228 bl_228 br_228 wl_159 vdd gnd cell_6t
Xbit_r160_c228 bl_228 br_228 wl_160 vdd gnd cell_6t
Xbit_r161_c228 bl_228 br_228 wl_161 vdd gnd cell_6t
Xbit_r162_c228 bl_228 br_228 wl_162 vdd gnd cell_6t
Xbit_r163_c228 bl_228 br_228 wl_163 vdd gnd cell_6t
Xbit_r164_c228 bl_228 br_228 wl_164 vdd gnd cell_6t
Xbit_r165_c228 bl_228 br_228 wl_165 vdd gnd cell_6t
Xbit_r166_c228 bl_228 br_228 wl_166 vdd gnd cell_6t
Xbit_r167_c228 bl_228 br_228 wl_167 vdd gnd cell_6t
Xbit_r168_c228 bl_228 br_228 wl_168 vdd gnd cell_6t
Xbit_r169_c228 bl_228 br_228 wl_169 vdd gnd cell_6t
Xbit_r170_c228 bl_228 br_228 wl_170 vdd gnd cell_6t
Xbit_r171_c228 bl_228 br_228 wl_171 vdd gnd cell_6t
Xbit_r172_c228 bl_228 br_228 wl_172 vdd gnd cell_6t
Xbit_r173_c228 bl_228 br_228 wl_173 vdd gnd cell_6t
Xbit_r174_c228 bl_228 br_228 wl_174 vdd gnd cell_6t
Xbit_r175_c228 bl_228 br_228 wl_175 vdd gnd cell_6t
Xbit_r176_c228 bl_228 br_228 wl_176 vdd gnd cell_6t
Xbit_r177_c228 bl_228 br_228 wl_177 vdd gnd cell_6t
Xbit_r178_c228 bl_228 br_228 wl_178 vdd gnd cell_6t
Xbit_r179_c228 bl_228 br_228 wl_179 vdd gnd cell_6t
Xbit_r180_c228 bl_228 br_228 wl_180 vdd gnd cell_6t
Xbit_r181_c228 bl_228 br_228 wl_181 vdd gnd cell_6t
Xbit_r182_c228 bl_228 br_228 wl_182 vdd gnd cell_6t
Xbit_r183_c228 bl_228 br_228 wl_183 vdd gnd cell_6t
Xbit_r184_c228 bl_228 br_228 wl_184 vdd gnd cell_6t
Xbit_r185_c228 bl_228 br_228 wl_185 vdd gnd cell_6t
Xbit_r186_c228 bl_228 br_228 wl_186 vdd gnd cell_6t
Xbit_r187_c228 bl_228 br_228 wl_187 vdd gnd cell_6t
Xbit_r188_c228 bl_228 br_228 wl_188 vdd gnd cell_6t
Xbit_r189_c228 bl_228 br_228 wl_189 vdd gnd cell_6t
Xbit_r190_c228 bl_228 br_228 wl_190 vdd gnd cell_6t
Xbit_r191_c228 bl_228 br_228 wl_191 vdd gnd cell_6t
Xbit_r192_c228 bl_228 br_228 wl_192 vdd gnd cell_6t
Xbit_r193_c228 bl_228 br_228 wl_193 vdd gnd cell_6t
Xbit_r194_c228 bl_228 br_228 wl_194 vdd gnd cell_6t
Xbit_r195_c228 bl_228 br_228 wl_195 vdd gnd cell_6t
Xbit_r196_c228 bl_228 br_228 wl_196 vdd gnd cell_6t
Xbit_r197_c228 bl_228 br_228 wl_197 vdd gnd cell_6t
Xbit_r198_c228 bl_228 br_228 wl_198 vdd gnd cell_6t
Xbit_r199_c228 bl_228 br_228 wl_199 vdd gnd cell_6t
Xbit_r200_c228 bl_228 br_228 wl_200 vdd gnd cell_6t
Xbit_r201_c228 bl_228 br_228 wl_201 vdd gnd cell_6t
Xbit_r202_c228 bl_228 br_228 wl_202 vdd gnd cell_6t
Xbit_r203_c228 bl_228 br_228 wl_203 vdd gnd cell_6t
Xbit_r204_c228 bl_228 br_228 wl_204 vdd gnd cell_6t
Xbit_r205_c228 bl_228 br_228 wl_205 vdd gnd cell_6t
Xbit_r206_c228 bl_228 br_228 wl_206 vdd gnd cell_6t
Xbit_r207_c228 bl_228 br_228 wl_207 vdd gnd cell_6t
Xbit_r208_c228 bl_228 br_228 wl_208 vdd gnd cell_6t
Xbit_r209_c228 bl_228 br_228 wl_209 vdd gnd cell_6t
Xbit_r210_c228 bl_228 br_228 wl_210 vdd gnd cell_6t
Xbit_r211_c228 bl_228 br_228 wl_211 vdd gnd cell_6t
Xbit_r212_c228 bl_228 br_228 wl_212 vdd gnd cell_6t
Xbit_r213_c228 bl_228 br_228 wl_213 vdd gnd cell_6t
Xbit_r214_c228 bl_228 br_228 wl_214 vdd gnd cell_6t
Xbit_r215_c228 bl_228 br_228 wl_215 vdd gnd cell_6t
Xbit_r216_c228 bl_228 br_228 wl_216 vdd gnd cell_6t
Xbit_r217_c228 bl_228 br_228 wl_217 vdd gnd cell_6t
Xbit_r218_c228 bl_228 br_228 wl_218 vdd gnd cell_6t
Xbit_r219_c228 bl_228 br_228 wl_219 vdd gnd cell_6t
Xbit_r220_c228 bl_228 br_228 wl_220 vdd gnd cell_6t
Xbit_r221_c228 bl_228 br_228 wl_221 vdd gnd cell_6t
Xbit_r222_c228 bl_228 br_228 wl_222 vdd gnd cell_6t
Xbit_r223_c228 bl_228 br_228 wl_223 vdd gnd cell_6t
Xbit_r224_c228 bl_228 br_228 wl_224 vdd gnd cell_6t
Xbit_r225_c228 bl_228 br_228 wl_225 vdd gnd cell_6t
Xbit_r226_c228 bl_228 br_228 wl_226 vdd gnd cell_6t
Xbit_r227_c228 bl_228 br_228 wl_227 vdd gnd cell_6t
Xbit_r228_c228 bl_228 br_228 wl_228 vdd gnd cell_6t
Xbit_r229_c228 bl_228 br_228 wl_229 vdd gnd cell_6t
Xbit_r230_c228 bl_228 br_228 wl_230 vdd gnd cell_6t
Xbit_r231_c228 bl_228 br_228 wl_231 vdd gnd cell_6t
Xbit_r232_c228 bl_228 br_228 wl_232 vdd gnd cell_6t
Xbit_r233_c228 bl_228 br_228 wl_233 vdd gnd cell_6t
Xbit_r234_c228 bl_228 br_228 wl_234 vdd gnd cell_6t
Xbit_r235_c228 bl_228 br_228 wl_235 vdd gnd cell_6t
Xbit_r236_c228 bl_228 br_228 wl_236 vdd gnd cell_6t
Xbit_r237_c228 bl_228 br_228 wl_237 vdd gnd cell_6t
Xbit_r238_c228 bl_228 br_228 wl_238 vdd gnd cell_6t
Xbit_r239_c228 bl_228 br_228 wl_239 vdd gnd cell_6t
Xbit_r240_c228 bl_228 br_228 wl_240 vdd gnd cell_6t
Xbit_r241_c228 bl_228 br_228 wl_241 vdd gnd cell_6t
Xbit_r242_c228 bl_228 br_228 wl_242 vdd gnd cell_6t
Xbit_r243_c228 bl_228 br_228 wl_243 vdd gnd cell_6t
Xbit_r244_c228 bl_228 br_228 wl_244 vdd gnd cell_6t
Xbit_r245_c228 bl_228 br_228 wl_245 vdd gnd cell_6t
Xbit_r246_c228 bl_228 br_228 wl_246 vdd gnd cell_6t
Xbit_r247_c228 bl_228 br_228 wl_247 vdd gnd cell_6t
Xbit_r248_c228 bl_228 br_228 wl_248 vdd gnd cell_6t
Xbit_r249_c228 bl_228 br_228 wl_249 vdd gnd cell_6t
Xbit_r250_c228 bl_228 br_228 wl_250 vdd gnd cell_6t
Xbit_r251_c228 bl_228 br_228 wl_251 vdd gnd cell_6t
Xbit_r252_c228 bl_228 br_228 wl_252 vdd gnd cell_6t
Xbit_r253_c228 bl_228 br_228 wl_253 vdd gnd cell_6t
Xbit_r254_c228 bl_228 br_228 wl_254 vdd gnd cell_6t
Xbit_r255_c228 bl_228 br_228 wl_255 vdd gnd cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd cell_6t
Xbit_r1_c229 bl_229 br_229 wl_1 vdd gnd cell_6t
Xbit_r2_c229 bl_229 br_229 wl_2 vdd gnd cell_6t
Xbit_r3_c229 bl_229 br_229 wl_3 vdd gnd cell_6t
Xbit_r4_c229 bl_229 br_229 wl_4 vdd gnd cell_6t
Xbit_r5_c229 bl_229 br_229 wl_5 vdd gnd cell_6t
Xbit_r6_c229 bl_229 br_229 wl_6 vdd gnd cell_6t
Xbit_r7_c229 bl_229 br_229 wl_7 vdd gnd cell_6t
Xbit_r8_c229 bl_229 br_229 wl_8 vdd gnd cell_6t
Xbit_r9_c229 bl_229 br_229 wl_9 vdd gnd cell_6t
Xbit_r10_c229 bl_229 br_229 wl_10 vdd gnd cell_6t
Xbit_r11_c229 bl_229 br_229 wl_11 vdd gnd cell_6t
Xbit_r12_c229 bl_229 br_229 wl_12 vdd gnd cell_6t
Xbit_r13_c229 bl_229 br_229 wl_13 vdd gnd cell_6t
Xbit_r14_c229 bl_229 br_229 wl_14 vdd gnd cell_6t
Xbit_r15_c229 bl_229 br_229 wl_15 vdd gnd cell_6t
Xbit_r16_c229 bl_229 br_229 wl_16 vdd gnd cell_6t
Xbit_r17_c229 bl_229 br_229 wl_17 vdd gnd cell_6t
Xbit_r18_c229 bl_229 br_229 wl_18 vdd gnd cell_6t
Xbit_r19_c229 bl_229 br_229 wl_19 vdd gnd cell_6t
Xbit_r20_c229 bl_229 br_229 wl_20 vdd gnd cell_6t
Xbit_r21_c229 bl_229 br_229 wl_21 vdd gnd cell_6t
Xbit_r22_c229 bl_229 br_229 wl_22 vdd gnd cell_6t
Xbit_r23_c229 bl_229 br_229 wl_23 vdd gnd cell_6t
Xbit_r24_c229 bl_229 br_229 wl_24 vdd gnd cell_6t
Xbit_r25_c229 bl_229 br_229 wl_25 vdd gnd cell_6t
Xbit_r26_c229 bl_229 br_229 wl_26 vdd gnd cell_6t
Xbit_r27_c229 bl_229 br_229 wl_27 vdd gnd cell_6t
Xbit_r28_c229 bl_229 br_229 wl_28 vdd gnd cell_6t
Xbit_r29_c229 bl_229 br_229 wl_29 vdd gnd cell_6t
Xbit_r30_c229 bl_229 br_229 wl_30 vdd gnd cell_6t
Xbit_r31_c229 bl_229 br_229 wl_31 vdd gnd cell_6t
Xbit_r32_c229 bl_229 br_229 wl_32 vdd gnd cell_6t
Xbit_r33_c229 bl_229 br_229 wl_33 vdd gnd cell_6t
Xbit_r34_c229 bl_229 br_229 wl_34 vdd gnd cell_6t
Xbit_r35_c229 bl_229 br_229 wl_35 vdd gnd cell_6t
Xbit_r36_c229 bl_229 br_229 wl_36 vdd gnd cell_6t
Xbit_r37_c229 bl_229 br_229 wl_37 vdd gnd cell_6t
Xbit_r38_c229 bl_229 br_229 wl_38 vdd gnd cell_6t
Xbit_r39_c229 bl_229 br_229 wl_39 vdd gnd cell_6t
Xbit_r40_c229 bl_229 br_229 wl_40 vdd gnd cell_6t
Xbit_r41_c229 bl_229 br_229 wl_41 vdd gnd cell_6t
Xbit_r42_c229 bl_229 br_229 wl_42 vdd gnd cell_6t
Xbit_r43_c229 bl_229 br_229 wl_43 vdd gnd cell_6t
Xbit_r44_c229 bl_229 br_229 wl_44 vdd gnd cell_6t
Xbit_r45_c229 bl_229 br_229 wl_45 vdd gnd cell_6t
Xbit_r46_c229 bl_229 br_229 wl_46 vdd gnd cell_6t
Xbit_r47_c229 bl_229 br_229 wl_47 vdd gnd cell_6t
Xbit_r48_c229 bl_229 br_229 wl_48 vdd gnd cell_6t
Xbit_r49_c229 bl_229 br_229 wl_49 vdd gnd cell_6t
Xbit_r50_c229 bl_229 br_229 wl_50 vdd gnd cell_6t
Xbit_r51_c229 bl_229 br_229 wl_51 vdd gnd cell_6t
Xbit_r52_c229 bl_229 br_229 wl_52 vdd gnd cell_6t
Xbit_r53_c229 bl_229 br_229 wl_53 vdd gnd cell_6t
Xbit_r54_c229 bl_229 br_229 wl_54 vdd gnd cell_6t
Xbit_r55_c229 bl_229 br_229 wl_55 vdd gnd cell_6t
Xbit_r56_c229 bl_229 br_229 wl_56 vdd gnd cell_6t
Xbit_r57_c229 bl_229 br_229 wl_57 vdd gnd cell_6t
Xbit_r58_c229 bl_229 br_229 wl_58 vdd gnd cell_6t
Xbit_r59_c229 bl_229 br_229 wl_59 vdd gnd cell_6t
Xbit_r60_c229 bl_229 br_229 wl_60 vdd gnd cell_6t
Xbit_r61_c229 bl_229 br_229 wl_61 vdd gnd cell_6t
Xbit_r62_c229 bl_229 br_229 wl_62 vdd gnd cell_6t
Xbit_r63_c229 bl_229 br_229 wl_63 vdd gnd cell_6t
Xbit_r64_c229 bl_229 br_229 wl_64 vdd gnd cell_6t
Xbit_r65_c229 bl_229 br_229 wl_65 vdd gnd cell_6t
Xbit_r66_c229 bl_229 br_229 wl_66 vdd gnd cell_6t
Xbit_r67_c229 bl_229 br_229 wl_67 vdd gnd cell_6t
Xbit_r68_c229 bl_229 br_229 wl_68 vdd gnd cell_6t
Xbit_r69_c229 bl_229 br_229 wl_69 vdd gnd cell_6t
Xbit_r70_c229 bl_229 br_229 wl_70 vdd gnd cell_6t
Xbit_r71_c229 bl_229 br_229 wl_71 vdd gnd cell_6t
Xbit_r72_c229 bl_229 br_229 wl_72 vdd gnd cell_6t
Xbit_r73_c229 bl_229 br_229 wl_73 vdd gnd cell_6t
Xbit_r74_c229 bl_229 br_229 wl_74 vdd gnd cell_6t
Xbit_r75_c229 bl_229 br_229 wl_75 vdd gnd cell_6t
Xbit_r76_c229 bl_229 br_229 wl_76 vdd gnd cell_6t
Xbit_r77_c229 bl_229 br_229 wl_77 vdd gnd cell_6t
Xbit_r78_c229 bl_229 br_229 wl_78 vdd gnd cell_6t
Xbit_r79_c229 bl_229 br_229 wl_79 vdd gnd cell_6t
Xbit_r80_c229 bl_229 br_229 wl_80 vdd gnd cell_6t
Xbit_r81_c229 bl_229 br_229 wl_81 vdd gnd cell_6t
Xbit_r82_c229 bl_229 br_229 wl_82 vdd gnd cell_6t
Xbit_r83_c229 bl_229 br_229 wl_83 vdd gnd cell_6t
Xbit_r84_c229 bl_229 br_229 wl_84 vdd gnd cell_6t
Xbit_r85_c229 bl_229 br_229 wl_85 vdd gnd cell_6t
Xbit_r86_c229 bl_229 br_229 wl_86 vdd gnd cell_6t
Xbit_r87_c229 bl_229 br_229 wl_87 vdd gnd cell_6t
Xbit_r88_c229 bl_229 br_229 wl_88 vdd gnd cell_6t
Xbit_r89_c229 bl_229 br_229 wl_89 vdd gnd cell_6t
Xbit_r90_c229 bl_229 br_229 wl_90 vdd gnd cell_6t
Xbit_r91_c229 bl_229 br_229 wl_91 vdd gnd cell_6t
Xbit_r92_c229 bl_229 br_229 wl_92 vdd gnd cell_6t
Xbit_r93_c229 bl_229 br_229 wl_93 vdd gnd cell_6t
Xbit_r94_c229 bl_229 br_229 wl_94 vdd gnd cell_6t
Xbit_r95_c229 bl_229 br_229 wl_95 vdd gnd cell_6t
Xbit_r96_c229 bl_229 br_229 wl_96 vdd gnd cell_6t
Xbit_r97_c229 bl_229 br_229 wl_97 vdd gnd cell_6t
Xbit_r98_c229 bl_229 br_229 wl_98 vdd gnd cell_6t
Xbit_r99_c229 bl_229 br_229 wl_99 vdd gnd cell_6t
Xbit_r100_c229 bl_229 br_229 wl_100 vdd gnd cell_6t
Xbit_r101_c229 bl_229 br_229 wl_101 vdd gnd cell_6t
Xbit_r102_c229 bl_229 br_229 wl_102 vdd gnd cell_6t
Xbit_r103_c229 bl_229 br_229 wl_103 vdd gnd cell_6t
Xbit_r104_c229 bl_229 br_229 wl_104 vdd gnd cell_6t
Xbit_r105_c229 bl_229 br_229 wl_105 vdd gnd cell_6t
Xbit_r106_c229 bl_229 br_229 wl_106 vdd gnd cell_6t
Xbit_r107_c229 bl_229 br_229 wl_107 vdd gnd cell_6t
Xbit_r108_c229 bl_229 br_229 wl_108 vdd gnd cell_6t
Xbit_r109_c229 bl_229 br_229 wl_109 vdd gnd cell_6t
Xbit_r110_c229 bl_229 br_229 wl_110 vdd gnd cell_6t
Xbit_r111_c229 bl_229 br_229 wl_111 vdd gnd cell_6t
Xbit_r112_c229 bl_229 br_229 wl_112 vdd gnd cell_6t
Xbit_r113_c229 bl_229 br_229 wl_113 vdd gnd cell_6t
Xbit_r114_c229 bl_229 br_229 wl_114 vdd gnd cell_6t
Xbit_r115_c229 bl_229 br_229 wl_115 vdd gnd cell_6t
Xbit_r116_c229 bl_229 br_229 wl_116 vdd gnd cell_6t
Xbit_r117_c229 bl_229 br_229 wl_117 vdd gnd cell_6t
Xbit_r118_c229 bl_229 br_229 wl_118 vdd gnd cell_6t
Xbit_r119_c229 bl_229 br_229 wl_119 vdd gnd cell_6t
Xbit_r120_c229 bl_229 br_229 wl_120 vdd gnd cell_6t
Xbit_r121_c229 bl_229 br_229 wl_121 vdd gnd cell_6t
Xbit_r122_c229 bl_229 br_229 wl_122 vdd gnd cell_6t
Xbit_r123_c229 bl_229 br_229 wl_123 vdd gnd cell_6t
Xbit_r124_c229 bl_229 br_229 wl_124 vdd gnd cell_6t
Xbit_r125_c229 bl_229 br_229 wl_125 vdd gnd cell_6t
Xbit_r126_c229 bl_229 br_229 wl_126 vdd gnd cell_6t
Xbit_r127_c229 bl_229 br_229 wl_127 vdd gnd cell_6t
Xbit_r128_c229 bl_229 br_229 wl_128 vdd gnd cell_6t
Xbit_r129_c229 bl_229 br_229 wl_129 vdd gnd cell_6t
Xbit_r130_c229 bl_229 br_229 wl_130 vdd gnd cell_6t
Xbit_r131_c229 bl_229 br_229 wl_131 vdd gnd cell_6t
Xbit_r132_c229 bl_229 br_229 wl_132 vdd gnd cell_6t
Xbit_r133_c229 bl_229 br_229 wl_133 vdd gnd cell_6t
Xbit_r134_c229 bl_229 br_229 wl_134 vdd gnd cell_6t
Xbit_r135_c229 bl_229 br_229 wl_135 vdd gnd cell_6t
Xbit_r136_c229 bl_229 br_229 wl_136 vdd gnd cell_6t
Xbit_r137_c229 bl_229 br_229 wl_137 vdd gnd cell_6t
Xbit_r138_c229 bl_229 br_229 wl_138 vdd gnd cell_6t
Xbit_r139_c229 bl_229 br_229 wl_139 vdd gnd cell_6t
Xbit_r140_c229 bl_229 br_229 wl_140 vdd gnd cell_6t
Xbit_r141_c229 bl_229 br_229 wl_141 vdd gnd cell_6t
Xbit_r142_c229 bl_229 br_229 wl_142 vdd gnd cell_6t
Xbit_r143_c229 bl_229 br_229 wl_143 vdd gnd cell_6t
Xbit_r144_c229 bl_229 br_229 wl_144 vdd gnd cell_6t
Xbit_r145_c229 bl_229 br_229 wl_145 vdd gnd cell_6t
Xbit_r146_c229 bl_229 br_229 wl_146 vdd gnd cell_6t
Xbit_r147_c229 bl_229 br_229 wl_147 vdd gnd cell_6t
Xbit_r148_c229 bl_229 br_229 wl_148 vdd gnd cell_6t
Xbit_r149_c229 bl_229 br_229 wl_149 vdd gnd cell_6t
Xbit_r150_c229 bl_229 br_229 wl_150 vdd gnd cell_6t
Xbit_r151_c229 bl_229 br_229 wl_151 vdd gnd cell_6t
Xbit_r152_c229 bl_229 br_229 wl_152 vdd gnd cell_6t
Xbit_r153_c229 bl_229 br_229 wl_153 vdd gnd cell_6t
Xbit_r154_c229 bl_229 br_229 wl_154 vdd gnd cell_6t
Xbit_r155_c229 bl_229 br_229 wl_155 vdd gnd cell_6t
Xbit_r156_c229 bl_229 br_229 wl_156 vdd gnd cell_6t
Xbit_r157_c229 bl_229 br_229 wl_157 vdd gnd cell_6t
Xbit_r158_c229 bl_229 br_229 wl_158 vdd gnd cell_6t
Xbit_r159_c229 bl_229 br_229 wl_159 vdd gnd cell_6t
Xbit_r160_c229 bl_229 br_229 wl_160 vdd gnd cell_6t
Xbit_r161_c229 bl_229 br_229 wl_161 vdd gnd cell_6t
Xbit_r162_c229 bl_229 br_229 wl_162 vdd gnd cell_6t
Xbit_r163_c229 bl_229 br_229 wl_163 vdd gnd cell_6t
Xbit_r164_c229 bl_229 br_229 wl_164 vdd gnd cell_6t
Xbit_r165_c229 bl_229 br_229 wl_165 vdd gnd cell_6t
Xbit_r166_c229 bl_229 br_229 wl_166 vdd gnd cell_6t
Xbit_r167_c229 bl_229 br_229 wl_167 vdd gnd cell_6t
Xbit_r168_c229 bl_229 br_229 wl_168 vdd gnd cell_6t
Xbit_r169_c229 bl_229 br_229 wl_169 vdd gnd cell_6t
Xbit_r170_c229 bl_229 br_229 wl_170 vdd gnd cell_6t
Xbit_r171_c229 bl_229 br_229 wl_171 vdd gnd cell_6t
Xbit_r172_c229 bl_229 br_229 wl_172 vdd gnd cell_6t
Xbit_r173_c229 bl_229 br_229 wl_173 vdd gnd cell_6t
Xbit_r174_c229 bl_229 br_229 wl_174 vdd gnd cell_6t
Xbit_r175_c229 bl_229 br_229 wl_175 vdd gnd cell_6t
Xbit_r176_c229 bl_229 br_229 wl_176 vdd gnd cell_6t
Xbit_r177_c229 bl_229 br_229 wl_177 vdd gnd cell_6t
Xbit_r178_c229 bl_229 br_229 wl_178 vdd gnd cell_6t
Xbit_r179_c229 bl_229 br_229 wl_179 vdd gnd cell_6t
Xbit_r180_c229 bl_229 br_229 wl_180 vdd gnd cell_6t
Xbit_r181_c229 bl_229 br_229 wl_181 vdd gnd cell_6t
Xbit_r182_c229 bl_229 br_229 wl_182 vdd gnd cell_6t
Xbit_r183_c229 bl_229 br_229 wl_183 vdd gnd cell_6t
Xbit_r184_c229 bl_229 br_229 wl_184 vdd gnd cell_6t
Xbit_r185_c229 bl_229 br_229 wl_185 vdd gnd cell_6t
Xbit_r186_c229 bl_229 br_229 wl_186 vdd gnd cell_6t
Xbit_r187_c229 bl_229 br_229 wl_187 vdd gnd cell_6t
Xbit_r188_c229 bl_229 br_229 wl_188 vdd gnd cell_6t
Xbit_r189_c229 bl_229 br_229 wl_189 vdd gnd cell_6t
Xbit_r190_c229 bl_229 br_229 wl_190 vdd gnd cell_6t
Xbit_r191_c229 bl_229 br_229 wl_191 vdd gnd cell_6t
Xbit_r192_c229 bl_229 br_229 wl_192 vdd gnd cell_6t
Xbit_r193_c229 bl_229 br_229 wl_193 vdd gnd cell_6t
Xbit_r194_c229 bl_229 br_229 wl_194 vdd gnd cell_6t
Xbit_r195_c229 bl_229 br_229 wl_195 vdd gnd cell_6t
Xbit_r196_c229 bl_229 br_229 wl_196 vdd gnd cell_6t
Xbit_r197_c229 bl_229 br_229 wl_197 vdd gnd cell_6t
Xbit_r198_c229 bl_229 br_229 wl_198 vdd gnd cell_6t
Xbit_r199_c229 bl_229 br_229 wl_199 vdd gnd cell_6t
Xbit_r200_c229 bl_229 br_229 wl_200 vdd gnd cell_6t
Xbit_r201_c229 bl_229 br_229 wl_201 vdd gnd cell_6t
Xbit_r202_c229 bl_229 br_229 wl_202 vdd gnd cell_6t
Xbit_r203_c229 bl_229 br_229 wl_203 vdd gnd cell_6t
Xbit_r204_c229 bl_229 br_229 wl_204 vdd gnd cell_6t
Xbit_r205_c229 bl_229 br_229 wl_205 vdd gnd cell_6t
Xbit_r206_c229 bl_229 br_229 wl_206 vdd gnd cell_6t
Xbit_r207_c229 bl_229 br_229 wl_207 vdd gnd cell_6t
Xbit_r208_c229 bl_229 br_229 wl_208 vdd gnd cell_6t
Xbit_r209_c229 bl_229 br_229 wl_209 vdd gnd cell_6t
Xbit_r210_c229 bl_229 br_229 wl_210 vdd gnd cell_6t
Xbit_r211_c229 bl_229 br_229 wl_211 vdd gnd cell_6t
Xbit_r212_c229 bl_229 br_229 wl_212 vdd gnd cell_6t
Xbit_r213_c229 bl_229 br_229 wl_213 vdd gnd cell_6t
Xbit_r214_c229 bl_229 br_229 wl_214 vdd gnd cell_6t
Xbit_r215_c229 bl_229 br_229 wl_215 vdd gnd cell_6t
Xbit_r216_c229 bl_229 br_229 wl_216 vdd gnd cell_6t
Xbit_r217_c229 bl_229 br_229 wl_217 vdd gnd cell_6t
Xbit_r218_c229 bl_229 br_229 wl_218 vdd gnd cell_6t
Xbit_r219_c229 bl_229 br_229 wl_219 vdd gnd cell_6t
Xbit_r220_c229 bl_229 br_229 wl_220 vdd gnd cell_6t
Xbit_r221_c229 bl_229 br_229 wl_221 vdd gnd cell_6t
Xbit_r222_c229 bl_229 br_229 wl_222 vdd gnd cell_6t
Xbit_r223_c229 bl_229 br_229 wl_223 vdd gnd cell_6t
Xbit_r224_c229 bl_229 br_229 wl_224 vdd gnd cell_6t
Xbit_r225_c229 bl_229 br_229 wl_225 vdd gnd cell_6t
Xbit_r226_c229 bl_229 br_229 wl_226 vdd gnd cell_6t
Xbit_r227_c229 bl_229 br_229 wl_227 vdd gnd cell_6t
Xbit_r228_c229 bl_229 br_229 wl_228 vdd gnd cell_6t
Xbit_r229_c229 bl_229 br_229 wl_229 vdd gnd cell_6t
Xbit_r230_c229 bl_229 br_229 wl_230 vdd gnd cell_6t
Xbit_r231_c229 bl_229 br_229 wl_231 vdd gnd cell_6t
Xbit_r232_c229 bl_229 br_229 wl_232 vdd gnd cell_6t
Xbit_r233_c229 bl_229 br_229 wl_233 vdd gnd cell_6t
Xbit_r234_c229 bl_229 br_229 wl_234 vdd gnd cell_6t
Xbit_r235_c229 bl_229 br_229 wl_235 vdd gnd cell_6t
Xbit_r236_c229 bl_229 br_229 wl_236 vdd gnd cell_6t
Xbit_r237_c229 bl_229 br_229 wl_237 vdd gnd cell_6t
Xbit_r238_c229 bl_229 br_229 wl_238 vdd gnd cell_6t
Xbit_r239_c229 bl_229 br_229 wl_239 vdd gnd cell_6t
Xbit_r240_c229 bl_229 br_229 wl_240 vdd gnd cell_6t
Xbit_r241_c229 bl_229 br_229 wl_241 vdd gnd cell_6t
Xbit_r242_c229 bl_229 br_229 wl_242 vdd gnd cell_6t
Xbit_r243_c229 bl_229 br_229 wl_243 vdd gnd cell_6t
Xbit_r244_c229 bl_229 br_229 wl_244 vdd gnd cell_6t
Xbit_r245_c229 bl_229 br_229 wl_245 vdd gnd cell_6t
Xbit_r246_c229 bl_229 br_229 wl_246 vdd gnd cell_6t
Xbit_r247_c229 bl_229 br_229 wl_247 vdd gnd cell_6t
Xbit_r248_c229 bl_229 br_229 wl_248 vdd gnd cell_6t
Xbit_r249_c229 bl_229 br_229 wl_249 vdd gnd cell_6t
Xbit_r250_c229 bl_229 br_229 wl_250 vdd gnd cell_6t
Xbit_r251_c229 bl_229 br_229 wl_251 vdd gnd cell_6t
Xbit_r252_c229 bl_229 br_229 wl_252 vdd gnd cell_6t
Xbit_r253_c229 bl_229 br_229 wl_253 vdd gnd cell_6t
Xbit_r254_c229 bl_229 br_229 wl_254 vdd gnd cell_6t
Xbit_r255_c229 bl_229 br_229 wl_255 vdd gnd cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd cell_6t
Xbit_r1_c230 bl_230 br_230 wl_1 vdd gnd cell_6t
Xbit_r2_c230 bl_230 br_230 wl_2 vdd gnd cell_6t
Xbit_r3_c230 bl_230 br_230 wl_3 vdd gnd cell_6t
Xbit_r4_c230 bl_230 br_230 wl_4 vdd gnd cell_6t
Xbit_r5_c230 bl_230 br_230 wl_5 vdd gnd cell_6t
Xbit_r6_c230 bl_230 br_230 wl_6 vdd gnd cell_6t
Xbit_r7_c230 bl_230 br_230 wl_7 vdd gnd cell_6t
Xbit_r8_c230 bl_230 br_230 wl_8 vdd gnd cell_6t
Xbit_r9_c230 bl_230 br_230 wl_9 vdd gnd cell_6t
Xbit_r10_c230 bl_230 br_230 wl_10 vdd gnd cell_6t
Xbit_r11_c230 bl_230 br_230 wl_11 vdd gnd cell_6t
Xbit_r12_c230 bl_230 br_230 wl_12 vdd gnd cell_6t
Xbit_r13_c230 bl_230 br_230 wl_13 vdd gnd cell_6t
Xbit_r14_c230 bl_230 br_230 wl_14 vdd gnd cell_6t
Xbit_r15_c230 bl_230 br_230 wl_15 vdd gnd cell_6t
Xbit_r16_c230 bl_230 br_230 wl_16 vdd gnd cell_6t
Xbit_r17_c230 bl_230 br_230 wl_17 vdd gnd cell_6t
Xbit_r18_c230 bl_230 br_230 wl_18 vdd gnd cell_6t
Xbit_r19_c230 bl_230 br_230 wl_19 vdd gnd cell_6t
Xbit_r20_c230 bl_230 br_230 wl_20 vdd gnd cell_6t
Xbit_r21_c230 bl_230 br_230 wl_21 vdd gnd cell_6t
Xbit_r22_c230 bl_230 br_230 wl_22 vdd gnd cell_6t
Xbit_r23_c230 bl_230 br_230 wl_23 vdd gnd cell_6t
Xbit_r24_c230 bl_230 br_230 wl_24 vdd gnd cell_6t
Xbit_r25_c230 bl_230 br_230 wl_25 vdd gnd cell_6t
Xbit_r26_c230 bl_230 br_230 wl_26 vdd gnd cell_6t
Xbit_r27_c230 bl_230 br_230 wl_27 vdd gnd cell_6t
Xbit_r28_c230 bl_230 br_230 wl_28 vdd gnd cell_6t
Xbit_r29_c230 bl_230 br_230 wl_29 vdd gnd cell_6t
Xbit_r30_c230 bl_230 br_230 wl_30 vdd gnd cell_6t
Xbit_r31_c230 bl_230 br_230 wl_31 vdd gnd cell_6t
Xbit_r32_c230 bl_230 br_230 wl_32 vdd gnd cell_6t
Xbit_r33_c230 bl_230 br_230 wl_33 vdd gnd cell_6t
Xbit_r34_c230 bl_230 br_230 wl_34 vdd gnd cell_6t
Xbit_r35_c230 bl_230 br_230 wl_35 vdd gnd cell_6t
Xbit_r36_c230 bl_230 br_230 wl_36 vdd gnd cell_6t
Xbit_r37_c230 bl_230 br_230 wl_37 vdd gnd cell_6t
Xbit_r38_c230 bl_230 br_230 wl_38 vdd gnd cell_6t
Xbit_r39_c230 bl_230 br_230 wl_39 vdd gnd cell_6t
Xbit_r40_c230 bl_230 br_230 wl_40 vdd gnd cell_6t
Xbit_r41_c230 bl_230 br_230 wl_41 vdd gnd cell_6t
Xbit_r42_c230 bl_230 br_230 wl_42 vdd gnd cell_6t
Xbit_r43_c230 bl_230 br_230 wl_43 vdd gnd cell_6t
Xbit_r44_c230 bl_230 br_230 wl_44 vdd gnd cell_6t
Xbit_r45_c230 bl_230 br_230 wl_45 vdd gnd cell_6t
Xbit_r46_c230 bl_230 br_230 wl_46 vdd gnd cell_6t
Xbit_r47_c230 bl_230 br_230 wl_47 vdd gnd cell_6t
Xbit_r48_c230 bl_230 br_230 wl_48 vdd gnd cell_6t
Xbit_r49_c230 bl_230 br_230 wl_49 vdd gnd cell_6t
Xbit_r50_c230 bl_230 br_230 wl_50 vdd gnd cell_6t
Xbit_r51_c230 bl_230 br_230 wl_51 vdd gnd cell_6t
Xbit_r52_c230 bl_230 br_230 wl_52 vdd gnd cell_6t
Xbit_r53_c230 bl_230 br_230 wl_53 vdd gnd cell_6t
Xbit_r54_c230 bl_230 br_230 wl_54 vdd gnd cell_6t
Xbit_r55_c230 bl_230 br_230 wl_55 vdd gnd cell_6t
Xbit_r56_c230 bl_230 br_230 wl_56 vdd gnd cell_6t
Xbit_r57_c230 bl_230 br_230 wl_57 vdd gnd cell_6t
Xbit_r58_c230 bl_230 br_230 wl_58 vdd gnd cell_6t
Xbit_r59_c230 bl_230 br_230 wl_59 vdd gnd cell_6t
Xbit_r60_c230 bl_230 br_230 wl_60 vdd gnd cell_6t
Xbit_r61_c230 bl_230 br_230 wl_61 vdd gnd cell_6t
Xbit_r62_c230 bl_230 br_230 wl_62 vdd gnd cell_6t
Xbit_r63_c230 bl_230 br_230 wl_63 vdd gnd cell_6t
Xbit_r64_c230 bl_230 br_230 wl_64 vdd gnd cell_6t
Xbit_r65_c230 bl_230 br_230 wl_65 vdd gnd cell_6t
Xbit_r66_c230 bl_230 br_230 wl_66 vdd gnd cell_6t
Xbit_r67_c230 bl_230 br_230 wl_67 vdd gnd cell_6t
Xbit_r68_c230 bl_230 br_230 wl_68 vdd gnd cell_6t
Xbit_r69_c230 bl_230 br_230 wl_69 vdd gnd cell_6t
Xbit_r70_c230 bl_230 br_230 wl_70 vdd gnd cell_6t
Xbit_r71_c230 bl_230 br_230 wl_71 vdd gnd cell_6t
Xbit_r72_c230 bl_230 br_230 wl_72 vdd gnd cell_6t
Xbit_r73_c230 bl_230 br_230 wl_73 vdd gnd cell_6t
Xbit_r74_c230 bl_230 br_230 wl_74 vdd gnd cell_6t
Xbit_r75_c230 bl_230 br_230 wl_75 vdd gnd cell_6t
Xbit_r76_c230 bl_230 br_230 wl_76 vdd gnd cell_6t
Xbit_r77_c230 bl_230 br_230 wl_77 vdd gnd cell_6t
Xbit_r78_c230 bl_230 br_230 wl_78 vdd gnd cell_6t
Xbit_r79_c230 bl_230 br_230 wl_79 vdd gnd cell_6t
Xbit_r80_c230 bl_230 br_230 wl_80 vdd gnd cell_6t
Xbit_r81_c230 bl_230 br_230 wl_81 vdd gnd cell_6t
Xbit_r82_c230 bl_230 br_230 wl_82 vdd gnd cell_6t
Xbit_r83_c230 bl_230 br_230 wl_83 vdd gnd cell_6t
Xbit_r84_c230 bl_230 br_230 wl_84 vdd gnd cell_6t
Xbit_r85_c230 bl_230 br_230 wl_85 vdd gnd cell_6t
Xbit_r86_c230 bl_230 br_230 wl_86 vdd gnd cell_6t
Xbit_r87_c230 bl_230 br_230 wl_87 vdd gnd cell_6t
Xbit_r88_c230 bl_230 br_230 wl_88 vdd gnd cell_6t
Xbit_r89_c230 bl_230 br_230 wl_89 vdd gnd cell_6t
Xbit_r90_c230 bl_230 br_230 wl_90 vdd gnd cell_6t
Xbit_r91_c230 bl_230 br_230 wl_91 vdd gnd cell_6t
Xbit_r92_c230 bl_230 br_230 wl_92 vdd gnd cell_6t
Xbit_r93_c230 bl_230 br_230 wl_93 vdd gnd cell_6t
Xbit_r94_c230 bl_230 br_230 wl_94 vdd gnd cell_6t
Xbit_r95_c230 bl_230 br_230 wl_95 vdd gnd cell_6t
Xbit_r96_c230 bl_230 br_230 wl_96 vdd gnd cell_6t
Xbit_r97_c230 bl_230 br_230 wl_97 vdd gnd cell_6t
Xbit_r98_c230 bl_230 br_230 wl_98 vdd gnd cell_6t
Xbit_r99_c230 bl_230 br_230 wl_99 vdd gnd cell_6t
Xbit_r100_c230 bl_230 br_230 wl_100 vdd gnd cell_6t
Xbit_r101_c230 bl_230 br_230 wl_101 vdd gnd cell_6t
Xbit_r102_c230 bl_230 br_230 wl_102 vdd gnd cell_6t
Xbit_r103_c230 bl_230 br_230 wl_103 vdd gnd cell_6t
Xbit_r104_c230 bl_230 br_230 wl_104 vdd gnd cell_6t
Xbit_r105_c230 bl_230 br_230 wl_105 vdd gnd cell_6t
Xbit_r106_c230 bl_230 br_230 wl_106 vdd gnd cell_6t
Xbit_r107_c230 bl_230 br_230 wl_107 vdd gnd cell_6t
Xbit_r108_c230 bl_230 br_230 wl_108 vdd gnd cell_6t
Xbit_r109_c230 bl_230 br_230 wl_109 vdd gnd cell_6t
Xbit_r110_c230 bl_230 br_230 wl_110 vdd gnd cell_6t
Xbit_r111_c230 bl_230 br_230 wl_111 vdd gnd cell_6t
Xbit_r112_c230 bl_230 br_230 wl_112 vdd gnd cell_6t
Xbit_r113_c230 bl_230 br_230 wl_113 vdd gnd cell_6t
Xbit_r114_c230 bl_230 br_230 wl_114 vdd gnd cell_6t
Xbit_r115_c230 bl_230 br_230 wl_115 vdd gnd cell_6t
Xbit_r116_c230 bl_230 br_230 wl_116 vdd gnd cell_6t
Xbit_r117_c230 bl_230 br_230 wl_117 vdd gnd cell_6t
Xbit_r118_c230 bl_230 br_230 wl_118 vdd gnd cell_6t
Xbit_r119_c230 bl_230 br_230 wl_119 vdd gnd cell_6t
Xbit_r120_c230 bl_230 br_230 wl_120 vdd gnd cell_6t
Xbit_r121_c230 bl_230 br_230 wl_121 vdd gnd cell_6t
Xbit_r122_c230 bl_230 br_230 wl_122 vdd gnd cell_6t
Xbit_r123_c230 bl_230 br_230 wl_123 vdd gnd cell_6t
Xbit_r124_c230 bl_230 br_230 wl_124 vdd gnd cell_6t
Xbit_r125_c230 bl_230 br_230 wl_125 vdd gnd cell_6t
Xbit_r126_c230 bl_230 br_230 wl_126 vdd gnd cell_6t
Xbit_r127_c230 bl_230 br_230 wl_127 vdd gnd cell_6t
Xbit_r128_c230 bl_230 br_230 wl_128 vdd gnd cell_6t
Xbit_r129_c230 bl_230 br_230 wl_129 vdd gnd cell_6t
Xbit_r130_c230 bl_230 br_230 wl_130 vdd gnd cell_6t
Xbit_r131_c230 bl_230 br_230 wl_131 vdd gnd cell_6t
Xbit_r132_c230 bl_230 br_230 wl_132 vdd gnd cell_6t
Xbit_r133_c230 bl_230 br_230 wl_133 vdd gnd cell_6t
Xbit_r134_c230 bl_230 br_230 wl_134 vdd gnd cell_6t
Xbit_r135_c230 bl_230 br_230 wl_135 vdd gnd cell_6t
Xbit_r136_c230 bl_230 br_230 wl_136 vdd gnd cell_6t
Xbit_r137_c230 bl_230 br_230 wl_137 vdd gnd cell_6t
Xbit_r138_c230 bl_230 br_230 wl_138 vdd gnd cell_6t
Xbit_r139_c230 bl_230 br_230 wl_139 vdd gnd cell_6t
Xbit_r140_c230 bl_230 br_230 wl_140 vdd gnd cell_6t
Xbit_r141_c230 bl_230 br_230 wl_141 vdd gnd cell_6t
Xbit_r142_c230 bl_230 br_230 wl_142 vdd gnd cell_6t
Xbit_r143_c230 bl_230 br_230 wl_143 vdd gnd cell_6t
Xbit_r144_c230 bl_230 br_230 wl_144 vdd gnd cell_6t
Xbit_r145_c230 bl_230 br_230 wl_145 vdd gnd cell_6t
Xbit_r146_c230 bl_230 br_230 wl_146 vdd gnd cell_6t
Xbit_r147_c230 bl_230 br_230 wl_147 vdd gnd cell_6t
Xbit_r148_c230 bl_230 br_230 wl_148 vdd gnd cell_6t
Xbit_r149_c230 bl_230 br_230 wl_149 vdd gnd cell_6t
Xbit_r150_c230 bl_230 br_230 wl_150 vdd gnd cell_6t
Xbit_r151_c230 bl_230 br_230 wl_151 vdd gnd cell_6t
Xbit_r152_c230 bl_230 br_230 wl_152 vdd gnd cell_6t
Xbit_r153_c230 bl_230 br_230 wl_153 vdd gnd cell_6t
Xbit_r154_c230 bl_230 br_230 wl_154 vdd gnd cell_6t
Xbit_r155_c230 bl_230 br_230 wl_155 vdd gnd cell_6t
Xbit_r156_c230 bl_230 br_230 wl_156 vdd gnd cell_6t
Xbit_r157_c230 bl_230 br_230 wl_157 vdd gnd cell_6t
Xbit_r158_c230 bl_230 br_230 wl_158 vdd gnd cell_6t
Xbit_r159_c230 bl_230 br_230 wl_159 vdd gnd cell_6t
Xbit_r160_c230 bl_230 br_230 wl_160 vdd gnd cell_6t
Xbit_r161_c230 bl_230 br_230 wl_161 vdd gnd cell_6t
Xbit_r162_c230 bl_230 br_230 wl_162 vdd gnd cell_6t
Xbit_r163_c230 bl_230 br_230 wl_163 vdd gnd cell_6t
Xbit_r164_c230 bl_230 br_230 wl_164 vdd gnd cell_6t
Xbit_r165_c230 bl_230 br_230 wl_165 vdd gnd cell_6t
Xbit_r166_c230 bl_230 br_230 wl_166 vdd gnd cell_6t
Xbit_r167_c230 bl_230 br_230 wl_167 vdd gnd cell_6t
Xbit_r168_c230 bl_230 br_230 wl_168 vdd gnd cell_6t
Xbit_r169_c230 bl_230 br_230 wl_169 vdd gnd cell_6t
Xbit_r170_c230 bl_230 br_230 wl_170 vdd gnd cell_6t
Xbit_r171_c230 bl_230 br_230 wl_171 vdd gnd cell_6t
Xbit_r172_c230 bl_230 br_230 wl_172 vdd gnd cell_6t
Xbit_r173_c230 bl_230 br_230 wl_173 vdd gnd cell_6t
Xbit_r174_c230 bl_230 br_230 wl_174 vdd gnd cell_6t
Xbit_r175_c230 bl_230 br_230 wl_175 vdd gnd cell_6t
Xbit_r176_c230 bl_230 br_230 wl_176 vdd gnd cell_6t
Xbit_r177_c230 bl_230 br_230 wl_177 vdd gnd cell_6t
Xbit_r178_c230 bl_230 br_230 wl_178 vdd gnd cell_6t
Xbit_r179_c230 bl_230 br_230 wl_179 vdd gnd cell_6t
Xbit_r180_c230 bl_230 br_230 wl_180 vdd gnd cell_6t
Xbit_r181_c230 bl_230 br_230 wl_181 vdd gnd cell_6t
Xbit_r182_c230 bl_230 br_230 wl_182 vdd gnd cell_6t
Xbit_r183_c230 bl_230 br_230 wl_183 vdd gnd cell_6t
Xbit_r184_c230 bl_230 br_230 wl_184 vdd gnd cell_6t
Xbit_r185_c230 bl_230 br_230 wl_185 vdd gnd cell_6t
Xbit_r186_c230 bl_230 br_230 wl_186 vdd gnd cell_6t
Xbit_r187_c230 bl_230 br_230 wl_187 vdd gnd cell_6t
Xbit_r188_c230 bl_230 br_230 wl_188 vdd gnd cell_6t
Xbit_r189_c230 bl_230 br_230 wl_189 vdd gnd cell_6t
Xbit_r190_c230 bl_230 br_230 wl_190 vdd gnd cell_6t
Xbit_r191_c230 bl_230 br_230 wl_191 vdd gnd cell_6t
Xbit_r192_c230 bl_230 br_230 wl_192 vdd gnd cell_6t
Xbit_r193_c230 bl_230 br_230 wl_193 vdd gnd cell_6t
Xbit_r194_c230 bl_230 br_230 wl_194 vdd gnd cell_6t
Xbit_r195_c230 bl_230 br_230 wl_195 vdd gnd cell_6t
Xbit_r196_c230 bl_230 br_230 wl_196 vdd gnd cell_6t
Xbit_r197_c230 bl_230 br_230 wl_197 vdd gnd cell_6t
Xbit_r198_c230 bl_230 br_230 wl_198 vdd gnd cell_6t
Xbit_r199_c230 bl_230 br_230 wl_199 vdd gnd cell_6t
Xbit_r200_c230 bl_230 br_230 wl_200 vdd gnd cell_6t
Xbit_r201_c230 bl_230 br_230 wl_201 vdd gnd cell_6t
Xbit_r202_c230 bl_230 br_230 wl_202 vdd gnd cell_6t
Xbit_r203_c230 bl_230 br_230 wl_203 vdd gnd cell_6t
Xbit_r204_c230 bl_230 br_230 wl_204 vdd gnd cell_6t
Xbit_r205_c230 bl_230 br_230 wl_205 vdd gnd cell_6t
Xbit_r206_c230 bl_230 br_230 wl_206 vdd gnd cell_6t
Xbit_r207_c230 bl_230 br_230 wl_207 vdd gnd cell_6t
Xbit_r208_c230 bl_230 br_230 wl_208 vdd gnd cell_6t
Xbit_r209_c230 bl_230 br_230 wl_209 vdd gnd cell_6t
Xbit_r210_c230 bl_230 br_230 wl_210 vdd gnd cell_6t
Xbit_r211_c230 bl_230 br_230 wl_211 vdd gnd cell_6t
Xbit_r212_c230 bl_230 br_230 wl_212 vdd gnd cell_6t
Xbit_r213_c230 bl_230 br_230 wl_213 vdd gnd cell_6t
Xbit_r214_c230 bl_230 br_230 wl_214 vdd gnd cell_6t
Xbit_r215_c230 bl_230 br_230 wl_215 vdd gnd cell_6t
Xbit_r216_c230 bl_230 br_230 wl_216 vdd gnd cell_6t
Xbit_r217_c230 bl_230 br_230 wl_217 vdd gnd cell_6t
Xbit_r218_c230 bl_230 br_230 wl_218 vdd gnd cell_6t
Xbit_r219_c230 bl_230 br_230 wl_219 vdd gnd cell_6t
Xbit_r220_c230 bl_230 br_230 wl_220 vdd gnd cell_6t
Xbit_r221_c230 bl_230 br_230 wl_221 vdd gnd cell_6t
Xbit_r222_c230 bl_230 br_230 wl_222 vdd gnd cell_6t
Xbit_r223_c230 bl_230 br_230 wl_223 vdd gnd cell_6t
Xbit_r224_c230 bl_230 br_230 wl_224 vdd gnd cell_6t
Xbit_r225_c230 bl_230 br_230 wl_225 vdd gnd cell_6t
Xbit_r226_c230 bl_230 br_230 wl_226 vdd gnd cell_6t
Xbit_r227_c230 bl_230 br_230 wl_227 vdd gnd cell_6t
Xbit_r228_c230 bl_230 br_230 wl_228 vdd gnd cell_6t
Xbit_r229_c230 bl_230 br_230 wl_229 vdd gnd cell_6t
Xbit_r230_c230 bl_230 br_230 wl_230 vdd gnd cell_6t
Xbit_r231_c230 bl_230 br_230 wl_231 vdd gnd cell_6t
Xbit_r232_c230 bl_230 br_230 wl_232 vdd gnd cell_6t
Xbit_r233_c230 bl_230 br_230 wl_233 vdd gnd cell_6t
Xbit_r234_c230 bl_230 br_230 wl_234 vdd gnd cell_6t
Xbit_r235_c230 bl_230 br_230 wl_235 vdd gnd cell_6t
Xbit_r236_c230 bl_230 br_230 wl_236 vdd gnd cell_6t
Xbit_r237_c230 bl_230 br_230 wl_237 vdd gnd cell_6t
Xbit_r238_c230 bl_230 br_230 wl_238 vdd gnd cell_6t
Xbit_r239_c230 bl_230 br_230 wl_239 vdd gnd cell_6t
Xbit_r240_c230 bl_230 br_230 wl_240 vdd gnd cell_6t
Xbit_r241_c230 bl_230 br_230 wl_241 vdd gnd cell_6t
Xbit_r242_c230 bl_230 br_230 wl_242 vdd gnd cell_6t
Xbit_r243_c230 bl_230 br_230 wl_243 vdd gnd cell_6t
Xbit_r244_c230 bl_230 br_230 wl_244 vdd gnd cell_6t
Xbit_r245_c230 bl_230 br_230 wl_245 vdd gnd cell_6t
Xbit_r246_c230 bl_230 br_230 wl_246 vdd gnd cell_6t
Xbit_r247_c230 bl_230 br_230 wl_247 vdd gnd cell_6t
Xbit_r248_c230 bl_230 br_230 wl_248 vdd gnd cell_6t
Xbit_r249_c230 bl_230 br_230 wl_249 vdd gnd cell_6t
Xbit_r250_c230 bl_230 br_230 wl_250 vdd gnd cell_6t
Xbit_r251_c230 bl_230 br_230 wl_251 vdd gnd cell_6t
Xbit_r252_c230 bl_230 br_230 wl_252 vdd gnd cell_6t
Xbit_r253_c230 bl_230 br_230 wl_253 vdd gnd cell_6t
Xbit_r254_c230 bl_230 br_230 wl_254 vdd gnd cell_6t
Xbit_r255_c230 bl_230 br_230 wl_255 vdd gnd cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd cell_6t
Xbit_r1_c231 bl_231 br_231 wl_1 vdd gnd cell_6t
Xbit_r2_c231 bl_231 br_231 wl_2 vdd gnd cell_6t
Xbit_r3_c231 bl_231 br_231 wl_3 vdd gnd cell_6t
Xbit_r4_c231 bl_231 br_231 wl_4 vdd gnd cell_6t
Xbit_r5_c231 bl_231 br_231 wl_5 vdd gnd cell_6t
Xbit_r6_c231 bl_231 br_231 wl_6 vdd gnd cell_6t
Xbit_r7_c231 bl_231 br_231 wl_7 vdd gnd cell_6t
Xbit_r8_c231 bl_231 br_231 wl_8 vdd gnd cell_6t
Xbit_r9_c231 bl_231 br_231 wl_9 vdd gnd cell_6t
Xbit_r10_c231 bl_231 br_231 wl_10 vdd gnd cell_6t
Xbit_r11_c231 bl_231 br_231 wl_11 vdd gnd cell_6t
Xbit_r12_c231 bl_231 br_231 wl_12 vdd gnd cell_6t
Xbit_r13_c231 bl_231 br_231 wl_13 vdd gnd cell_6t
Xbit_r14_c231 bl_231 br_231 wl_14 vdd gnd cell_6t
Xbit_r15_c231 bl_231 br_231 wl_15 vdd gnd cell_6t
Xbit_r16_c231 bl_231 br_231 wl_16 vdd gnd cell_6t
Xbit_r17_c231 bl_231 br_231 wl_17 vdd gnd cell_6t
Xbit_r18_c231 bl_231 br_231 wl_18 vdd gnd cell_6t
Xbit_r19_c231 bl_231 br_231 wl_19 vdd gnd cell_6t
Xbit_r20_c231 bl_231 br_231 wl_20 vdd gnd cell_6t
Xbit_r21_c231 bl_231 br_231 wl_21 vdd gnd cell_6t
Xbit_r22_c231 bl_231 br_231 wl_22 vdd gnd cell_6t
Xbit_r23_c231 bl_231 br_231 wl_23 vdd gnd cell_6t
Xbit_r24_c231 bl_231 br_231 wl_24 vdd gnd cell_6t
Xbit_r25_c231 bl_231 br_231 wl_25 vdd gnd cell_6t
Xbit_r26_c231 bl_231 br_231 wl_26 vdd gnd cell_6t
Xbit_r27_c231 bl_231 br_231 wl_27 vdd gnd cell_6t
Xbit_r28_c231 bl_231 br_231 wl_28 vdd gnd cell_6t
Xbit_r29_c231 bl_231 br_231 wl_29 vdd gnd cell_6t
Xbit_r30_c231 bl_231 br_231 wl_30 vdd gnd cell_6t
Xbit_r31_c231 bl_231 br_231 wl_31 vdd gnd cell_6t
Xbit_r32_c231 bl_231 br_231 wl_32 vdd gnd cell_6t
Xbit_r33_c231 bl_231 br_231 wl_33 vdd gnd cell_6t
Xbit_r34_c231 bl_231 br_231 wl_34 vdd gnd cell_6t
Xbit_r35_c231 bl_231 br_231 wl_35 vdd gnd cell_6t
Xbit_r36_c231 bl_231 br_231 wl_36 vdd gnd cell_6t
Xbit_r37_c231 bl_231 br_231 wl_37 vdd gnd cell_6t
Xbit_r38_c231 bl_231 br_231 wl_38 vdd gnd cell_6t
Xbit_r39_c231 bl_231 br_231 wl_39 vdd gnd cell_6t
Xbit_r40_c231 bl_231 br_231 wl_40 vdd gnd cell_6t
Xbit_r41_c231 bl_231 br_231 wl_41 vdd gnd cell_6t
Xbit_r42_c231 bl_231 br_231 wl_42 vdd gnd cell_6t
Xbit_r43_c231 bl_231 br_231 wl_43 vdd gnd cell_6t
Xbit_r44_c231 bl_231 br_231 wl_44 vdd gnd cell_6t
Xbit_r45_c231 bl_231 br_231 wl_45 vdd gnd cell_6t
Xbit_r46_c231 bl_231 br_231 wl_46 vdd gnd cell_6t
Xbit_r47_c231 bl_231 br_231 wl_47 vdd gnd cell_6t
Xbit_r48_c231 bl_231 br_231 wl_48 vdd gnd cell_6t
Xbit_r49_c231 bl_231 br_231 wl_49 vdd gnd cell_6t
Xbit_r50_c231 bl_231 br_231 wl_50 vdd gnd cell_6t
Xbit_r51_c231 bl_231 br_231 wl_51 vdd gnd cell_6t
Xbit_r52_c231 bl_231 br_231 wl_52 vdd gnd cell_6t
Xbit_r53_c231 bl_231 br_231 wl_53 vdd gnd cell_6t
Xbit_r54_c231 bl_231 br_231 wl_54 vdd gnd cell_6t
Xbit_r55_c231 bl_231 br_231 wl_55 vdd gnd cell_6t
Xbit_r56_c231 bl_231 br_231 wl_56 vdd gnd cell_6t
Xbit_r57_c231 bl_231 br_231 wl_57 vdd gnd cell_6t
Xbit_r58_c231 bl_231 br_231 wl_58 vdd gnd cell_6t
Xbit_r59_c231 bl_231 br_231 wl_59 vdd gnd cell_6t
Xbit_r60_c231 bl_231 br_231 wl_60 vdd gnd cell_6t
Xbit_r61_c231 bl_231 br_231 wl_61 vdd gnd cell_6t
Xbit_r62_c231 bl_231 br_231 wl_62 vdd gnd cell_6t
Xbit_r63_c231 bl_231 br_231 wl_63 vdd gnd cell_6t
Xbit_r64_c231 bl_231 br_231 wl_64 vdd gnd cell_6t
Xbit_r65_c231 bl_231 br_231 wl_65 vdd gnd cell_6t
Xbit_r66_c231 bl_231 br_231 wl_66 vdd gnd cell_6t
Xbit_r67_c231 bl_231 br_231 wl_67 vdd gnd cell_6t
Xbit_r68_c231 bl_231 br_231 wl_68 vdd gnd cell_6t
Xbit_r69_c231 bl_231 br_231 wl_69 vdd gnd cell_6t
Xbit_r70_c231 bl_231 br_231 wl_70 vdd gnd cell_6t
Xbit_r71_c231 bl_231 br_231 wl_71 vdd gnd cell_6t
Xbit_r72_c231 bl_231 br_231 wl_72 vdd gnd cell_6t
Xbit_r73_c231 bl_231 br_231 wl_73 vdd gnd cell_6t
Xbit_r74_c231 bl_231 br_231 wl_74 vdd gnd cell_6t
Xbit_r75_c231 bl_231 br_231 wl_75 vdd gnd cell_6t
Xbit_r76_c231 bl_231 br_231 wl_76 vdd gnd cell_6t
Xbit_r77_c231 bl_231 br_231 wl_77 vdd gnd cell_6t
Xbit_r78_c231 bl_231 br_231 wl_78 vdd gnd cell_6t
Xbit_r79_c231 bl_231 br_231 wl_79 vdd gnd cell_6t
Xbit_r80_c231 bl_231 br_231 wl_80 vdd gnd cell_6t
Xbit_r81_c231 bl_231 br_231 wl_81 vdd gnd cell_6t
Xbit_r82_c231 bl_231 br_231 wl_82 vdd gnd cell_6t
Xbit_r83_c231 bl_231 br_231 wl_83 vdd gnd cell_6t
Xbit_r84_c231 bl_231 br_231 wl_84 vdd gnd cell_6t
Xbit_r85_c231 bl_231 br_231 wl_85 vdd gnd cell_6t
Xbit_r86_c231 bl_231 br_231 wl_86 vdd gnd cell_6t
Xbit_r87_c231 bl_231 br_231 wl_87 vdd gnd cell_6t
Xbit_r88_c231 bl_231 br_231 wl_88 vdd gnd cell_6t
Xbit_r89_c231 bl_231 br_231 wl_89 vdd gnd cell_6t
Xbit_r90_c231 bl_231 br_231 wl_90 vdd gnd cell_6t
Xbit_r91_c231 bl_231 br_231 wl_91 vdd gnd cell_6t
Xbit_r92_c231 bl_231 br_231 wl_92 vdd gnd cell_6t
Xbit_r93_c231 bl_231 br_231 wl_93 vdd gnd cell_6t
Xbit_r94_c231 bl_231 br_231 wl_94 vdd gnd cell_6t
Xbit_r95_c231 bl_231 br_231 wl_95 vdd gnd cell_6t
Xbit_r96_c231 bl_231 br_231 wl_96 vdd gnd cell_6t
Xbit_r97_c231 bl_231 br_231 wl_97 vdd gnd cell_6t
Xbit_r98_c231 bl_231 br_231 wl_98 vdd gnd cell_6t
Xbit_r99_c231 bl_231 br_231 wl_99 vdd gnd cell_6t
Xbit_r100_c231 bl_231 br_231 wl_100 vdd gnd cell_6t
Xbit_r101_c231 bl_231 br_231 wl_101 vdd gnd cell_6t
Xbit_r102_c231 bl_231 br_231 wl_102 vdd gnd cell_6t
Xbit_r103_c231 bl_231 br_231 wl_103 vdd gnd cell_6t
Xbit_r104_c231 bl_231 br_231 wl_104 vdd gnd cell_6t
Xbit_r105_c231 bl_231 br_231 wl_105 vdd gnd cell_6t
Xbit_r106_c231 bl_231 br_231 wl_106 vdd gnd cell_6t
Xbit_r107_c231 bl_231 br_231 wl_107 vdd gnd cell_6t
Xbit_r108_c231 bl_231 br_231 wl_108 vdd gnd cell_6t
Xbit_r109_c231 bl_231 br_231 wl_109 vdd gnd cell_6t
Xbit_r110_c231 bl_231 br_231 wl_110 vdd gnd cell_6t
Xbit_r111_c231 bl_231 br_231 wl_111 vdd gnd cell_6t
Xbit_r112_c231 bl_231 br_231 wl_112 vdd gnd cell_6t
Xbit_r113_c231 bl_231 br_231 wl_113 vdd gnd cell_6t
Xbit_r114_c231 bl_231 br_231 wl_114 vdd gnd cell_6t
Xbit_r115_c231 bl_231 br_231 wl_115 vdd gnd cell_6t
Xbit_r116_c231 bl_231 br_231 wl_116 vdd gnd cell_6t
Xbit_r117_c231 bl_231 br_231 wl_117 vdd gnd cell_6t
Xbit_r118_c231 bl_231 br_231 wl_118 vdd gnd cell_6t
Xbit_r119_c231 bl_231 br_231 wl_119 vdd gnd cell_6t
Xbit_r120_c231 bl_231 br_231 wl_120 vdd gnd cell_6t
Xbit_r121_c231 bl_231 br_231 wl_121 vdd gnd cell_6t
Xbit_r122_c231 bl_231 br_231 wl_122 vdd gnd cell_6t
Xbit_r123_c231 bl_231 br_231 wl_123 vdd gnd cell_6t
Xbit_r124_c231 bl_231 br_231 wl_124 vdd gnd cell_6t
Xbit_r125_c231 bl_231 br_231 wl_125 vdd gnd cell_6t
Xbit_r126_c231 bl_231 br_231 wl_126 vdd gnd cell_6t
Xbit_r127_c231 bl_231 br_231 wl_127 vdd gnd cell_6t
Xbit_r128_c231 bl_231 br_231 wl_128 vdd gnd cell_6t
Xbit_r129_c231 bl_231 br_231 wl_129 vdd gnd cell_6t
Xbit_r130_c231 bl_231 br_231 wl_130 vdd gnd cell_6t
Xbit_r131_c231 bl_231 br_231 wl_131 vdd gnd cell_6t
Xbit_r132_c231 bl_231 br_231 wl_132 vdd gnd cell_6t
Xbit_r133_c231 bl_231 br_231 wl_133 vdd gnd cell_6t
Xbit_r134_c231 bl_231 br_231 wl_134 vdd gnd cell_6t
Xbit_r135_c231 bl_231 br_231 wl_135 vdd gnd cell_6t
Xbit_r136_c231 bl_231 br_231 wl_136 vdd gnd cell_6t
Xbit_r137_c231 bl_231 br_231 wl_137 vdd gnd cell_6t
Xbit_r138_c231 bl_231 br_231 wl_138 vdd gnd cell_6t
Xbit_r139_c231 bl_231 br_231 wl_139 vdd gnd cell_6t
Xbit_r140_c231 bl_231 br_231 wl_140 vdd gnd cell_6t
Xbit_r141_c231 bl_231 br_231 wl_141 vdd gnd cell_6t
Xbit_r142_c231 bl_231 br_231 wl_142 vdd gnd cell_6t
Xbit_r143_c231 bl_231 br_231 wl_143 vdd gnd cell_6t
Xbit_r144_c231 bl_231 br_231 wl_144 vdd gnd cell_6t
Xbit_r145_c231 bl_231 br_231 wl_145 vdd gnd cell_6t
Xbit_r146_c231 bl_231 br_231 wl_146 vdd gnd cell_6t
Xbit_r147_c231 bl_231 br_231 wl_147 vdd gnd cell_6t
Xbit_r148_c231 bl_231 br_231 wl_148 vdd gnd cell_6t
Xbit_r149_c231 bl_231 br_231 wl_149 vdd gnd cell_6t
Xbit_r150_c231 bl_231 br_231 wl_150 vdd gnd cell_6t
Xbit_r151_c231 bl_231 br_231 wl_151 vdd gnd cell_6t
Xbit_r152_c231 bl_231 br_231 wl_152 vdd gnd cell_6t
Xbit_r153_c231 bl_231 br_231 wl_153 vdd gnd cell_6t
Xbit_r154_c231 bl_231 br_231 wl_154 vdd gnd cell_6t
Xbit_r155_c231 bl_231 br_231 wl_155 vdd gnd cell_6t
Xbit_r156_c231 bl_231 br_231 wl_156 vdd gnd cell_6t
Xbit_r157_c231 bl_231 br_231 wl_157 vdd gnd cell_6t
Xbit_r158_c231 bl_231 br_231 wl_158 vdd gnd cell_6t
Xbit_r159_c231 bl_231 br_231 wl_159 vdd gnd cell_6t
Xbit_r160_c231 bl_231 br_231 wl_160 vdd gnd cell_6t
Xbit_r161_c231 bl_231 br_231 wl_161 vdd gnd cell_6t
Xbit_r162_c231 bl_231 br_231 wl_162 vdd gnd cell_6t
Xbit_r163_c231 bl_231 br_231 wl_163 vdd gnd cell_6t
Xbit_r164_c231 bl_231 br_231 wl_164 vdd gnd cell_6t
Xbit_r165_c231 bl_231 br_231 wl_165 vdd gnd cell_6t
Xbit_r166_c231 bl_231 br_231 wl_166 vdd gnd cell_6t
Xbit_r167_c231 bl_231 br_231 wl_167 vdd gnd cell_6t
Xbit_r168_c231 bl_231 br_231 wl_168 vdd gnd cell_6t
Xbit_r169_c231 bl_231 br_231 wl_169 vdd gnd cell_6t
Xbit_r170_c231 bl_231 br_231 wl_170 vdd gnd cell_6t
Xbit_r171_c231 bl_231 br_231 wl_171 vdd gnd cell_6t
Xbit_r172_c231 bl_231 br_231 wl_172 vdd gnd cell_6t
Xbit_r173_c231 bl_231 br_231 wl_173 vdd gnd cell_6t
Xbit_r174_c231 bl_231 br_231 wl_174 vdd gnd cell_6t
Xbit_r175_c231 bl_231 br_231 wl_175 vdd gnd cell_6t
Xbit_r176_c231 bl_231 br_231 wl_176 vdd gnd cell_6t
Xbit_r177_c231 bl_231 br_231 wl_177 vdd gnd cell_6t
Xbit_r178_c231 bl_231 br_231 wl_178 vdd gnd cell_6t
Xbit_r179_c231 bl_231 br_231 wl_179 vdd gnd cell_6t
Xbit_r180_c231 bl_231 br_231 wl_180 vdd gnd cell_6t
Xbit_r181_c231 bl_231 br_231 wl_181 vdd gnd cell_6t
Xbit_r182_c231 bl_231 br_231 wl_182 vdd gnd cell_6t
Xbit_r183_c231 bl_231 br_231 wl_183 vdd gnd cell_6t
Xbit_r184_c231 bl_231 br_231 wl_184 vdd gnd cell_6t
Xbit_r185_c231 bl_231 br_231 wl_185 vdd gnd cell_6t
Xbit_r186_c231 bl_231 br_231 wl_186 vdd gnd cell_6t
Xbit_r187_c231 bl_231 br_231 wl_187 vdd gnd cell_6t
Xbit_r188_c231 bl_231 br_231 wl_188 vdd gnd cell_6t
Xbit_r189_c231 bl_231 br_231 wl_189 vdd gnd cell_6t
Xbit_r190_c231 bl_231 br_231 wl_190 vdd gnd cell_6t
Xbit_r191_c231 bl_231 br_231 wl_191 vdd gnd cell_6t
Xbit_r192_c231 bl_231 br_231 wl_192 vdd gnd cell_6t
Xbit_r193_c231 bl_231 br_231 wl_193 vdd gnd cell_6t
Xbit_r194_c231 bl_231 br_231 wl_194 vdd gnd cell_6t
Xbit_r195_c231 bl_231 br_231 wl_195 vdd gnd cell_6t
Xbit_r196_c231 bl_231 br_231 wl_196 vdd gnd cell_6t
Xbit_r197_c231 bl_231 br_231 wl_197 vdd gnd cell_6t
Xbit_r198_c231 bl_231 br_231 wl_198 vdd gnd cell_6t
Xbit_r199_c231 bl_231 br_231 wl_199 vdd gnd cell_6t
Xbit_r200_c231 bl_231 br_231 wl_200 vdd gnd cell_6t
Xbit_r201_c231 bl_231 br_231 wl_201 vdd gnd cell_6t
Xbit_r202_c231 bl_231 br_231 wl_202 vdd gnd cell_6t
Xbit_r203_c231 bl_231 br_231 wl_203 vdd gnd cell_6t
Xbit_r204_c231 bl_231 br_231 wl_204 vdd gnd cell_6t
Xbit_r205_c231 bl_231 br_231 wl_205 vdd gnd cell_6t
Xbit_r206_c231 bl_231 br_231 wl_206 vdd gnd cell_6t
Xbit_r207_c231 bl_231 br_231 wl_207 vdd gnd cell_6t
Xbit_r208_c231 bl_231 br_231 wl_208 vdd gnd cell_6t
Xbit_r209_c231 bl_231 br_231 wl_209 vdd gnd cell_6t
Xbit_r210_c231 bl_231 br_231 wl_210 vdd gnd cell_6t
Xbit_r211_c231 bl_231 br_231 wl_211 vdd gnd cell_6t
Xbit_r212_c231 bl_231 br_231 wl_212 vdd gnd cell_6t
Xbit_r213_c231 bl_231 br_231 wl_213 vdd gnd cell_6t
Xbit_r214_c231 bl_231 br_231 wl_214 vdd gnd cell_6t
Xbit_r215_c231 bl_231 br_231 wl_215 vdd gnd cell_6t
Xbit_r216_c231 bl_231 br_231 wl_216 vdd gnd cell_6t
Xbit_r217_c231 bl_231 br_231 wl_217 vdd gnd cell_6t
Xbit_r218_c231 bl_231 br_231 wl_218 vdd gnd cell_6t
Xbit_r219_c231 bl_231 br_231 wl_219 vdd gnd cell_6t
Xbit_r220_c231 bl_231 br_231 wl_220 vdd gnd cell_6t
Xbit_r221_c231 bl_231 br_231 wl_221 vdd gnd cell_6t
Xbit_r222_c231 bl_231 br_231 wl_222 vdd gnd cell_6t
Xbit_r223_c231 bl_231 br_231 wl_223 vdd gnd cell_6t
Xbit_r224_c231 bl_231 br_231 wl_224 vdd gnd cell_6t
Xbit_r225_c231 bl_231 br_231 wl_225 vdd gnd cell_6t
Xbit_r226_c231 bl_231 br_231 wl_226 vdd gnd cell_6t
Xbit_r227_c231 bl_231 br_231 wl_227 vdd gnd cell_6t
Xbit_r228_c231 bl_231 br_231 wl_228 vdd gnd cell_6t
Xbit_r229_c231 bl_231 br_231 wl_229 vdd gnd cell_6t
Xbit_r230_c231 bl_231 br_231 wl_230 vdd gnd cell_6t
Xbit_r231_c231 bl_231 br_231 wl_231 vdd gnd cell_6t
Xbit_r232_c231 bl_231 br_231 wl_232 vdd gnd cell_6t
Xbit_r233_c231 bl_231 br_231 wl_233 vdd gnd cell_6t
Xbit_r234_c231 bl_231 br_231 wl_234 vdd gnd cell_6t
Xbit_r235_c231 bl_231 br_231 wl_235 vdd gnd cell_6t
Xbit_r236_c231 bl_231 br_231 wl_236 vdd gnd cell_6t
Xbit_r237_c231 bl_231 br_231 wl_237 vdd gnd cell_6t
Xbit_r238_c231 bl_231 br_231 wl_238 vdd gnd cell_6t
Xbit_r239_c231 bl_231 br_231 wl_239 vdd gnd cell_6t
Xbit_r240_c231 bl_231 br_231 wl_240 vdd gnd cell_6t
Xbit_r241_c231 bl_231 br_231 wl_241 vdd gnd cell_6t
Xbit_r242_c231 bl_231 br_231 wl_242 vdd gnd cell_6t
Xbit_r243_c231 bl_231 br_231 wl_243 vdd gnd cell_6t
Xbit_r244_c231 bl_231 br_231 wl_244 vdd gnd cell_6t
Xbit_r245_c231 bl_231 br_231 wl_245 vdd gnd cell_6t
Xbit_r246_c231 bl_231 br_231 wl_246 vdd gnd cell_6t
Xbit_r247_c231 bl_231 br_231 wl_247 vdd gnd cell_6t
Xbit_r248_c231 bl_231 br_231 wl_248 vdd gnd cell_6t
Xbit_r249_c231 bl_231 br_231 wl_249 vdd gnd cell_6t
Xbit_r250_c231 bl_231 br_231 wl_250 vdd gnd cell_6t
Xbit_r251_c231 bl_231 br_231 wl_251 vdd gnd cell_6t
Xbit_r252_c231 bl_231 br_231 wl_252 vdd gnd cell_6t
Xbit_r253_c231 bl_231 br_231 wl_253 vdd gnd cell_6t
Xbit_r254_c231 bl_231 br_231 wl_254 vdd gnd cell_6t
Xbit_r255_c231 bl_231 br_231 wl_255 vdd gnd cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd cell_6t
Xbit_r1_c232 bl_232 br_232 wl_1 vdd gnd cell_6t
Xbit_r2_c232 bl_232 br_232 wl_2 vdd gnd cell_6t
Xbit_r3_c232 bl_232 br_232 wl_3 vdd gnd cell_6t
Xbit_r4_c232 bl_232 br_232 wl_4 vdd gnd cell_6t
Xbit_r5_c232 bl_232 br_232 wl_5 vdd gnd cell_6t
Xbit_r6_c232 bl_232 br_232 wl_6 vdd gnd cell_6t
Xbit_r7_c232 bl_232 br_232 wl_7 vdd gnd cell_6t
Xbit_r8_c232 bl_232 br_232 wl_8 vdd gnd cell_6t
Xbit_r9_c232 bl_232 br_232 wl_9 vdd gnd cell_6t
Xbit_r10_c232 bl_232 br_232 wl_10 vdd gnd cell_6t
Xbit_r11_c232 bl_232 br_232 wl_11 vdd gnd cell_6t
Xbit_r12_c232 bl_232 br_232 wl_12 vdd gnd cell_6t
Xbit_r13_c232 bl_232 br_232 wl_13 vdd gnd cell_6t
Xbit_r14_c232 bl_232 br_232 wl_14 vdd gnd cell_6t
Xbit_r15_c232 bl_232 br_232 wl_15 vdd gnd cell_6t
Xbit_r16_c232 bl_232 br_232 wl_16 vdd gnd cell_6t
Xbit_r17_c232 bl_232 br_232 wl_17 vdd gnd cell_6t
Xbit_r18_c232 bl_232 br_232 wl_18 vdd gnd cell_6t
Xbit_r19_c232 bl_232 br_232 wl_19 vdd gnd cell_6t
Xbit_r20_c232 bl_232 br_232 wl_20 vdd gnd cell_6t
Xbit_r21_c232 bl_232 br_232 wl_21 vdd gnd cell_6t
Xbit_r22_c232 bl_232 br_232 wl_22 vdd gnd cell_6t
Xbit_r23_c232 bl_232 br_232 wl_23 vdd gnd cell_6t
Xbit_r24_c232 bl_232 br_232 wl_24 vdd gnd cell_6t
Xbit_r25_c232 bl_232 br_232 wl_25 vdd gnd cell_6t
Xbit_r26_c232 bl_232 br_232 wl_26 vdd gnd cell_6t
Xbit_r27_c232 bl_232 br_232 wl_27 vdd gnd cell_6t
Xbit_r28_c232 bl_232 br_232 wl_28 vdd gnd cell_6t
Xbit_r29_c232 bl_232 br_232 wl_29 vdd gnd cell_6t
Xbit_r30_c232 bl_232 br_232 wl_30 vdd gnd cell_6t
Xbit_r31_c232 bl_232 br_232 wl_31 vdd gnd cell_6t
Xbit_r32_c232 bl_232 br_232 wl_32 vdd gnd cell_6t
Xbit_r33_c232 bl_232 br_232 wl_33 vdd gnd cell_6t
Xbit_r34_c232 bl_232 br_232 wl_34 vdd gnd cell_6t
Xbit_r35_c232 bl_232 br_232 wl_35 vdd gnd cell_6t
Xbit_r36_c232 bl_232 br_232 wl_36 vdd gnd cell_6t
Xbit_r37_c232 bl_232 br_232 wl_37 vdd gnd cell_6t
Xbit_r38_c232 bl_232 br_232 wl_38 vdd gnd cell_6t
Xbit_r39_c232 bl_232 br_232 wl_39 vdd gnd cell_6t
Xbit_r40_c232 bl_232 br_232 wl_40 vdd gnd cell_6t
Xbit_r41_c232 bl_232 br_232 wl_41 vdd gnd cell_6t
Xbit_r42_c232 bl_232 br_232 wl_42 vdd gnd cell_6t
Xbit_r43_c232 bl_232 br_232 wl_43 vdd gnd cell_6t
Xbit_r44_c232 bl_232 br_232 wl_44 vdd gnd cell_6t
Xbit_r45_c232 bl_232 br_232 wl_45 vdd gnd cell_6t
Xbit_r46_c232 bl_232 br_232 wl_46 vdd gnd cell_6t
Xbit_r47_c232 bl_232 br_232 wl_47 vdd gnd cell_6t
Xbit_r48_c232 bl_232 br_232 wl_48 vdd gnd cell_6t
Xbit_r49_c232 bl_232 br_232 wl_49 vdd gnd cell_6t
Xbit_r50_c232 bl_232 br_232 wl_50 vdd gnd cell_6t
Xbit_r51_c232 bl_232 br_232 wl_51 vdd gnd cell_6t
Xbit_r52_c232 bl_232 br_232 wl_52 vdd gnd cell_6t
Xbit_r53_c232 bl_232 br_232 wl_53 vdd gnd cell_6t
Xbit_r54_c232 bl_232 br_232 wl_54 vdd gnd cell_6t
Xbit_r55_c232 bl_232 br_232 wl_55 vdd gnd cell_6t
Xbit_r56_c232 bl_232 br_232 wl_56 vdd gnd cell_6t
Xbit_r57_c232 bl_232 br_232 wl_57 vdd gnd cell_6t
Xbit_r58_c232 bl_232 br_232 wl_58 vdd gnd cell_6t
Xbit_r59_c232 bl_232 br_232 wl_59 vdd gnd cell_6t
Xbit_r60_c232 bl_232 br_232 wl_60 vdd gnd cell_6t
Xbit_r61_c232 bl_232 br_232 wl_61 vdd gnd cell_6t
Xbit_r62_c232 bl_232 br_232 wl_62 vdd gnd cell_6t
Xbit_r63_c232 bl_232 br_232 wl_63 vdd gnd cell_6t
Xbit_r64_c232 bl_232 br_232 wl_64 vdd gnd cell_6t
Xbit_r65_c232 bl_232 br_232 wl_65 vdd gnd cell_6t
Xbit_r66_c232 bl_232 br_232 wl_66 vdd gnd cell_6t
Xbit_r67_c232 bl_232 br_232 wl_67 vdd gnd cell_6t
Xbit_r68_c232 bl_232 br_232 wl_68 vdd gnd cell_6t
Xbit_r69_c232 bl_232 br_232 wl_69 vdd gnd cell_6t
Xbit_r70_c232 bl_232 br_232 wl_70 vdd gnd cell_6t
Xbit_r71_c232 bl_232 br_232 wl_71 vdd gnd cell_6t
Xbit_r72_c232 bl_232 br_232 wl_72 vdd gnd cell_6t
Xbit_r73_c232 bl_232 br_232 wl_73 vdd gnd cell_6t
Xbit_r74_c232 bl_232 br_232 wl_74 vdd gnd cell_6t
Xbit_r75_c232 bl_232 br_232 wl_75 vdd gnd cell_6t
Xbit_r76_c232 bl_232 br_232 wl_76 vdd gnd cell_6t
Xbit_r77_c232 bl_232 br_232 wl_77 vdd gnd cell_6t
Xbit_r78_c232 bl_232 br_232 wl_78 vdd gnd cell_6t
Xbit_r79_c232 bl_232 br_232 wl_79 vdd gnd cell_6t
Xbit_r80_c232 bl_232 br_232 wl_80 vdd gnd cell_6t
Xbit_r81_c232 bl_232 br_232 wl_81 vdd gnd cell_6t
Xbit_r82_c232 bl_232 br_232 wl_82 vdd gnd cell_6t
Xbit_r83_c232 bl_232 br_232 wl_83 vdd gnd cell_6t
Xbit_r84_c232 bl_232 br_232 wl_84 vdd gnd cell_6t
Xbit_r85_c232 bl_232 br_232 wl_85 vdd gnd cell_6t
Xbit_r86_c232 bl_232 br_232 wl_86 vdd gnd cell_6t
Xbit_r87_c232 bl_232 br_232 wl_87 vdd gnd cell_6t
Xbit_r88_c232 bl_232 br_232 wl_88 vdd gnd cell_6t
Xbit_r89_c232 bl_232 br_232 wl_89 vdd gnd cell_6t
Xbit_r90_c232 bl_232 br_232 wl_90 vdd gnd cell_6t
Xbit_r91_c232 bl_232 br_232 wl_91 vdd gnd cell_6t
Xbit_r92_c232 bl_232 br_232 wl_92 vdd gnd cell_6t
Xbit_r93_c232 bl_232 br_232 wl_93 vdd gnd cell_6t
Xbit_r94_c232 bl_232 br_232 wl_94 vdd gnd cell_6t
Xbit_r95_c232 bl_232 br_232 wl_95 vdd gnd cell_6t
Xbit_r96_c232 bl_232 br_232 wl_96 vdd gnd cell_6t
Xbit_r97_c232 bl_232 br_232 wl_97 vdd gnd cell_6t
Xbit_r98_c232 bl_232 br_232 wl_98 vdd gnd cell_6t
Xbit_r99_c232 bl_232 br_232 wl_99 vdd gnd cell_6t
Xbit_r100_c232 bl_232 br_232 wl_100 vdd gnd cell_6t
Xbit_r101_c232 bl_232 br_232 wl_101 vdd gnd cell_6t
Xbit_r102_c232 bl_232 br_232 wl_102 vdd gnd cell_6t
Xbit_r103_c232 bl_232 br_232 wl_103 vdd gnd cell_6t
Xbit_r104_c232 bl_232 br_232 wl_104 vdd gnd cell_6t
Xbit_r105_c232 bl_232 br_232 wl_105 vdd gnd cell_6t
Xbit_r106_c232 bl_232 br_232 wl_106 vdd gnd cell_6t
Xbit_r107_c232 bl_232 br_232 wl_107 vdd gnd cell_6t
Xbit_r108_c232 bl_232 br_232 wl_108 vdd gnd cell_6t
Xbit_r109_c232 bl_232 br_232 wl_109 vdd gnd cell_6t
Xbit_r110_c232 bl_232 br_232 wl_110 vdd gnd cell_6t
Xbit_r111_c232 bl_232 br_232 wl_111 vdd gnd cell_6t
Xbit_r112_c232 bl_232 br_232 wl_112 vdd gnd cell_6t
Xbit_r113_c232 bl_232 br_232 wl_113 vdd gnd cell_6t
Xbit_r114_c232 bl_232 br_232 wl_114 vdd gnd cell_6t
Xbit_r115_c232 bl_232 br_232 wl_115 vdd gnd cell_6t
Xbit_r116_c232 bl_232 br_232 wl_116 vdd gnd cell_6t
Xbit_r117_c232 bl_232 br_232 wl_117 vdd gnd cell_6t
Xbit_r118_c232 bl_232 br_232 wl_118 vdd gnd cell_6t
Xbit_r119_c232 bl_232 br_232 wl_119 vdd gnd cell_6t
Xbit_r120_c232 bl_232 br_232 wl_120 vdd gnd cell_6t
Xbit_r121_c232 bl_232 br_232 wl_121 vdd gnd cell_6t
Xbit_r122_c232 bl_232 br_232 wl_122 vdd gnd cell_6t
Xbit_r123_c232 bl_232 br_232 wl_123 vdd gnd cell_6t
Xbit_r124_c232 bl_232 br_232 wl_124 vdd gnd cell_6t
Xbit_r125_c232 bl_232 br_232 wl_125 vdd gnd cell_6t
Xbit_r126_c232 bl_232 br_232 wl_126 vdd gnd cell_6t
Xbit_r127_c232 bl_232 br_232 wl_127 vdd gnd cell_6t
Xbit_r128_c232 bl_232 br_232 wl_128 vdd gnd cell_6t
Xbit_r129_c232 bl_232 br_232 wl_129 vdd gnd cell_6t
Xbit_r130_c232 bl_232 br_232 wl_130 vdd gnd cell_6t
Xbit_r131_c232 bl_232 br_232 wl_131 vdd gnd cell_6t
Xbit_r132_c232 bl_232 br_232 wl_132 vdd gnd cell_6t
Xbit_r133_c232 bl_232 br_232 wl_133 vdd gnd cell_6t
Xbit_r134_c232 bl_232 br_232 wl_134 vdd gnd cell_6t
Xbit_r135_c232 bl_232 br_232 wl_135 vdd gnd cell_6t
Xbit_r136_c232 bl_232 br_232 wl_136 vdd gnd cell_6t
Xbit_r137_c232 bl_232 br_232 wl_137 vdd gnd cell_6t
Xbit_r138_c232 bl_232 br_232 wl_138 vdd gnd cell_6t
Xbit_r139_c232 bl_232 br_232 wl_139 vdd gnd cell_6t
Xbit_r140_c232 bl_232 br_232 wl_140 vdd gnd cell_6t
Xbit_r141_c232 bl_232 br_232 wl_141 vdd gnd cell_6t
Xbit_r142_c232 bl_232 br_232 wl_142 vdd gnd cell_6t
Xbit_r143_c232 bl_232 br_232 wl_143 vdd gnd cell_6t
Xbit_r144_c232 bl_232 br_232 wl_144 vdd gnd cell_6t
Xbit_r145_c232 bl_232 br_232 wl_145 vdd gnd cell_6t
Xbit_r146_c232 bl_232 br_232 wl_146 vdd gnd cell_6t
Xbit_r147_c232 bl_232 br_232 wl_147 vdd gnd cell_6t
Xbit_r148_c232 bl_232 br_232 wl_148 vdd gnd cell_6t
Xbit_r149_c232 bl_232 br_232 wl_149 vdd gnd cell_6t
Xbit_r150_c232 bl_232 br_232 wl_150 vdd gnd cell_6t
Xbit_r151_c232 bl_232 br_232 wl_151 vdd gnd cell_6t
Xbit_r152_c232 bl_232 br_232 wl_152 vdd gnd cell_6t
Xbit_r153_c232 bl_232 br_232 wl_153 vdd gnd cell_6t
Xbit_r154_c232 bl_232 br_232 wl_154 vdd gnd cell_6t
Xbit_r155_c232 bl_232 br_232 wl_155 vdd gnd cell_6t
Xbit_r156_c232 bl_232 br_232 wl_156 vdd gnd cell_6t
Xbit_r157_c232 bl_232 br_232 wl_157 vdd gnd cell_6t
Xbit_r158_c232 bl_232 br_232 wl_158 vdd gnd cell_6t
Xbit_r159_c232 bl_232 br_232 wl_159 vdd gnd cell_6t
Xbit_r160_c232 bl_232 br_232 wl_160 vdd gnd cell_6t
Xbit_r161_c232 bl_232 br_232 wl_161 vdd gnd cell_6t
Xbit_r162_c232 bl_232 br_232 wl_162 vdd gnd cell_6t
Xbit_r163_c232 bl_232 br_232 wl_163 vdd gnd cell_6t
Xbit_r164_c232 bl_232 br_232 wl_164 vdd gnd cell_6t
Xbit_r165_c232 bl_232 br_232 wl_165 vdd gnd cell_6t
Xbit_r166_c232 bl_232 br_232 wl_166 vdd gnd cell_6t
Xbit_r167_c232 bl_232 br_232 wl_167 vdd gnd cell_6t
Xbit_r168_c232 bl_232 br_232 wl_168 vdd gnd cell_6t
Xbit_r169_c232 bl_232 br_232 wl_169 vdd gnd cell_6t
Xbit_r170_c232 bl_232 br_232 wl_170 vdd gnd cell_6t
Xbit_r171_c232 bl_232 br_232 wl_171 vdd gnd cell_6t
Xbit_r172_c232 bl_232 br_232 wl_172 vdd gnd cell_6t
Xbit_r173_c232 bl_232 br_232 wl_173 vdd gnd cell_6t
Xbit_r174_c232 bl_232 br_232 wl_174 vdd gnd cell_6t
Xbit_r175_c232 bl_232 br_232 wl_175 vdd gnd cell_6t
Xbit_r176_c232 bl_232 br_232 wl_176 vdd gnd cell_6t
Xbit_r177_c232 bl_232 br_232 wl_177 vdd gnd cell_6t
Xbit_r178_c232 bl_232 br_232 wl_178 vdd gnd cell_6t
Xbit_r179_c232 bl_232 br_232 wl_179 vdd gnd cell_6t
Xbit_r180_c232 bl_232 br_232 wl_180 vdd gnd cell_6t
Xbit_r181_c232 bl_232 br_232 wl_181 vdd gnd cell_6t
Xbit_r182_c232 bl_232 br_232 wl_182 vdd gnd cell_6t
Xbit_r183_c232 bl_232 br_232 wl_183 vdd gnd cell_6t
Xbit_r184_c232 bl_232 br_232 wl_184 vdd gnd cell_6t
Xbit_r185_c232 bl_232 br_232 wl_185 vdd gnd cell_6t
Xbit_r186_c232 bl_232 br_232 wl_186 vdd gnd cell_6t
Xbit_r187_c232 bl_232 br_232 wl_187 vdd gnd cell_6t
Xbit_r188_c232 bl_232 br_232 wl_188 vdd gnd cell_6t
Xbit_r189_c232 bl_232 br_232 wl_189 vdd gnd cell_6t
Xbit_r190_c232 bl_232 br_232 wl_190 vdd gnd cell_6t
Xbit_r191_c232 bl_232 br_232 wl_191 vdd gnd cell_6t
Xbit_r192_c232 bl_232 br_232 wl_192 vdd gnd cell_6t
Xbit_r193_c232 bl_232 br_232 wl_193 vdd gnd cell_6t
Xbit_r194_c232 bl_232 br_232 wl_194 vdd gnd cell_6t
Xbit_r195_c232 bl_232 br_232 wl_195 vdd gnd cell_6t
Xbit_r196_c232 bl_232 br_232 wl_196 vdd gnd cell_6t
Xbit_r197_c232 bl_232 br_232 wl_197 vdd gnd cell_6t
Xbit_r198_c232 bl_232 br_232 wl_198 vdd gnd cell_6t
Xbit_r199_c232 bl_232 br_232 wl_199 vdd gnd cell_6t
Xbit_r200_c232 bl_232 br_232 wl_200 vdd gnd cell_6t
Xbit_r201_c232 bl_232 br_232 wl_201 vdd gnd cell_6t
Xbit_r202_c232 bl_232 br_232 wl_202 vdd gnd cell_6t
Xbit_r203_c232 bl_232 br_232 wl_203 vdd gnd cell_6t
Xbit_r204_c232 bl_232 br_232 wl_204 vdd gnd cell_6t
Xbit_r205_c232 bl_232 br_232 wl_205 vdd gnd cell_6t
Xbit_r206_c232 bl_232 br_232 wl_206 vdd gnd cell_6t
Xbit_r207_c232 bl_232 br_232 wl_207 vdd gnd cell_6t
Xbit_r208_c232 bl_232 br_232 wl_208 vdd gnd cell_6t
Xbit_r209_c232 bl_232 br_232 wl_209 vdd gnd cell_6t
Xbit_r210_c232 bl_232 br_232 wl_210 vdd gnd cell_6t
Xbit_r211_c232 bl_232 br_232 wl_211 vdd gnd cell_6t
Xbit_r212_c232 bl_232 br_232 wl_212 vdd gnd cell_6t
Xbit_r213_c232 bl_232 br_232 wl_213 vdd gnd cell_6t
Xbit_r214_c232 bl_232 br_232 wl_214 vdd gnd cell_6t
Xbit_r215_c232 bl_232 br_232 wl_215 vdd gnd cell_6t
Xbit_r216_c232 bl_232 br_232 wl_216 vdd gnd cell_6t
Xbit_r217_c232 bl_232 br_232 wl_217 vdd gnd cell_6t
Xbit_r218_c232 bl_232 br_232 wl_218 vdd gnd cell_6t
Xbit_r219_c232 bl_232 br_232 wl_219 vdd gnd cell_6t
Xbit_r220_c232 bl_232 br_232 wl_220 vdd gnd cell_6t
Xbit_r221_c232 bl_232 br_232 wl_221 vdd gnd cell_6t
Xbit_r222_c232 bl_232 br_232 wl_222 vdd gnd cell_6t
Xbit_r223_c232 bl_232 br_232 wl_223 vdd gnd cell_6t
Xbit_r224_c232 bl_232 br_232 wl_224 vdd gnd cell_6t
Xbit_r225_c232 bl_232 br_232 wl_225 vdd gnd cell_6t
Xbit_r226_c232 bl_232 br_232 wl_226 vdd gnd cell_6t
Xbit_r227_c232 bl_232 br_232 wl_227 vdd gnd cell_6t
Xbit_r228_c232 bl_232 br_232 wl_228 vdd gnd cell_6t
Xbit_r229_c232 bl_232 br_232 wl_229 vdd gnd cell_6t
Xbit_r230_c232 bl_232 br_232 wl_230 vdd gnd cell_6t
Xbit_r231_c232 bl_232 br_232 wl_231 vdd gnd cell_6t
Xbit_r232_c232 bl_232 br_232 wl_232 vdd gnd cell_6t
Xbit_r233_c232 bl_232 br_232 wl_233 vdd gnd cell_6t
Xbit_r234_c232 bl_232 br_232 wl_234 vdd gnd cell_6t
Xbit_r235_c232 bl_232 br_232 wl_235 vdd gnd cell_6t
Xbit_r236_c232 bl_232 br_232 wl_236 vdd gnd cell_6t
Xbit_r237_c232 bl_232 br_232 wl_237 vdd gnd cell_6t
Xbit_r238_c232 bl_232 br_232 wl_238 vdd gnd cell_6t
Xbit_r239_c232 bl_232 br_232 wl_239 vdd gnd cell_6t
Xbit_r240_c232 bl_232 br_232 wl_240 vdd gnd cell_6t
Xbit_r241_c232 bl_232 br_232 wl_241 vdd gnd cell_6t
Xbit_r242_c232 bl_232 br_232 wl_242 vdd gnd cell_6t
Xbit_r243_c232 bl_232 br_232 wl_243 vdd gnd cell_6t
Xbit_r244_c232 bl_232 br_232 wl_244 vdd gnd cell_6t
Xbit_r245_c232 bl_232 br_232 wl_245 vdd gnd cell_6t
Xbit_r246_c232 bl_232 br_232 wl_246 vdd gnd cell_6t
Xbit_r247_c232 bl_232 br_232 wl_247 vdd gnd cell_6t
Xbit_r248_c232 bl_232 br_232 wl_248 vdd gnd cell_6t
Xbit_r249_c232 bl_232 br_232 wl_249 vdd gnd cell_6t
Xbit_r250_c232 bl_232 br_232 wl_250 vdd gnd cell_6t
Xbit_r251_c232 bl_232 br_232 wl_251 vdd gnd cell_6t
Xbit_r252_c232 bl_232 br_232 wl_252 vdd gnd cell_6t
Xbit_r253_c232 bl_232 br_232 wl_253 vdd gnd cell_6t
Xbit_r254_c232 bl_232 br_232 wl_254 vdd gnd cell_6t
Xbit_r255_c232 bl_232 br_232 wl_255 vdd gnd cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd cell_6t
Xbit_r1_c233 bl_233 br_233 wl_1 vdd gnd cell_6t
Xbit_r2_c233 bl_233 br_233 wl_2 vdd gnd cell_6t
Xbit_r3_c233 bl_233 br_233 wl_3 vdd gnd cell_6t
Xbit_r4_c233 bl_233 br_233 wl_4 vdd gnd cell_6t
Xbit_r5_c233 bl_233 br_233 wl_5 vdd gnd cell_6t
Xbit_r6_c233 bl_233 br_233 wl_6 vdd gnd cell_6t
Xbit_r7_c233 bl_233 br_233 wl_7 vdd gnd cell_6t
Xbit_r8_c233 bl_233 br_233 wl_8 vdd gnd cell_6t
Xbit_r9_c233 bl_233 br_233 wl_9 vdd gnd cell_6t
Xbit_r10_c233 bl_233 br_233 wl_10 vdd gnd cell_6t
Xbit_r11_c233 bl_233 br_233 wl_11 vdd gnd cell_6t
Xbit_r12_c233 bl_233 br_233 wl_12 vdd gnd cell_6t
Xbit_r13_c233 bl_233 br_233 wl_13 vdd gnd cell_6t
Xbit_r14_c233 bl_233 br_233 wl_14 vdd gnd cell_6t
Xbit_r15_c233 bl_233 br_233 wl_15 vdd gnd cell_6t
Xbit_r16_c233 bl_233 br_233 wl_16 vdd gnd cell_6t
Xbit_r17_c233 bl_233 br_233 wl_17 vdd gnd cell_6t
Xbit_r18_c233 bl_233 br_233 wl_18 vdd gnd cell_6t
Xbit_r19_c233 bl_233 br_233 wl_19 vdd gnd cell_6t
Xbit_r20_c233 bl_233 br_233 wl_20 vdd gnd cell_6t
Xbit_r21_c233 bl_233 br_233 wl_21 vdd gnd cell_6t
Xbit_r22_c233 bl_233 br_233 wl_22 vdd gnd cell_6t
Xbit_r23_c233 bl_233 br_233 wl_23 vdd gnd cell_6t
Xbit_r24_c233 bl_233 br_233 wl_24 vdd gnd cell_6t
Xbit_r25_c233 bl_233 br_233 wl_25 vdd gnd cell_6t
Xbit_r26_c233 bl_233 br_233 wl_26 vdd gnd cell_6t
Xbit_r27_c233 bl_233 br_233 wl_27 vdd gnd cell_6t
Xbit_r28_c233 bl_233 br_233 wl_28 vdd gnd cell_6t
Xbit_r29_c233 bl_233 br_233 wl_29 vdd gnd cell_6t
Xbit_r30_c233 bl_233 br_233 wl_30 vdd gnd cell_6t
Xbit_r31_c233 bl_233 br_233 wl_31 vdd gnd cell_6t
Xbit_r32_c233 bl_233 br_233 wl_32 vdd gnd cell_6t
Xbit_r33_c233 bl_233 br_233 wl_33 vdd gnd cell_6t
Xbit_r34_c233 bl_233 br_233 wl_34 vdd gnd cell_6t
Xbit_r35_c233 bl_233 br_233 wl_35 vdd gnd cell_6t
Xbit_r36_c233 bl_233 br_233 wl_36 vdd gnd cell_6t
Xbit_r37_c233 bl_233 br_233 wl_37 vdd gnd cell_6t
Xbit_r38_c233 bl_233 br_233 wl_38 vdd gnd cell_6t
Xbit_r39_c233 bl_233 br_233 wl_39 vdd gnd cell_6t
Xbit_r40_c233 bl_233 br_233 wl_40 vdd gnd cell_6t
Xbit_r41_c233 bl_233 br_233 wl_41 vdd gnd cell_6t
Xbit_r42_c233 bl_233 br_233 wl_42 vdd gnd cell_6t
Xbit_r43_c233 bl_233 br_233 wl_43 vdd gnd cell_6t
Xbit_r44_c233 bl_233 br_233 wl_44 vdd gnd cell_6t
Xbit_r45_c233 bl_233 br_233 wl_45 vdd gnd cell_6t
Xbit_r46_c233 bl_233 br_233 wl_46 vdd gnd cell_6t
Xbit_r47_c233 bl_233 br_233 wl_47 vdd gnd cell_6t
Xbit_r48_c233 bl_233 br_233 wl_48 vdd gnd cell_6t
Xbit_r49_c233 bl_233 br_233 wl_49 vdd gnd cell_6t
Xbit_r50_c233 bl_233 br_233 wl_50 vdd gnd cell_6t
Xbit_r51_c233 bl_233 br_233 wl_51 vdd gnd cell_6t
Xbit_r52_c233 bl_233 br_233 wl_52 vdd gnd cell_6t
Xbit_r53_c233 bl_233 br_233 wl_53 vdd gnd cell_6t
Xbit_r54_c233 bl_233 br_233 wl_54 vdd gnd cell_6t
Xbit_r55_c233 bl_233 br_233 wl_55 vdd gnd cell_6t
Xbit_r56_c233 bl_233 br_233 wl_56 vdd gnd cell_6t
Xbit_r57_c233 bl_233 br_233 wl_57 vdd gnd cell_6t
Xbit_r58_c233 bl_233 br_233 wl_58 vdd gnd cell_6t
Xbit_r59_c233 bl_233 br_233 wl_59 vdd gnd cell_6t
Xbit_r60_c233 bl_233 br_233 wl_60 vdd gnd cell_6t
Xbit_r61_c233 bl_233 br_233 wl_61 vdd gnd cell_6t
Xbit_r62_c233 bl_233 br_233 wl_62 vdd gnd cell_6t
Xbit_r63_c233 bl_233 br_233 wl_63 vdd gnd cell_6t
Xbit_r64_c233 bl_233 br_233 wl_64 vdd gnd cell_6t
Xbit_r65_c233 bl_233 br_233 wl_65 vdd gnd cell_6t
Xbit_r66_c233 bl_233 br_233 wl_66 vdd gnd cell_6t
Xbit_r67_c233 bl_233 br_233 wl_67 vdd gnd cell_6t
Xbit_r68_c233 bl_233 br_233 wl_68 vdd gnd cell_6t
Xbit_r69_c233 bl_233 br_233 wl_69 vdd gnd cell_6t
Xbit_r70_c233 bl_233 br_233 wl_70 vdd gnd cell_6t
Xbit_r71_c233 bl_233 br_233 wl_71 vdd gnd cell_6t
Xbit_r72_c233 bl_233 br_233 wl_72 vdd gnd cell_6t
Xbit_r73_c233 bl_233 br_233 wl_73 vdd gnd cell_6t
Xbit_r74_c233 bl_233 br_233 wl_74 vdd gnd cell_6t
Xbit_r75_c233 bl_233 br_233 wl_75 vdd gnd cell_6t
Xbit_r76_c233 bl_233 br_233 wl_76 vdd gnd cell_6t
Xbit_r77_c233 bl_233 br_233 wl_77 vdd gnd cell_6t
Xbit_r78_c233 bl_233 br_233 wl_78 vdd gnd cell_6t
Xbit_r79_c233 bl_233 br_233 wl_79 vdd gnd cell_6t
Xbit_r80_c233 bl_233 br_233 wl_80 vdd gnd cell_6t
Xbit_r81_c233 bl_233 br_233 wl_81 vdd gnd cell_6t
Xbit_r82_c233 bl_233 br_233 wl_82 vdd gnd cell_6t
Xbit_r83_c233 bl_233 br_233 wl_83 vdd gnd cell_6t
Xbit_r84_c233 bl_233 br_233 wl_84 vdd gnd cell_6t
Xbit_r85_c233 bl_233 br_233 wl_85 vdd gnd cell_6t
Xbit_r86_c233 bl_233 br_233 wl_86 vdd gnd cell_6t
Xbit_r87_c233 bl_233 br_233 wl_87 vdd gnd cell_6t
Xbit_r88_c233 bl_233 br_233 wl_88 vdd gnd cell_6t
Xbit_r89_c233 bl_233 br_233 wl_89 vdd gnd cell_6t
Xbit_r90_c233 bl_233 br_233 wl_90 vdd gnd cell_6t
Xbit_r91_c233 bl_233 br_233 wl_91 vdd gnd cell_6t
Xbit_r92_c233 bl_233 br_233 wl_92 vdd gnd cell_6t
Xbit_r93_c233 bl_233 br_233 wl_93 vdd gnd cell_6t
Xbit_r94_c233 bl_233 br_233 wl_94 vdd gnd cell_6t
Xbit_r95_c233 bl_233 br_233 wl_95 vdd gnd cell_6t
Xbit_r96_c233 bl_233 br_233 wl_96 vdd gnd cell_6t
Xbit_r97_c233 bl_233 br_233 wl_97 vdd gnd cell_6t
Xbit_r98_c233 bl_233 br_233 wl_98 vdd gnd cell_6t
Xbit_r99_c233 bl_233 br_233 wl_99 vdd gnd cell_6t
Xbit_r100_c233 bl_233 br_233 wl_100 vdd gnd cell_6t
Xbit_r101_c233 bl_233 br_233 wl_101 vdd gnd cell_6t
Xbit_r102_c233 bl_233 br_233 wl_102 vdd gnd cell_6t
Xbit_r103_c233 bl_233 br_233 wl_103 vdd gnd cell_6t
Xbit_r104_c233 bl_233 br_233 wl_104 vdd gnd cell_6t
Xbit_r105_c233 bl_233 br_233 wl_105 vdd gnd cell_6t
Xbit_r106_c233 bl_233 br_233 wl_106 vdd gnd cell_6t
Xbit_r107_c233 bl_233 br_233 wl_107 vdd gnd cell_6t
Xbit_r108_c233 bl_233 br_233 wl_108 vdd gnd cell_6t
Xbit_r109_c233 bl_233 br_233 wl_109 vdd gnd cell_6t
Xbit_r110_c233 bl_233 br_233 wl_110 vdd gnd cell_6t
Xbit_r111_c233 bl_233 br_233 wl_111 vdd gnd cell_6t
Xbit_r112_c233 bl_233 br_233 wl_112 vdd gnd cell_6t
Xbit_r113_c233 bl_233 br_233 wl_113 vdd gnd cell_6t
Xbit_r114_c233 bl_233 br_233 wl_114 vdd gnd cell_6t
Xbit_r115_c233 bl_233 br_233 wl_115 vdd gnd cell_6t
Xbit_r116_c233 bl_233 br_233 wl_116 vdd gnd cell_6t
Xbit_r117_c233 bl_233 br_233 wl_117 vdd gnd cell_6t
Xbit_r118_c233 bl_233 br_233 wl_118 vdd gnd cell_6t
Xbit_r119_c233 bl_233 br_233 wl_119 vdd gnd cell_6t
Xbit_r120_c233 bl_233 br_233 wl_120 vdd gnd cell_6t
Xbit_r121_c233 bl_233 br_233 wl_121 vdd gnd cell_6t
Xbit_r122_c233 bl_233 br_233 wl_122 vdd gnd cell_6t
Xbit_r123_c233 bl_233 br_233 wl_123 vdd gnd cell_6t
Xbit_r124_c233 bl_233 br_233 wl_124 vdd gnd cell_6t
Xbit_r125_c233 bl_233 br_233 wl_125 vdd gnd cell_6t
Xbit_r126_c233 bl_233 br_233 wl_126 vdd gnd cell_6t
Xbit_r127_c233 bl_233 br_233 wl_127 vdd gnd cell_6t
Xbit_r128_c233 bl_233 br_233 wl_128 vdd gnd cell_6t
Xbit_r129_c233 bl_233 br_233 wl_129 vdd gnd cell_6t
Xbit_r130_c233 bl_233 br_233 wl_130 vdd gnd cell_6t
Xbit_r131_c233 bl_233 br_233 wl_131 vdd gnd cell_6t
Xbit_r132_c233 bl_233 br_233 wl_132 vdd gnd cell_6t
Xbit_r133_c233 bl_233 br_233 wl_133 vdd gnd cell_6t
Xbit_r134_c233 bl_233 br_233 wl_134 vdd gnd cell_6t
Xbit_r135_c233 bl_233 br_233 wl_135 vdd gnd cell_6t
Xbit_r136_c233 bl_233 br_233 wl_136 vdd gnd cell_6t
Xbit_r137_c233 bl_233 br_233 wl_137 vdd gnd cell_6t
Xbit_r138_c233 bl_233 br_233 wl_138 vdd gnd cell_6t
Xbit_r139_c233 bl_233 br_233 wl_139 vdd gnd cell_6t
Xbit_r140_c233 bl_233 br_233 wl_140 vdd gnd cell_6t
Xbit_r141_c233 bl_233 br_233 wl_141 vdd gnd cell_6t
Xbit_r142_c233 bl_233 br_233 wl_142 vdd gnd cell_6t
Xbit_r143_c233 bl_233 br_233 wl_143 vdd gnd cell_6t
Xbit_r144_c233 bl_233 br_233 wl_144 vdd gnd cell_6t
Xbit_r145_c233 bl_233 br_233 wl_145 vdd gnd cell_6t
Xbit_r146_c233 bl_233 br_233 wl_146 vdd gnd cell_6t
Xbit_r147_c233 bl_233 br_233 wl_147 vdd gnd cell_6t
Xbit_r148_c233 bl_233 br_233 wl_148 vdd gnd cell_6t
Xbit_r149_c233 bl_233 br_233 wl_149 vdd gnd cell_6t
Xbit_r150_c233 bl_233 br_233 wl_150 vdd gnd cell_6t
Xbit_r151_c233 bl_233 br_233 wl_151 vdd gnd cell_6t
Xbit_r152_c233 bl_233 br_233 wl_152 vdd gnd cell_6t
Xbit_r153_c233 bl_233 br_233 wl_153 vdd gnd cell_6t
Xbit_r154_c233 bl_233 br_233 wl_154 vdd gnd cell_6t
Xbit_r155_c233 bl_233 br_233 wl_155 vdd gnd cell_6t
Xbit_r156_c233 bl_233 br_233 wl_156 vdd gnd cell_6t
Xbit_r157_c233 bl_233 br_233 wl_157 vdd gnd cell_6t
Xbit_r158_c233 bl_233 br_233 wl_158 vdd gnd cell_6t
Xbit_r159_c233 bl_233 br_233 wl_159 vdd gnd cell_6t
Xbit_r160_c233 bl_233 br_233 wl_160 vdd gnd cell_6t
Xbit_r161_c233 bl_233 br_233 wl_161 vdd gnd cell_6t
Xbit_r162_c233 bl_233 br_233 wl_162 vdd gnd cell_6t
Xbit_r163_c233 bl_233 br_233 wl_163 vdd gnd cell_6t
Xbit_r164_c233 bl_233 br_233 wl_164 vdd gnd cell_6t
Xbit_r165_c233 bl_233 br_233 wl_165 vdd gnd cell_6t
Xbit_r166_c233 bl_233 br_233 wl_166 vdd gnd cell_6t
Xbit_r167_c233 bl_233 br_233 wl_167 vdd gnd cell_6t
Xbit_r168_c233 bl_233 br_233 wl_168 vdd gnd cell_6t
Xbit_r169_c233 bl_233 br_233 wl_169 vdd gnd cell_6t
Xbit_r170_c233 bl_233 br_233 wl_170 vdd gnd cell_6t
Xbit_r171_c233 bl_233 br_233 wl_171 vdd gnd cell_6t
Xbit_r172_c233 bl_233 br_233 wl_172 vdd gnd cell_6t
Xbit_r173_c233 bl_233 br_233 wl_173 vdd gnd cell_6t
Xbit_r174_c233 bl_233 br_233 wl_174 vdd gnd cell_6t
Xbit_r175_c233 bl_233 br_233 wl_175 vdd gnd cell_6t
Xbit_r176_c233 bl_233 br_233 wl_176 vdd gnd cell_6t
Xbit_r177_c233 bl_233 br_233 wl_177 vdd gnd cell_6t
Xbit_r178_c233 bl_233 br_233 wl_178 vdd gnd cell_6t
Xbit_r179_c233 bl_233 br_233 wl_179 vdd gnd cell_6t
Xbit_r180_c233 bl_233 br_233 wl_180 vdd gnd cell_6t
Xbit_r181_c233 bl_233 br_233 wl_181 vdd gnd cell_6t
Xbit_r182_c233 bl_233 br_233 wl_182 vdd gnd cell_6t
Xbit_r183_c233 bl_233 br_233 wl_183 vdd gnd cell_6t
Xbit_r184_c233 bl_233 br_233 wl_184 vdd gnd cell_6t
Xbit_r185_c233 bl_233 br_233 wl_185 vdd gnd cell_6t
Xbit_r186_c233 bl_233 br_233 wl_186 vdd gnd cell_6t
Xbit_r187_c233 bl_233 br_233 wl_187 vdd gnd cell_6t
Xbit_r188_c233 bl_233 br_233 wl_188 vdd gnd cell_6t
Xbit_r189_c233 bl_233 br_233 wl_189 vdd gnd cell_6t
Xbit_r190_c233 bl_233 br_233 wl_190 vdd gnd cell_6t
Xbit_r191_c233 bl_233 br_233 wl_191 vdd gnd cell_6t
Xbit_r192_c233 bl_233 br_233 wl_192 vdd gnd cell_6t
Xbit_r193_c233 bl_233 br_233 wl_193 vdd gnd cell_6t
Xbit_r194_c233 bl_233 br_233 wl_194 vdd gnd cell_6t
Xbit_r195_c233 bl_233 br_233 wl_195 vdd gnd cell_6t
Xbit_r196_c233 bl_233 br_233 wl_196 vdd gnd cell_6t
Xbit_r197_c233 bl_233 br_233 wl_197 vdd gnd cell_6t
Xbit_r198_c233 bl_233 br_233 wl_198 vdd gnd cell_6t
Xbit_r199_c233 bl_233 br_233 wl_199 vdd gnd cell_6t
Xbit_r200_c233 bl_233 br_233 wl_200 vdd gnd cell_6t
Xbit_r201_c233 bl_233 br_233 wl_201 vdd gnd cell_6t
Xbit_r202_c233 bl_233 br_233 wl_202 vdd gnd cell_6t
Xbit_r203_c233 bl_233 br_233 wl_203 vdd gnd cell_6t
Xbit_r204_c233 bl_233 br_233 wl_204 vdd gnd cell_6t
Xbit_r205_c233 bl_233 br_233 wl_205 vdd gnd cell_6t
Xbit_r206_c233 bl_233 br_233 wl_206 vdd gnd cell_6t
Xbit_r207_c233 bl_233 br_233 wl_207 vdd gnd cell_6t
Xbit_r208_c233 bl_233 br_233 wl_208 vdd gnd cell_6t
Xbit_r209_c233 bl_233 br_233 wl_209 vdd gnd cell_6t
Xbit_r210_c233 bl_233 br_233 wl_210 vdd gnd cell_6t
Xbit_r211_c233 bl_233 br_233 wl_211 vdd gnd cell_6t
Xbit_r212_c233 bl_233 br_233 wl_212 vdd gnd cell_6t
Xbit_r213_c233 bl_233 br_233 wl_213 vdd gnd cell_6t
Xbit_r214_c233 bl_233 br_233 wl_214 vdd gnd cell_6t
Xbit_r215_c233 bl_233 br_233 wl_215 vdd gnd cell_6t
Xbit_r216_c233 bl_233 br_233 wl_216 vdd gnd cell_6t
Xbit_r217_c233 bl_233 br_233 wl_217 vdd gnd cell_6t
Xbit_r218_c233 bl_233 br_233 wl_218 vdd gnd cell_6t
Xbit_r219_c233 bl_233 br_233 wl_219 vdd gnd cell_6t
Xbit_r220_c233 bl_233 br_233 wl_220 vdd gnd cell_6t
Xbit_r221_c233 bl_233 br_233 wl_221 vdd gnd cell_6t
Xbit_r222_c233 bl_233 br_233 wl_222 vdd gnd cell_6t
Xbit_r223_c233 bl_233 br_233 wl_223 vdd gnd cell_6t
Xbit_r224_c233 bl_233 br_233 wl_224 vdd gnd cell_6t
Xbit_r225_c233 bl_233 br_233 wl_225 vdd gnd cell_6t
Xbit_r226_c233 bl_233 br_233 wl_226 vdd gnd cell_6t
Xbit_r227_c233 bl_233 br_233 wl_227 vdd gnd cell_6t
Xbit_r228_c233 bl_233 br_233 wl_228 vdd gnd cell_6t
Xbit_r229_c233 bl_233 br_233 wl_229 vdd gnd cell_6t
Xbit_r230_c233 bl_233 br_233 wl_230 vdd gnd cell_6t
Xbit_r231_c233 bl_233 br_233 wl_231 vdd gnd cell_6t
Xbit_r232_c233 bl_233 br_233 wl_232 vdd gnd cell_6t
Xbit_r233_c233 bl_233 br_233 wl_233 vdd gnd cell_6t
Xbit_r234_c233 bl_233 br_233 wl_234 vdd gnd cell_6t
Xbit_r235_c233 bl_233 br_233 wl_235 vdd gnd cell_6t
Xbit_r236_c233 bl_233 br_233 wl_236 vdd gnd cell_6t
Xbit_r237_c233 bl_233 br_233 wl_237 vdd gnd cell_6t
Xbit_r238_c233 bl_233 br_233 wl_238 vdd gnd cell_6t
Xbit_r239_c233 bl_233 br_233 wl_239 vdd gnd cell_6t
Xbit_r240_c233 bl_233 br_233 wl_240 vdd gnd cell_6t
Xbit_r241_c233 bl_233 br_233 wl_241 vdd gnd cell_6t
Xbit_r242_c233 bl_233 br_233 wl_242 vdd gnd cell_6t
Xbit_r243_c233 bl_233 br_233 wl_243 vdd gnd cell_6t
Xbit_r244_c233 bl_233 br_233 wl_244 vdd gnd cell_6t
Xbit_r245_c233 bl_233 br_233 wl_245 vdd gnd cell_6t
Xbit_r246_c233 bl_233 br_233 wl_246 vdd gnd cell_6t
Xbit_r247_c233 bl_233 br_233 wl_247 vdd gnd cell_6t
Xbit_r248_c233 bl_233 br_233 wl_248 vdd gnd cell_6t
Xbit_r249_c233 bl_233 br_233 wl_249 vdd gnd cell_6t
Xbit_r250_c233 bl_233 br_233 wl_250 vdd gnd cell_6t
Xbit_r251_c233 bl_233 br_233 wl_251 vdd gnd cell_6t
Xbit_r252_c233 bl_233 br_233 wl_252 vdd gnd cell_6t
Xbit_r253_c233 bl_233 br_233 wl_253 vdd gnd cell_6t
Xbit_r254_c233 bl_233 br_233 wl_254 vdd gnd cell_6t
Xbit_r255_c233 bl_233 br_233 wl_255 vdd gnd cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd cell_6t
Xbit_r1_c234 bl_234 br_234 wl_1 vdd gnd cell_6t
Xbit_r2_c234 bl_234 br_234 wl_2 vdd gnd cell_6t
Xbit_r3_c234 bl_234 br_234 wl_3 vdd gnd cell_6t
Xbit_r4_c234 bl_234 br_234 wl_4 vdd gnd cell_6t
Xbit_r5_c234 bl_234 br_234 wl_5 vdd gnd cell_6t
Xbit_r6_c234 bl_234 br_234 wl_6 vdd gnd cell_6t
Xbit_r7_c234 bl_234 br_234 wl_7 vdd gnd cell_6t
Xbit_r8_c234 bl_234 br_234 wl_8 vdd gnd cell_6t
Xbit_r9_c234 bl_234 br_234 wl_9 vdd gnd cell_6t
Xbit_r10_c234 bl_234 br_234 wl_10 vdd gnd cell_6t
Xbit_r11_c234 bl_234 br_234 wl_11 vdd gnd cell_6t
Xbit_r12_c234 bl_234 br_234 wl_12 vdd gnd cell_6t
Xbit_r13_c234 bl_234 br_234 wl_13 vdd gnd cell_6t
Xbit_r14_c234 bl_234 br_234 wl_14 vdd gnd cell_6t
Xbit_r15_c234 bl_234 br_234 wl_15 vdd gnd cell_6t
Xbit_r16_c234 bl_234 br_234 wl_16 vdd gnd cell_6t
Xbit_r17_c234 bl_234 br_234 wl_17 vdd gnd cell_6t
Xbit_r18_c234 bl_234 br_234 wl_18 vdd gnd cell_6t
Xbit_r19_c234 bl_234 br_234 wl_19 vdd gnd cell_6t
Xbit_r20_c234 bl_234 br_234 wl_20 vdd gnd cell_6t
Xbit_r21_c234 bl_234 br_234 wl_21 vdd gnd cell_6t
Xbit_r22_c234 bl_234 br_234 wl_22 vdd gnd cell_6t
Xbit_r23_c234 bl_234 br_234 wl_23 vdd gnd cell_6t
Xbit_r24_c234 bl_234 br_234 wl_24 vdd gnd cell_6t
Xbit_r25_c234 bl_234 br_234 wl_25 vdd gnd cell_6t
Xbit_r26_c234 bl_234 br_234 wl_26 vdd gnd cell_6t
Xbit_r27_c234 bl_234 br_234 wl_27 vdd gnd cell_6t
Xbit_r28_c234 bl_234 br_234 wl_28 vdd gnd cell_6t
Xbit_r29_c234 bl_234 br_234 wl_29 vdd gnd cell_6t
Xbit_r30_c234 bl_234 br_234 wl_30 vdd gnd cell_6t
Xbit_r31_c234 bl_234 br_234 wl_31 vdd gnd cell_6t
Xbit_r32_c234 bl_234 br_234 wl_32 vdd gnd cell_6t
Xbit_r33_c234 bl_234 br_234 wl_33 vdd gnd cell_6t
Xbit_r34_c234 bl_234 br_234 wl_34 vdd gnd cell_6t
Xbit_r35_c234 bl_234 br_234 wl_35 vdd gnd cell_6t
Xbit_r36_c234 bl_234 br_234 wl_36 vdd gnd cell_6t
Xbit_r37_c234 bl_234 br_234 wl_37 vdd gnd cell_6t
Xbit_r38_c234 bl_234 br_234 wl_38 vdd gnd cell_6t
Xbit_r39_c234 bl_234 br_234 wl_39 vdd gnd cell_6t
Xbit_r40_c234 bl_234 br_234 wl_40 vdd gnd cell_6t
Xbit_r41_c234 bl_234 br_234 wl_41 vdd gnd cell_6t
Xbit_r42_c234 bl_234 br_234 wl_42 vdd gnd cell_6t
Xbit_r43_c234 bl_234 br_234 wl_43 vdd gnd cell_6t
Xbit_r44_c234 bl_234 br_234 wl_44 vdd gnd cell_6t
Xbit_r45_c234 bl_234 br_234 wl_45 vdd gnd cell_6t
Xbit_r46_c234 bl_234 br_234 wl_46 vdd gnd cell_6t
Xbit_r47_c234 bl_234 br_234 wl_47 vdd gnd cell_6t
Xbit_r48_c234 bl_234 br_234 wl_48 vdd gnd cell_6t
Xbit_r49_c234 bl_234 br_234 wl_49 vdd gnd cell_6t
Xbit_r50_c234 bl_234 br_234 wl_50 vdd gnd cell_6t
Xbit_r51_c234 bl_234 br_234 wl_51 vdd gnd cell_6t
Xbit_r52_c234 bl_234 br_234 wl_52 vdd gnd cell_6t
Xbit_r53_c234 bl_234 br_234 wl_53 vdd gnd cell_6t
Xbit_r54_c234 bl_234 br_234 wl_54 vdd gnd cell_6t
Xbit_r55_c234 bl_234 br_234 wl_55 vdd gnd cell_6t
Xbit_r56_c234 bl_234 br_234 wl_56 vdd gnd cell_6t
Xbit_r57_c234 bl_234 br_234 wl_57 vdd gnd cell_6t
Xbit_r58_c234 bl_234 br_234 wl_58 vdd gnd cell_6t
Xbit_r59_c234 bl_234 br_234 wl_59 vdd gnd cell_6t
Xbit_r60_c234 bl_234 br_234 wl_60 vdd gnd cell_6t
Xbit_r61_c234 bl_234 br_234 wl_61 vdd gnd cell_6t
Xbit_r62_c234 bl_234 br_234 wl_62 vdd gnd cell_6t
Xbit_r63_c234 bl_234 br_234 wl_63 vdd gnd cell_6t
Xbit_r64_c234 bl_234 br_234 wl_64 vdd gnd cell_6t
Xbit_r65_c234 bl_234 br_234 wl_65 vdd gnd cell_6t
Xbit_r66_c234 bl_234 br_234 wl_66 vdd gnd cell_6t
Xbit_r67_c234 bl_234 br_234 wl_67 vdd gnd cell_6t
Xbit_r68_c234 bl_234 br_234 wl_68 vdd gnd cell_6t
Xbit_r69_c234 bl_234 br_234 wl_69 vdd gnd cell_6t
Xbit_r70_c234 bl_234 br_234 wl_70 vdd gnd cell_6t
Xbit_r71_c234 bl_234 br_234 wl_71 vdd gnd cell_6t
Xbit_r72_c234 bl_234 br_234 wl_72 vdd gnd cell_6t
Xbit_r73_c234 bl_234 br_234 wl_73 vdd gnd cell_6t
Xbit_r74_c234 bl_234 br_234 wl_74 vdd gnd cell_6t
Xbit_r75_c234 bl_234 br_234 wl_75 vdd gnd cell_6t
Xbit_r76_c234 bl_234 br_234 wl_76 vdd gnd cell_6t
Xbit_r77_c234 bl_234 br_234 wl_77 vdd gnd cell_6t
Xbit_r78_c234 bl_234 br_234 wl_78 vdd gnd cell_6t
Xbit_r79_c234 bl_234 br_234 wl_79 vdd gnd cell_6t
Xbit_r80_c234 bl_234 br_234 wl_80 vdd gnd cell_6t
Xbit_r81_c234 bl_234 br_234 wl_81 vdd gnd cell_6t
Xbit_r82_c234 bl_234 br_234 wl_82 vdd gnd cell_6t
Xbit_r83_c234 bl_234 br_234 wl_83 vdd gnd cell_6t
Xbit_r84_c234 bl_234 br_234 wl_84 vdd gnd cell_6t
Xbit_r85_c234 bl_234 br_234 wl_85 vdd gnd cell_6t
Xbit_r86_c234 bl_234 br_234 wl_86 vdd gnd cell_6t
Xbit_r87_c234 bl_234 br_234 wl_87 vdd gnd cell_6t
Xbit_r88_c234 bl_234 br_234 wl_88 vdd gnd cell_6t
Xbit_r89_c234 bl_234 br_234 wl_89 vdd gnd cell_6t
Xbit_r90_c234 bl_234 br_234 wl_90 vdd gnd cell_6t
Xbit_r91_c234 bl_234 br_234 wl_91 vdd gnd cell_6t
Xbit_r92_c234 bl_234 br_234 wl_92 vdd gnd cell_6t
Xbit_r93_c234 bl_234 br_234 wl_93 vdd gnd cell_6t
Xbit_r94_c234 bl_234 br_234 wl_94 vdd gnd cell_6t
Xbit_r95_c234 bl_234 br_234 wl_95 vdd gnd cell_6t
Xbit_r96_c234 bl_234 br_234 wl_96 vdd gnd cell_6t
Xbit_r97_c234 bl_234 br_234 wl_97 vdd gnd cell_6t
Xbit_r98_c234 bl_234 br_234 wl_98 vdd gnd cell_6t
Xbit_r99_c234 bl_234 br_234 wl_99 vdd gnd cell_6t
Xbit_r100_c234 bl_234 br_234 wl_100 vdd gnd cell_6t
Xbit_r101_c234 bl_234 br_234 wl_101 vdd gnd cell_6t
Xbit_r102_c234 bl_234 br_234 wl_102 vdd gnd cell_6t
Xbit_r103_c234 bl_234 br_234 wl_103 vdd gnd cell_6t
Xbit_r104_c234 bl_234 br_234 wl_104 vdd gnd cell_6t
Xbit_r105_c234 bl_234 br_234 wl_105 vdd gnd cell_6t
Xbit_r106_c234 bl_234 br_234 wl_106 vdd gnd cell_6t
Xbit_r107_c234 bl_234 br_234 wl_107 vdd gnd cell_6t
Xbit_r108_c234 bl_234 br_234 wl_108 vdd gnd cell_6t
Xbit_r109_c234 bl_234 br_234 wl_109 vdd gnd cell_6t
Xbit_r110_c234 bl_234 br_234 wl_110 vdd gnd cell_6t
Xbit_r111_c234 bl_234 br_234 wl_111 vdd gnd cell_6t
Xbit_r112_c234 bl_234 br_234 wl_112 vdd gnd cell_6t
Xbit_r113_c234 bl_234 br_234 wl_113 vdd gnd cell_6t
Xbit_r114_c234 bl_234 br_234 wl_114 vdd gnd cell_6t
Xbit_r115_c234 bl_234 br_234 wl_115 vdd gnd cell_6t
Xbit_r116_c234 bl_234 br_234 wl_116 vdd gnd cell_6t
Xbit_r117_c234 bl_234 br_234 wl_117 vdd gnd cell_6t
Xbit_r118_c234 bl_234 br_234 wl_118 vdd gnd cell_6t
Xbit_r119_c234 bl_234 br_234 wl_119 vdd gnd cell_6t
Xbit_r120_c234 bl_234 br_234 wl_120 vdd gnd cell_6t
Xbit_r121_c234 bl_234 br_234 wl_121 vdd gnd cell_6t
Xbit_r122_c234 bl_234 br_234 wl_122 vdd gnd cell_6t
Xbit_r123_c234 bl_234 br_234 wl_123 vdd gnd cell_6t
Xbit_r124_c234 bl_234 br_234 wl_124 vdd gnd cell_6t
Xbit_r125_c234 bl_234 br_234 wl_125 vdd gnd cell_6t
Xbit_r126_c234 bl_234 br_234 wl_126 vdd gnd cell_6t
Xbit_r127_c234 bl_234 br_234 wl_127 vdd gnd cell_6t
Xbit_r128_c234 bl_234 br_234 wl_128 vdd gnd cell_6t
Xbit_r129_c234 bl_234 br_234 wl_129 vdd gnd cell_6t
Xbit_r130_c234 bl_234 br_234 wl_130 vdd gnd cell_6t
Xbit_r131_c234 bl_234 br_234 wl_131 vdd gnd cell_6t
Xbit_r132_c234 bl_234 br_234 wl_132 vdd gnd cell_6t
Xbit_r133_c234 bl_234 br_234 wl_133 vdd gnd cell_6t
Xbit_r134_c234 bl_234 br_234 wl_134 vdd gnd cell_6t
Xbit_r135_c234 bl_234 br_234 wl_135 vdd gnd cell_6t
Xbit_r136_c234 bl_234 br_234 wl_136 vdd gnd cell_6t
Xbit_r137_c234 bl_234 br_234 wl_137 vdd gnd cell_6t
Xbit_r138_c234 bl_234 br_234 wl_138 vdd gnd cell_6t
Xbit_r139_c234 bl_234 br_234 wl_139 vdd gnd cell_6t
Xbit_r140_c234 bl_234 br_234 wl_140 vdd gnd cell_6t
Xbit_r141_c234 bl_234 br_234 wl_141 vdd gnd cell_6t
Xbit_r142_c234 bl_234 br_234 wl_142 vdd gnd cell_6t
Xbit_r143_c234 bl_234 br_234 wl_143 vdd gnd cell_6t
Xbit_r144_c234 bl_234 br_234 wl_144 vdd gnd cell_6t
Xbit_r145_c234 bl_234 br_234 wl_145 vdd gnd cell_6t
Xbit_r146_c234 bl_234 br_234 wl_146 vdd gnd cell_6t
Xbit_r147_c234 bl_234 br_234 wl_147 vdd gnd cell_6t
Xbit_r148_c234 bl_234 br_234 wl_148 vdd gnd cell_6t
Xbit_r149_c234 bl_234 br_234 wl_149 vdd gnd cell_6t
Xbit_r150_c234 bl_234 br_234 wl_150 vdd gnd cell_6t
Xbit_r151_c234 bl_234 br_234 wl_151 vdd gnd cell_6t
Xbit_r152_c234 bl_234 br_234 wl_152 vdd gnd cell_6t
Xbit_r153_c234 bl_234 br_234 wl_153 vdd gnd cell_6t
Xbit_r154_c234 bl_234 br_234 wl_154 vdd gnd cell_6t
Xbit_r155_c234 bl_234 br_234 wl_155 vdd gnd cell_6t
Xbit_r156_c234 bl_234 br_234 wl_156 vdd gnd cell_6t
Xbit_r157_c234 bl_234 br_234 wl_157 vdd gnd cell_6t
Xbit_r158_c234 bl_234 br_234 wl_158 vdd gnd cell_6t
Xbit_r159_c234 bl_234 br_234 wl_159 vdd gnd cell_6t
Xbit_r160_c234 bl_234 br_234 wl_160 vdd gnd cell_6t
Xbit_r161_c234 bl_234 br_234 wl_161 vdd gnd cell_6t
Xbit_r162_c234 bl_234 br_234 wl_162 vdd gnd cell_6t
Xbit_r163_c234 bl_234 br_234 wl_163 vdd gnd cell_6t
Xbit_r164_c234 bl_234 br_234 wl_164 vdd gnd cell_6t
Xbit_r165_c234 bl_234 br_234 wl_165 vdd gnd cell_6t
Xbit_r166_c234 bl_234 br_234 wl_166 vdd gnd cell_6t
Xbit_r167_c234 bl_234 br_234 wl_167 vdd gnd cell_6t
Xbit_r168_c234 bl_234 br_234 wl_168 vdd gnd cell_6t
Xbit_r169_c234 bl_234 br_234 wl_169 vdd gnd cell_6t
Xbit_r170_c234 bl_234 br_234 wl_170 vdd gnd cell_6t
Xbit_r171_c234 bl_234 br_234 wl_171 vdd gnd cell_6t
Xbit_r172_c234 bl_234 br_234 wl_172 vdd gnd cell_6t
Xbit_r173_c234 bl_234 br_234 wl_173 vdd gnd cell_6t
Xbit_r174_c234 bl_234 br_234 wl_174 vdd gnd cell_6t
Xbit_r175_c234 bl_234 br_234 wl_175 vdd gnd cell_6t
Xbit_r176_c234 bl_234 br_234 wl_176 vdd gnd cell_6t
Xbit_r177_c234 bl_234 br_234 wl_177 vdd gnd cell_6t
Xbit_r178_c234 bl_234 br_234 wl_178 vdd gnd cell_6t
Xbit_r179_c234 bl_234 br_234 wl_179 vdd gnd cell_6t
Xbit_r180_c234 bl_234 br_234 wl_180 vdd gnd cell_6t
Xbit_r181_c234 bl_234 br_234 wl_181 vdd gnd cell_6t
Xbit_r182_c234 bl_234 br_234 wl_182 vdd gnd cell_6t
Xbit_r183_c234 bl_234 br_234 wl_183 vdd gnd cell_6t
Xbit_r184_c234 bl_234 br_234 wl_184 vdd gnd cell_6t
Xbit_r185_c234 bl_234 br_234 wl_185 vdd gnd cell_6t
Xbit_r186_c234 bl_234 br_234 wl_186 vdd gnd cell_6t
Xbit_r187_c234 bl_234 br_234 wl_187 vdd gnd cell_6t
Xbit_r188_c234 bl_234 br_234 wl_188 vdd gnd cell_6t
Xbit_r189_c234 bl_234 br_234 wl_189 vdd gnd cell_6t
Xbit_r190_c234 bl_234 br_234 wl_190 vdd gnd cell_6t
Xbit_r191_c234 bl_234 br_234 wl_191 vdd gnd cell_6t
Xbit_r192_c234 bl_234 br_234 wl_192 vdd gnd cell_6t
Xbit_r193_c234 bl_234 br_234 wl_193 vdd gnd cell_6t
Xbit_r194_c234 bl_234 br_234 wl_194 vdd gnd cell_6t
Xbit_r195_c234 bl_234 br_234 wl_195 vdd gnd cell_6t
Xbit_r196_c234 bl_234 br_234 wl_196 vdd gnd cell_6t
Xbit_r197_c234 bl_234 br_234 wl_197 vdd gnd cell_6t
Xbit_r198_c234 bl_234 br_234 wl_198 vdd gnd cell_6t
Xbit_r199_c234 bl_234 br_234 wl_199 vdd gnd cell_6t
Xbit_r200_c234 bl_234 br_234 wl_200 vdd gnd cell_6t
Xbit_r201_c234 bl_234 br_234 wl_201 vdd gnd cell_6t
Xbit_r202_c234 bl_234 br_234 wl_202 vdd gnd cell_6t
Xbit_r203_c234 bl_234 br_234 wl_203 vdd gnd cell_6t
Xbit_r204_c234 bl_234 br_234 wl_204 vdd gnd cell_6t
Xbit_r205_c234 bl_234 br_234 wl_205 vdd gnd cell_6t
Xbit_r206_c234 bl_234 br_234 wl_206 vdd gnd cell_6t
Xbit_r207_c234 bl_234 br_234 wl_207 vdd gnd cell_6t
Xbit_r208_c234 bl_234 br_234 wl_208 vdd gnd cell_6t
Xbit_r209_c234 bl_234 br_234 wl_209 vdd gnd cell_6t
Xbit_r210_c234 bl_234 br_234 wl_210 vdd gnd cell_6t
Xbit_r211_c234 bl_234 br_234 wl_211 vdd gnd cell_6t
Xbit_r212_c234 bl_234 br_234 wl_212 vdd gnd cell_6t
Xbit_r213_c234 bl_234 br_234 wl_213 vdd gnd cell_6t
Xbit_r214_c234 bl_234 br_234 wl_214 vdd gnd cell_6t
Xbit_r215_c234 bl_234 br_234 wl_215 vdd gnd cell_6t
Xbit_r216_c234 bl_234 br_234 wl_216 vdd gnd cell_6t
Xbit_r217_c234 bl_234 br_234 wl_217 vdd gnd cell_6t
Xbit_r218_c234 bl_234 br_234 wl_218 vdd gnd cell_6t
Xbit_r219_c234 bl_234 br_234 wl_219 vdd gnd cell_6t
Xbit_r220_c234 bl_234 br_234 wl_220 vdd gnd cell_6t
Xbit_r221_c234 bl_234 br_234 wl_221 vdd gnd cell_6t
Xbit_r222_c234 bl_234 br_234 wl_222 vdd gnd cell_6t
Xbit_r223_c234 bl_234 br_234 wl_223 vdd gnd cell_6t
Xbit_r224_c234 bl_234 br_234 wl_224 vdd gnd cell_6t
Xbit_r225_c234 bl_234 br_234 wl_225 vdd gnd cell_6t
Xbit_r226_c234 bl_234 br_234 wl_226 vdd gnd cell_6t
Xbit_r227_c234 bl_234 br_234 wl_227 vdd gnd cell_6t
Xbit_r228_c234 bl_234 br_234 wl_228 vdd gnd cell_6t
Xbit_r229_c234 bl_234 br_234 wl_229 vdd gnd cell_6t
Xbit_r230_c234 bl_234 br_234 wl_230 vdd gnd cell_6t
Xbit_r231_c234 bl_234 br_234 wl_231 vdd gnd cell_6t
Xbit_r232_c234 bl_234 br_234 wl_232 vdd gnd cell_6t
Xbit_r233_c234 bl_234 br_234 wl_233 vdd gnd cell_6t
Xbit_r234_c234 bl_234 br_234 wl_234 vdd gnd cell_6t
Xbit_r235_c234 bl_234 br_234 wl_235 vdd gnd cell_6t
Xbit_r236_c234 bl_234 br_234 wl_236 vdd gnd cell_6t
Xbit_r237_c234 bl_234 br_234 wl_237 vdd gnd cell_6t
Xbit_r238_c234 bl_234 br_234 wl_238 vdd gnd cell_6t
Xbit_r239_c234 bl_234 br_234 wl_239 vdd gnd cell_6t
Xbit_r240_c234 bl_234 br_234 wl_240 vdd gnd cell_6t
Xbit_r241_c234 bl_234 br_234 wl_241 vdd gnd cell_6t
Xbit_r242_c234 bl_234 br_234 wl_242 vdd gnd cell_6t
Xbit_r243_c234 bl_234 br_234 wl_243 vdd gnd cell_6t
Xbit_r244_c234 bl_234 br_234 wl_244 vdd gnd cell_6t
Xbit_r245_c234 bl_234 br_234 wl_245 vdd gnd cell_6t
Xbit_r246_c234 bl_234 br_234 wl_246 vdd gnd cell_6t
Xbit_r247_c234 bl_234 br_234 wl_247 vdd gnd cell_6t
Xbit_r248_c234 bl_234 br_234 wl_248 vdd gnd cell_6t
Xbit_r249_c234 bl_234 br_234 wl_249 vdd gnd cell_6t
Xbit_r250_c234 bl_234 br_234 wl_250 vdd gnd cell_6t
Xbit_r251_c234 bl_234 br_234 wl_251 vdd gnd cell_6t
Xbit_r252_c234 bl_234 br_234 wl_252 vdd gnd cell_6t
Xbit_r253_c234 bl_234 br_234 wl_253 vdd gnd cell_6t
Xbit_r254_c234 bl_234 br_234 wl_254 vdd gnd cell_6t
Xbit_r255_c234 bl_234 br_234 wl_255 vdd gnd cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd cell_6t
Xbit_r1_c235 bl_235 br_235 wl_1 vdd gnd cell_6t
Xbit_r2_c235 bl_235 br_235 wl_2 vdd gnd cell_6t
Xbit_r3_c235 bl_235 br_235 wl_3 vdd gnd cell_6t
Xbit_r4_c235 bl_235 br_235 wl_4 vdd gnd cell_6t
Xbit_r5_c235 bl_235 br_235 wl_5 vdd gnd cell_6t
Xbit_r6_c235 bl_235 br_235 wl_6 vdd gnd cell_6t
Xbit_r7_c235 bl_235 br_235 wl_7 vdd gnd cell_6t
Xbit_r8_c235 bl_235 br_235 wl_8 vdd gnd cell_6t
Xbit_r9_c235 bl_235 br_235 wl_9 vdd gnd cell_6t
Xbit_r10_c235 bl_235 br_235 wl_10 vdd gnd cell_6t
Xbit_r11_c235 bl_235 br_235 wl_11 vdd gnd cell_6t
Xbit_r12_c235 bl_235 br_235 wl_12 vdd gnd cell_6t
Xbit_r13_c235 bl_235 br_235 wl_13 vdd gnd cell_6t
Xbit_r14_c235 bl_235 br_235 wl_14 vdd gnd cell_6t
Xbit_r15_c235 bl_235 br_235 wl_15 vdd gnd cell_6t
Xbit_r16_c235 bl_235 br_235 wl_16 vdd gnd cell_6t
Xbit_r17_c235 bl_235 br_235 wl_17 vdd gnd cell_6t
Xbit_r18_c235 bl_235 br_235 wl_18 vdd gnd cell_6t
Xbit_r19_c235 bl_235 br_235 wl_19 vdd gnd cell_6t
Xbit_r20_c235 bl_235 br_235 wl_20 vdd gnd cell_6t
Xbit_r21_c235 bl_235 br_235 wl_21 vdd gnd cell_6t
Xbit_r22_c235 bl_235 br_235 wl_22 vdd gnd cell_6t
Xbit_r23_c235 bl_235 br_235 wl_23 vdd gnd cell_6t
Xbit_r24_c235 bl_235 br_235 wl_24 vdd gnd cell_6t
Xbit_r25_c235 bl_235 br_235 wl_25 vdd gnd cell_6t
Xbit_r26_c235 bl_235 br_235 wl_26 vdd gnd cell_6t
Xbit_r27_c235 bl_235 br_235 wl_27 vdd gnd cell_6t
Xbit_r28_c235 bl_235 br_235 wl_28 vdd gnd cell_6t
Xbit_r29_c235 bl_235 br_235 wl_29 vdd gnd cell_6t
Xbit_r30_c235 bl_235 br_235 wl_30 vdd gnd cell_6t
Xbit_r31_c235 bl_235 br_235 wl_31 vdd gnd cell_6t
Xbit_r32_c235 bl_235 br_235 wl_32 vdd gnd cell_6t
Xbit_r33_c235 bl_235 br_235 wl_33 vdd gnd cell_6t
Xbit_r34_c235 bl_235 br_235 wl_34 vdd gnd cell_6t
Xbit_r35_c235 bl_235 br_235 wl_35 vdd gnd cell_6t
Xbit_r36_c235 bl_235 br_235 wl_36 vdd gnd cell_6t
Xbit_r37_c235 bl_235 br_235 wl_37 vdd gnd cell_6t
Xbit_r38_c235 bl_235 br_235 wl_38 vdd gnd cell_6t
Xbit_r39_c235 bl_235 br_235 wl_39 vdd gnd cell_6t
Xbit_r40_c235 bl_235 br_235 wl_40 vdd gnd cell_6t
Xbit_r41_c235 bl_235 br_235 wl_41 vdd gnd cell_6t
Xbit_r42_c235 bl_235 br_235 wl_42 vdd gnd cell_6t
Xbit_r43_c235 bl_235 br_235 wl_43 vdd gnd cell_6t
Xbit_r44_c235 bl_235 br_235 wl_44 vdd gnd cell_6t
Xbit_r45_c235 bl_235 br_235 wl_45 vdd gnd cell_6t
Xbit_r46_c235 bl_235 br_235 wl_46 vdd gnd cell_6t
Xbit_r47_c235 bl_235 br_235 wl_47 vdd gnd cell_6t
Xbit_r48_c235 bl_235 br_235 wl_48 vdd gnd cell_6t
Xbit_r49_c235 bl_235 br_235 wl_49 vdd gnd cell_6t
Xbit_r50_c235 bl_235 br_235 wl_50 vdd gnd cell_6t
Xbit_r51_c235 bl_235 br_235 wl_51 vdd gnd cell_6t
Xbit_r52_c235 bl_235 br_235 wl_52 vdd gnd cell_6t
Xbit_r53_c235 bl_235 br_235 wl_53 vdd gnd cell_6t
Xbit_r54_c235 bl_235 br_235 wl_54 vdd gnd cell_6t
Xbit_r55_c235 bl_235 br_235 wl_55 vdd gnd cell_6t
Xbit_r56_c235 bl_235 br_235 wl_56 vdd gnd cell_6t
Xbit_r57_c235 bl_235 br_235 wl_57 vdd gnd cell_6t
Xbit_r58_c235 bl_235 br_235 wl_58 vdd gnd cell_6t
Xbit_r59_c235 bl_235 br_235 wl_59 vdd gnd cell_6t
Xbit_r60_c235 bl_235 br_235 wl_60 vdd gnd cell_6t
Xbit_r61_c235 bl_235 br_235 wl_61 vdd gnd cell_6t
Xbit_r62_c235 bl_235 br_235 wl_62 vdd gnd cell_6t
Xbit_r63_c235 bl_235 br_235 wl_63 vdd gnd cell_6t
Xbit_r64_c235 bl_235 br_235 wl_64 vdd gnd cell_6t
Xbit_r65_c235 bl_235 br_235 wl_65 vdd gnd cell_6t
Xbit_r66_c235 bl_235 br_235 wl_66 vdd gnd cell_6t
Xbit_r67_c235 bl_235 br_235 wl_67 vdd gnd cell_6t
Xbit_r68_c235 bl_235 br_235 wl_68 vdd gnd cell_6t
Xbit_r69_c235 bl_235 br_235 wl_69 vdd gnd cell_6t
Xbit_r70_c235 bl_235 br_235 wl_70 vdd gnd cell_6t
Xbit_r71_c235 bl_235 br_235 wl_71 vdd gnd cell_6t
Xbit_r72_c235 bl_235 br_235 wl_72 vdd gnd cell_6t
Xbit_r73_c235 bl_235 br_235 wl_73 vdd gnd cell_6t
Xbit_r74_c235 bl_235 br_235 wl_74 vdd gnd cell_6t
Xbit_r75_c235 bl_235 br_235 wl_75 vdd gnd cell_6t
Xbit_r76_c235 bl_235 br_235 wl_76 vdd gnd cell_6t
Xbit_r77_c235 bl_235 br_235 wl_77 vdd gnd cell_6t
Xbit_r78_c235 bl_235 br_235 wl_78 vdd gnd cell_6t
Xbit_r79_c235 bl_235 br_235 wl_79 vdd gnd cell_6t
Xbit_r80_c235 bl_235 br_235 wl_80 vdd gnd cell_6t
Xbit_r81_c235 bl_235 br_235 wl_81 vdd gnd cell_6t
Xbit_r82_c235 bl_235 br_235 wl_82 vdd gnd cell_6t
Xbit_r83_c235 bl_235 br_235 wl_83 vdd gnd cell_6t
Xbit_r84_c235 bl_235 br_235 wl_84 vdd gnd cell_6t
Xbit_r85_c235 bl_235 br_235 wl_85 vdd gnd cell_6t
Xbit_r86_c235 bl_235 br_235 wl_86 vdd gnd cell_6t
Xbit_r87_c235 bl_235 br_235 wl_87 vdd gnd cell_6t
Xbit_r88_c235 bl_235 br_235 wl_88 vdd gnd cell_6t
Xbit_r89_c235 bl_235 br_235 wl_89 vdd gnd cell_6t
Xbit_r90_c235 bl_235 br_235 wl_90 vdd gnd cell_6t
Xbit_r91_c235 bl_235 br_235 wl_91 vdd gnd cell_6t
Xbit_r92_c235 bl_235 br_235 wl_92 vdd gnd cell_6t
Xbit_r93_c235 bl_235 br_235 wl_93 vdd gnd cell_6t
Xbit_r94_c235 bl_235 br_235 wl_94 vdd gnd cell_6t
Xbit_r95_c235 bl_235 br_235 wl_95 vdd gnd cell_6t
Xbit_r96_c235 bl_235 br_235 wl_96 vdd gnd cell_6t
Xbit_r97_c235 bl_235 br_235 wl_97 vdd gnd cell_6t
Xbit_r98_c235 bl_235 br_235 wl_98 vdd gnd cell_6t
Xbit_r99_c235 bl_235 br_235 wl_99 vdd gnd cell_6t
Xbit_r100_c235 bl_235 br_235 wl_100 vdd gnd cell_6t
Xbit_r101_c235 bl_235 br_235 wl_101 vdd gnd cell_6t
Xbit_r102_c235 bl_235 br_235 wl_102 vdd gnd cell_6t
Xbit_r103_c235 bl_235 br_235 wl_103 vdd gnd cell_6t
Xbit_r104_c235 bl_235 br_235 wl_104 vdd gnd cell_6t
Xbit_r105_c235 bl_235 br_235 wl_105 vdd gnd cell_6t
Xbit_r106_c235 bl_235 br_235 wl_106 vdd gnd cell_6t
Xbit_r107_c235 bl_235 br_235 wl_107 vdd gnd cell_6t
Xbit_r108_c235 bl_235 br_235 wl_108 vdd gnd cell_6t
Xbit_r109_c235 bl_235 br_235 wl_109 vdd gnd cell_6t
Xbit_r110_c235 bl_235 br_235 wl_110 vdd gnd cell_6t
Xbit_r111_c235 bl_235 br_235 wl_111 vdd gnd cell_6t
Xbit_r112_c235 bl_235 br_235 wl_112 vdd gnd cell_6t
Xbit_r113_c235 bl_235 br_235 wl_113 vdd gnd cell_6t
Xbit_r114_c235 bl_235 br_235 wl_114 vdd gnd cell_6t
Xbit_r115_c235 bl_235 br_235 wl_115 vdd gnd cell_6t
Xbit_r116_c235 bl_235 br_235 wl_116 vdd gnd cell_6t
Xbit_r117_c235 bl_235 br_235 wl_117 vdd gnd cell_6t
Xbit_r118_c235 bl_235 br_235 wl_118 vdd gnd cell_6t
Xbit_r119_c235 bl_235 br_235 wl_119 vdd gnd cell_6t
Xbit_r120_c235 bl_235 br_235 wl_120 vdd gnd cell_6t
Xbit_r121_c235 bl_235 br_235 wl_121 vdd gnd cell_6t
Xbit_r122_c235 bl_235 br_235 wl_122 vdd gnd cell_6t
Xbit_r123_c235 bl_235 br_235 wl_123 vdd gnd cell_6t
Xbit_r124_c235 bl_235 br_235 wl_124 vdd gnd cell_6t
Xbit_r125_c235 bl_235 br_235 wl_125 vdd gnd cell_6t
Xbit_r126_c235 bl_235 br_235 wl_126 vdd gnd cell_6t
Xbit_r127_c235 bl_235 br_235 wl_127 vdd gnd cell_6t
Xbit_r128_c235 bl_235 br_235 wl_128 vdd gnd cell_6t
Xbit_r129_c235 bl_235 br_235 wl_129 vdd gnd cell_6t
Xbit_r130_c235 bl_235 br_235 wl_130 vdd gnd cell_6t
Xbit_r131_c235 bl_235 br_235 wl_131 vdd gnd cell_6t
Xbit_r132_c235 bl_235 br_235 wl_132 vdd gnd cell_6t
Xbit_r133_c235 bl_235 br_235 wl_133 vdd gnd cell_6t
Xbit_r134_c235 bl_235 br_235 wl_134 vdd gnd cell_6t
Xbit_r135_c235 bl_235 br_235 wl_135 vdd gnd cell_6t
Xbit_r136_c235 bl_235 br_235 wl_136 vdd gnd cell_6t
Xbit_r137_c235 bl_235 br_235 wl_137 vdd gnd cell_6t
Xbit_r138_c235 bl_235 br_235 wl_138 vdd gnd cell_6t
Xbit_r139_c235 bl_235 br_235 wl_139 vdd gnd cell_6t
Xbit_r140_c235 bl_235 br_235 wl_140 vdd gnd cell_6t
Xbit_r141_c235 bl_235 br_235 wl_141 vdd gnd cell_6t
Xbit_r142_c235 bl_235 br_235 wl_142 vdd gnd cell_6t
Xbit_r143_c235 bl_235 br_235 wl_143 vdd gnd cell_6t
Xbit_r144_c235 bl_235 br_235 wl_144 vdd gnd cell_6t
Xbit_r145_c235 bl_235 br_235 wl_145 vdd gnd cell_6t
Xbit_r146_c235 bl_235 br_235 wl_146 vdd gnd cell_6t
Xbit_r147_c235 bl_235 br_235 wl_147 vdd gnd cell_6t
Xbit_r148_c235 bl_235 br_235 wl_148 vdd gnd cell_6t
Xbit_r149_c235 bl_235 br_235 wl_149 vdd gnd cell_6t
Xbit_r150_c235 bl_235 br_235 wl_150 vdd gnd cell_6t
Xbit_r151_c235 bl_235 br_235 wl_151 vdd gnd cell_6t
Xbit_r152_c235 bl_235 br_235 wl_152 vdd gnd cell_6t
Xbit_r153_c235 bl_235 br_235 wl_153 vdd gnd cell_6t
Xbit_r154_c235 bl_235 br_235 wl_154 vdd gnd cell_6t
Xbit_r155_c235 bl_235 br_235 wl_155 vdd gnd cell_6t
Xbit_r156_c235 bl_235 br_235 wl_156 vdd gnd cell_6t
Xbit_r157_c235 bl_235 br_235 wl_157 vdd gnd cell_6t
Xbit_r158_c235 bl_235 br_235 wl_158 vdd gnd cell_6t
Xbit_r159_c235 bl_235 br_235 wl_159 vdd gnd cell_6t
Xbit_r160_c235 bl_235 br_235 wl_160 vdd gnd cell_6t
Xbit_r161_c235 bl_235 br_235 wl_161 vdd gnd cell_6t
Xbit_r162_c235 bl_235 br_235 wl_162 vdd gnd cell_6t
Xbit_r163_c235 bl_235 br_235 wl_163 vdd gnd cell_6t
Xbit_r164_c235 bl_235 br_235 wl_164 vdd gnd cell_6t
Xbit_r165_c235 bl_235 br_235 wl_165 vdd gnd cell_6t
Xbit_r166_c235 bl_235 br_235 wl_166 vdd gnd cell_6t
Xbit_r167_c235 bl_235 br_235 wl_167 vdd gnd cell_6t
Xbit_r168_c235 bl_235 br_235 wl_168 vdd gnd cell_6t
Xbit_r169_c235 bl_235 br_235 wl_169 vdd gnd cell_6t
Xbit_r170_c235 bl_235 br_235 wl_170 vdd gnd cell_6t
Xbit_r171_c235 bl_235 br_235 wl_171 vdd gnd cell_6t
Xbit_r172_c235 bl_235 br_235 wl_172 vdd gnd cell_6t
Xbit_r173_c235 bl_235 br_235 wl_173 vdd gnd cell_6t
Xbit_r174_c235 bl_235 br_235 wl_174 vdd gnd cell_6t
Xbit_r175_c235 bl_235 br_235 wl_175 vdd gnd cell_6t
Xbit_r176_c235 bl_235 br_235 wl_176 vdd gnd cell_6t
Xbit_r177_c235 bl_235 br_235 wl_177 vdd gnd cell_6t
Xbit_r178_c235 bl_235 br_235 wl_178 vdd gnd cell_6t
Xbit_r179_c235 bl_235 br_235 wl_179 vdd gnd cell_6t
Xbit_r180_c235 bl_235 br_235 wl_180 vdd gnd cell_6t
Xbit_r181_c235 bl_235 br_235 wl_181 vdd gnd cell_6t
Xbit_r182_c235 bl_235 br_235 wl_182 vdd gnd cell_6t
Xbit_r183_c235 bl_235 br_235 wl_183 vdd gnd cell_6t
Xbit_r184_c235 bl_235 br_235 wl_184 vdd gnd cell_6t
Xbit_r185_c235 bl_235 br_235 wl_185 vdd gnd cell_6t
Xbit_r186_c235 bl_235 br_235 wl_186 vdd gnd cell_6t
Xbit_r187_c235 bl_235 br_235 wl_187 vdd gnd cell_6t
Xbit_r188_c235 bl_235 br_235 wl_188 vdd gnd cell_6t
Xbit_r189_c235 bl_235 br_235 wl_189 vdd gnd cell_6t
Xbit_r190_c235 bl_235 br_235 wl_190 vdd gnd cell_6t
Xbit_r191_c235 bl_235 br_235 wl_191 vdd gnd cell_6t
Xbit_r192_c235 bl_235 br_235 wl_192 vdd gnd cell_6t
Xbit_r193_c235 bl_235 br_235 wl_193 vdd gnd cell_6t
Xbit_r194_c235 bl_235 br_235 wl_194 vdd gnd cell_6t
Xbit_r195_c235 bl_235 br_235 wl_195 vdd gnd cell_6t
Xbit_r196_c235 bl_235 br_235 wl_196 vdd gnd cell_6t
Xbit_r197_c235 bl_235 br_235 wl_197 vdd gnd cell_6t
Xbit_r198_c235 bl_235 br_235 wl_198 vdd gnd cell_6t
Xbit_r199_c235 bl_235 br_235 wl_199 vdd gnd cell_6t
Xbit_r200_c235 bl_235 br_235 wl_200 vdd gnd cell_6t
Xbit_r201_c235 bl_235 br_235 wl_201 vdd gnd cell_6t
Xbit_r202_c235 bl_235 br_235 wl_202 vdd gnd cell_6t
Xbit_r203_c235 bl_235 br_235 wl_203 vdd gnd cell_6t
Xbit_r204_c235 bl_235 br_235 wl_204 vdd gnd cell_6t
Xbit_r205_c235 bl_235 br_235 wl_205 vdd gnd cell_6t
Xbit_r206_c235 bl_235 br_235 wl_206 vdd gnd cell_6t
Xbit_r207_c235 bl_235 br_235 wl_207 vdd gnd cell_6t
Xbit_r208_c235 bl_235 br_235 wl_208 vdd gnd cell_6t
Xbit_r209_c235 bl_235 br_235 wl_209 vdd gnd cell_6t
Xbit_r210_c235 bl_235 br_235 wl_210 vdd gnd cell_6t
Xbit_r211_c235 bl_235 br_235 wl_211 vdd gnd cell_6t
Xbit_r212_c235 bl_235 br_235 wl_212 vdd gnd cell_6t
Xbit_r213_c235 bl_235 br_235 wl_213 vdd gnd cell_6t
Xbit_r214_c235 bl_235 br_235 wl_214 vdd gnd cell_6t
Xbit_r215_c235 bl_235 br_235 wl_215 vdd gnd cell_6t
Xbit_r216_c235 bl_235 br_235 wl_216 vdd gnd cell_6t
Xbit_r217_c235 bl_235 br_235 wl_217 vdd gnd cell_6t
Xbit_r218_c235 bl_235 br_235 wl_218 vdd gnd cell_6t
Xbit_r219_c235 bl_235 br_235 wl_219 vdd gnd cell_6t
Xbit_r220_c235 bl_235 br_235 wl_220 vdd gnd cell_6t
Xbit_r221_c235 bl_235 br_235 wl_221 vdd gnd cell_6t
Xbit_r222_c235 bl_235 br_235 wl_222 vdd gnd cell_6t
Xbit_r223_c235 bl_235 br_235 wl_223 vdd gnd cell_6t
Xbit_r224_c235 bl_235 br_235 wl_224 vdd gnd cell_6t
Xbit_r225_c235 bl_235 br_235 wl_225 vdd gnd cell_6t
Xbit_r226_c235 bl_235 br_235 wl_226 vdd gnd cell_6t
Xbit_r227_c235 bl_235 br_235 wl_227 vdd gnd cell_6t
Xbit_r228_c235 bl_235 br_235 wl_228 vdd gnd cell_6t
Xbit_r229_c235 bl_235 br_235 wl_229 vdd gnd cell_6t
Xbit_r230_c235 bl_235 br_235 wl_230 vdd gnd cell_6t
Xbit_r231_c235 bl_235 br_235 wl_231 vdd gnd cell_6t
Xbit_r232_c235 bl_235 br_235 wl_232 vdd gnd cell_6t
Xbit_r233_c235 bl_235 br_235 wl_233 vdd gnd cell_6t
Xbit_r234_c235 bl_235 br_235 wl_234 vdd gnd cell_6t
Xbit_r235_c235 bl_235 br_235 wl_235 vdd gnd cell_6t
Xbit_r236_c235 bl_235 br_235 wl_236 vdd gnd cell_6t
Xbit_r237_c235 bl_235 br_235 wl_237 vdd gnd cell_6t
Xbit_r238_c235 bl_235 br_235 wl_238 vdd gnd cell_6t
Xbit_r239_c235 bl_235 br_235 wl_239 vdd gnd cell_6t
Xbit_r240_c235 bl_235 br_235 wl_240 vdd gnd cell_6t
Xbit_r241_c235 bl_235 br_235 wl_241 vdd gnd cell_6t
Xbit_r242_c235 bl_235 br_235 wl_242 vdd gnd cell_6t
Xbit_r243_c235 bl_235 br_235 wl_243 vdd gnd cell_6t
Xbit_r244_c235 bl_235 br_235 wl_244 vdd gnd cell_6t
Xbit_r245_c235 bl_235 br_235 wl_245 vdd gnd cell_6t
Xbit_r246_c235 bl_235 br_235 wl_246 vdd gnd cell_6t
Xbit_r247_c235 bl_235 br_235 wl_247 vdd gnd cell_6t
Xbit_r248_c235 bl_235 br_235 wl_248 vdd gnd cell_6t
Xbit_r249_c235 bl_235 br_235 wl_249 vdd gnd cell_6t
Xbit_r250_c235 bl_235 br_235 wl_250 vdd gnd cell_6t
Xbit_r251_c235 bl_235 br_235 wl_251 vdd gnd cell_6t
Xbit_r252_c235 bl_235 br_235 wl_252 vdd gnd cell_6t
Xbit_r253_c235 bl_235 br_235 wl_253 vdd gnd cell_6t
Xbit_r254_c235 bl_235 br_235 wl_254 vdd gnd cell_6t
Xbit_r255_c235 bl_235 br_235 wl_255 vdd gnd cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd cell_6t
Xbit_r1_c236 bl_236 br_236 wl_1 vdd gnd cell_6t
Xbit_r2_c236 bl_236 br_236 wl_2 vdd gnd cell_6t
Xbit_r3_c236 bl_236 br_236 wl_3 vdd gnd cell_6t
Xbit_r4_c236 bl_236 br_236 wl_4 vdd gnd cell_6t
Xbit_r5_c236 bl_236 br_236 wl_5 vdd gnd cell_6t
Xbit_r6_c236 bl_236 br_236 wl_6 vdd gnd cell_6t
Xbit_r7_c236 bl_236 br_236 wl_7 vdd gnd cell_6t
Xbit_r8_c236 bl_236 br_236 wl_8 vdd gnd cell_6t
Xbit_r9_c236 bl_236 br_236 wl_9 vdd gnd cell_6t
Xbit_r10_c236 bl_236 br_236 wl_10 vdd gnd cell_6t
Xbit_r11_c236 bl_236 br_236 wl_11 vdd gnd cell_6t
Xbit_r12_c236 bl_236 br_236 wl_12 vdd gnd cell_6t
Xbit_r13_c236 bl_236 br_236 wl_13 vdd gnd cell_6t
Xbit_r14_c236 bl_236 br_236 wl_14 vdd gnd cell_6t
Xbit_r15_c236 bl_236 br_236 wl_15 vdd gnd cell_6t
Xbit_r16_c236 bl_236 br_236 wl_16 vdd gnd cell_6t
Xbit_r17_c236 bl_236 br_236 wl_17 vdd gnd cell_6t
Xbit_r18_c236 bl_236 br_236 wl_18 vdd gnd cell_6t
Xbit_r19_c236 bl_236 br_236 wl_19 vdd gnd cell_6t
Xbit_r20_c236 bl_236 br_236 wl_20 vdd gnd cell_6t
Xbit_r21_c236 bl_236 br_236 wl_21 vdd gnd cell_6t
Xbit_r22_c236 bl_236 br_236 wl_22 vdd gnd cell_6t
Xbit_r23_c236 bl_236 br_236 wl_23 vdd gnd cell_6t
Xbit_r24_c236 bl_236 br_236 wl_24 vdd gnd cell_6t
Xbit_r25_c236 bl_236 br_236 wl_25 vdd gnd cell_6t
Xbit_r26_c236 bl_236 br_236 wl_26 vdd gnd cell_6t
Xbit_r27_c236 bl_236 br_236 wl_27 vdd gnd cell_6t
Xbit_r28_c236 bl_236 br_236 wl_28 vdd gnd cell_6t
Xbit_r29_c236 bl_236 br_236 wl_29 vdd gnd cell_6t
Xbit_r30_c236 bl_236 br_236 wl_30 vdd gnd cell_6t
Xbit_r31_c236 bl_236 br_236 wl_31 vdd gnd cell_6t
Xbit_r32_c236 bl_236 br_236 wl_32 vdd gnd cell_6t
Xbit_r33_c236 bl_236 br_236 wl_33 vdd gnd cell_6t
Xbit_r34_c236 bl_236 br_236 wl_34 vdd gnd cell_6t
Xbit_r35_c236 bl_236 br_236 wl_35 vdd gnd cell_6t
Xbit_r36_c236 bl_236 br_236 wl_36 vdd gnd cell_6t
Xbit_r37_c236 bl_236 br_236 wl_37 vdd gnd cell_6t
Xbit_r38_c236 bl_236 br_236 wl_38 vdd gnd cell_6t
Xbit_r39_c236 bl_236 br_236 wl_39 vdd gnd cell_6t
Xbit_r40_c236 bl_236 br_236 wl_40 vdd gnd cell_6t
Xbit_r41_c236 bl_236 br_236 wl_41 vdd gnd cell_6t
Xbit_r42_c236 bl_236 br_236 wl_42 vdd gnd cell_6t
Xbit_r43_c236 bl_236 br_236 wl_43 vdd gnd cell_6t
Xbit_r44_c236 bl_236 br_236 wl_44 vdd gnd cell_6t
Xbit_r45_c236 bl_236 br_236 wl_45 vdd gnd cell_6t
Xbit_r46_c236 bl_236 br_236 wl_46 vdd gnd cell_6t
Xbit_r47_c236 bl_236 br_236 wl_47 vdd gnd cell_6t
Xbit_r48_c236 bl_236 br_236 wl_48 vdd gnd cell_6t
Xbit_r49_c236 bl_236 br_236 wl_49 vdd gnd cell_6t
Xbit_r50_c236 bl_236 br_236 wl_50 vdd gnd cell_6t
Xbit_r51_c236 bl_236 br_236 wl_51 vdd gnd cell_6t
Xbit_r52_c236 bl_236 br_236 wl_52 vdd gnd cell_6t
Xbit_r53_c236 bl_236 br_236 wl_53 vdd gnd cell_6t
Xbit_r54_c236 bl_236 br_236 wl_54 vdd gnd cell_6t
Xbit_r55_c236 bl_236 br_236 wl_55 vdd gnd cell_6t
Xbit_r56_c236 bl_236 br_236 wl_56 vdd gnd cell_6t
Xbit_r57_c236 bl_236 br_236 wl_57 vdd gnd cell_6t
Xbit_r58_c236 bl_236 br_236 wl_58 vdd gnd cell_6t
Xbit_r59_c236 bl_236 br_236 wl_59 vdd gnd cell_6t
Xbit_r60_c236 bl_236 br_236 wl_60 vdd gnd cell_6t
Xbit_r61_c236 bl_236 br_236 wl_61 vdd gnd cell_6t
Xbit_r62_c236 bl_236 br_236 wl_62 vdd gnd cell_6t
Xbit_r63_c236 bl_236 br_236 wl_63 vdd gnd cell_6t
Xbit_r64_c236 bl_236 br_236 wl_64 vdd gnd cell_6t
Xbit_r65_c236 bl_236 br_236 wl_65 vdd gnd cell_6t
Xbit_r66_c236 bl_236 br_236 wl_66 vdd gnd cell_6t
Xbit_r67_c236 bl_236 br_236 wl_67 vdd gnd cell_6t
Xbit_r68_c236 bl_236 br_236 wl_68 vdd gnd cell_6t
Xbit_r69_c236 bl_236 br_236 wl_69 vdd gnd cell_6t
Xbit_r70_c236 bl_236 br_236 wl_70 vdd gnd cell_6t
Xbit_r71_c236 bl_236 br_236 wl_71 vdd gnd cell_6t
Xbit_r72_c236 bl_236 br_236 wl_72 vdd gnd cell_6t
Xbit_r73_c236 bl_236 br_236 wl_73 vdd gnd cell_6t
Xbit_r74_c236 bl_236 br_236 wl_74 vdd gnd cell_6t
Xbit_r75_c236 bl_236 br_236 wl_75 vdd gnd cell_6t
Xbit_r76_c236 bl_236 br_236 wl_76 vdd gnd cell_6t
Xbit_r77_c236 bl_236 br_236 wl_77 vdd gnd cell_6t
Xbit_r78_c236 bl_236 br_236 wl_78 vdd gnd cell_6t
Xbit_r79_c236 bl_236 br_236 wl_79 vdd gnd cell_6t
Xbit_r80_c236 bl_236 br_236 wl_80 vdd gnd cell_6t
Xbit_r81_c236 bl_236 br_236 wl_81 vdd gnd cell_6t
Xbit_r82_c236 bl_236 br_236 wl_82 vdd gnd cell_6t
Xbit_r83_c236 bl_236 br_236 wl_83 vdd gnd cell_6t
Xbit_r84_c236 bl_236 br_236 wl_84 vdd gnd cell_6t
Xbit_r85_c236 bl_236 br_236 wl_85 vdd gnd cell_6t
Xbit_r86_c236 bl_236 br_236 wl_86 vdd gnd cell_6t
Xbit_r87_c236 bl_236 br_236 wl_87 vdd gnd cell_6t
Xbit_r88_c236 bl_236 br_236 wl_88 vdd gnd cell_6t
Xbit_r89_c236 bl_236 br_236 wl_89 vdd gnd cell_6t
Xbit_r90_c236 bl_236 br_236 wl_90 vdd gnd cell_6t
Xbit_r91_c236 bl_236 br_236 wl_91 vdd gnd cell_6t
Xbit_r92_c236 bl_236 br_236 wl_92 vdd gnd cell_6t
Xbit_r93_c236 bl_236 br_236 wl_93 vdd gnd cell_6t
Xbit_r94_c236 bl_236 br_236 wl_94 vdd gnd cell_6t
Xbit_r95_c236 bl_236 br_236 wl_95 vdd gnd cell_6t
Xbit_r96_c236 bl_236 br_236 wl_96 vdd gnd cell_6t
Xbit_r97_c236 bl_236 br_236 wl_97 vdd gnd cell_6t
Xbit_r98_c236 bl_236 br_236 wl_98 vdd gnd cell_6t
Xbit_r99_c236 bl_236 br_236 wl_99 vdd gnd cell_6t
Xbit_r100_c236 bl_236 br_236 wl_100 vdd gnd cell_6t
Xbit_r101_c236 bl_236 br_236 wl_101 vdd gnd cell_6t
Xbit_r102_c236 bl_236 br_236 wl_102 vdd gnd cell_6t
Xbit_r103_c236 bl_236 br_236 wl_103 vdd gnd cell_6t
Xbit_r104_c236 bl_236 br_236 wl_104 vdd gnd cell_6t
Xbit_r105_c236 bl_236 br_236 wl_105 vdd gnd cell_6t
Xbit_r106_c236 bl_236 br_236 wl_106 vdd gnd cell_6t
Xbit_r107_c236 bl_236 br_236 wl_107 vdd gnd cell_6t
Xbit_r108_c236 bl_236 br_236 wl_108 vdd gnd cell_6t
Xbit_r109_c236 bl_236 br_236 wl_109 vdd gnd cell_6t
Xbit_r110_c236 bl_236 br_236 wl_110 vdd gnd cell_6t
Xbit_r111_c236 bl_236 br_236 wl_111 vdd gnd cell_6t
Xbit_r112_c236 bl_236 br_236 wl_112 vdd gnd cell_6t
Xbit_r113_c236 bl_236 br_236 wl_113 vdd gnd cell_6t
Xbit_r114_c236 bl_236 br_236 wl_114 vdd gnd cell_6t
Xbit_r115_c236 bl_236 br_236 wl_115 vdd gnd cell_6t
Xbit_r116_c236 bl_236 br_236 wl_116 vdd gnd cell_6t
Xbit_r117_c236 bl_236 br_236 wl_117 vdd gnd cell_6t
Xbit_r118_c236 bl_236 br_236 wl_118 vdd gnd cell_6t
Xbit_r119_c236 bl_236 br_236 wl_119 vdd gnd cell_6t
Xbit_r120_c236 bl_236 br_236 wl_120 vdd gnd cell_6t
Xbit_r121_c236 bl_236 br_236 wl_121 vdd gnd cell_6t
Xbit_r122_c236 bl_236 br_236 wl_122 vdd gnd cell_6t
Xbit_r123_c236 bl_236 br_236 wl_123 vdd gnd cell_6t
Xbit_r124_c236 bl_236 br_236 wl_124 vdd gnd cell_6t
Xbit_r125_c236 bl_236 br_236 wl_125 vdd gnd cell_6t
Xbit_r126_c236 bl_236 br_236 wl_126 vdd gnd cell_6t
Xbit_r127_c236 bl_236 br_236 wl_127 vdd gnd cell_6t
Xbit_r128_c236 bl_236 br_236 wl_128 vdd gnd cell_6t
Xbit_r129_c236 bl_236 br_236 wl_129 vdd gnd cell_6t
Xbit_r130_c236 bl_236 br_236 wl_130 vdd gnd cell_6t
Xbit_r131_c236 bl_236 br_236 wl_131 vdd gnd cell_6t
Xbit_r132_c236 bl_236 br_236 wl_132 vdd gnd cell_6t
Xbit_r133_c236 bl_236 br_236 wl_133 vdd gnd cell_6t
Xbit_r134_c236 bl_236 br_236 wl_134 vdd gnd cell_6t
Xbit_r135_c236 bl_236 br_236 wl_135 vdd gnd cell_6t
Xbit_r136_c236 bl_236 br_236 wl_136 vdd gnd cell_6t
Xbit_r137_c236 bl_236 br_236 wl_137 vdd gnd cell_6t
Xbit_r138_c236 bl_236 br_236 wl_138 vdd gnd cell_6t
Xbit_r139_c236 bl_236 br_236 wl_139 vdd gnd cell_6t
Xbit_r140_c236 bl_236 br_236 wl_140 vdd gnd cell_6t
Xbit_r141_c236 bl_236 br_236 wl_141 vdd gnd cell_6t
Xbit_r142_c236 bl_236 br_236 wl_142 vdd gnd cell_6t
Xbit_r143_c236 bl_236 br_236 wl_143 vdd gnd cell_6t
Xbit_r144_c236 bl_236 br_236 wl_144 vdd gnd cell_6t
Xbit_r145_c236 bl_236 br_236 wl_145 vdd gnd cell_6t
Xbit_r146_c236 bl_236 br_236 wl_146 vdd gnd cell_6t
Xbit_r147_c236 bl_236 br_236 wl_147 vdd gnd cell_6t
Xbit_r148_c236 bl_236 br_236 wl_148 vdd gnd cell_6t
Xbit_r149_c236 bl_236 br_236 wl_149 vdd gnd cell_6t
Xbit_r150_c236 bl_236 br_236 wl_150 vdd gnd cell_6t
Xbit_r151_c236 bl_236 br_236 wl_151 vdd gnd cell_6t
Xbit_r152_c236 bl_236 br_236 wl_152 vdd gnd cell_6t
Xbit_r153_c236 bl_236 br_236 wl_153 vdd gnd cell_6t
Xbit_r154_c236 bl_236 br_236 wl_154 vdd gnd cell_6t
Xbit_r155_c236 bl_236 br_236 wl_155 vdd gnd cell_6t
Xbit_r156_c236 bl_236 br_236 wl_156 vdd gnd cell_6t
Xbit_r157_c236 bl_236 br_236 wl_157 vdd gnd cell_6t
Xbit_r158_c236 bl_236 br_236 wl_158 vdd gnd cell_6t
Xbit_r159_c236 bl_236 br_236 wl_159 vdd gnd cell_6t
Xbit_r160_c236 bl_236 br_236 wl_160 vdd gnd cell_6t
Xbit_r161_c236 bl_236 br_236 wl_161 vdd gnd cell_6t
Xbit_r162_c236 bl_236 br_236 wl_162 vdd gnd cell_6t
Xbit_r163_c236 bl_236 br_236 wl_163 vdd gnd cell_6t
Xbit_r164_c236 bl_236 br_236 wl_164 vdd gnd cell_6t
Xbit_r165_c236 bl_236 br_236 wl_165 vdd gnd cell_6t
Xbit_r166_c236 bl_236 br_236 wl_166 vdd gnd cell_6t
Xbit_r167_c236 bl_236 br_236 wl_167 vdd gnd cell_6t
Xbit_r168_c236 bl_236 br_236 wl_168 vdd gnd cell_6t
Xbit_r169_c236 bl_236 br_236 wl_169 vdd gnd cell_6t
Xbit_r170_c236 bl_236 br_236 wl_170 vdd gnd cell_6t
Xbit_r171_c236 bl_236 br_236 wl_171 vdd gnd cell_6t
Xbit_r172_c236 bl_236 br_236 wl_172 vdd gnd cell_6t
Xbit_r173_c236 bl_236 br_236 wl_173 vdd gnd cell_6t
Xbit_r174_c236 bl_236 br_236 wl_174 vdd gnd cell_6t
Xbit_r175_c236 bl_236 br_236 wl_175 vdd gnd cell_6t
Xbit_r176_c236 bl_236 br_236 wl_176 vdd gnd cell_6t
Xbit_r177_c236 bl_236 br_236 wl_177 vdd gnd cell_6t
Xbit_r178_c236 bl_236 br_236 wl_178 vdd gnd cell_6t
Xbit_r179_c236 bl_236 br_236 wl_179 vdd gnd cell_6t
Xbit_r180_c236 bl_236 br_236 wl_180 vdd gnd cell_6t
Xbit_r181_c236 bl_236 br_236 wl_181 vdd gnd cell_6t
Xbit_r182_c236 bl_236 br_236 wl_182 vdd gnd cell_6t
Xbit_r183_c236 bl_236 br_236 wl_183 vdd gnd cell_6t
Xbit_r184_c236 bl_236 br_236 wl_184 vdd gnd cell_6t
Xbit_r185_c236 bl_236 br_236 wl_185 vdd gnd cell_6t
Xbit_r186_c236 bl_236 br_236 wl_186 vdd gnd cell_6t
Xbit_r187_c236 bl_236 br_236 wl_187 vdd gnd cell_6t
Xbit_r188_c236 bl_236 br_236 wl_188 vdd gnd cell_6t
Xbit_r189_c236 bl_236 br_236 wl_189 vdd gnd cell_6t
Xbit_r190_c236 bl_236 br_236 wl_190 vdd gnd cell_6t
Xbit_r191_c236 bl_236 br_236 wl_191 vdd gnd cell_6t
Xbit_r192_c236 bl_236 br_236 wl_192 vdd gnd cell_6t
Xbit_r193_c236 bl_236 br_236 wl_193 vdd gnd cell_6t
Xbit_r194_c236 bl_236 br_236 wl_194 vdd gnd cell_6t
Xbit_r195_c236 bl_236 br_236 wl_195 vdd gnd cell_6t
Xbit_r196_c236 bl_236 br_236 wl_196 vdd gnd cell_6t
Xbit_r197_c236 bl_236 br_236 wl_197 vdd gnd cell_6t
Xbit_r198_c236 bl_236 br_236 wl_198 vdd gnd cell_6t
Xbit_r199_c236 bl_236 br_236 wl_199 vdd gnd cell_6t
Xbit_r200_c236 bl_236 br_236 wl_200 vdd gnd cell_6t
Xbit_r201_c236 bl_236 br_236 wl_201 vdd gnd cell_6t
Xbit_r202_c236 bl_236 br_236 wl_202 vdd gnd cell_6t
Xbit_r203_c236 bl_236 br_236 wl_203 vdd gnd cell_6t
Xbit_r204_c236 bl_236 br_236 wl_204 vdd gnd cell_6t
Xbit_r205_c236 bl_236 br_236 wl_205 vdd gnd cell_6t
Xbit_r206_c236 bl_236 br_236 wl_206 vdd gnd cell_6t
Xbit_r207_c236 bl_236 br_236 wl_207 vdd gnd cell_6t
Xbit_r208_c236 bl_236 br_236 wl_208 vdd gnd cell_6t
Xbit_r209_c236 bl_236 br_236 wl_209 vdd gnd cell_6t
Xbit_r210_c236 bl_236 br_236 wl_210 vdd gnd cell_6t
Xbit_r211_c236 bl_236 br_236 wl_211 vdd gnd cell_6t
Xbit_r212_c236 bl_236 br_236 wl_212 vdd gnd cell_6t
Xbit_r213_c236 bl_236 br_236 wl_213 vdd gnd cell_6t
Xbit_r214_c236 bl_236 br_236 wl_214 vdd gnd cell_6t
Xbit_r215_c236 bl_236 br_236 wl_215 vdd gnd cell_6t
Xbit_r216_c236 bl_236 br_236 wl_216 vdd gnd cell_6t
Xbit_r217_c236 bl_236 br_236 wl_217 vdd gnd cell_6t
Xbit_r218_c236 bl_236 br_236 wl_218 vdd gnd cell_6t
Xbit_r219_c236 bl_236 br_236 wl_219 vdd gnd cell_6t
Xbit_r220_c236 bl_236 br_236 wl_220 vdd gnd cell_6t
Xbit_r221_c236 bl_236 br_236 wl_221 vdd gnd cell_6t
Xbit_r222_c236 bl_236 br_236 wl_222 vdd gnd cell_6t
Xbit_r223_c236 bl_236 br_236 wl_223 vdd gnd cell_6t
Xbit_r224_c236 bl_236 br_236 wl_224 vdd gnd cell_6t
Xbit_r225_c236 bl_236 br_236 wl_225 vdd gnd cell_6t
Xbit_r226_c236 bl_236 br_236 wl_226 vdd gnd cell_6t
Xbit_r227_c236 bl_236 br_236 wl_227 vdd gnd cell_6t
Xbit_r228_c236 bl_236 br_236 wl_228 vdd gnd cell_6t
Xbit_r229_c236 bl_236 br_236 wl_229 vdd gnd cell_6t
Xbit_r230_c236 bl_236 br_236 wl_230 vdd gnd cell_6t
Xbit_r231_c236 bl_236 br_236 wl_231 vdd gnd cell_6t
Xbit_r232_c236 bl_236 br_236 wl_232 vdd gnd cell_6t
Xbit_r233_c236 bl_236 br_236 wl_233 vdd gnd cell_6t
Xbit_r234_c236 bl_236 br_236 wl_234 vdd gnd cell_6t
Xbit_r235_c236 bl_236 br_236 wl_235 vdd gnd cell_6t
Xbit_r236_c236 bl_236 br_236 wl_236 vdd gnd cell_6t
Xbit_r237_c236 bl_236 br_236 wl_237 vdd gnd cell_6t
Xbit_r238_c236 bl_236 br_236 wl_238 vdd gnd cell_6t
Xbit_r239_c236 bl_236 br_236 wl_239 vdd gnd cell_6t
Xbit_r240_c236 bl_236 br_236 wl_240 vdd gnd cell_6t
Xbit_r241_c236 bl_236 br_236 wl_241 vdd gnd cell_6t
Xbit_r242_c236 bl_236 br_236 wl_242 vdd gnd cell_6t
Xbit_r243_c236 bl_236 br_236 wl_243 vdd gnd cell_6t
Xbit_r244_c236 bl_236 br_236 wl_244 vdd gnd cell_6t
Xbit_r245_c236 bl_236 br_236 wl_245 vdd gnd cell_6t
Xbit_r246_c236 bl_236 br_236 wl_246 vdd gnd cell_6t
Xbit_r247_c236 bl_236 br_236 wl_247 vdd gnd cell_6t
Xbit_r248_c236 bl_236 br_236 wl_248 vdd gnd cell_6t
Xbit_r249_c236 bl_236 br_236 wl_249 vdd gnd cell_6t
Xbit_r250_c236 bl_236 br_236 wl_250 vdd gnd cell_6t
Xbit_r251_c236 bl_236 br_236 wl_251 vdd gnd cell_6t
Xbit_r252_c236 bl_236 br_236 wl_252 vdd gnd cell_6t
Xbit_r253_c236 bl_236 br_236 wl_253 vdd gnd cell_6t
Xbit_r254_c236 bl_236 br_236 wl_254 vdd gnd cell_6t
Xbit_r255_c236 bl_236 br_236 wl_255 vdd gnd cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd cell_6t
Xbit_r1_c237 bl_237 br_237 wl_1 vdd gnd cell_6t
Xbit_r2_c237 bl_237 br_237 wl_2 vdd gnd cell_6t
Xbit_r3_c237 bl_237 br_237 wl_3 vdd gnd cell_6t
Xbit_r4_c237 bl_237 br_237 wl_4 vdd gnd cell_6t
Xbit_r5_c237 bl_237 br_237 wl_5 vdd gnd cell_6t
Xbit_r6_c237 bl_237 br_237 wl_6 vdd gnd cell_6t
Xbit_r7_c237 bl_237 br_237 wl_7 vdd gnd cell_6t
Xbit_r8_c237 bl_237 br_237 wl_8 vdd gnd cell_6t
Xbit_r9_c237 bl_237 br_237 wl_9 vdd gnd cell_6t
Xbit_r10_c237 bl_237 br_237 wl_10 vdd gnd cell_6t
Xbit_r11_c237 bl_237 br_237 wl_11 vdd gnd cell_6t
Xbit_r12_c237 bl_237 br_237 wl_12 vdd gnd cell_6t
Xbit_r13_c237 bl_237 br_237 wl_13 vdd gnd cell_6t
Xbit_r14_c237 bl_237 br_237 wl_14 vdd gnd cell_6t
Xbit_r15_c237 bl_237 br_237 wl_15 vdd gnd cell_6t
Xbit_r16_c237 bl_237 br_237 wl_16 vdd gnd cell_6t
Xbit_r17_c237 bl_237 br_237 wl_17 vdd gnd cell_6t
Xbit_r18_c237 bl_237 br_237 wl_18 vdd gnd cell_6t
Xbit_r19_c237 bl_237 br_237 wl_19 vdd gnd cell_6t
Xbit_r20_c237 bl_237 br_237 wl_20 vdd gnd cell_6t
Xbit_r21_c237 bl_237 br_237 wl_21 vdd gnd cell_6t
Xbit_r22_c237 bl_237 br_237 wl_22 vdd gnd cell_6t
Xbit_r23_c237 bl_237 br_237 wl_23 vdd gnd cell_6t
Xbit_r24_c237 bl_237 br_237 wl_24 vdd gnd cell_6t
Xbit_r25_c237 bl_237 br_237 wl_25 vdd gnd cell_6t
Xbit_r26_c237 bl_237 br_237 wl_26 vdd gnd cell_6t
Xbit_r27_c237 bl_237 br_237 wl_27 vdd gnd cell_6t
Xbit_r28_c237 bl_237 br_237 wl_28 vdd gnd cell_6t
Xbit_r29_c237 bl_237 br_237 wl_29 vdd gnd cell_6t
Xbit_r30_c237 bl_237 br_237 wl_30 vdd gnd cell_6t
Xbit_r31_c237 bl_237 br_237 wl_31 vdd gnd cell_6t
Xbit_r32_c237 bl_237 br_237 wl_32 vdd gnd cell_6t
Xbit_r33_c237 bl_237 br_237 wl_33 vdd gnd cell_6t
Xbit_r34_c237 bl_237 br_237 wl_34 vdd gnd cell_6t
Xbit_r35_c237 bl_237 br_237 wl_35 vdd gnd cell_6t
Xbit_r36_c237 bl_237 br_237 wl_36 vdd gnd cell_6t
Xbit_r37_c237 bl_237 br_237 wl_37 vdd gnd cell_6t
Xbit_r38_c237 bl_237 br_237 wl_38 vdd gnd cell_6t
Xbit_r39_c237 bl_237 br_237 wl_39 vdd gnd cell_6t
Xbit_r40_c237 bl_237 br_237 wl_40 vdd gnd cell_6t
Xbit_r41_c237 bl_237 br_237 wl_41 vdd gnd cell_6t
Xbit_r42_c237 bl_237 br_237 wl_42 vdd gnd cell_6t
Xbit_r43_c237 bl_237 br_237 wl_43 vdd gnd cell_6t
Xbit_r44_c237 bl_237 br_237 wl_44 vdd gnd cell_6t
Xbit_r45_c237 bl_237 br_237 wl_45 vdd gnd cell_6t
Xbit_r46_c237 bl_237 br_237 wl_46 vdd gnd cell_6t
Xbit_r47_c237 bl_237 br_237 wl_47 vdd gnd cell_6t
Xbit_r48_c237 bl_237 br_237 wl_48 vdd gnd cell_6t
Xbit_r49_c237 bl_237 br_237 wl_49 vdd gnd cell_6t
Xbit_r50_c237 bl_237 br_237 wl_50 vdd gnd cell_6t
Xbit_r51_c237 bl_237 br_237 wl_51 vdd gnd cell_6t
Xbit_r52_c237 bl_237 br_237 wl_52 vdd gnd cell_6t
Xbit_r53_c237 bl_237 br_237 wl_53 vdd gnd cell_6t
Xbit_r54_c237 bl_237 br_237 wl_54 vdd gnd cell_6t
Xbit_r55_c237 bl_237 br_237 wl_55 vdd gnd cell_6t
Xbit_r56_c237 bl_237 br_237 wl_56 vdd gnd cell_6t
Xbit_r57_c237 bl_237 br_237 wl_57 vdd gnd cell_6t
Xbit_r58_c237 bl_237 br_237 wl_58 vdd gnd cell_6t
Xbit_r59_c237 bl_237 br_237 wl_59 vdd gnd cell_6t
Xbit_r60_c237 bl_237 br_237 wl_60 vdd gnd cell_6t
Xbit_r61_c237 bl_237 br_237 wl_61 vdd gnd cell_6t
Xbit_r62_c237 bl_237 br_237 wl_62 vdd gnd cell_6t
Xbit_r63_c237 bl_237 br_237 wl_63 vdd gnd cell_6t
Xbit_r64_c237 bl_237 br_237 wl_64 vdd gnd cell_6t
Xbit_r65_c237 bl_237 br_237 wl_65 vdd gnd cell_6t
Xbit_r66_c237 bl_237 br_237 wl_66 vdd gnd cell_6t
Xbit_r67_c237 bl_237 br_237 wl_67 vdd gnd cell_6t
Xbit_r68_c237 bl_237 br_237 wl_68 vdd gnd cell_6t
Xbit_r69_c237 bl_237 br_237 wl_69 vdd gnd cell_6t
Xbit_r70_c237 bl_237 br_237 wl_70 vdd gnd cell_6t
Xbit_r71_c237 bl_237 br_237 wl_71 vdd gnd cell_6t
Xbit_r72_c237 bl_237 br_237 wl_72 vdd gnd cell_6t
Xbit_r73_c237 bl_237 br_237 wl_73 vdd gnd cell_6t
Xbit_r74_c237 bl_237 br_237 wl_74 vdd gnd cell_6t
Xbit_r75_c237 bl_237 br_237 wl_75 vdd gnd cell_6t
Xbit_r76_c237 bl_237 br_237 wl_76 vdd gnd cell_6t
Xbit_r77_c237 bl_237 br_237 wl_77 vdd gnd cell_6t
Xbit_r78_c237 bl_237 br_237 wl_78 vdd gnd cell_6t
Xbit_r79_c237 bl_237 br_237 wl_79 vdd gnd cell_6t
Xbit_r80_c237 bl_237 br_237 wl_80 vdd gnd cell_6t
Xbit_r81_c237 bl_237 br_237 wl_81 vdd gnd cell_6t
Xbit_r82_c237 bl_237 br_237 wl_82 vdd gnd cell_6t
Xbit_r83_c237 bl_237 br_237 wl_83 vdd gnd cell_6t
Xbit_r84_c237 bl_237 br_237 wl_84 vdd gnd cell_6t
Xbit_r85_c237 bl_237 br_237 wl_85 vdd gnd cell_6t
Xbit_r86_c237 bl_237 br_237 wl_86 vdd gnd cell_6t
Xbit_r87_c237 bl_237 br_237 wl_87 vdd gnd cell_6t
Xbit_r88_c237 bl_237 br_237 wl_88 vdd gnd cell_6t
Xbit_r89_c237 bl_237 br_237 wl_89 vdd gnd cell_6t
Xbit_r90_c237 bl_237 br_237 wl_90 vdd gnd cell_6t
Xbit_r91_c237 bl_237 br_237 wl_91 vdd gnd cell_6t
Xbit_r92_c237 bl_237 br_237 wl_92 vdd gnd cell_6t
Xbit_r93_c237 bl_237 br_237 wl_93 vdd gnd cell_6t
Xbit_r94_c237 bl_237 br_237 wl_94 vdd gnd cell_6t
Xbit_r95_c237 bl_237 br_237 wl_95 vdd gnd cell_6t
Xbit_r96_c237 bl_237 br_237 wl_96 vdd gnd cell_6t
Xbit_r97_c237 bl_237 br_237 wl_97 vdd gnd cell_6t
Xbit_r98_c237 bl_237 br_237 wl_98 vdd gnd cell_6t
Xbit_r99_c237 bl_237 br_237 wl_99 vdd gnd cell_6t
Xbit_r100_c237 bl_237 br_237 wl_100 vdd gnd cell_6t
Xbit_r101_c237 bl_237 br_237 wl_101 vdd gnd cell_6t
Xbit_r102_c237 bl_237 br_237 wl_102 vdd gnd cell_6t
Xbit_r103_c237 bl_237 br_237 wl_103 vdd gnd cell_6t
Xbit_r104_c237 bl_237 br_237 wl_104 vdd gnd cell_6t
Xbit_r105_c237 bl_237 br_237 wl_105 vdd gnd cell_6t
Xbit_r106_c237 bl_237 br_237 wl_106 vdd gnd cell_6t
Xbit_r107_c237 bl_237 br_237 wl_107 vdd gnd cell_6t
Xbit_r108_c237 bl_237 br_237 wl_108 vdd gnd cell_6t
Xbit_r109_c237 bl_237 br_237 wl_109 vdd gnd cell_6t
Xbit_r110_c237 bl_237 br_237 wl_110 vdd gnd cell_6t
Xbit_r111_c237 bl_237 br_237 wl_111 vdd gnd cell_6t
Xbit_r112_c237 bl_237 br_237 wl_112 vdd gnd cell_6t
Xbit_r113_c237 bl_237 br_237 wl_113 vdd gnd cell_6t
Xbit_r114_c237 bl_237 br_237 wl_114 vdd gnd cell_6t
Xbit_r115_c237 bl_237 br_237 wl_115 vdd gnd cell_6t
Xbit_r116_c237 bl_237 br_237 wl_116 vdd gnd cell_6t
Xbit_r117_c237 bl_237 br_237 wl_117 vdd gnd cell_6t
Xbit_r118_c237 bl_237 br_237 wl_118 vdd gnd cell_6t
Xbit_r119_c237 bl_237 br_237 wl_119 vdd gnd cell_6t
Xbit_r120_c237 bl_237 br_237 wl_120 vdd gnd cell_6t
Xbit_r121_c237 bl_237 br_237 wl_121 vdd gnd cell_6t
Xbit_r122_c237 bl_237 br_237 wl_122 vdd gnd cell_6t
Xbit_r123_c237 bl_237 br_237 wl_123 vdd gnd cell_6t
Xbit_r124_c237 bl_237 br_237 wl_124 vdd gnd cell_6t
Xbit_r125_c237 bl_237 br_237 wl_125 vdd gnd cell_6t
Xbit_r126_c237 bl_237 br_237 wl_126 vdd gnd cell_6t
Xbit_r127_c237 bl_237 br_237 wl_127 vdd gnd cell_6t
Xbit_r128_c237 bl_237 br_237 wl_128 vdd gnd cell_6t
Xbit_r129_c237 bl_237 br_237 wl_129 vdd gnd cell_6t
Xbit_r130_c237 bl_237 br_237 wl_130 vdd gnd cell_6t
Xbit_r131_c237 bl_237 br_237 wl_131 vdd gnd cell_6t
Xbit_r132_c237 bl_237 br_237 wl_132 vdd gnd cell_6t
Xbit_r133_c237 bl_237 br_237 wl_133 vdd gnd cell_6t
Xbit_r134_c237 bl_237 br_237 wl_134 vdd gnd cell_6t
Xbit_r135_c237 bl_237 br_237 wl_135 vdd gnd cell_6t
Xbit_r136_c237 bl_237 br_237 wl_136 vdd gnd cell_6t
Xbit_r137_c237 bl_237 br_237 wl_137 vdd gnd cell_6t
Xbit_r138_c237 bl_237 br_237 wl_138 vdd gnd cell_6t
Xbit_r139_c237 bl_237 br_237 wl_139 vdd gnd cell_6t
Xbit_r140_c237 bl_237 br_237 wl_140 vdd gnd cell_6t
Xbit_r141_c237 bl_237 br_237 wl_141 vdd gnd cell_6t
Xbit_r142_c237 bl_237 br_237 wl_142 vdd gnd cell_6t
Xbit_r143_c237 bl_237 br_237 wl_143 vdd gnd cell_6t
Xbit_r144_c237 bl_237 br_237 wl_144 vdd gnd cell_6t
Xbit_r145_c237 bl_237 br_237 wl_145 vdd gnd cell_6t
Xbit_r146_c237 bl_237 br_237 wl_146 vdd gnd cell_6t
Xbit_r147_c237 bl_237 br_237 wl_147 vdd gnd cell_6t
Xbit_r148_c237 bl_237 br_237 wl_148 vdd gnd cell_6t
Xbit_r149_c237 bl_237 br_237 wl_149 vdd gnd cell_6t
Xbit_r150_c237 bl_237 br_237 wl_150 vdd gnd cell_6t
Xbit_r151_c237 bl_237 br_237 wl_151 vdd gnd cell_6t
Xbit_r152_c237 bl_237 br_237 wl_152 vdd gnd cell_6t
Xbit_r153_c237 bl_237 br_237 wl_153 vdd gnd cell_6t
Xbit_r154_c237 bl_237 br_237 wl_154 vdd gnd cell_6t
Xbit_r155_c237 bl_237 br_237 wl_155 vdd gnd cell_6t
Xbit_r156_c237 bl_237 br_237 wl_156 vdd gnd cell_6t
Xbit_r157_c237 bl_237 br_237 wl_157 vdd gnd cell_6t
Xbit_r158_c237 bl_237 br_237 wl_158 vdd gnd cell_6t
Xbit_r159_c237 bl_237 br_237 wl_159 vdd gnd cell_6t
Xbit_r160_c237 bl_237 br_237 wl_160 vdd gnd cell_6t
Xbit_r161_c237 bl_237 br_237 wl_161 vdd gnd cell_6t
Xbit_r162_c237 bl_237 br_237 wl_162 vdd gnd cell_6t
Xbit_r163_c237 bl_237 br_237 wl_163 vdd gnd cell_6t
Xbit_r164_c237 bl_237 br_237 wl_164 vdd gnd cell_6t
Xbit_r165_c237 bl_237 br_237 wl_165 vdd gnd cell_6t
Xbit_r166_c237 bl_237 br_237 wl_166 vdd gnd cell_6t
Xbit_r167_c237 bl_237 br_237 wl_167 vdd gnd cell_6t
Xbit_r168_c237 bl_237 br_237 wl_168 vdd gnd cell_6t
Xbit_r169_c237 bl_237 br_237 wl_169 vdd gnd cell_6t
Xbit_r170_c237 bl_237 br_237 wl_170 vdd gnd cell_6t
Xbit_r171_c237 bl_237 br_237 wl_171 vdd gnd cell_6t
Xbit_r172_c237 bl_237 br_237 wl_172 vdd gnd cell_6t
Xbit_r173_c237 bl_237 br_237 wl_173 vdd gnd cell_6t
Xbit_r174_c237 bl_237 br_237 wl_174 vdd gnd cell_6t
Xbit_r175_c237 bl_237 br_237 wl_175 vdd gnd cell_6t
Xbit_r176_c237 bl_237 br_237 wl_176 vdd gnd cell_6t
Xbit_r177_c237 bl_237 br_237 wl_177 vdd gnd cell_6t
Xbit_r178_c237 bl_237 br_237 wl_178 vdd gnd cell_6t
Xbit_r179_c237 bl_237 br_237 wl_179 vdd gnd cell_6t
Xbit_r180_c237 bl_237 br_237 wl_180 vdd gnd cell_6t
Xbit_r181_c237 bl_237 br_237 wl_181 vdd gnd cell_6t
Xbit_r182_c237 bl_237 br_237 wl_182 vdd gnd cell_6t
Xbit_r183_c237 bl_237 br_237 wl_183 vdd gnd cell_6t
Xbit_r184_c237 bl_237 br_237 wl_184 vdd gnd cell_6t
Xbit_r185_c237 bl_237 br_237 wl_185 vdd gnd cell_6t
Xbit_r186_c237 bl_237 br_237 wl_186 vdd gnd cell_6t
Xbit_r187_c237 bl_237 br_237 wl_187 vdd gnd cell_6t
Xbit_r188_c237 bl_237 br_237 wl_188 vdd gnd cell_6t
Xbit_r189_c237 bl_237 br_237 wl_189 vdd gnd cell_6t
Xbit_r190_c237 bl_237 br_237 wl_190 vdd gnd cell_6t
Xbit_r191_c237 bl_237 br_237 wl_191 vdd gnd cell_6t
Xbit_r192_c237 bl_237 br_237 wl_192 vdd gnd cell_6t
Xbit_r193_c237 bl_237 br_237 wl_193 vdd gnd cell_6t
Xbit_r194_c237 bl_237 br_237 wl_194 vdd gnd cell_6t
Xbit_r195_c237 bl_237 br_237 wl_195 vdd gnd cell_6t
Xbit_r196_c237 bl_237 br_237 wl_196 vdd gnd cell_6t
Xbit_r197_c237 bl_237 br_237 wl_197 vdd gnd cell_6t
Xbit_r198_c237 bl_237 br_237 wl_198 vdd gnd cell_6t
Xbit_r199_c237 bl_237 br_237 wl_199 vdd gnd cell_6t
Xbit_r200_c237 bl_237 br_237 wl_200 vdd gnd cell_6t
Xbit_r201_c237 bl_237 br_237 wl_201 vdd gnd cell_6t
Xbit_r202_c237 bl_237 br_237 wl_202 vdd gnd cell_6t
Xbit_r203_c237 bl_237 br_237 wl_203 vdd gnd cell_6t
Xbit_r204_c237 bl_237 br_237 wl_204 vdd gnd cell_6t
Xbit_r205_c237 bl_237 br_237 wl_205 vdd gnd cell_6t
Xbit_r206_c237 bl_237 br_237 wl_206 vdd gnd cell_6t
Xbit_r207_c237 bl_237 br_237 wl_207 vdd gnd cell_6t
Xbit_r208_c237 bl_237 br_237 wl_208 vdd gnd cell_6t
Xbit_r209_c237 bl_237 br_237 wl_209 vdd gnd cell_6t
Xbit_r210_c237 bl_237 br_237 wl_210 vdd gnd cell_6t
Xbit_r211_c237 bl_237 br_237 wl_211 vdd gnd cell_6t
Xbit_r212_c237 bl_237 br_237 wl_212 vdd gnd cell_6t
Xbit_r213_c237 bl_237 br_237 wl_213 vdd gnd cell_6t
Xbit_r214_c237 bl_237 br_237 wl_214 vdd gnd cell_6t
Xbit_r215_c237 bl_237 br_237 wl_215 vdd gnd cell_6t
Xbit_r216_c237 bl_237 br_237 wl_216 vdd gnd cell_6t
Xbit_r217_c237 bl_237 br_237 wl_217 vdd gnd cell_6t
Xbit_r218_c237 bl_237 br_237 wl_218 vdd gnd cell_6t
Xbit_r219_c237 bl_237 br_237 wl_219 vdd gnd cell_6t
Xbit_r220_c237 bl_237 br_237 wl_220 vdd gnd cell_6t
Xbit_r221_c237 bl_237 br_237 wl_221 vdd gnd cell_6t
Xbit_r222_c237 bl_237 br_237 wl_222 vdd gnd cell_6t
Xbit_r223_c237 bl_237 br_237 wl_223 vdd gnd cell_6t
Xbit_r224_c237 bl_237 br_237 wl_224 vdd gnd cell_6t
Xbit_r225_c237 bl_237 br_237 wl_225 vdd gnd cell_6t
Xbit_r226_c237 bl_237 br_237 wl_226 vdd gnd cell_6t
Xbit_r227_c237 bl_237 br_237 wl_227 vdd gnd cell_6t
Xbit_r228_c237 bl_237 br_237 wl_228 vdd gnd cell_6t
Xbit_r229_c237 bl_237 br_237 wl_229 vdd gnd cell_6t
Xbit_r230_c237 bl_237 br_237 wl_230 vdd gnd cell_6t
Xbit_r231_c237 bl_237 br_237 wl_231 vdd gnd cell_6t
Xbit_r232_c237 bl_237 br_237 wl_232 vdd gnd cell_6t
Xbit_r233_c237 bl_237 br_237 wl_233 vdd gnd cell_6t
Xbit_r234_c237 bl_237 br_237 wl_234 vdd gnd cell_6t
Xbit_r235_c237 bl_237 br_237 wl_235 vdd gnd cell_6t
Xbit_r236_c237 bl_237 br_237 wl_236 vdd gnd cell_6t
Xbit_r237_c237 bl_237 br_237 wl_237 vdd gnd cell_6t
Xbit_r238_c237 bl_237 br_237 wl_238 vdd gnd cell_6t
Xbit_r239_c237 bl_237 br_237 wl_239 vdd gnd cell_6t
Xbit_r240_c237 bl_237 br_237 wl_240 vdd gnd cell_6t
Xbit_r241_c237 bl_237 br_237 wl_241 vdd gnd cell_6t
Xbit_r242_c237 bl_237 br_237 wl_242 vdd gnd cell_6t
Xbit_r243_c237 bl_237 br_237 wl_243 vdd gnd cell_6t
Xbit_r244_c237 bl_237 br_237 wl_244 vdd gnd cell_6t
Xbit_r245_c237 bl_237 br_237 wl_245 vdd gnd cell_6t
Xbit_r246_c237 bl_237 br_237 wl_246 vdd gnd cell_6t
Xbit_r247_c237 bl_237 br_237 wl_247 vdd gnd cell_6t
Xbit_r248_c237 bl_237 br_237 wl_248 vdd gnd cell_6t
Xbit_r249_c237 bl_237 br_237 wl_249 vdd gnd cell_6t
Xbit_r250_c237 bl_237 br_237 wl_250 vdd gnd cell_6t
Xbit_r251_c237 bl_237 br_237 wl_251 vdd gnd cell_6t
Xbit_r252_c237 bl_237 br_237 wl_252 vdd gnd cell_6t
Xbit_r253_c237 bl_237 br_237 wl_253 vdd gnd cell_6t
Xbit_r254_c237 bl_237 br_237 wl_254 vdd gnd cell_6t
Xbit_r255_c237 bl_237 br_237 wl_255 vdd gnd cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd cell_6t
Xbit_r1_c238 bl_238 br_238 wl_1 vdd gnd cell_6t
Xbit_r2_c238 bl_238 br_238 wl_2 vdd gnd cell_6t
Xbit_r3_c238 bl_238 br_238 wl_3 vdd gnd cell_6t
Xbit_r4_c238 bl_238 br_238 wl_4 vdd gnd cell_6t
Xbit_r5_c238 bl_238 br_238 wl_5 vdd gnd cell_6t
Xbit_r6_c238 bl_238 br_238 wl_6 vdd gnd cell_6t
Xbit_r7_c238 bl_238 br_238 wl_7 vdd gnd cell_6t
Xbit_r8_c238 bl_238 br_238 wl_8 vdd gnd cell_6t
Xbit_r9_c238 bl_238 br_238 wl_9 vdd gnd cell_6t
Xbit_r10_c238 bl_238 br_238 wl_10 vdd gnd cell_6t
Xbit_r11_c238 bl_238 br_238 wl_11 vdd gnd cell_6t
Xbit_r12_c238 bl_238 br_238 wl_12 vdd gnd cell_6t
Xbit_r13_c238 bl_238 br_238 wl_13 vdd gnd cell_6t
Xbit_r14_c238 bl_238 br_238 wl_14 vdd gnd cell_6t
Xbit_r15_c238 bl_238 br_238 wl_15 vdd gnd cell_6t
Xbit_r16_c238 bl_238 br_238 wl_16 vdd gnd cell_6t
Xbit_r17_c238 bl_238 br_238 wl_17 vdd gnd cell_6t
Xbit_r18_c238 bl_238 br_238 wl_18 vdd gnd cell_6t
Xbit_r19_c238 bl_238 br_238 wl_19 vdd gnd cell_6t
Xbit_r20_c238 bl_238 br_238 wl_20 vdd gnd cell_6t
Xbit_r21_c238 bl_238 br_238 wl_21 vdd gnd cell_6t
Xbit_r22_c238 bl_238 br_238 wl_22 vdd gnd cell_6t
Xbit_r23_c238 bl_238 br_238 wl_23 vdd gnd cell_6t
Xbit_r24_c238 bl_238 br_238 wl_24 vdd gnd cell_6t
Xbit_r25_c238 bl_238 br_238 wl_25 vdd gnd cell_6t
Xbit_r26_c238 bl_238 br_238 wl_26 vdd gnd cell_6t
Xbit_r27_c238 bl_238 br_238 wl_27 vdd gnd cell_6t
Xbit_r28_c238 bl_238 br_238 wl_28 vdd gnd cell_6t
Xbit_r29_c238 bl_238 br_238 wl_29 vdd gnd cell_6t
Xbit_r30_c238 bl_238 br_238 wl_30 vdd gnd cell_6t
Xbit_r31_c238 bl_238 br_238 wl_31 vdd gnd cell_6t
Xbit_r32_c238 bl_238 br_238 wl_32 vdd gnd cell_6t
Xbit_r33_c238 bl_238 br_238 wl_33 vdd gnd cell_6t
Xbit_r34_c238 bl_238 br_238 wl_34 vdd gnd cell_6t
Xbit_r35_c238 bl_238 br_238 wl_35 vdd gnd cell_6t
Xbit_r36_c238 bl_238 br_238 wl_36 vdd gnd cell_6t
Xbit_r37_c238 bl_238 br_238 wl_37 vdd gnd cell_6t
Xbit_r38_c238 bl_238 br_238 wl_38 vdd gnd cell_6t
Xbit_r39_c238 bl_238 br_238 wl_39 vdd gnd cell_6t
Xbit_r40_c238 bl_238 br_238 wl_40 vdd gnd cell_6t
Xbit_r41_c238 bl_238 br_238 wl_41 vdd gnd cell_6t
Xbit_r42_c238 bl_238 br_238 wl_42 vdd gnd cell_6t
Xbit_r43_c238 bl_238 br_238 wl_43 vdd gnd cell_6t
Xbit_r44_c238 bl_238 br_238 wl_44 vdd gnd cell_6t
Xbit_r45_c238 bl_238 br_238 wl_45 vdd gnd cell_6t
Xbit_r46_c238 bl_238 br_238 wl_46 vdd gnd cell_6t
Xbit_r47_c238 bl_238 br_238 wl_47 vdd gnd cell_6t
Xbit_r48_c238 bl_238 br_238 wl_48 vdd gnd cell_6t
Xbit_r49_c238 bl_238 br_238 wl_49 vdd gnd cell_6t
Xbit_r50_c238 bl_238 br_238 wl_50 vdd gnd cell_6t
Xbit_r51_c238 bl_238 br_238 wl_51 vdd gnd cell_6t
Xbit_r52_c238 bl_238 br_238 wl_52 vdd gnd cell_6t
Xbit_r53_c238 bl_238 br_238 wl_53 vdd gnd cell_6t
Xbit_r54_c238 bl_238 br_238 wl_54 vdd gnd cell_6t
Xbit_r55_c238 bl_238 br_238 wl_55 vdd gnd cell_6t
Xbit_r56_c238 bl_238 br_238 wl_56 vdd gnd cell_6t
Xbit_r57_c238 bl_238 br_238 wl_57 vdd gnd cell_6t
Xbit_r58_c238 bl_238 br_238 wl_58 vdd gnd cell_6t
Xbit_r59_c238 bl_238 br_238 wl_59 vdd gnd cell_6t
Xbit_r60_c238 bl_238 br_238 wl_60 vdd gnd cell_6t
Xbit_r61_c238 bl_238 br_238 wl_61 vdd gnd cell_6t
Xbit_r62_c238 bl_238 br_238 wl_62 vdd gnd cell_6t
Xbit_r63_c238 bl_238 br_238 wl_63 vdd gnd cell_6t
Xbit_r64_c238 bl_238 br_238 wl_64 vdd gnd cell_6t
Xbit_r65_c238 bl_238 br_238 wl_65 vdd gnd cell_6t
Xbit_r66_c238 bl_238 br_238 wl_66 vdd gnd cell_6t
Xbit_r67_c238 bl_238 br_238 wl_67 vdd gnd cell_6t
Xbit_r68_c238 bl_238 br_238 wl_68 vdd gnd cell_6t
Xbit_r69_c238 bl_238 br_238 wl_69 vdd gnd cell_6t
Xbit_r70_c238 bl_238 br_238 wl_70 vdd gnd cell_6t
Xbit_r71_c238 bl_238 br_238 wl_71 vdd gnd cell_6t
Xbit_r72_c238 bl_238 br_238 wl_72 vdd gnd cell_6t
Xbit_r73_c238 bl_238 br_238 wl_73 vdd gnd cell_6t
Xbit_r74_c238 bl_238 br_238 wl_74 vdd gnd cell_6t
Xbit_r75_c238 bl_238 br_238 wl_75 vdd gnd cell_6t
Xbit_r76_c238 bl_238 br_238 wl_76 vdd gnd cell_6t
Xbit_r77_c238 bl_238 br_238 wl_77 vdd gnd cell_6t
Xbit_r78_c238 bl_238 br_238 wl_78 vdd gnd cell_6t
Xbit_r79_c238 bl_238 br_238 wl_79 vdd gnd cell_6t
Xbit_r80_c238 bl_238 br_238 wl_80 vdd gnd cell_6t
Xbit_r81_c238 bl_238 br_238 wl_81 vdd gnd cell_6t
Xbit_r82_c238 bl_238 br_238 wl_82 vdd gnd cell_6t
Xbit_r83_c238 bl_238 br_238 wl_83 vdd gnd cell_6t
Xbit_r84_c238 bl_238 br_238 wl_84 vdd gnd cell_6t
Xbit_r85_c238 bl_238 br_238 wl_85 vdd gnd cell_6t
Xbit_r86_c238 bl_238 br_238 wl_86 vdd gnd cell_6t
Xbit_r87_c238 bl_238 br_238 wl_87 vdd gnd cell_6t
Xbit_r88_c238 bl_238 br_238 wl_88 vdd gnd cell_6t
Xbit_r89_c238 bl_238 br_238 wl_89 vdd gnd cell_6t
Xbit_r90_c238 bl_238 br_238 wl_90 vdd gnd cell_6t
Xbit_r91_c238 bl_238 br_238 wl_91 vdd gnd cell_6t
Xbit_r92_c238 bl_238 br_238 wl_92 vdd gnd cell_6t
Xbit_r93_c238 bl_238 br_238 wl_93 vdd gnd cell_6t
Xbit_r94_c238 bl_238 br_238 wl_94 vdd gnd cell_6t
Xbit_r95_c238 bl_238 br_238 wl_95 vdd gnd cell_6t
Xbit_r96_c238 bl_238 br_238 wl_96 vdd gnd cell_6t
Xbit_r97_c238 bl_238 br_238 wl_97 vdd gnd cell_6t
Xbit_r98_c238 bl_238 br_238 wl_98 vdd gnd cell_6t
Xbit_r99_c238 bl_238 br_238 wl_99 vdd gnd cell_6t
Xbit_r100_c238 bl_238 br_238 wl_100 vdd gnd cell_6t
Xbit_r101_c238 bl_238 br_238 wl_101 vdd gnd cell_6t
Xbit_r102_c238 bl_238 br_238 wl_102 vdd gnd cell_6t
Xbit_r103_c238 bl_238 br_238 wl_103 vdd gnd cell_6t
Xbit_r104_c238 bl_238 br_238 wl_104 vdd gnd cell_6t
Xbit_r105_c238 bl_238 br_238 wl_105 vdd gnd cell_6t
Xbit_r106_c238 bl_238 br_238 wl_106 vdd gnd cell_6t
Xbit_r107_c238 bl_238 br_238 wl_107 vdd gnd cell_6t
Xbit_r108_c238 bl_238 br_238 wl_108 vdd gnd cell_6t
Xbit_r109_c238 bl_238 br_238 wl_109 vdd gnd cell_6t
Xbit_r110_c238 bl_238 br_238 wl_110 vdd gnd cell_6t
Xbit_r111_c238 bl_238 br_238 wl_111 vdd gnd cell_6t
Xbit_r112_c238 bl_238 br_238 wl_112 vdd gnd cell_6t
Xbit_r113_c238 bl_238 br_238 wl_113 vdd gnd cell_6t
Xbit_r114_c238 bl_238 br_238 wl_114 vdd gnd cell_6t
Xbit_r115_c238 bl_238 br_238 wl_115 vdd gnd cell_6t
Xbit_r116_c238 bl_238 br_238 wl_116 vdd gnd cell_6t
Xbit_r117_c238 bl_238 br_238 wl_117 vdd gnd cell_6t
Xbit_r118_c238 bl_238 br_238 wl_118 vdd gnd cell_6t
Xbit_r119_c238 bl_238 br_238 wl_119 vdd gnd cell_6t
Xbit_r120_c238 bl_238 br_238 wl_120 vdd gnd cell_6t
Xbit_r121_c238 bl_238 br_238 wl_121 vdd gnd cell_6t
Xbit_r122_c238 bl_238 br_238 wl_122 vdd gnd cell_6t
Xbit_r123_c238 bl_238 br_238 wl_123 vdd gnd cell_6t
Xbit_r124_c238 bl_238 br_238 wl_124 vdd gnd cell_6t
Xbit_r125_c238 bl_238 br_238 wl_125 vdd gnd cell_6t
Xbit_r126_c238 bl_238 br_238 wl_126 vdd gnd cell_6t
Xbit_r127_c238 bl_238 br_238 wl_127 vdd gnd cell_6t
Xbit_r128_c238 bl_238 br_238 wl_128 vdd gnd cell_6t
Xbit_r129_c238 bl_238 br_238 wl_129 vdd gnd cell_6t
Xbit_r130_c238 bl_238 br_238 wl_130 vdd gnd cell_6t
Xbit_r131_c238 bl_238 br_238 wl_131 vdd gnd cell_6t
Xbit_r132_c238 bl_238 br_238 wl_132 vdd gnd cell_6t
Xbit_r133_c238 bl_238 br_238 wl_133 vdd gnd cell_6t
Xbit_r134_c238 bl_238 br_238 wl_134 vdd gnd cell_6t
Xbit_r135_c238 bl_238 br_238 wl_135 vdd gnd cell_6t
Xbit_r136_c238 bl_238 br_238 wl_136 vdd gnd cell_6t
Xbit_r137_c238 bl_238 br_238 wl_137 vdd gnd cell_6t
Xbit_r138_c238 bl_238 br_238 wl_138 vdd gnd cell_6t
Xbit_r139_c238 bl_238 br_238 wl_139 vdd gnd cell_6t
Xbit_r140_c238 bl_238 br_238 wl_140 vdd gnd cell_6t
Xbit_r141_c238 bl_238 br_238 wl_141 vdd gnd cell_6t
Xbit_r142_c238 bl_238 br_238 wl_142 vdd gnd cell_6t
Xbit_r143_c238 bl_238 br_238 wl_143 vdd gnd cell_6t
Xbit_r144_c238 bl_238 br_238 wl_144 vdd gnd cell_6t
Xbit_r145_c238 bl_238 br_238 wl_145 vdd gnd cell_6t
Xbit_r146_c238 bl_238 br_238 wl_146 vdd gnd cell_6t
Xbit_r147_c238 bl_238 br_238 wl_147 vdd gnd cell_6t
Xbit_r148_c238 bl_238 br_238 wl_148 vdd gnd cell_6t
Xbit_r149_c238 bl_238 br_238 wl_149 vdd gnd cell_6t
Xbit_r150_c238 bl_238 br_238 wl_150 vdd gnd cell_6t
Xbit_r151_c238 bl_238 br_238 wl_151 vdd gnd cell_6t
Xbit_r152_c238 bl_238 br_238 wl_152 vdd gnd cell_6t
Xbit_r153_c238 bl_238 br_238 wl_153 vdd gnd cell_6t
Xbit_r154_c238 bl_238 br_238 wl_154 vdd gnd cell_6t
Xbit_r155_c238 bl_238 br_238 wl_155 vdd gnd cell_6t
Xbit_r156_c238 bl_238 br_238 wl_156 vdd gnd cell_6t
Xbit_r157_c238 bl_238 br_238 wl_157 vdd gnd cell_6t
Xbit_r158_c238 bl_238 br_238 wl_158 vdd gnd cell_6t
Xbit_r159_c238 bl_238 br_238 wl_159 vdd gnd cell_6t
Xbit_r160_c238 bl_238 br_238 wl_160 vdd gnd cell_6t
Xbit_r161_c238 bl_238 br_238 wl_161 vdd gnd cell_6t
Xbit_r162_c238 bl_238 br_238 wl_162 vdd gnd cell_6t
Xbit_r163_c238 bl_238 br_238 wl_163 vdd gnd cell_6t
Xbit_r164_c238 bl_238 br_238 wl_164 vdd gnd cell_6t
Xbit_r165_c238 bl_238 br_238 wl_165 vdd gnd cell_6t
Xbit_r166_c238 bl_238 br_238 wl_166 vdd gnd cell_6t
Xbit_r167_c238 bl_238 br_238 wl_167 vdd gnd cell_6t
Xbit_r168_c238 bl_238 br_238 wl_168 vdd gnd cell_6t
Xbit_r169_c238 bl_238 br_238 wl_169 vdd gnd cell_6t
Xbit_r170_c238 bl_238 br_238 wl_170 vdd gnd cell_6t
Xbit_r171_c238 bl_238 br_238 wl_171 vdd gnd cell_6t
Xbit_r172_c238 bl_238 br_238 wl_172 vdd gnd cell_6t
Xbit_r173_c238 bl_238 br_238 wl_173 vdd gnd cell_6t
Xbit_r174_c238 bl_238 br_238 wl_174 vdd gnd cell_6t
Xbit_r175_c238 bl_238 br_238 wl_175 vdd gnd cell_6t
Xbit_r176_c238 bl_238 br_238 wl_176 vdd gnd cell_6t
Xbit_r177_c238 bl_238 br_238 wl_177 vdd gnd cell_6t
Xbit_r178_c238 bl_238 br_238 wl_178 vdd gnd cell_6t
Xbit_r179_c238 bl_238 br_238 wl_179 vdd gnd cell_6t
Xbit_r180_c238 bl_238 br_238 wl_180 vdd gnd cell_6t
Xbit_r181_c238 bl_238 br_238 wl_181 vdd gnd cell_6t
Xbit_r182_c238 bl_238 br_238 wl_182 vdd gnd cell_6t
Xbit_r183_c238 bl_238 br_238 wl_183 vdd gnd cell_6t
Xbit_r184_c238 bl_238 br_238 wl_184 vdd gnd cell_6t
Xbit_r185_c238 bl_238 br_238 wl_185 vdd gnd cell_6t
Xbit_r186_c238 bl_238 br_238 wl_186 vdd gnd cell_6t
Xbit_r187_c238 bl_238 br_238 wl_187 vdd gnd cell_6t
Xbit_r188_c238 bl_238 br_238 wl_188 vdd gnd cell_6t
Xbit_r189_c238 bl_238 br_238 wl_189 vdd gnd cell_6t
Xbit_r190_c238 bl_238 br_238 wl_190 vdd gnd cell_6t
Xbit_r191_c238 bl_238 br_238 wl_191 vdd gnd cell_6t
Xbit_r192_c238 bl_238 br_238 wl_192 vdd gnd cell_6t
Xbit_r193_c238 bl_238 br_238 wl_193 vdd gnd cell_6t
Xbit_r194_c238 bl_238 br_238 wl_194 vdd gnd cell_6t
Xbit_r195_c238 bl_238 br_238 wl_195 vdd gnd cell_6t
Xbit_r196_c238 bl_238 br_238 wl_196 vdd gnd cell_6t
Xbit_r197_c238 bl_238 br_238 wl_197 vdd gnd cell_6t
Xbit_r198_c238 bl_238 br_238 wl_198 vdd gnd cell_6t
Xbit_r199_c238 bl_238 br_238 wl_199 vdd gnd cell_6t
Xbit_r200_c238 bl_238 br_238 wl_200 vdd gnd cell_6t
Xbit_r201_c238 bl_238 br_238 wl_201 vdd gnd cell_6t
Xbit_r202_c238 bl_238 br_238 wl_202 vdd gnd cell_6t
Xbit_r203_c238 bl_238 br_238 wl_203 vdd gnd cell_6t
Xbit_r204_c238 bl_238 br_238 wl_204 vdd gnd cell_6t
Xbit_r205_c238 bl_238 br_238 wl_205 vdd gnd cell_6t
Xbit_r206_c238 bl_238 br_238 wl_206 vdd gnd cell_6t
Xbit_r207_c238 bl_238 br_238 wl_207 vdd gnd cell_6t
Xbit_r208_c238 bl_238 br_238 wl_208 vdd gnd cell_6t
Xbit_r209_c238 bl_238 br_238 wl_209 vdd gnd cell_6t
Xbit_r210_c238 bl_238 br_238 wl_210 vdd gnd cell_6t
Xbit_r211_c238 bl_238 br_238 wl_211 vdd gnd cell_6t
Xbit_r212_c238 bl_238 br_238 wl_212 vdd gnd cell_6t
Xbit_r213_c238 bl_238 br_238 wl_213 vdd gnd cell_6t
Xbit_r214_c238 bl_238 br_238 wl_214 vdd gnd cell_6t
Xbit_r215_c238 bl_238 br_238 wl_215 vdd gnd cell_6t
Xbit_r216_c238 bl_238 br_238 wl_216 vdd gnd cell_6t
Xbit_r217_c238 bl_238 br_238 wl_217 vdd gnd cell_6t
Xbit_r218_c238 bl_238 br_238 wl_218 vdd gnd cell_6t
Xbit_r219_c238 bl_238 br_238 wl_219 vdd gnd cell_6t
Xbit_r220_c238 bl_238 br_238 wl_220 vdd gnd cell_6t
Xbit_r221_c238 bl_238 br_238 wl_221 vdd gnd cell_6t
Xbit_r222_c238 bl_238 br_238 wl_222 vdd gnd cell_6t
Xbit_r223_c238 bl_238 br_238 wl_223 vdd gnd cell_6t
Xbit_r224_c238 bl_238 br_238 wl_224 vdd gnd cell_6t
Xbit_r225_c238 bl_238 br_238 wl_225 vdd gnd cell_6t
Xbit_r226_c238 bl_238 br_238 wl_226 vdd gnd cell_6t
Xbit_r227_c238 bl_238 br_238 wl_227 vdd gnd cell_6t
Xbit_r228_c238 bl_238 br_238 wl_228 vdd gnd cell_6t
Xbit_r229_c238 bl_238 br_238 wl_229 vdd gnd cell_6t
Xbit_r230_c238 bl_238 br_238 wl_230 vdd gnd cell_6t
Xbit_r231_c238 bl_238 br_238 wl_231 vdd gnd cell_6t
Xbit_r232_c238 bl_238 br_238 wl_232 vdd gnd cell_6t
Xbit_r233_c238 bl_238 br_238 wl_233 vdd gnd cell_6t
Xbit_r234_c238 bl_238 br_238 wl_234 vdd gnd cell_6t
Xbit_r235_c238 bl_238 br_238 wl_235 vdd gnd cell_6t
Xbit_r236_c238 bl_238 br_238 wl_236 vdd gnd cell_6t
Xbit_r237_c238 bl_238 br_238 wl_237 vdd gnd cell_6t
Xbit_r238_c238 bl_238 br_238 wl_238 vdd gnd cell_6t
Xbit_r239_c238 bl_238 br_238 wl_239 vdd gnd cell_6t
Xbit_r240_c238 bl_238 br_238 wl_240 vdd gnd cell_6t
Xbit_r241_c238 bl_238 br_238 wl_241 vdd gnd cell_6t
Xbit_r242_c238 bl_238 br_238 wl_242 vdd gnd cell_6t
Xbit_r243_c238 bl_238 br_238 wl_243 vdd gnd cell_6t
Xbit_r244_c238 bl_238 br_238 wl_244 vdd gnd cell_6t
Xbit_r245_c238 bl_238 br_238 wl_245 vdd gnd cell_6t
Xbit_r246_c238 bl_238 br_238 wl_246 vdd gnd cell_6t
Xbit_r247_c238 bl_238 br_238 wl_247 vdd gnd cell_6t
Xbit_r248_c238 bl_238 br_238 wl_248 vdd gnd cell_6t
Xbit_r249_c238 bl_238 br_238 wl_249 vdd gnd cell_6t
Xbit_r250_c238 bl_238 br_238 wl_250 vdd gnd cell_6t
Xbit_r251_c238 bl_238 br_238 wl_251 vdd gnd cell_6t
Xbit_r252_c238 bl_238 br_238 wl_252 vdd gnd cell_6t
Xbit_r253_c238 bl_238 br_238 wl_253 vdd gnd cell_6t
Xbit_r254_c238 bl_238 br_238 wl_254 vdd gnd cell_6t
Xbit_r255_c238 bl_238 br_238 wl_255 vdd gnd cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd cell_6t
Xbit_r1_c239 bl_239 br_239 wl_1 vdd gnd cell_6t
Xbit_r2_c239 bl_239 br_239 wl_2 vdd gnd cell_6t
Xbit_r3_c239 bl_239 br_239 wl_3 vdd gnd cell_6t
Xbit_r4_c239 bl_239 br_239 wl_4 vdd gnd cell_6t
Xbit_r5_c239 bl_239 br_239 wl_5 vdd gnd cell_6t
Xbit_r6_c239 bl_239 br_239 wl_6 vdd gnd cell_6t
Xbit_r7_c239 bl_239 br_239 wl_7 vdd gnd cell_6t
Xbit_r8_c239 bl_239 br_239 wl_8 vdd gnd cell_6t
Xbit_r9_c239 bl_239 br_239 wl_9 vdd gnd cell_6t
Xbit_r10_c239 bl_239 br_239 wl_10 vdd gnd cell_6t
Xbit_r11_c239 bl_239 br_239 wl_11 vdd gnd cell_6t
Xbit_r12_c239 bl_239 br_239 wl_12 vdd gnd cell_6t
Xbit_r13_c239 bl_239 br_239 wl_13 vdd gnd cell_6t
Xbit_r14_c239 bl_239 br_239 wl_14 vdd gnd cell_6t
Xbit_r15_c239 bl_239 br_239 wl_15 vdd gnd cell_6t
Xbit_r16_c239 bl_239 br_239 wl_16 vdd gnd cell_6t
Xbit_r17_c239 bl_239 br_239 wl_17 vdd gnd cell_6t
Xbit_r18_c239 bl_239 br_239 wl_18 vdd gnd cell_6t
Xbit_r19_c239 bl_239 br_239 wl_19 vdd gnd cell_6t
Xbit_r20_c239 bl_239 br_239 wl_20 vdd gnd cell_6t
Xbit_r21_c239 bl_239 br_239 wl_21 vdd gnd cell_6t
Xbit_r22_c239 bl_239 br_239 wl_22 vdd gnd cell_6t
Xbit_r23_c239 bl_239 br_239 wl_23 vdd gnd cell_6t
Xbit_r24_c239 bl_239 br_239 wl_24 vdd gnd cell_6t
Xbit_r25_c239 bl_239 br_239 wl_25 vdd gnd cell_6t
Xbit_r26_c239 bl_239 br_239 wl_26 vdd gnd cell_6t
Xbit_r27_c239 bl_239 br_239 wl_27 vdd gnd cell_6t
Xbit_r28_c239 bl_239 br_239 wl_28 vdd gnd cell_6t
Xbit_r29_c239 bl_239 br_239 wl_29 vdd gnd cell_6t
Xbit_r30_c239 bl_239 br_239 wl_30 vdd gnd cell_6t
Xbit_r31_c239 bl_239 br_239 wl_31 vdd gnd cell_6t
Xbit_r32_c239 bl_239 br_239 wl_32 vdd gnd cell_6t
Xbit_r33_c239 bl_239 br_239 wl_33 vdd gnd cell_6t
Xbit_r34_c239 bl_239 br_239 wl_34 vdd gnd cell_6t
Xbit_r35_c239 bl_239 br_239 wl_35 vdd gnd cell_6t
Xbit_r36_c239 bl_239 br_239 wl_36 vdd gnd cell_6t
Xbit_r37_c239 bl_239 br_239 wl_37 vdd gnd cell_6t
Xbit_r38_c239 bl_239 br_239 wl_38 vdd gnd cell_6t
Xbit_r39_c239 bl_239 br_239 wl_39 vdd gnd cell_6t
Xbit_r40_c239 bl_239 br_239 wl_40 vdd gnd cell_6t
Xbit_r41_c239 bl_239 br_239 wl_41 vdd gnd cell_6t
Xbit_r42_c239 bl_239 br_239 wl_42 vdd gnd cell_6t
Xbit_r43_c239 bl_239 br_239 wl_43 vdd gnd cell_6t
Xbit_r44_c239 bl_239 br_239 wl_44 vdd gnd cell_6t
Xbit_r45_c239 bl_239 br_239 wl_45 vdd gnd cell_6t
Xbit_r46_c239 bl_239 br_239 wl_46 vdd gnd cell_6t
Xbit_r47_c239 bl_239 br_239 wl_47 vdd gnd cell_6t
Xbit_r48_c239 bl_239 br_239 wl_48 vdd gnd cell_6t
Xbit_r49_c239 bl_239 br_239 wl_49 vdd gnd cell_6t
Xbit_r50_c239 bl_239 br_239 wl_50 vdd gnd cell_6t
Xbit_r51_c239 bl_239 br_239 wl_51 vdd gnd cell_6t
Xbit_r52_c239 bl_239 br_239 wl_52 vdd gnd cell_6t
Xbit_r53_c239 bl_239 br_239 wl_53 vdd gnd cell_6t
Xbit_r54_c239 bl_239 br_239 wl_54 vdd gnd cell_6t
Xbit_r55_c239 bl_239 br_239 wl_55 vdd gnd cell_6t
Xbit_r56_c239 bl_239 br_239 wl_56 vdd gnd cell_6t
Xbit_r57_c239 bl_239 br_239 wl_57 vdd gnd cell_6t
Xbit_r58_c239 bl_239 br_239 wl_58 vdd gnd cell_6t
Xbit_r59_c239 bl_239 br_239 wl_59 vdd gnd cell_6t
Xbit_r60_c239 bl_239 br_239 wl_60 vdd gnd cell_6t
Xbit_r61_c239 bl_239 br_239 wl_61 vdd gnd cell_6t
Xbit_r62_c239 bl_239 br_239 wl_62 vdd gnd cell_6t
Xbit_r63_c239 bl_239 br_239 wl_63 vdd gnd cell_6t
Xbit_r64_c239 bl_239 br_239 wl_64 vdd gnd cell_6t
Xbit_r65_c239 bl_239 br_239 wl_65 vdd gnd cell_6t
Xbit_r66_c239 bl_239 br_239 wl_66 vdd gnd cell_6t
Xbit_r67_c239 bl_239 br_239 wl_67 vdd gnd cell_6t
Xbit_r68_c239 bl_239 br_239 wl_68 vdd gnd cell_6t
Xbit_r69_c239 bl_239 br_239 wl_69 vdd gnd cell_6t
Xbit_r70_c239 bl_239 br_239 wl_70 vdd gnd cell_6t
Xbit_r71_c239 bl_239 br_239 wl_71 vdd gnd cell_6t
Xbit_r72_c239 bl_239 br_239 wl_72 vdd gnd cell_6t
Xbit_r73_c239 bl_239 br_239 wl_73 vdd gnd cell_6t
Xbit_r74_c239 bl_239 br_239 wl_74 vdd gnd cell_6t
Xbit_r75_c239 bl_239 br_239 wl_75 vdd gnd cell_6t
Xbit_r76_c239 bl_239 br_239 wl_76 vdd gnd cell_6t
Xbit_r77_c239 bl_239 br_239 wl_77 vdd gnd cell_6t
Xbit_r78_c239 bl_239 br_239 wl_78 vdd gnd cell_6t
Xbit_r79_c239 bl_239 br_239 wl_79 vdd gnd cell_6t
Xbit_r80_c239 bl_239 br_239 wl_80 vdd gnd cell_6t
Xbit_r81_c239 bl_239 br_239 wl_81 vdd gnd cell_6t
Xbit_r82_c239 bl_239 br_239 wl_82 vdd gnd cell_6t
Xbit_r83_c239 bl_239 br_239 wl_83 vdd gnd cell_6t
Xbit_r84_c239 bl_239 br_239 wl_84 vdd gnd cell_6t
Xbit_r85_c239 bl_239 br_239 wl_85 vdd gnd cell_6t
Xbit_r86_c239 bl_239 br_239 wl_86 vdd gnd cell_6t
Xbit_r87_c239 bl_239 br_239 wl_87 vdd gnd cell_6t
Xbit_r88_c239 bl_239 br_239 wl_88 vdd gnd cell_6t
Xbit_r89_c239 bl_239 br_239 wl_89 vdd gnd cell_6t
Xbit_r90_c239 bl_239 br_239 wl_90 vdd gnd cell_6t
Xbit_r91_c239 bl_239 br_239 wl_91 vdd gnd cell_6t
Xbit_r92_c239 bl_239 br_239 wl_92 vdd gnd cell_6t
Xbit_r93_c239 bl_239 br_239 wl_93 vdd gnd cell_6t
Xbit_r94_c239 bl_239 br_239 wl_94 vdd gnd cell_6t
Xbit_r95_c239 bl_239 br_239 wl_95 vdd gnd cell_6t
Xbit_r96_c239 bl_239 br_239 wl_96 vdd gnd cell_6t
Xbit_r97_c239 bl_239 br_239 wl_97 vdd gnd cell_6t
Xbit_r98_c239 bl_239 br_239 wl_98 vdd gnd cell_6t
Xbit_r99_c239 bl_239 br_239 wl_99 vdd gnd cell_6t
Xbit_r100_c239 bl_239 br_239 wl_100 vdd gnd cell_6t
Xbit_r101_c239 bl_239 br_239 wl_101 vdd gnd cell_6t
Xbit_r102_c239 bl_239 br_239 wl_102 vdd gnd cell_6t
Xbit_r103_c239 bl_239 br_239 wl_103 vdd gnd cell_6t
Xbit_r104_c239 bl_239 br_239 wl_104 vdd gnd cell_6t
Xbit_r105_c239 bl_239 br_239 wl_105 vdd gnd cell_6t
Xbit_r106_c239 bl_239 br_239 wl_106 vdd gnd cell_6t
Xbit_r107_c239 bl_239 br_239 wl_107 vdd gnd cell_6t
Xbit_r108_c239 bl_239 br_239 wl_108 vdd gnd cell_6t
Xbit_r109_c239 bl_239 br_239 wl_109 vdd gnd cell_6t
Xbit_r110_c239 bl_239 br_239 wl_110 vdd gnd cell_6t
Xbit_r111_c239 bl_239 br_239 wl_111 vdd gnd cell_6t
Xbit_r112_c239 bl_239 br_239 wl_112 vdd gnd cell_6t
Xbit_r113_c239 bl_239 br_239 wl_113 vdd gnd cell_6t
Xbit_r114_c239 bl_239 br_239 wl_114 vdd gnd cell_6t
Xbit_r115_c239 bl_239 br_239 wl_115 vdd gnd cell_6t
Xbit_r116_c239 bl_239 br_239 wl_116 vdd gnd cell_6t
Xbit_r117_c239 bl_239 br_239 wl_117 vdd gnd cell_6t
Xbit_r118_c239 bl_239 br_239 wl_118 vdd gnd cell_6t
Xbit_r119_c239 bl_239 br_239 wl_119 vdd gnd cell_6t
Xbit_r120_c239 bl_239 br_239 wl_120 vdd gnd cell_6t
Xbit_r121_c239 bl_239 br_239 wl_121 vdd gnd cell_6t
Xbit_r122_c239 bl_239 br_239 wl_122 vdd gnd cell_6t
Xbit_r123_c239 bl_239 br_239 wl_123 vdd gnd cell_6t
Xbit_r124_c239 bl_239 br_239 wl_124 vdd gnd cell_6t
Xbit_r125_c239 bl_239 br_239 wl_125 vdd gnd cell_6t
Xbit_r126_c239 bl_239 br_239 wl_126 vdd gnd cell_6t
Xbit_r127_c239 bl_239 br_239 wl_127 vdd gnd cell_6t
Xbit_r128_c239 bl_239 br_239 wl_128 vdd gnd cell_6t
Xbit_r129_c239 bl_239 br_239 wl_129 vdd gnd cell_6t
Xbit_r130_c239 bl_239 br_239 wl_130 vdd gnd cell_6t
Xbit_r131_c239 bl_239 br_239 wl_131 vdd gnd cell_6t
Xbit_r132_c239 bl_239 br_239 wl_132 vdd gnd cell_6t
Xbit_r133_c239 bl_239 br_239 wl_133 vdd gnd cell_6t
Xbit_r134_c239 bl_239 br_239 wl_134 vdd gnd cell_6t
Xbit_r135_c239 bl_239 br_239 wl_135 vdd gnd cell_6t
Xbit_r136_c239 bl_239 br_239 wl_136 vdd gnd cell_6t
Xbit_r137_c239 bl_239 br_239 wl_137 vdd gnd cell_6t
Xbit_r138_c239 bl_239 br_239 wl_138 vdd gnd cell_6t
Xbit_r139_c239 bl_239 br_239 wl_139 vdd gnd cell_6t
Xbit_r140_c239 bl_239 br_239 wl_140 vdd gnd cell_6t
Xbit_r141_c239 bl_239 br_239 wl_141 vdd gnd cell_6t
Xbit_r142_c239 bl_239 br_239 wl_142 vdd gnd cell_6t
Xbit_r143_c239 bl_239 br_239 wl_143 vdd gnd cell_6t
Xbit_r144_c239 bl_239 br_239 wl_144 vdd gnd cell_6t
Xbit_r145_c239 bl_239 br_239 wl_145 vdd gnd cell_6t
Xbit_r146_c239 bl_239 br_239 wl_146 vdd gnd cell_6t
Xbit_r147_c239 bl_239 br_239 wl_147 vdd gnd cell_6t
Xbit_r148_c239 bl_239 br_239 wl_148 vdd gnd cell_6t
Xbit_r149_c239 bl_239 br_239 wl_149 vdd gnd cell_6t
Xbit_r150_c239 bl_239 br_239 wl_150 vdd gnd cell_6t
Xbit_r151_c239 bl_239 br_239 wl_151 vdd gnd cell_6t
Xbit_r152_c239 bl_239 br_239 wl_152 vdd gnd cell_6t
Xbit_r153_c239 bl_239 br_239 wl_153 vdd gnd cell_6t
Xbit_r154_c239 bl_239 br_239 wl_154 vdd gnd cell_6t
Xbit_r155_c239 bl_239 br_239 wl_155 vdd gnd cell_6t
Xbit_r156_c239 bl_239 br_239 wl_156 vdd gnd cell_6t
Xbit_r157_c239 bl_239 br_239 wl_157 vdd gnd cell_6t
Xbit_r158_c239 bl_239 br_239 wl_158 vdd gnd cell_6t
Xbit_r159_c239 bl_239 br_239 wl_159 vdd gnd cell_6t
Xbit_r160_c239 bl_239 br_239 wl_160 vdd gnd cell_6t
Xbit_r161_c239 bl_239 br_239 wl_161 vdd gnd cell_6t
Xbit_r162_c239 bl_239 br_239 wl_162 vdd gnd cell_6t
Xbit_r163_c239 bl_239 br_239 wl_163 vdd gnd cell_6t
Xbit_r164_c239 bl_239 br_239 wl_164 vdd gnd cell_6t
Xbit_r165_c239 bl_239 br_239 wl_165 vdd gnd cell_6t
Xbit_r166_c239 bl_239 br_239 wl_166 vdd gnd cell_6t
Xbit_r167_c239 bl_239 br_239 wl_167 vdd gnd cell_6t
Xbit_r168_c239 bl_239 br_239 wl_168 vdd gnd cell_6t
Xbit_r169_c239 bl_239 br_239 wl_169 vdd gnd cell_6t
Xbit_r170_c239 bl_239 br_239 wl_170 vdd gnd cell_6t
Xbit_r171_c239 bl_239 br_239 wl_171 vdd gnd cell_6t
Xbit_r172_c239 bl_239 br_239 wl_172 vdd gnd cell_6t
Xbit_r173_c239 bl_239 br_239 wl_173 vdd gnd cell_6t
Xbit_r174_c239 bl_239 br_239 wl_174 vdd gnd cell_6t
Xbit_r175_c239 bl_239 br_239 wl_175 vdd gnd cell_6t
Xbit_r176_c239 bl_239 br_239 wl_176 vdd gnd cell_6t
Xbit_r177_c239 bl_239 br_239 wl_177 vdd gnd cell_6t
Xbit_r178_c239 bl_239 br_239 wl_178 vdd gnd cell_6t
Xbit_r179_c239 bl_239 br_239 wl_179 vdd gnd cell_6t
Xbit_r180_c239 bl_239 br_239 wl_180 vdd gnd cell_6t
Xbit_r181_c239 bl_239 br_239 wl_181 vdd gnd cell_6t
Xbit_r182_c239 bl_239 br_239 wl_182 vdd gnd cell_6t
Xbit_r183_c239 bl_239 br_239 wl_183 vdd gnd cell_6t
Xbit_r184_c239 bl_239 br_239 wl_184 vdd gnd cell_6t
Xbit_r185_c239 bl_239 br_239 wl_185 vdd gnd cell_6t
Xbit_r186_c239 bl_239 br_239 wl_186 vdd gnd cell_6t
Xbit_r187_c239 bl_239 br_239 wl_187 vdd gnd cell_6t
Xbit_r188_c239 bl_239 br_239 wl_188 vdd gnd cell_6t
Xbit_r189_c239 bl_239 br_239 wl_189 vdd gnd cell_6t
Xbit_r190_c239 bl_239 br_239 wl_190 vdd gnd cell_6t
Xbit_r191_c239 bl_239 br_239 wl_191 vdd gnd cell_6t
Xbit_r192_c239 bl_239 br_239 wl_192 vdd gnd cell_6t
Xbit_r193_c239 bl_239 br_239 wl_193 vdd gnd cell_6t
Xbit_r194_c239 bl_239 br_239 wl_194 vdd gnd cell_6t
Xbit_r195_c239 bl_239 br_239 wl_195 vdd gnd cell_6t
Xbit_r196_c239 bl_239 br_239 wl_196 vdd gnd cell_6t
Xbit_r197_c239 bl_239 br_239 wl_197 vdd gnd cell_6t
Xbit_r198_c239 bl_239 br_239 wl_198 vdd gnd cell_6t
Xbit_r199_c239 bl_239 br_239 wl_199 vdd gnd cell_6t
Xbit_r200_c239 bl_239 br_239 wl_200 vdd gnd cell_6t
Xbit_r201_c239 bl_239 br_239 wl_201 vdd gnd cell_6t
Xbit_r202_c239 bl_239 br_239 wl_202 vdd gnd cell_6t
Xbit_r203_c239 bl_239 br_239 wl_203 vdd gnd cell_6t
Xbit_r204_c239 bl_239 br_239 wl_204 vdd gnd cell_6t
Xbit_r205_c239 bl_239 br_239 wl_205 vdd gnd cell_6t
Xbit_r206_c239 bl_239 br_239 wl_206 vdd gnd cell_6t
Xbit_r207_c239 bl_239 br_239 wl_207 vdd gnd cell_6t
Xbit_r208_c239 bl_239 br_239 wl_208 vdd gnd cell_6t
Xbit_r209_c239 bl_239 br_239 wl_209 vdd gnd cell_6t
Xbit_r210_c239 bl_239 br_239 wl_210 vdd gnd cell_6t
Xbit_r211_c239 bl_239 br_239 wl_211 vdd gnd cell_6t
Xbit_r212_c239 bl_239 br_239 wl_212 vdd gnd cell_6t
Xbit_r213_c239 bl_239 br_239 wl_213 vdd gnd cell_6t
Xbit_r214_c239 bl_239 br_239 wl_214 vdd gnd cell_6t
Xbit_r215_c239 bl_239 br_239 wl_215 vdd gnd cell_6t
Xbit_r216_c239 bl_239 br_239 wl_216 vdd gnd cell_6t
Xbit_r217_c239 bl_239 br_239 wl_217 vdd gnd cell_6t
Xbit_r218_c239 bl_239 br_239 wl_218 vdd gnd cell_6t
Xbit_r219_c239 bl_239 br_239 wl_219 vdd gnd cell_6t
Xbit_r220_c239 bl_239 br_239 wl_220 vdd gnd cell_6t
Xbit_r221_c239 bl_239 br_239 wl_221 vdd gnd cell_6t
Xbit_r222_c239 bl_239 br_239 wl_222 vdd gnd cell_6t
Xbit_r223_c239 bl_239 br_239 wl_223 vdd gnd cell_6t
Xbit_r224_c239 bl_239 br_239 wl_224 vdd gnd cell_6t
Xbit_r225_c239 bl_239 br_239 wl_225 vdd gnd cell_6t
Xbit_r226_c239 bl_239 br_239 wl_226 vdd gnd cell_6t
Xbit_r227_c239 bl_239 br_239 wl_227 vdd gnd cell_6t
Xbit_r228_c239 bl_239 br_239 wl_228 vdd gnd cell_6t
Xbit_r229_c239 bl_239 br_239 wl_229 vdd gnd cell_6t
Xbit_r230_c239 bl_239 br_239 wl_230 vdd gnd cell_6t
Xbit_r231_c239 bl_239 br_239 wl_231 vdd gnd cell_6t
Xbit_r232_c239 bl_239 br_239 wl_232 vdd gnd cell_6t
Xbit_r233_c239 bl_239 br_239 wl_233 vdd gnd cell_6t
Xbit_r234_c239 bl_239 br_239 wl_234 vdd gnd cell_6t
Xbit_r235_c239 bl_239 br_239 wl_235 vdd gnd cell_6t
Xbit_r236_c239 bl_239 br_239 wl_236 vdd gnd cell_6t
Xbit_r237_c239 bl_239 br_239 wl_237 vdd gnd cell_6t
Xbit_r238_c239 bl_239 br_239 wl_238 vdd gnd cell_6t
Xbit_r239_c239 bl_239 br_239 wl_239 vdd gnd cell_6t
Xbit_r240_c239 bl_239 br_239 wl_240 vdd gnd cell_6t
Xbit_r241_c239 bl_239 br_239 wl_241 vdd gnd cell_6t
Xbit_r242_c239 bl_239 br_239 wl_242 vdd gnd cell_6t
Xbit_r243_c239 bl_239 br_239 wl_243 vdd gnd cell_6t
Xbit_r244_c239 bl_239 br_239 wl_244 vdd gnd cell_6t
Xbit_r245_c239 bl_239 br_239 wl_245 vdd gnd cell_6t
Xbit_r246_c239 bl_239 br_239 wl_246 vdd gnd cell_6t
Xbit_r247_c239 bl_239 br_239 wl_247 vdd gnd cell_6t
Xbit_r248_c239 bl_239 br_239 wl_248 vdd gnd cell_6t
Xbit_r249_c239 bl_239 br_239 wl_249 vdd gnd cell_6t
Xbit_r250_c239 bl_239 br_239 wl_250 vdd gnd cell_6t
Xbit_r251_c239 bl_239 br_239 wl_251 vdd gnd cell_6t
Xbit_r252_c239 bl_239 br_239 wl_252 vdd gnd cell_6t
Xbit_r253_c239 bl_239 br_239 wl_253 vdd gnd cell_6t
Xbit_r254_c239 bl_239 br_239 wl_254 vdd gnd cell_6t
Xbit_r255_c239 bl_239 br_239 wl_255 vdd gnd cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd cell_6t
Xbit_r1_c240 bl_240 br_240 wl_1 vdd gnd cell_6t
Xbit_r2_c240 bl_240 br_240 wl_2 vdd gnd cell_6t
Xbit_r3_c240 bl_240 br_240 wl_3 vdd gnd cell_6t
Xbit_r4_c240 bl_240 br_240 wl_4 vdd gnd cell_6t
Xbit_r5_c240 bl_240 br_240 wl_5 vdd gnd cell_6t
Xbit_r6_c240 bl_240 br_240 wl_6 vdd gnd cell_6t
Xbit_r7_c240 bl_240 br_240 wl_7 vdd gnd cell_6t
Xbit_r8_c240 bl_240 br_240 wl_8 vdd gnd cell_6t
Xbit_r9_c240 bl_240 br_240 wl_9 vdd gnd cell_6t
Xbit_r10_c240 bl_240 br_240 wl_10 vdd gnd cell_6t
Xbit_r11_c240 bl_240 br_240 wl_11 vdd gnd cell_6t
Xbit_r12_c240 bl_240 br_240 wl_12 vdd gnd cell_6t
Xbit_r13_c240 bl_240 br_240 wl_13 vdd gnd cell_6t
Xbit_r14_c240 bl_240 br_240 wl_14 vdd gnd cell_6t
Xbit_r15_c240 bl_240 br_240 wl_15 vdd gnd cell_6t
Xbit_r16_c240 bl_240 br_240 wl_16 vdd gnd cell_6t
Xbit_r17_c240 bl_240 br_240 wl_17 vdd gnd cell_6t
Xbit_r18_c240 bl_240 br_240 wl_18 vdd gnd cell_6t
Xbit_r19_c240 bl_240 br_240 wl_19 vdd gnd cell_6t
Xbit_r20_c240 bl_240 br_240 wl_20 vdd gnd cell_6t
Xbit_r21_c240 bl_240 br_240 wl_21 vdd gnd cell_6t
Xbit_r22_c240 bl_240 br_240 wl_22 vdd gnd cell_6t
Xbit_r23_c240 bl_240 br_240 wl_23 vdd gnd cell_6t
Xbit_r24_c240 bl_240 br_240 wl_24 vdd gnd cell_6t
Xbit_r25_c240 bl_240 br_240 wl_25 vdd gnd cell_6t
Xbit_r26_c240 bl_240 br_240 wl_26 vdd gnd cell_6t
Xbit_r27_c240 bl_240 br_240 wl_27 vdd gnd cell_6t
Xbit_r28_c240 bl_240 br_240 wl_28 vdd gnd cell_6t
Xbit_r29_c240 bl_240 br_240 wl_29 vdd gnd cell_6t
Xbit_r30_c240 bl_240 br_240 wl_30 vdd gnd cell_6t
Xbit_r31_c240 bl_240 br_240 wl_31 vdd gnd cell_6t
Xbit_r32_c240 bl_240 br_240 wl_32 vdd gnd cell_6t
Xbit_r33_c240 bl_240 br_240 wl_33 vdd gnd cell_6t
Xbit_r34_c240 bl_240 br_240 wl_34 vdd gnd cell_6t
Xbit_r35_c240 bl_240 br_240 wl_35 vdd gnd cell_6t
Xbit_r36_c240 bl_240 br_240 wl_36 vdd gnd cell_6t
Xbit_r37_c240 bl_240 br_240 wl_37 vdd gnd cell_6t
Xbit_r38_c240 bl_240 br_240 wl_38 vdd gnd cell_6t
Xbit_r39_c240 bl_240 br_240 wl_39 vdd gnd cell_6t
Xbit_r40_c240 bl_240 br_240 wl_40 vdd gnd cell_6t
Xbit_r41_c240 bl_240 br_240 wl_41 vdd gnd cell_6t
Xbit_r42_c240 bl_240 br_240 wl_42 vdd gnd cell_6t
Xbit_r43_c240 bl_240 br_240 wl_43 vdd gnd cell_6t
Xbit_r44_c240 bl_240 br_240 wl_44 vdd gnd cell_6t
Xbit_r45_c240 bl_240 br_240 wl_45 vdd gnd cell_6t
Xbit_r46_c240 bl_240 br_240 wl_46 vdd gnd cell_6t
Xbit_r47_c240 bl_240 br_240 wl_47 vdd gnd cell_6t
Xbit_r48_c240 bl_240 br_240 wl_48 vdd gnd cell_6t
Xbit_r49_c240 bl_240 br_240 wl_49 vdd gnd cell_6t
Xbit_r50_c240 bl_240 br_240 wl_50 vdd gnd cell_6t
Xbit_r51_c240 bl_240 br_240 wl_51 vdd gnd cell_6t
Xbit_r52_c240 bl_240 br_240 wl_52 vdd gnd cell_6t
Xbit_r53_c240 bl_240 br_240 wl_53 vdd gnd cell_6t
Xbit_r54_c240 bl_240 br_240 wl_54 vdd gnd cell_6t
Xbit_r55_c240 bl_240 br_240 wl_55 vdd gnd cell_6t
Xbit_r56_c240 bl_240 br_240 wl_56 vdd gnd cell_6t
Xbit_r57_c240 bl_240 br_240 wl_57 vdd gnd cell_6t
Xbit_r58_c240 bl_240 br_240 wl_58 vdd gnd cell_6t
Xbit_r59_c240 bl_240 br_240 wl_59 vdd gnd cell_6t
Xbit_r60_c240 bl_240 br_240 wl_60 vdd gnd cell_6t
Xbit_r61_c240 bl_240 br_240 wl_61 vdd gnd cell_6t
Xbit_r62_c240 bl_240 br_240 wl_62 vdd gnd cell_6t
Xbit_r63_c240 bl_240 br_240 wl_63 vdd gnd cell_6t
Xbit_r64_c240 bl_240 br_240 wl_64 vdd gnd cell_6t
Xbit_r65_c240 bl_240 br_240 wl_65 vdd gnd cell_6t
Xbit_r66_c240 bl_240 br_240 wl_66 vdd gnd cell_6t
Xbit_r67_c240 bl_240 br_240 wl_67 vdd gnd cell_6t
Xbit_r68_c240 bl_240 br_240 wl_68 vdd gnd cell_6t
Xbit_r69_c240 bl_240 br_240 wl_69 vdd gnd cell_6t
Xbit_r70_c240 bl_240 br_240 wl_70 vdd gnd cell_6t
Xbit_r71_c240 bl_240 br_240 wl_71 vdd gnd cell_6t
Xbit_r72_c240 bl_240 br_240 wl_72 vdd gnd cell_6t
Xbit_r73_c240 bl_240 br_240 wl_73 vdd gnd cell_6t
Xbit_r74_c240 bl_240 br_240 wl_74 vdd gnd cell_6t
Xbit_r75_c240 bl_240 br_240 wl_75 vdd gnd cell_6t
Xbit_r76_c240 bl_240 br_240 wl_76 vdd gnd cell_6t
Xbit_r77_c240 bl_240 br_240 wl_77 vdd gnd cell_6t
Xbit_r78_c240 bl_240 br_240 wl_78 vdd gnd cell_6t
Xbit_r79_c240 bl_240 br_240 wl_79 vdd gnd cell_6t
Xbit_r80_c240 bl_240 br_240 wl_80 vdd gnd cell_6t
Xbit_r81_c240 bl_240 br_240 wl_81 vdd gnd cell_6t
Xbit_r82_c240 bl_240 br_240 wl_82 vdd gnd cell_6t
Xbit_r83_c240 bl_240 br_240 wl_83 vdd gnd cell_6t
Xbit_r84_c240 bl_240 br_240 wl_84 vdd gnd cell_6t
Xbit_r85_c240 bl_240 br_240 wl_85 vdd gnd cell_6t
Xbit_r86_c240 bl_240 br_240 wl_86 vdd gnd cell_6t
Xbit_r87_c240 bl_240 br_240 wl_87 vdd gnd cell_6t
Xbit_r88_c240 bl_240 br_240 wl_88 vdd gnd cell_6t
Xbit_r89_c240 bl_240 br_240 wl_89 vdd gnd cell_6t
Xbit_r90_c240 bl_240 br_240 wl_90 vdd gnd cell_6t
Xbit_r91_c240 bl_240 br_240 wl_91 vdd gnd cell_6t
Xbit_r92_c240 bl_240 br_240 wl_92 vdd gnd cell_6t
Xbit_r93_c240 bl_240 br_240 wl_93 vdd gnd cell_6t
Xbit_r94_c240 bl_240 br_240 wl_94 vdd gnd cell_6t
Xbit_r95_c240 bl_240 br_240 wl_95 vdd gnd cell_6t
Xbit_r96_c240 bl_240 br_240 wl_96 vdd gnd cell_6t
Xbit_r97_c240 bl_240 br_240 wl_97 vdd gnd cell_6t
Xbit_r98_c240 bl_240 br_240 wl_98 vdd gnd cell_6t
Xbit_r99_c240 bl_240 br_240 wl_99 vdd gnd cell_6t
Xbit_r100_c240 bl_240 br_240 wl_100 vdd gnd cell_6t
Xbit_r101_c240 bl_240 br_240 wl_101 vdd gnd cell_6t
Xbit_r102_c240 bl_240 br_240 wl_102 vdd gnd cell_6t
Xbit_r103_c240 bl_240 br_240 wl_103 vdd gnd cell_6t
Xbit_r104_c240 bl_240 br_240 wl_104 vdd gnd cell_6t
Xbit_r105_c240 bl_240 br_240 wl_105 vdd gnd cell_6t
Xbit_r106_c240 bl_240 br_240 wl_106 vdd gnd cell_6t
Xbit_r107_c240 bl_240 br_240 wl_107 vdd gnd cell_6t
Xbit_r108_c240 bl_240 br_240 wl_108 vdd gnd cell_6t
Xbit_r109_c240 bl_240 br_240 wl_109 vdd gnd cell_6t
Xbit_r110_c240 bl_240 br_240 wl_110 vdd gnd cell_6t
Xbit_r111_c240 bl_240 br_240 wl_111 vdd gnd cell_6t
Xbit_r112_c240 bl_240 br_240 wl_112 vdd gnd cell_6t
Xbit_r113_c240 bl_240 br_240 wl_113 vdd gnd cell_6t
Xbit_r114_c240 bl_240 br_240 wl_114 vdd gnd cell_6t
Xbit_r115_c240 bl_240 br_240 wl_115 vdd gnd cell_6t
Xbit_r116_c240 bl_240 br_240 wl_116 vdd gnd cell_6t
Xbit_r117_c240 bl_240 br_240 wl_117 vdd gnd cell_6t
Xbit_r118_c240 bl_240 br_240 wl_118 vdd gnd cell_6t
Xbit_r119_c240 bl_240 br_240 wl_119 vdd gnd cell_6t
Xbit_r120_c240 bl_240 br_240 wl_120 vdd gnd cell_6t
Xbit_r121_c240 bl_240 br_240 wl_121 vdd gnd cell_6t
Xbit_r122_c240 bl_240 br_240 wl_122 vdd gnd cell_6t
Xbit_r123_c240 bl_240 br_240 wl_123 vdd gnd cell_6t
Xbit_r124_c240 bl_240 br_240 wl_124 vdd gnd cell_6t
Xbit_r125_c240 bl_240 br_240 wl_125 vdd gnd cell_6t
Xbit_r126_c240 bl_240 br_240 wl_126 vdd gnd cell_6t
Xbit_r127_c240 bl_240 br_240 wl_127 vdd gnd cell_6t
Xbit_r128_c240 bl_240 br_240 wl_128 vdd gnd cell_6t
Xbit_r129_c240 bl_240 br_240 wl_129 vdd gnd cell_6t
Xbit_r130_c240 bl_240 br_240 wl_130 vdd gnd cell_6t
Xbit_r131_c240 bl_240 br_240 wl_131 vdd gnd cell_6t
Xbit_r132_c240 bl_240 br_240 wl_132 vdd gnd cell_6t
Xbit_r133_c240 bl_240 br_240 wl_133 vdd gnd cell_6t
Xbit_r134_c240 bl_240 br_240 wl_134 vdd gnd cell_6t
Xbit_r135_c240 bl_240 br_240 wl_135 vdd gnd cell_6t
Xbit_r136_c240 bl_240 br_240 wl_136 vdd gnd cell_6t
Xbit_r137_c240 bl_240 br_240 wl_137 vdd gnd cell_6t
Xbit_r138_c240 bl_240 br_240 wl_138 vdd gnd cell_6t
Xbit_r139_c240 bl_240 br_240 wl_139 vdd gnd cell_6t
Xbit_r140_c240 bl_240 br_240 wl_140 vdd gnd cell_6t
Xbit_r141_c240 bl_240 br_240 wl_141 vdd gnd cell_6t
Xbit_r142_c240 bl_240 br_240 wl_142 vdd gnd cell_6t
Xbit_r143_c240 bl_240 br_240 wl_143 vdd gnd cell_6t
Xbit_r144_c240 bl_240 br_240 wl_144 vdd gnd cell_6t
Xbit_r145_c240 bl_240 br_240 wl_145 vdd gnd cell_6t
Xbit_r146_c240 bl_240 br_240 wl_146 vdd gnd cell_6t
Xbit_r147_c240 bl_240 br_240 wl_147 vdd gnd cell_6t
Xbit_r148_c240 bl_240 br_240 wl_148 vdd gnd cell_6t
Xbit_r149_c240 bl_240 br_240 wl_149 vdd gnd cell_6t
Xbit_r150_c240 bl_240 br_240 wl_150 vdd gnd cell_6t
Xbit_r151_c240 bl_240 br_240 wl_151 vdd gnd cell_6t
Xbit_r152_c240 bl_240 br_240 wl_152 vdd gnd cell_6t
Xbit_r153_c240 bl_240 br_240 wl_153 vdd gnd cell_6t
Xbit_r154_c240 bl_240 br_240 wl_154 vdd gnd cell_6t
Xbit_r155_c240 bl_240 br_240 wl_155 vdd gnd cell_6t
Xbit_r156_c240 bl_240 br_240 wl_156 vdd gnd cell_6t
Xbit_r157_c240 bl_240 br_240 wl_157 vdd gnd cell_6t
Xbit_r158_c240 bl_240 br_240 wl_158 vdd gnd cell_6t
Xbit_r159_c240 bl_240 br_240 wl_159 vdd gnd cell_6t
Xbit_r160_c240 bl_240 br_240 wl_160 vdd gnd cell_6t
Xbit_r161_c240 bl_240 br_240 wl_161 vdd gnd cell_6t
Xbit_r162_c240 bl_240 br_240 wl_162 vdd gnd cell_6t
Xbit_r163_c240 bl_240 br_240 wl_163 vdd gnd cell_6t
Xbit_r164_c240 bl_240 br_240 wl_164 vdd gnd cell_6t
Xbit_r165_c240 bl_240 br_240 wl_165 vdd gnd cell_6t
Xbit_r166_c240 bl_240 br_240 wl_166 vdd gnd cell_6t
Xbit_r167_c240 bl_240 br_240 wl_167 vdd gnd cell_6t
Xbit_r168_c240 bl_240 br_240 wl_168 vdd gnd cell_6t
Xbit_r169_c240 bl_240 br_240 wl_169 vdd gnd cell_6t
Xbit_r170_c240 bl_240 br_240 wl_170 vdd gnd cell_6t
Xbit_r171_c240 bl_240 br_240 wl_171 vdd gnd cell_6t
Xbit_r172_c240 bl_240 br_240 wl_172 vdd gnd cell_6t
Xbit_r173_c240 bl_240 br_240 wl_173 vdd gnd cell_6t
Xbit_r174_c240 bl_240 br_240 wl_174 vdd gnd cell_6t
Xbit_r175_c240 bl_240 br_240 wl_175 vdd gnd cell_6t
Xbit_r176_c240 bl_240 br_240 wl_176 vdd gnd cell_6t
Xbit_r177_c240 bl_240 br_240 wl_177 vdd gnd cell_6t
Xbit_r178_c240 bl_240 br_240 wl_178 vdd gnd cell_6t
Xbit_r179_c240 bl_240 br_240 wl_179 vdd gnd cell_6t
Xbit_r180_c240 bl_240 br_240 wl_180 vdd gnd cell_6t
Xbit_r181_c240 bl_240 br_240 wl_181 vdd gnd cell_6t
Xbit_r182_c240 bl_240 br_240 wl_182 vdd gnd cell_6t
Xbit_r183_c240 bl_240 br_240 wl_183 vdd gnd cell_6t
Xbit_r184_c240 bl_240 br_240 wl_184 vdd gnd cell_6t
Xbit_r185_c240 bl_240 br_240 wl_185 vdd gnd cell_6t
Xbit_r186_c240 bl_240 br_240 wl_186 vdd gnd cell_6t
Xbit_r187_c240 bl_240 br_240 wl_187 vdd gnd cell_6t
Xbit_r188_c240 bl_240 br_240 wl_188 vdd gnd cell_6t
Xbit_r189_c240 bl_240 br_240 wl_189 vdd gnd cell_6t
Xbit_r190_c240 bl_240 br_240 wl_190 vdd gnd cell_6t
Xbit_r191_c240 bl_240 br_240 wl_191 vdd gnd cell_6t
Xbit_r192_c240 bl_240 br_240 wl_192 vdd gnd cell_6t
Xbit_r193_c240 bl_240 br_240 wl_193 vdd gnd cell_6t
Xbit_r194_c240 bl_240 br_240 wl_194 vdd gnd cell_6t
Xbit_r195_c240 bl_240 br_240 wl_195 vdd gnd cell_6t
Xbit_r196_c240 bl_240 br_240 wl_196 vdd gnd cell_6t
Xbit_r197_c240 bl_240 br_240 wl_197 vdd gnd cell_6t
Xbit_r198_c240 bl_240 br_240 wl_198 vdd gnd cell_6t
Xbit_r199_c240 bl_240 br_240 wl_199 vdd gnd cell_6t
Xbit_r200_c240 bl_240 br_240 wl_200 vdd gnd cell_6t
Xbit_r201_c240 bl_240 br_240 wl_201 vdd gnd cell_6t
Xbit_r202_c240 bl_240 br_240 wl_202 vdd gnd cell_6t
Xbit_r203_c240 bl_240 br_240 wl_203 vdd gnd cell_6t
Xbit_r204_c240 bl_240 br_240 wl_204 vdd gnd cell_6t
Xbit_r205_c240 bl_240 br_240 wl_205 vdd gnd cell_6t
Xbit_r206_c240 bl_240 br_240 wl_206 vdd gnd cell_6t
Xbit_r207_c240 bl_240 br_240 wl_207 vdd gnd cell_6t
Xbit_r208_c240 bl_240 br_240 wl_208 vdd gnd cell_6t
Xbit_r209_c240 bl_240 br_240 wl_209 vdd gnd cell_6t
Xbit_r210_c240 bl_240 br_240 wl_210 vdd gnd cell_6t
Xbit_r211_c240 bl_240 br_240 wl_211 vdd gnd cell_6t
Xbit_r212_c240 bl_240 br_240 wl_212 vdd gnd cell_6t
Xbit_r213_c240 bl_240 br_240 wl_213 vdd gnd cell_6t
Xbit_r214_c240 bl_240 br_240 wl_214 vdd gnd cell_6t
Xbit_r215_c240 bl_240 br_240 wl_215 vdd gnd cell_6t
Xbit_r216_c240 bl_240 br_240 wl_216 vdd gnd cell_6t
Xbit_r217_c240 bl_240 br_240 wl_217 vdd gnd cell_6t
Xbit_r218_c240 bl_240 br_240 wl_218 vdd gnd cell_6t
Xbit_r219_c240 bl_240 br_240 wl_219 vdd gnd cell_6t
Xbit_r220_c240 bl_240 br_240 wl_220 vdd gnd cell_6t
Xbit_r221_c240 bl_240 br_240 wl_221 vdd gnd cell_6t
Xbit_r222_c240 bl_240 br_240 wl_222 vdd gnd cell_6t
Xbit_r223_c240 bl_240 br_240 wl_223 vdd gnd cell_6t
Xbit_r224_c240 bl_240 br_240 wl_224 vdd gnd cell_6t
Xbit_r225_c240 bl_240 br_240 wl_225 vdd gnd cell_6t
Xbit_r226_c240 bl_240 br_240 wl_226 vdd gnd cell_6t
Xbit_r227_c240 bl_240 br_240 wl_227 vdd gnd cell_6t
Xbit_r228_c240 bl_240 br_240 wl_228 vdd gnd cell_6t
Xbit_r229_c240 bl_240 br_240 wl_229 vdd gnd cell_6t
Xbit_r230_c240 bl_240 br_240 wl_230 vdd gnd cell_6t
Xbit_r231_c240 bl_240 br_240 wl_231 vdd gnd cell_6t
Xbit_r232_c240 bl_240 br_240 wl_232 vdd gnd cell_6t
Xbit_r233_c240 bl_240 br_240 wl_233 vdd gnd cell_6t
Xbit_r234_c240 bl_240 br_240 wl_234 vdd gnd cell_6t
Xbit_r235_c240 bl_240 br_240 wl_235 vdd gnd cell_6t
Xbit_r236_c240 bl_240 br_240 wl_236 vdd gnd cell_6t
Xbit_r237_c240 bl_240 br_240 wl_237 vdd gnd cell_6t
Xbit_r238_c240 bl_240 br_240 wl_238 vdd gnd cell_6t
Xbit_r239_c240 bl_240 br_240 wl_239 vdd gnd cell_6t
Xbit_r240_c240 bl_240 br_240 wl_240 vdd gnd cell_6t
Xbit_r241_c240 bl_240 br_240 wl_241 vdd gnd cell_6t
Xbit_r242_c240 bl_240 br_240 wl_242 vdd gnd cell_6t
Xbit_r243_c240 bl_240 br_240 wl_243 vdd gnd cell_6t
Xbit_r244_c240 bl_240 br_240 wl_244 vdd gnd cell_6t
Xbit_r245_c240 bl_240 br_240 wl_245 vdd gnd cell_6t
Xbit_r246_c240 bl_240 br_240 wl_246 vdd gnd cell_6t
Xbit_r247_c240 bl_240 br_240 wl_247 vdd gnd cell_6t
Xbit_r248_c240 bl_240 br_240 wl_248 vdd gnd cell_6t
Xbit_r249_c240 bl_240 br_240 wl_249 vdd gnd cell_6t
Xbit_r250_c240 bl_240 br_240 wl_250 vdd gnd cell_6t
Xbit_r251_c240 bl_240 br_240 wl_251 vdd gnd cell_6t
Xbit_r252_c240 bl_240 br_240 wl_252 vdd gnd cell_6t
Xbit_r253_c240 bl_240 br_240 wl_253 vdd gnd cell_6t
Xbit_r254_c240 bl_240 br_240 wl_254 vdd gnd cell_6t
Xbit_r255_c240 bl_240 br_240 wl_255 vdd gnd cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd cell_6t
Xbit_r1_c241 bl_241 br_241 wl_1 vdd gnd cell_6t
Xbit_r2_c241 bl_241 br_241 wl_2 vdd gnd cell_6t
Xbit_r3_c241 bl_241 br_241 wl_3 vdd gnd cell_6t
Xbit_r4_c241 bl_241 br_241 wl_4 vdd gnd cell_6t
Xbit_r5_c241 bl_241 br_241 wl_5 vdd gnd cell_6t
Xbit_r6_c241 bl_241 br_241 wl_6 vdd gnd cell_6t
Xbit_r7_c241 bl_241 br_241 wl_7 vdd gnd cell_6t
Xbit_r8_c241 bl_241 br_241 wl_8 vdd gnd cell_6t
Xbit_r9_c241 bl_241 br_241 wl_9 vdd gnd cell_6t
Xbit_r10_c241 bl_241 br_241 wl_10 vdd gnd cell_6t
Xbit_r11_c241 bl_241 br_241 wl_11 vdd gnd cell_6t
Xbit_r12_c241 bl_241 br_241 wl_12 vdd gnd cell_6t
Xbit_r13_c241 bl_241 br_241 wl_13 vdd gnd cell_6t
Xbit_r14_c241 bl_241 br_241 wl_14 vdd gnd cell_6t
Xbit_r15_c241 bl_241 br_241 wl_15 vdd gnd cell_6t
Xbit_r16_c241 bl_241 br_241 wl_16 vdd gnd cell_6t
Xbit_r17_c241 bl_241 br_241 wl_17 vdd gnd cell_6t
Xbit_r18_c241 bl_241 br_241 wl_18 vdd gnd cell_6t
Xbit_r19_c241 bl_241 br_241 wl_19 vdd gnd cell_6t
Xbit_r20_c241 bl_241 br_241 wl_20 vdd gnd cell_6t
Xbit_r21_c241 bl_241 br_241 wl_21 vdd gnd cell_6t
Xbit_r22_c241 bl_241 br_241 wl_22 vdd gnd cell_6t
Xbit_r23_c241 bl_241 br_241 wl_23 vdd gnd cell_6t
Xbit_r24_c241 bl_241 br_241 wl_24 vdd gnd cell_6t
Xbit_r25_c241 bl_241 br_241 wl_25 vdd gnd cell_6t
Xbit_r26_c241 bl_241 br_241 wl_26 vdd gnd cell_6t
Xbit_r27_c241 bl_241 br_241 wl_27 vdd gnd cell_6t
Xbit_r28_c241 bl_241 br_241 wl_28 vdd gnd cell_6t
Xbit_r29_c241 bl_241 br_241 wl_29 vdd gnd cell_6t
Xbit_r30_c241 bl_241 br_241 wl_30 vdd gnd cell_6t
Xbit_r31_c241 bl_241 br_241 wl_31 vdd gnd cell_6t
Xbit_r32_c241 bl_241 br_241 wl_32 vdd gnd cell_6t
Xbit_r33_c241 bl_241 br_241 wl_33 vdd gnd cell_6t
Xbit_r34_c241 bl_241 br_241 wl_34 vdd gnd cell_6t
Xbit_r35_c241 bl_241 br_241 wl_35 vdd gnd cell_6t
Xbit_r36_c241 bl_241 br_241 wl_36 vdd gnd cell_6t
Xbit_r37_c241 bl_241 br_241 wl_37 vdd gnd cell_6t
Xbit_r38_c241 bl_241 br_241 wl_38 vdd gnd cell_6t
Xbit_r39_c241 bl_241 br_241 wl_39 vdd gnd cell_6t
Xbit_r40_c241 bl_241 br_241 wl_40 vdd gnd cell_6t
Xbit_r41_c241 bl_241 br_241 wl_41 vdd gnd cell_6t
Xbit_r42_c241 bl_241 br_241 wl_42 vdd gnd cell_6t
Xbit_r43_c241 bl_241 br_241 wl_43 vdd gnd cell_6t
Xbit_r44_c241 bl_241 br_241 wl_44 vdd gnd cell_6t
Xbit_r45_c241 bl_241 br_241 wl_45 vdd gnd cell_6t
Xbit_r46_c241 bl_241 br_241 wl_46 vdd gnd cell_6t
Xbit_r47_c241 bl_241 br_241 wl_47 vdd gnd cell_6t
Xbit_r48_c241 bl_241 br_241 wl_48 vdd gnd cell_6t
Xbit_r49_c241 bl_241 br_241 wl_49 vdd gnd cell_6t
Xbit_r50_c241 bl_241 br_241 wl_50 vdd gnd cell_6t
Xbit_r51_c241 bl_241 br_241 wl_51 vdd gnd cell_6t
Xbit_r52_c241 bl_241 br_241 wl_52 vdd gnd cell_6t
Xbit_r53_c241 bl_241 br_241 wl_53 vdd gnd cell_6t
Xbit_r54_c241 bl_241 br_241 wl_54 vdd gnd cell_6t
Xbit_r55_c241 bl_241 br_241 wl_55 vdd gnd cell_6t
Xbit_r56_c241 bl_241 br_241 wl_56 vdd gnd cell_6t
Xbit_r57_c241 bl_241 br_241 wl_57 vdd gnd cell_6t
Xbit_r58_c241 bl_241 br_241 wl_58 vdd gnd cell_6t
Xbit_r59_c241 bl_241 br_241 wl_59 vdd gnd cell_6t
Xbit_r60_c241 bl_241 br_241 wl_60 vdd gnd cell_6t
Xbit_r61_c241 bl_241 br_241 wl_61 vdd gnd cell_6t
Xbit_r62_c241 bl_241 br_241 wl_62 vdd gnd cell_6t
Xbit_r63_c241 bl_241 br_241 wl_63 vdd gnd cell_6t
Xbit_r64_c241 bl_241 br_241 wl_64 vdd gnd cell_6t
Xbit_r65_c241 bl_241 br_241 wl_65 vdd gnd cell_6t
Xbit_r66_c241 bl_241 br_241 wl_66 vdd gnd cell_6t
Xbit_r67_c241 bl_241 br_241 wl_67 vdd gnd cell_6t
Xbit_r68_c241 bl_241 br_241 wl_68 vdd gnd cell_6t
Xbit_r69_c241 bl_241 br_241 wl_69 vdd gnd cell_6t
Xbit_r70_c241 bl_241 br_241 wl_70 vdd gnd cell_6t
Xbit_r71_c241 bl_241 br_241 wl_71 vdd gnd cell_6t
Xbit_r72_c241 bl_241 br_241 wl_72 vdd gnd cell_6t
Xbit_r73_c241 bl_241 br_241 wl_73 vdd gnd cell_6t
Xbit_r74_c241 bl_241 br_241 wl_74 vdd gnd cell_6t
Xbit_r75_c241 bl_241 br_241 wl_75 vdd gnd cell_6t
Xbit_r76_c241 bl_241 br_241 wl_76 vdd gnd cell_6t
Xbit_r77_c241 bl_241 br_241 wl_77 vdd gnd cell_6t
Xbit_r78_c241 bl_241 br_241 wl_78 vdd gnd cell_6t
Xbit_r79_c241 bl_241 br_241 wl_79 vdd gnd cell_6t
Xbit_r80_c241 bl_241 br_241 wl_80 vdd gnd cell_6t
Xbit_r81_c241 bl_241 br_241 wl_81 vdd gnd cell_6t
Xbit_r82_c241 bl_241 br_241 wl_82 vdd gnd cell_6t
Xbit_r83_c241 bl_241 br_241 wl_83 vdd gnd cell_6t
Xbit_r84_c241 bl_241 br_241 wl_84 vdd gnd cell_6t
Xbit_r85_c241 bl_241 br_241 wl_85 vdd gnd cell_6t
Xbit_r86_c241 bl_241 br_241 wl_86 vdd gnd cell_6t
Xbit_r87_c241 bl_241 br_241 wl_87 vdd gnd cell_6t
Xbit_r88_c241 bl_241 br_241 wl_88 vdd gnd cell_6t
Xbit_r89_c241 bl_241 br_241 wl_89 vdd gnd cell_6t
Xbit_r90_c241 bl_241 br_241 wl_90 vdd gnd cell_6t
Xbit_r91_c241 bl_241 br_241 wl_91 vdd gnd cell_6t
Xbit_r92_c241 bl_241 br_241 wl_92 vdd gnd cell_6t
Xbit_r93_c241 bl_241 br_241 wl_93 vdd gnd cell_6t
Xbit_r94_c241 bl_241 br_241 wl_94 vdd gnd cell_6t
Xbit_r95_c241 bl_241 br_241 wl_95 vdd gnd cell_6t
Xbit_r96_c241 bl_241 br_241 wl_96 vdd gnd cell_6t
Xbit_r97_c241 bl_241 br_241 wl_97 vdd gnd cell_6t
Xbit_r98_c241 bl_241 br_241 wl_98 vdd gnd cell_6t
Xbit_r99_c241 bl_241 br_241 wl_99 vdd gnd cell_6t
Xbit_r100_c241 bl_241 br_241 wl_100 vdd gnd cell_6t
Xbit_r101_c241 bl_241 br_241 wl_101 vdd gnd cell_6t
Xbit_r102_c241 bl_241 br_241 wl_102 vdd gnd cell_6t
Xbit_r103_c241 bl_241 br_241 wl_103 vdd gnd cell_6t
Xbit_r104_c241 bl_241 br_241 wl_104 vdd gnd cell_6t
Xbit_r105_c241 bl_241 br_241 wl_105 vdd gnd cell_6t
Xbit_r106_c241 bl_241 br_241 wl_106 vdd gnd cell_6t
Xbit_r107_c241 bl_241 br_241 wl_107 vdd gnd cell_6t
Xbit_r108_c241 bl_241 br_241 wl_108 vdd gnd cell_6t
Xbit_r109_c241 bl_241 br_241 wl_109 vdd gnd cell_6t
Xbit_r110_c241 bl_241 br_241 wl_110 vdd gnd cell_6t
Xbit_r111_c241 bl_241 br_241 wl_111 vdd gnd cell_6t
Xbit_r112_c241 bl_241 br_241 wl_112 vdd gnd cell_6t
Xbit_r113_c241 bl_241 br_241 wl_113 vdd gnd cell_6t
Xbit_r114_c241 bl_241 br_241 wl_114 vdd gnd cell_6t
Xbit_r115_c241 bl_241 br_241 wl_115 vdd gnd cell_6t
Xbit_r116_c241 bl_241 br_241 wl_116 vdd gnd cell_6t
Xbit_r117_c241 bl_241 br_241 wl_117 vdd gnd cell_6t
Xbit_r118_c241 bl_241 br_241 wl_118 vdd gnd cell_6t
Xbit_r119_c241 bl_241 br_241 wl_119 vdd gnd cell_6t
Xbit_r120_c241 bl_241 br_241 wl_120 vdd gnd cell_6t
Xbit_r121_c241 bl_241 br_241 wl_121 vdd gnd cell_6t
Xbit_r122_c241 bl_241 br_241 wl_122 vdd gnd cell_6t
Xbit_r123_c241 bl_241 br_241 wl_123 vdd gnd cell_6t
Xbit_r124_c241 bl_241 br_241 wl_124 vdd gnd cell_6t
Xbit_r125_c241 bl_241 br_241 wl_125 vdd gnd cell_6t
Xbit_r126_c241 bl_241 br_241 wl_126 vdd gnd cell_6t
Xbit_r127_c241 bl_241 br_241 wl_127 vdd gnd cell_6t
Xbit_r128_c241 bl_241 br_241 wl_128 vdd gnd cell_6t
Xbit_r129_c241 bl_241 br_241 wl_129 vdd gnd cell_6t
Xbit_r130_c241 bl_241 br_241 wl_130 vdd gnd cell_6t
Xbit_r131_c241 bl_241 br_241 wl_131 vdd gnd cell_6t
Xbit_r132_c241 bl_241 br_241 wl_132 vdd gnd cell_6t
Xbit_r133_c241 bl_241 br_241 wl_133 vdd gnd cell_6t
Xbit_r134_c241 bl_241 br_241 wl_134 vdd gnd cell_6t
Xbit_r135_c241 bl_241 br_241 wl_135 vdd gnd cell_6t
Xbit_r136_c241 bl_241 br_241 wl_136 vdd gnd cell_6t
Xbit_r137_c241 bl_241 br_241 wl_137 vdd gnd cell_6t
Xbit_r138_c241 bl_241 br_241 wl_138 vdd gnd cell_6t
Xbit_r139_c241 bl_241 br_241 wl_139 vdd gnd cell_6t
Xbit_r140_c241 bl_241 br_241 wl_140 vdd gnd cell_6t
Xbit_r141_c241 bl_241 br_241 wl_141 vdd gnd cell_6t
Xbit_r142_c241 bl_241 br_241 wl_142 vdd gnd cell_6t
Xbit_r143_c241 bl_241 br_241 wl_143 vdd gnd cell_6t
Xbit_r144_c241 bl_241 br_241 wl_144 vdd gnd cell_6t
Xbit_r145_c241 bl_241 br_241 wl_145 vdd gnd cell_6t
Xbit_r146_c241 bl_241 br_241 wl_146 vdd gnd cell_6t
Xbit_r147_c241 bl_241 br_241 wl_147 vdd gnd cell_6t
Xbit_r148_c241 bl_241 br_241 wl_148 vdd gnd cell_6t
Xbit_r149_c241 bl_241 br_241 wl_149 vdd gnd cell_6t
Xbit_r150_c241 bl_241 br_241 wl_150 vdd gnd cell_6t
Xbit_r151_c241 bl_241 br_241 wl_151 vdd gnd cell_6t
Xbit_r152_c241 bl_241 br_241 wl_152 vdd gnd cell_6t
Xbit_r153_c241 bl_241 br_241 wl_153 vdd gnd cell_6t
Xbit_r154_c241 bl_241 br_241 wl_154 vdd gnd cell_6t
Xbit_r155_c241 bl_241 br_241 wl_155 vdd gnd cell_6t
Xbit_r156_c241 bl_241 br_241 wl_156 vdd gnd cell_6t
Xbit_r157_c241 bl_241 br_241 wl_157 vdd gnd cell_6t
Xbit_r158_c241 bl_241 br_241 wl_158 vdd gnd cell_6t
Xbit_r159_c241 bl_241 br_241 wl_159 vdd gnd cell_6t
Xbit_r160_c241 bl_241 br_241 wl_160 vdd gnd cell_6t
Xbit_r161_c241 bl_241 br_241 wl_161 vdd gnd cell_6t
Xbit_r162_c241 bl_241 br_241 wl_162 vdd gnd cell_6t
Xbit_r163_c241 bl_241 br_241 wl_163 vdd gnd cell_6t
Xbit_r164_c241 bl_241 br_241 wl_164 vdd gnd cell_6t
Xbit_r165_c241 bl_241 br_241 wl_165 vdd gnd cell_6t
Xbit_r166_c241 bl_241 br_241 wl_166 vdd gnd cell_6t
Xbit_r167_c241 bl_241 br_241 wl_167 vdd gnd cell_6t
Xbit_r168_c241 bl_241 br_241 wl_168 vdd gnd cell_6t
Xbit_r169_c241 bl_241 br_241 wl_169 vdd gnd cell_6t
Xbit_r170_c241 bl_241 br_241 wl_170 vdd gnd cell_6t
Xbit_r171_c241 bl_241 br_241 wl_171 vdd gnd cell_6t
Xbit_r172_c241 bl_241 br_241 wl_172 vdd gnd cell_6t
Xbit_r173_c241 bl_241 br_241 wl_173 vdd gnd cell_6t
Xbit_r174_c241 bl_241 br_241 wl_174 vdd gnd cell_6t
Xbit_r175_c241 bl_241 br_241 wl_175 vdd gnd cell_6t
Xbit_r176_c241 bl_241 br_241 wl_176 vdd gnd cell_6t
Xbit_r177_c241 bl_241 br_241 wl_177 vdd gnd cell_6t
Xbit_r178_c241 bl_241 br_241 wl_178 vdd gnd cell_6t
Xbit_r179_c241 bl_241 br_241 wl_179 vdd gnd cell_6t
Xbit_r180_c241 bl_241 br_241 wl_180 vdd gnd cell_6t
Xbit_r181_c241 bl_241 br_241 wl_181 vdd gnd cell_6t
Xbit_r182_c241 bl_241 br_241 wl_182 vdd gnd cell_6t
Xbit_r183_c241 bl_241 br_241 wl_183 vdd gnd cell_6t
Xbit_r184_c241 bl_241 br_241 wl_184 vdd gnd cell_6t
Xbit_r185_c241 bl_241 br_241 wl_185 vdd gnd cell_6t
Xbit_r186_c241 bl_241 br_241 wl_186 vdd gnd cell_6t
Xbit_r187_c241 bl_241 br_241 wl_187 vdd gnd cell_6t
Xbit_r188_c241 bl_241 br_241 wl_188 vdd gnd cell_6t
Xbit_r189_c241 bl_241 br_241 wl_189 vdd gnd cell_6t
Xbit_r190_c241 bl_241 br_241 wl_190 vdd gnd cell_6t
Xbit_r191_c241 bl_241 br_241 wl_191 vdd gnd cell_6t
Xbit_r192_c241 bl_241 br_241 wl_192 vdd gnd cell_6t
Xbit_r193_c241 bl_241 br_241 wl_193 vdd gnd cell_6t
Xbit_r194_c241 bl_241 br_241 wl_194 vdd gnd cell_6t
Xbit_r195_c241 bl_241 br_241 wl_195 vdd gnd cell_6t
Xbit_r196_c241 bl_241 br_241 wl_196 vdd gnd cell_6t
Xbit_r197_c241 bl_241 br_241 wl_197 vdd gnd cell_6t
Xbit_r198_c241 bl_241 br_241 wl_198 vdd gnd cell_6t
Xbit_r199_c241 bl_241 br_241 wl_199 vdd gnd cell_6t
Xbit_r200_c241 bl_241 br_241 wl_200 vdd gnd cell_6t
Xbit_r201_c241 bl_241 br_241 wl_201 vdd gnd cell_6t
Xbit_r202_c241 bl_241 br_241 wl_202 vdd gnd cell_6t
Xbit_r203_c241 bl_241 br_241 wl_203 vdd gnd cell_6t
Xbit_r204_c241 bl_241 br_241 wl_204 vdd gnd cell_6t
Xbit_r205_c241 bl_241 br_241 wl_205 vdd gnd cell_6t
Xbit_r206_c241 bl_241 br_241 wl_206 vdd gnd cell_6t
Xbit_r207_c241 bl_241 br_241 wl_207 vdd gnd cell_6t
Xbit_r208_c241 bl_241 br_241 wl_208 vdd gnd cell_6t
Xbit_r209_c241 bl_241 br_241 wl_209 vdd gnd cell_6t
Xbit_r210_c241 bl_241 br_241 wl_210 vdd gnd cell_6t
Xbit_r211_c241 bl_241 br_241 wl_211 vdd gnd cell_6t
Xbit_r212_c241 bl_241 br_241 wl_212 vdd gnd cell_6t
Xbit_r213_c241 bl_241 br_241 wl_213 vdd gnd cell_6t
Xbit_r214_c241 bl_241 br_241 wl_214 vdd gnd cell_6t
Xbit_r215_c241 bl_241 br_241 wl_215 vdd gnd cell_6t
Xbit_r216_c241 bl_241 br_241 wl_216 vdd gnd cell_6t
Xbit_r217_c241 bl_241 br_241 wl_217 vdd gnd cell_6t
Xbit_r218_c241 bl_241 br_241 wl_218 vdd gnd cell_6t
Xbit_r219_c241 bl_241 br_241 wl_219 vdd gnd cell_6t
Xbit_r220_c241 bl_241 br_241 wl_220 vdd gnd cell_6t
Xbit_r221_c241 bl_241 br_241 wl_221 vdd gnd cell_6t
Xbit_r222_c241 bl_241 br_241 wl_222 vdd gnd cell_6t
Xbit_r223_c241 bl_241 br_241 wl_223 vdd gnd cell_6t
Xbit_r224_c241 bl_241 br_241 wl_224 vdd gnd cell_6t
Xbit_r225_c241 bl_241 br_241 wl_225 vdd gnd cell_6t
Xbit_r226_c241 bl_241 br_241 wl_226 vdd gnd cell_6t
Xbit_r227_c241 bl_241 br_241 wl_227 vdd gnd cell_6t
Xbit_r228_c241 bl_241 br_241 wl_228 vdd gnd cell_6t
Xbit_r229_c241 bl_241 br_241 wl_229 vdd gnd cell_6t
Xbit_r230_c241 bl_241 br_241 wl_230 vdd gnd cell_6t
Xbit_r231_c241 bl_241 br_241 wl_231 vdd gnd cell_6t
Xbit_r232_c241 bl_241 br_241 wl_232 vdd gnd cell_6t
Xbit_r233_c241 bl_241 br_241 wl_233 vdd gnd cell_6t
Xbit_r234_c241 bl_241 br_241 wl_234 vdd gnd cell_6t
Xbit_r235_c241 bl_241 br_241 wl_235 vdd gnd cell_6t
Xbit_r236_c241 bl_241 br_241 wl_236 vdd gnd cell_6t
Xbit_r237_c241 bl_241 br_241 wl_237 vdd gnd cell_6t
Xbit_r238_c241 bl_241 br_241 wl_238 vdd gnd cell_6t
Xbit_r239_c241 bl_241 br_241 wl_239 vdd gnd cell_6t
Xbit_r240_c241 bl_241 br_241 wl_240 vdd gnd cell_6t
Xbit_r241_c241 bl_241 br_241 wl_241 vdd gnd cell_6t
Xbit_r242_c241 bl_241 br_241 wl_242 vdd gnd cell_6t
Xbit_r243_c241 bl_241 br_241 wl_243 vdd gnd cell_6t
Xbit_r244_c241 bl_241 br_241 wl_244 vdd gnd cell_6t
Xbit_r245_c241 bl_241 br_241 wl_245 vdd gnd cell_6t
Xbit_r246_c241 bl_241 br_241 wl_246 vdd gnd cell_6t
Xbit_r247_c241 bl_241 br_241 wl_247 vdd gnd cell_6t
Xbit_r248_c241 bl_241 br_241 wl_248 vdd gnd cell_6t
Xbit_r249_c241 bl_241 br_241 wl_249 vdd gnd cell_6t
Xbit_r250_c241 bl_241 br_241 wl_250 vdd gnd cell_6t
Xbit_r251_c241 bl_241 br_241 wl_251 vdd gnd cell_6t
Xbit_r252_c241 bl_241 br_241 wl_252 vdd gnd cell_6t
Xbit_r253_c241 bl_241 br_241 wl_253 vdd gnd cell_6t
Xbit_r254_c241 bl_241 br_241 wl_254 vdd gnd cell_6t
Xbit_r255_c241 bl_241 br_241 wl_255 vdd gnd cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd cell_6t
Xbit_r1_c242 bl_242 br_242 wl_1 vdd gnd cell_6t
Xbit_r2_c242 bl_242 br_242 wl_2 vdd gnd cell_6t
Xbit_r3_c242 bl_242 br_242 wl_3 vdd gnd cell_6t
Xbit_r4_c242 bl_242 br_242 wl_4 vdd gnd cell_6t
Xbit_r5_c242 bl_242 br_242 wl_5 vdd gnd cell_6t
Xbit_r6_c242 bl_242 br_242 wl_6 vdd gnd cell_6t
Xbit_r7_c242 bl_242 br_242 wl_7 vdd gnd cell_6t
Xbit_r8_c242 bl_242 br_242 wl_8 vdd gnd cell_6t
Xbit_r9_c242 bl_242 br_242 wl_9 vdd gnd cell_6t
Xbit_r10_c242 bl_242 br_242 wl_10 vdd gnd cell_6t
Xbit_r11_c242 bl_242 br_242 wl_11 vdd gnd cell_6t
Xbit_r12_c242 bl_242 br_242 wl_12 vdd gnd cell_6t
Xbit_r13_c242 bl_242 br_242 wl_13 vdd gnd cell_6t
Xbit_r14_c242 bl_242 br_242 wl_14 vdd gnd cell_6t
Xbit_r15_c242 bl_242 br_242 wl_15 vdd gnd cell_6t
Xbit_r16_c242 bl_242 br_242 wl_16 vdd gnd cell_6t
Xbit_r17_c242 bl_242 br_242 wl_17 vdd gnd cell_6t
Xbit_r18_c242 bl_242 br_242 wl_18 vdd gnd cell_6t
Xbit_r19_c242 bl_242 br_242 wl_19 vdd gnd cell_6t
Xbit_r20_c242 bl_242 br_242 wl_20 vdd gnd cell_6t
Xbit_r21_c242 bl_242 br_242 wl_21 vdd gnd cell_6t
Xbit_r22_c242 bl_242 br_242 wl_22 vdd gnd cell_6t
Xbit_r23_c242 bl_242 br_242 wl_23 vdd gnd cell_6t
Xbit_r24_c242 bl_242 br_242 wl_24 vdd gnd cell_6t
Xbit_r25_c242 bl_242 br_242 wl_25 vdd gnd cell_6t
Xbit_r26_c242 bl_242 br_242 wl_26 vdd gnd cell_6t
Xbit_r27_c242 bl_242 br_242 wl_27 vdd gnd cell_6t
Xbit_r28_c242 bl_242 br_242 wl_28 vdd gnd cell_6t
Xbit_r29_c242 bl_242 br_242 wl_29 vdd gnd cell_6t
Xbit_r30_c242 bl_242 br_242 wl_30 vdd gnd cell_6t
Xbit_r31_c242 bl_242 br_242 wl_31 vdd gnd cell_6t
Xbit_r32_c242 bl_242 br_242 wl_32 vdd gnd cell_6t
Xbit_r33_c242 bl_242 br_242 wl_33 vdd gnd cell_6t
Xbit_r34_c242 bl_242 br_242 wl_34 vdd gnd cell_6t
Xbit_r35_c242 bl_242 br_242 wl_35 vdd gnd cell_6t
Xbit_r36_c242 bl_242 br_242 wl_36 vdd gnd cell_6t
Xbit_r37_c242 bl_242 br_242 wl_37 vdd gnd cell_6t
Xbit_r38_c242 bl_242 br_242 wl_38 vdd gnd cell_6t
Xbit_r39_c242 bl_242 br_242 wl_39 vdd gnd cell_6t
Xbit_r40_c242 bl_242 br_242 wl_40 vdd gnd cell_6t
Xbit_r41_c242 bl_242 br_242 wl_41 vdd gnd cell_6t
Xbit_r42_c242 bl_242 br_242 wl_42 vdd gnd cell_6t
Xbit_r43_c242 bl_242 br_242 wl_43 vdd gnd cell_6t
Xbit_r44_c242 bl_242 br_242 wl_44 vdd gnd cell_6t
Xbit_r45_c242 bl_242 br_242 wl_45 vdd gnd cell_6t
Xbit_r46_c242 bl_242 br_242 wl_46 vdd gnd cell_6t
Xbit_r47_c242 bl_242 br_242 wl_47 vdd gnd cell_6t
Xbit_r48_c242 bl_242 br_242 wl_48 vdd gnd cell_6t
Xbit_r49_c242 bl_242 br_242 wl_49 vdd gnd cell_6t
Xbit_r50_c242 bl_242 br_242 wl_50 vdd gnd cell_6t
Xbit_r51_c242 bl_242 br_242 wl_51 vdd gnd cell_6t
Xbit_r52_c242 bl_242 br_242 wl_52 vdd gnd cell_6t
Xbit_r53_c242 bl_242 br_242 wl_53 vdd gnd cell_6t
Xbit_r54_c242 bl_242 br_242 wl_54 vdd gnd cell_6t
Xbit_r55_c242 bl_242 br_242 wl_55 vdd gnd cell_6t
Xbit_r56_c242 bl_242 br_242 wl_56 vdd gnd cell_6t
Xbit_r57_c242 bl_242 br_242 wl_57 vdd gnd cell_6t
Xbit_r58_c242 bl_242 br_242 wl_58 vdd gnd cell_6t
Xbit_r59_c242 bl_242 br_242 wl_59 vdd gnd cell_6t
Xbit_r60_c242 bl_242 br_242 wl_60 vdd gnd cell_6t
Xbit_r61_c242 bl_242 br_242 wl_61 vdd gnd cell_6t
Xbit_r62_c242 bl_242 br_242 wl_62 vdd gnd cell_6t
Xbit_r63_c242 bl_242 br_242 wl_63 vdd gnd cell_6t
Xbit_r64_c242 bl_242 br_242 wl_64 vdd gnd cell_6t
Xbit_r65_c242 bl_242 br_242 wl_65 vdd gnd cell_6t
Xbit_r66_c242 bl_242 br_242 wl_66 vdd gnd cell_6t
Xbit_r67_c242 bl_242 br_242 wl_67 vdd gnd cell_6t
Xbit_r68_c242 bl_242 br_242 wl_68 vdd gnd cell_6t
Xbit_r69_c242 bl_242 br_242 wl_69 vdd gnd cell_6t
Xbit_r70_c242 bl_242 br_242 wl_70 vdd gnd cell_6t
Xbit_r71_c242 bl_242 br_242 wl_71 vdd gnd cell_6t
Xbit_r72_c242 bl_242 br_242 wl_72 vdd gnd cell_6t
Xbit_r73_c242 bl_242 br_242 wl_73 vdd gnd cell_6t
Xbit_r74_c242 bl_242 br_242 wl_74 vdd gnd cell_6t
Xbit_r75_c242 bl_242 br_242 wl_75 vdd gnd cell_6t
Xbit_r76_c242 bl_242 br_242 wl_76 vdd gnd cell_6t
Xbit_r77_c242 bl_242 br_242 wl_77 vdd gnd cell_6t
Xbit_r78_c242 bl_242 br_242 wl_78 vdd gnd cell_6t
Xbit_r79_c242 bl_242 br_242 wl_79 vdd gnd cell_6t
Xbit_r80_c242 bl_242 br_242 wl_80 vdd gnd cell_6t
Xbit_r81_c242 bl_242 br_242 wl_81 vdd gnd cell_6t
Xbit_r82_c242 bl_242 br_242 wl_82 vdd gnd cell_6t
Xbit_r83_c242 bl_242 br_242 wl_83 vdd gnd cell_6t
Xbit_r84_c242 bl_242 br_242 wl_84 vdd gnd cell_6t
Xbit_r85_c242 bl_242 br_242 wl_85 vdd gnd cell_6t
Xbit_r86_c242 bl_242 br_242 wl_86 vdd gnd cell_6t
Xbit_r87_c242 bl_242 br_242 wl_87 vdd gnd cell_6t
Xbit_r88_c242 bl_242 br_242 wl_88 vdd gnd cell_6t
Xbit_r89_c242 bl_242 br_242 wl_89 vdd gnd cell_6t
Xbit_r90_c242 bl_242 br_242 wl_90 vdd gnd cell_6t
Xbit_r91_c242 bl_242 br_242 wl_91 vdd gnd cell_6t
Xbit_r92_c242 bl_242 br_242 wl_92 vdd gnd cell_6t
Xbit_r93_c242 bl_242 br_242 wl_93 vdd gnd cell_6t
Xbit_r94_c242 bl_242 br_242 wl_94 vdd gnd cell_6t
Xbit_r95_c242 bl_242 br_242 wl_95 vdd gnd cell_6t
Xbit_r96_c242 bl_242 br_242 wl_96 vdd gnd cell_6t
Xbit_r97_c242 bl_242 br_242 wl_97 vdd gnd cell_6t
Xbit_r98_c242 bl_242 br_242 wl_98 vdd gnd cell_6t
Xbit_r99_c242 bl_242 br_242 wl_99 vdd gnd cell_6t
Xbit_r100_c242 bl_242 br_242 wl_100 vdd gnd cell_6t
Xbit_r101_c242 bl_242 br_242 wl_101 vdd gnd cell_6t
Xbit_r102_c242 bl_242 br_242 wl_102 vdd gnd cell_6t
Xbit_r103_c242 bl_242 br_242 wl_103 vdd gnd cell_6t
Xbit_r104_c242 bl_242 br_242 wl_104 vdd gnd cell_6t
Xbit_r105_c242 bl_242 br_242 wl_105 vdd gnd cell_6t
Xbit_r106_c242 bl_242 br_242 wl_106 vdd gnd cell_6t
Xbit_r107_c242 bl_242 br_242 wl_107 vdd gnd cell_6t
Xbit_r108_c242 bl_242 br_242 wl_108 vdd gnd cell_6t
Xbit_r109_c242 bl_242 br_242 wl_109 vdd gnd cell_6t
Xbit_r110_c242 bl_242 br_242 wl_110 vdd gnd cell_6t
Xbit_r111_c242 bl_242 br_242 wl_111 vdd gnd cell_6t
Xbit_r112_c242 bl_242 br_242 wl_112 vdd gnd cell_6t
Xbit_r113_c242 bl_242 br_242 wl_113 vdd gnd cell_6t
Xbit_r114_c242 bl_242 br_242 wl_114 vdd gnd cell_6t
Xbit_r115_c242 bl_242 br_242 wl_115 vdd gnd cell_6t
Xbit_r116_c242 bl_242 br_242 wl_116 vdd gnd cell_6t
Xbit_r117_c242 bl_242 br_242 wl_117 vdd gnd cell_6t
Xbit_r118_c242 bl_242 br_242 wl_118 vdd gnd cell_6t
Xbit_r119_c242 bl_242 br_242 wl_119 vdd gnd cell_6t
Xbit_r120_c242 bl_242 br_242 wl_120 vdd gnd cell_6t
Xbit_r121_c242 bl_242 br_242 wl_121 vdd gnd cell_6t
Xbit_r122_c242 bl_242 br_242 wl_122 vdd gnd cell_6t
Xbit_r123_c242 bl_242 br_242 wl_123 vdd gnd cell_6t
Xbit_r124_c242 bl_242 br_242 wl_124 vdd gnd cell_6t
Xbit_r125_c242 bl_242 br_242 wl_125 vdd gnd cell_6t
Xbit_r126_c242 bl_242 br_242 wl_126 vdd gnd cell_6t
Xbit_r127_c242 bl_242 br_242 wl_127 vdd gnd cell_6t
Xbit_r128_c242 bl_242 br_242 wl_128 vdd gnd cell_6t
Xbit_r129_c242 bl_242 br_242 wl_129 vdd gnd cell_6t
Xbit_r130_c242 bl_242 br_242 wl_130 vdd gnd cell_6t
Xbit_r131_c242 bl_242 br_242 wl_131 vdd gnd cell_6t
Xbit_r132_c242 bl_242 br_242 wl_132 vdd gnd cell_6t
Xbit_r133_c242 bl_242 br_242 wl_133 vdd gnd cell_6t
Xbit_r134_c242 bl_242 br_242 wl_134 vdd gnd cell_6t
Xbit_r135_c242 bl_242 br_242 wl_135 vdd gnd cell_6t
Xbit_r136_c242 bl_242 br_242 wl_136 vdd gnd cell_6t
Xbit_r137_c242 bl_242 br_242 wl_137 vdd gnd cell_6t
Xbit_r138_c242 bl_242 br_242 wl_138 vdd gnd cell_6t
Xbit_r139_c242 bl_242 br_242 wl_139 vdd gnd cell_6t
Xbit_r140_c242 bl_242 br_242 wl_140 vdd gnd cell_6t
Xbit_r141_c242 bl_242 br_242 wl_141 vdd gnd cell_6t
Xbit_r142_c242 bl_242 br_242 wl_142 vdd gnd cell_6t
Xbit_r143_c242 bl_242 br_242 wl_143 vdd gnd cell_6t
Xbit_r144_c242 bl_242 br_242 wl_144 vdd gnd cell_6t
Xbit_r145_c242 bl_242 br_242 wl_145 vdd gnd cell_6t
Xbit_r146_c242 bl_242 br_242 wl_146 vdd gnd cell_6t
Xbit_r147_c242 bl_242 br_242 wl_147 vdd gnd cell_6t
Xbit_r148_c242 bl_242 br_242 wl_148 vdd gnd cell_6t
Xbit_r149_c242 bl_242 br_242 wl_149 vdd gnd cell_6t
Xbit_r150_c242 bl_242 br_242 wl_150 vdd gnd cell_6t
Xbit_r151_c242 bl_242 br_242 wl_151 vdd gnd cell_6t
Xbit_r152_c242 bl_242 br_242 wl_152 vdd gnd cell_6t
Xbit_r153_c242 bl_242 br_242 wl_153 vdd gnd cell_6t
Xbit_r154_c242 bl_242 br_242 wl_154 vdd gnd cell_6t
Xbit_r155_c242 bl_242 br_242 wl_155 vdd gnd cell_6t
Xbit_r156_c242 bl_242 br_242 wl_156 vdd gnd cell_6t
Xbit_r157_c242 bl_242 br_242 wl_157 vdd gnd cell_6t
Xbit_r158_c242 bl_242 br_242 wl_158 vdd gnd cell_6t
Xbit_r159_c242 bl_242 br_242 wl_159 vdd gnd cell_6t
Xbit_r160_c242 bl_242 br_242 wl_160 vdd gnd cell_6t
Xbit_r161_c242 bl_242 br_242 wl_161 vdd gnd cell_6t
Xbit_r162_c242 bl_242 br_242 wl_162 vdd gnd cell_6t
Xbit_r163_c242 bl_242 br_242 wl_163 vdd gnd cell_6t
Xbit_r164_c242 bl_242 br_242 wl_164 vdd gnd cell_6t
Xbit_r165_c242 bl_242 br_242 wl_165 vdd gnd cell_6t
Xbit_r166_c242 bl_242 br_242 wl_166 vdd gnd cell_6t
Xbit_r167_c242 bl_242 br_242 wl_167 vdd gnd cell_6t
Xbit_r168_c242 bl_242 br_242 wl_168 vdd gnd cell_6t
Xbit_r169_c242 bl_242 br_242 wl_169 vdd gnd cell_6t
Xbit_r170_c242 bl_242 br_242 wl_170 vdd gnd cell_6t
Xbit_r171_c242 bl_242 br_242 wl_171 vdd gnd cell_6t
Xbit_r172_c242 bl_242 br_242 wl_172 vdd gnd cell_6t
Xbit_r173_c242 bl_242 br_242 wl_173 vdd gnd cell_6t
Xbit_r174_c242 bl_242 br_242 wl_174 vdd gnd cell_6t
Xbit_r175_c242 bl_242 br_242 wl_175 vdd gnd cell_6t
Xbit_r176_c242 bl_242 br_242 wl_176 vdd gnd cell_6t
Xbit_r177_c242 bl_242 br_242 wl_177 vdd gnd cell_6t
Xbit_r178_c242 bl_242 br_242 wl_178 vdd gnd cell_6t
Xbit_r179_c242 bl_242 br_242 wl_179 vdd gnd cell_6t
Xbit_r180_c242 bl_242 br_242 wl_180 vdd gnd cell_6t
Xbit_r181_c242 bl_242 br_242 wl_181 vdd gnd cell_6t
Xbit_r182_c242 bl_242 br_242 wl_182 vdd gnd cell_6t
Xbit_r183_c242 bl_242 br_242 wl_183 vdd gnd cell_6t
Xbit_r184_c242 bl_242 br_242 wl_184 vdd gnd cell_6t
Xbit_r185_c242 bl_242 br_242 wl_185 vdd gnd cell_6t
Xbit_r186_c242 bl_242 br_242 wl_186 vdd gnd cell_6t
Xbit_r187_c242 bl_242 br_242 wl_187 vdd gnd cell_6t
Xbit_r188_c242 bl_242 br_242 wl_188 vdd gnd cell_6t
Xbit_r189_c242 bl_242 br_242 wl_189 vdd gnd cell_6t
Xbit_r190_c242 bl_242 br_242 wl_190 vdd gnd cell_6t
Xbit_r191_c242 bl_242 br_242 wl_191 vdd gnd cell_6t
Xbit_r192_c242 bl_242 br_242 wl_192 vdd gnd cell_6t
Xbit_r193_c242 bl_242 br_242 wl_193 vdd gnd cell_6t
Xbit_r194_c242 bl_242 br_242 wl_194 vdd gnd cell_6t
Xbit_r195_c242 bl_242 br_242 wl_195 vdd gnd cell_6t
Xbit_r196_c242 bl_242 br_242 wl_196 vdd gnd cell_6t
Xbit_r197_c242 bl_242 br_242 wl_197 vdd gnd cell_6t
Xbit_r198_c242 bl_242 br_242 wl_198 vdd gnd cell_6t
Xbit_r199_c242 bl_242 br_242 wl_199 vdd gnd cell_6t
Xbit_r200_c242 bl_242 br_242 wl_200 vdd gnd cell_6t
Xbit_r201_c242 bl_242 br_242 wl_201 vdd gnd cell_6t
Xbit_r202_c242 bl_242 br_242 wl_202 vdd gnd cell_6t
Xbit_r203_c242 bl_242 br_242 wl_203 vdd gnd cell_6t
Xbit_r204_c242 bl_242 br_242 wl_204 vdd gnd cell_6t
Xbit_r205_c242 bl_242 br_242 wl_205 vdd gnd cell_6t
Xbit_r206_c242 bl_242 br_242 wl_206 vdd gnd cell_6t
Xbit_r207_c242 bl_242 br_242 wl_207 vdd gnd cell_6t
Xbit_r208_c242 bl_242 br_242 wl_208 vdd gnd cell_6t
Xbit_r209_c242 bl_242 br_242 wl_209 vdd gnd cell_6t
Xbit_r210_c242 bl_242 br_242 wl_210 vdd gnd cell_6t
Xbit_r211_c242 bl_242 br_242 wl_211 vdd gnd cell_6t
Xbit_r212_c242 bl_242 br_242 wl_212 vdd gnd cell_6t
Xbit_r213_c242 bl_242 br_242 wl_213 vdd gnd cell_6t
Xbit_r214_c242 bl_242 br_242 wl_214 vdd gnd cell_6t
Xbit_r215_c242 bl_242 br_242 wl_215 vdd gnd cell_6t
Xbit_r216_c242 bl_242 br_242 wl_216 vdd gnd cell_6t
Xbit_r217_c242 bl_242 br_242 wl_217 vdd gnd cell_6t
Xbit_r218_c242 bl_242 br_242 wl_218 vdd gnd cell_6t
Xbit_r219_c242 bl_242 br_242 wl_219 vdd gnd cell_6t
Xbit_r220_c242 bl_242 br_242 wl_220 vdd gnd cell_6t
Xbit_r221_c242 bl_242 br_242 wl_221 vdd gnd cell_6t
Xbit_r222_c242 bl_242 br_242 wl_222 vdd gnd cell_6t
Xbit_r223_c242 bl_242 br_242 wl_223 vdd gnd cell_6t
Xbit_r224_c242 bl_242 br_242 wl_224 vdd gnd cell_6t
Xbit_r225_c242 bl_242 br_242 wl_225 vdd gnd cell_6t
Xbit_r226_c242 bl_242 br_242 wl_226 vdd gnd cell_6t
Xbit_r227_c242 bl_242 br_242 wl_227 vdd gnd cell_6t
Xbit_r228_c242 bl_242 br_242 wl_228 vdd gnd cell_6t
Xbit_r229_c242 bl_242 br_242 wl_229 vdd gnd cell_6t
Xbit_r230_c242 bl_242 br_242 wl_230 vdd gnd cell_6t
Xbit_r231_c242 bl_242 br_242 wl_231 vdd gnd cell_6t
Xbit_r232_c242 bl_242 br_242 wl_232 vdd gnd cell_6t
Xbit_r233_c242 bl_242 br_242 wl_233 vdd gnd cell_6t
Xbit_r234_c242 bl_242 br_242 wl_234 vdd gnd cell_6t
Xbit_r235_c242 bl_242 br_242 wl_235 vdd gnd cell_6t
Xbit_r236_c242 bl_242 br_242 wl_236 vdd gnd cell_6t
Xbit_r237_c242 bl_242 br_242 wl_237 vdd gnd cell_6t
Xbit_r238_c242 bl_242 br_242 wl_238 vdd gnd cell_6t
Xbit_r239_c242 bl_242 br_242 wl_239 vdd gnd cell_6t
Xbit_r240_c242 bl_242 br_242 wl_240 vdd gnd cell_6t
Xbit_r241_c242 bl_242 br_242 wl_241 vdd gnd cell_6t
Xbit_r242_c242 bl_242 br_242 wl_242 vdd gnd cell_6t
Xbit_r243_c242 bl_242 br_242 wl_243 vdd gnd cell_6t
Xbit_r244_c242 bl_242 br_242 wl_244 vdd gnd cell_6t
Xbit_r245_c242 bl_242 br_242 wl_245 vdd gnd cell_6t
Xbit_r246_c242 bl_242 br_242 wl_246 vdd gnd cell_6t
Xbit_r247_c242 bl_242 br_242 wl_247 vdd gnd cell_6t
Xbit_r248_c242 bl_242 br_242 wl_248 vdd gnd cell_6t
Xbit_r249_c242 bl_242 br_242 wl_249 vdd gnd cell_6t
Xbit_r250_c242 bl_242 br_242 wl_250 vdd gnd cell_6t
Xbit_r251_c242 bl_242 br_242 wl_251 vdd gnd cell_6t
Xbit_r252_c242 bl_242 br_242 wl_252 vdd gnd cell_6t
Xbit_r253_c242 bl_242 br_242 wl_253 vdd gnd cell_6t
Xbit_r254_c242 bl_242 br_242 wl_254 vdd gnd cell_6t
Xbit_r255_c242 bl_242 br_242 wl_255 vdd gnd cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd cell_6t
Xbit_r1_c243 bl_243 br_243 wl_1 vdd gnd cell_6t
Xbit_r2_c243 bl_243 br_243 wl_2 vdd gnd cell_6t
Xbit_r3_c243 bl_243 br_243 wl_3 vdd gnd cell_6t
Xbit_r4_c243 bl_243 br_243 wl_4 vdd gnd cell_6t
Xbit_r5_c243 bl_243 br_243 wl_5 vdd gnd cell_6t
Xbit_r6_c243 bl_243 br_243 wl_6 vdd gnd cell_6t
Xbit_r7_c243 bl_243 br_243 wl_7 vdd gnd cell_6t
Xbit_r8_c243 bl_243 br_243 wl_8 vdd gnd cell_6t
Xbit_r9_c243 bl_243 br_243 wl_9 vdd gnd cell_6t
Xbit_r10_c243 bl_243 br_243 wl_10 vdd gnd cell_6t
Xbit_r11_c243 bl_243 br_243 wl_11 vdd gnd cell_6t
Xbit_r12_c243 bl_243 br_243 wl_12 vdd gnd cell_6t
Xbit_r13_c243 bl_243 br_243 wl_13 vdd gnd cell_6t
Xbit_r14_c243 bl_243 br_243 wl_14 vdd gnd cell_6t
Xbit_r15_c243 bl_243 br_243 wl_15 vdd gnd cell_6t
Xbit_r16_c243 bl_243 br_243 wl_16 vdd gnd cell_6t
Xbit_r17_c243 bl_243 br_243 wl_17 vdd gnd cell_6t
Xbit_r18_c243 bl_243 br_243 wl_18 vdd gnd cell_6t
Xbit_r19_c243 bl_243 br_243 wl_19 vdd gnd cell_6t
Xbit_r20_c243 bl_243 br_243 wl_20 vdd gnd cell_6t
Xbit_r21_c243 bl_243 br_243 wl_21 vdd gnd cell_6t
Xbit_r22_c243 bl_243 br_243 wl_22 vdd gnd cell_6t
Xbit_r23_c243 bl_243 br_243 wl_23 vdd gnd cell_6t
Xbit_r24_c243 bl_243 br_243 wl_24 vdd gnd cell_6t
Xbit_r25_c243 bl_243 br_243 wl_25 vdd gnd cell_6t
Xbit_r26_c243 bl_243 br_243 wl_26 vdd gnd cell_6t
Xbit_r27_c243 bl_243 br_243 wl_27 vdd gnd cell_6t
Xbit_r28_c243 bl_243 br_243 wl_28 vdd gnd cell_6t
Xbit_r29_c243 bl_243 br_243 wl_29 vdd gnd cell_6t
Xbit_r30_c243 bl_243 br_243 wl_30 vdd gnd cell_6t
Xbit_r31_c243 bl_243 br_243 wl_31 vdd gnd cell_6t
Xbit_r32_c243 bl_243 br_243 wl_32 vdd gnd cell_6t
Xbit_r33_c243 bl_243 br_243 wl_33 vdd gnd cell_6t
Xbit_r34_c243 bl_243 br_243 wl_34 vdd gnd cell_6t
Xbit_r35_c243 bl_243 br_243 wl_35 vdd gnd cell_6t
Xbit_r36_c243 bl_243 br_243 wl_36 vdd gnd cell_6t
Xbit_r37_c243 bl_243 br_243 wl_37 vdd gnd cell_6t
Xbit_r38_c243 bl_243 br_243 wl_38 vdd gnd cell_6t
Xbit_r39_c243 bl_243 br_243 wl_39 vdd gnd cell_6t
Xbit_r40_c243 bl_243 br_243 wl_40 vdd gnd cell_6t
Xbit_r41_c243 bl_243 br_243 wl_41 vdd gnd cell_6t
Xbit_r42_c243 bl_243 br_243 wl_42 vdd gnd cell_6t
Xbit_r43_c243 bl_243 br_243 wl_43 vdd gnd cell_6t
Xbit_r44_c243 bl_243 br_243 wl_44 vdd gnd cell_6t
Xbit_r45_c243 bl_243 br_243 wl_45 vdd gnd cell_6t
Xbit_r46_c243 bl_243 br_243 wl_46 vdd gnd cell_6t
Xbit_r47_c243 bl_243 br_243 wl_47 vdd gnd cell_6t
Xbit_r48_c243 bl_243 br_243 wl_48 vdd gnd cell_6t
Xbit_r49_c243 bl_243 br_243 wl_49 vdd gnd cell_6t
Xbit_r50_c243 bl_243 br_243 wl_50 vdd gnd cell_6t
Xbit_r51_c243 bl_243 br_243 wl_51 vdd gnd cell_6t
Xbit_r52_c243 bl_243 br_243 wl_52 vdd gnd cell_6t
Xbit_r53_c243 bl_243 br_243 wl_53 vdd gnd cell_6t
Xbit_r54_c243 bl_243 br_243 wl_54 vdd gnd cell_6t
Xbit_r55_c243 bl_243 br_243 wl_55 vdd gnd cell_6t
Xbit_r56_c243 bl_243 br_243 wl_56 vdd gnd cell_6t
Xbit_r57_c243 bl_243 br_243 wl_57 vdd gnd cell_6t
Xbit_r58_c243 bl_243 br_243 wl_58 vdd gnd cell_6t
Xbit_r59_c243 bl_243 br_243 wl_59 vdd gnd cell_6t
Xbit_r60_c243 bl_243 br_243 wl_60 vdd gnd cell_6t
Xbit_r61_c243 bl_243 br_243 wl_61 vdd gnd cell_6t
Xbit_r62_c243 bl_243 br_243 wl_62 vdd gnd cell_6t
Xbit_r63_c243 bl_243 br_243 wl_63 vdd gnd cell_6t
Xbit_r64_c243 bl_243 br_243 wl_64 vdd gnd cell_6t
Xbit_r65_c243 bl_243 br_243 wl_65 vdd gnd cell_6t
Xbit_r66_c243 bl_243 br_243 wl_66 vdd gnd cell_6t
Xbit_r67_c243 bl_243 br_243 wl_67 vdd gnd cell_6t
Xbit_r68_c243 bl_243 br_243 wl_68 vdd gnd cell_6t
Xbit_r69_c243 bl_243 br_243 wl_69 vdd gnd cell_6t
Xbit_r70_c243 bl_243 br_243 wl_70 vdd gnd cell_6t
Xbit_r71_c243 bl_243 br_243 wl_71 vdd gnd cell_6t
Xbit_r72_c243 bl_243 br_243 wl_72 vdd gnd cell_6t
Xbit_r73_c243 bl_243 br_243 wl_73 vdd gnd cell_6t
Xbit_r74_c243 bl_243 br_243 wl_74 vdd gnd cell_6t
Xbit_r75_c243 bl_243 br_243 wl_75 vdd gnd cell_6t
Xbit_r76_c243 bl_243 br_243 wl_76 vdd gnd cell_6t
Xbit_r77_c243 bl_243 br_243 wl_77 vdd gnd cell_6t
Xbit_r78_c243 bl_243 br_243 wl_78 vdd gnd cell_6t
Xbit_r79_c243 bl_243 br_243 wl_79 vdd gnd cell_6t
Xbit_r80_c243 bl_243 br_243 wl_80 vdd gnd cell_6t
Xbit_r81_c243 bl_243 br_243 wl_81 vdd gnd cell_6t
Xbit_r82_c243 bl_243 br_243 wl_82 vdd gnd cell_6t
Xbit_r83_c243 bl_243 br_243 wl_83 vdd gnd cell_6t
Xbit_r84_c243 bl_243 br_243 wl_84 vdd gnd cell_6t
Xbit_r85_c243 bl_243 br_243 wl_85 vdd gnd cell_6t
Xbit_r86_c243 bl_243 br_243 wl_86 vdd gnd cell_6t
Xbit_r87_c243 bl_243 br_243 wl_87 vdd gnd cell_6t
Xbit_r88_c243 bl_243 br_243 wl_88 vdd gnd cell_6t
Xbit_r89_c243 bl_243 br_243 wl_89 vdd gnd cell_6t
Xbit_r90_c243 bl_243 br_243 wl_90 vdd gnd cell_6t
Xbit_r91_c243 bl_243 br_243 wl_91 vdd gnd cell_6t
Xbit_r92_c243 bl_243 br_243 wl_92 vdd gnd cell_6t
Xbit_r93_c243 bl_243 br_243 wl_93 vdd gnd cell_6t
Xbit_r94_c243 bl_243 br_243 wl_94 vdd gnd cell_6t
Xbit_r95_c243 bl_243 br_243 wl_95 vdd gnd cell_6t
Xbit_r96_c243 bl_243 br_243 wl_96 vdd gnd cell_6t
Xbit_r97_c243 bl_243 br_243 wl_97 vdd gnd cell_6t
Xbit_r98_c243 bl_243 br_243 wl_98 vdd gnd cell_6t
Xbit_r99_c243 bl_243 br_243 wl_99 vdd gnd cell_6t
Xbit_r100_c243 bl_243 br_243 wl_100 vdd gnd cell_6t
Xbit_r101_c243 bl_243 br_243 wl_101 vdd gnd cell_6t
Xbit_r102_c243 bl_243 br_243 wl_102 vdd gnd cell_6t
Xbit_r103_c243 bl_243 br_243 wl_103 vdd gnd cell_6t
Xbit_r104_c243 bl_243 br_243 wl_104 vdd gnd cell_6t
Xbit_r105_c243 bl_243 br_243 wl_105 vdd gnd cell_6t
Xbit_r106_c243 bl_243 br_243 wl_106 vdd gnd cell_6t
Xbit_r107_c243 bl_243 br_243 wl_107 vdd gnd cell_6t
Xbit_r108_c243 bl_243 br_243 wl_108 vdd gnd cell_6t
Xbit_r109_c243 bl_243 br_243 wl_109 vdd gnd cell_6t
Xbit_r110_c243 bl_243 br_243 wl_110 vdd gnd cell_6t
Xbit_r111_c243 bl_243 br_243 wl_111 vdd gnd cell_6t
Xbit_r112_c243 bl_243 br_243 wl_112 vdd gnd cell_6t
Xbit_r113_c243 bl_243 br_243 wl_113 vdd gnd cell_6t
Xbit_r114_c243 bl_243 br_243 wl_114 vdd gnd cell_6t
Xbit_r115_c243 bl_243 br_243 wl_115 vdd gnd cell_6t
Xbit_r116_c243 bl_243 br_243 wl_116 vdd gnd cell_6t
Xbit_r117_c243 bl_243 br_243 wl_117 vdd gnd cell_6t
Xbit_r118_c243 bl_243 br_243 wl_118 vdd gnd cell_6t
Xbit_r119_c243 bl_243 br_243 wl_119 vdd gnd cell_6t
Xbit_r120_c243 bl_243 br_243 wl_120 vdd gnd cell_6t
Xbit_r121_c243 bl_243 br_243 wl_121 vdd gnd cell_6t
Xbit_r122_c243 bl_243 br_243 wl_122 vdd gnd cell_6t
Xbit_r123_c243 bl_243 br_243 wl_123 vdd gnd cell_6t
Xbit_r124_c243 bl_243 br_243 wl_124 vdd gnd cell_6t
Xbit_r125_c243 bl_243 br_243 wl_125 vdd gnd cell_6t
Xbit_r126_c243 bl_243 br_243 wl_126 vdd gnd cell_6t
Xbit_r127_c243 bl_243 br_243 wl_127 vdd gnd cell_6t
Xbit_r128_c243 bl_243 br_243 wl_128 vdd gnd cell_6t
Xbit_r129_c243 bl_243 br_243 wl_129 vdd gnd cell_6t
Xbit_r130_c243 bl_243 br_243 wl_130 vdd gnd cell_6t
Xbit_r131_c243 bl_243 br_243 wl_131 vdd gnd cell_6t
Xbit_r132_c243 bl_243 br_243 wl_132 vdd gnd cell_6t
Xbit_r133_c243 bl_243 br_243 wl_133 vdd gnd cell_6t
Xbit_r134_c243 bl_243 br_243 wl_134 vdd gnd cell_6t
Xbit_r135_c243 bl_243 br_243 wl_135 vdd gnd cell_6t
Xbit_r136_c243 bl_243 br_243 wl_136 vdd gnd cell_6t
Xbit_r137_c243 bl_243 br_243 wl_137 vdd gnd cell_6t
Xbit_r138_c243 bl_243 br_243 wl_138 vdd gnd cell_6t
Xbit_r139_c243 bl_243 br_243 wl_139 vdd gnd cell_6t
Xbit_r140_c243 bl_243 br_243 wl_140 vdd gnd cell_6t
Xbit_r141_c243 bl_243 br_243 wl_141 vdd gnd cell_6t
Xbit_r142_c243 bl_243 br_243 wl_142 vdd gnd cell_6t
Xbit_r143_c243 bl_243 br_243 wl_143 vdd gnd cell_6t
Xbit_r144_c243 bl_243 br_243 wl_144 vdd gnd cell_6t
Xbit_r145_c243 bl_243 br_243 wl_145 vdd gnd cell_6t
Xbit_r146_c243 bl_243 br_243 wl_146 vdd gnd cell_6t
Xbit_r147_c243 bl_243 br_243 wl_147 vdd gnd cell_6t
Xbit_r148_c243 bl_243 br_243 wl_148 vdd gnd cell_6t
Xbit_r149_c243 bl_243 br_243 wl_149 vdd gnd cell_6t
Xbit_r150_c243 bl_243 br_243 wl_150 vdd gnd cell_6t
Xbit_r151_c243 bl_243 br_243 wl_151 vdd gnd cell_6t
Xbit_r152_c243 bl_243 br_243 wl_152 vdd gnd cell_6t
Xbit_r153_c243 bl_243 br_243 wl_153 vdd gnd cell_6t
Xbit_r154_c243 bl_243 br_243 wl_154 vdd gnd cell_6t
Xbit_r155_c243 bl_243 br_243 wl_155 vdd gnd cell_6t
Xbit_r156_c243 bl_243 br_243 wl_156 vdd gnd cell_6t
Xbit_r157_c243 bl_243 br_243 wl_157 vdd gnd cell_6t
Xbit_r158_c243 bl_243 br_243 wl_158 vdd gnd cell_6t
Xbit_r159_c243 bl_243 br_243 wl_159 vdd gnd cell_6t
Xbit_r160_c243 bl_243 br_243 wl_160 vdd gnd cell_6t
Xbit_r161_c243 bl_243 br_243 wl_161 vdd gnd cell_6t
Xbit_r162_c243 bl_243 br_243 wl_162 vdd gnd cell_6t
Xbit_r163_c243 bl_243 br_243 wl_163 vdd gnd cell_6t
Xbit_r164_c243 bl_243 br_243 wl_164 vdd gnd cell_6t
Xbit_r165_c243 bl_243 br_243 wl_165 vdd gnd cell_6t
Xbit_r166_c243 bl_243 br_243 wl_166 vdd gnd cell_6t
Xbit_r167_c243 bl_243 br_243 wl_167 vdd gnd cell_6t
Xbit_r168_c243 bl_243 br_243 wl_168 vdd gnd cell_6t
Xbit_r169_c243 bl_243 br_243 wl_169 vdd gnd cell_6t
Xbit_r170_c243 bl_243 br_243 wl_170 vdd gnd cell_6t
Xbit_r171_c243 bl_243 br_243 wl_171 vdd gnd cell_6t
Xbit_r172_c243 bl_243 br_243 wl_172 vdd gnd cell_6t
Xbit_r173_c243 bl_243 br_243 wl_173 vdd gnd cell_6t
Xbit_r174_c243 bl_243 br_243 wl_174 vdd gnd cell_6t
Xbit_r175_c243 bl_243 br_243 wl_175 vdd gnd cell_6t
Xbit_r176_c243 bl_243 br_243 wl_176 vdd gnd cell_6t
Xbit_r177_c243 bl_243 br_243 wl_177 vdd gnd cell_6t
Xbit_r178_c243 bl_243 br_243 wl_178 vdd gnd cell_6t
Xbit_r179_c243 bl_243 br_243 wl_179 vdd gnd cell_6t
Xbit_r180_c243 bl_243 br_243 wl_180 vdd gnd cell_6t
Xbit_r181_c243 bl_243 br_243 wl_181 vdd gnd cell_6t
Xbit_r182_c243 bl_243 br_243 wl_182 vdd gnd cell_6t
Xbit_r183_c243 bl_243 br_243 wl_183 vdd gnd cell_6t
Xbit_r184_c243 bl_243 br_243 wl_184 vdd gnd cell_6t
Xbit_r185_c243 bl_243 br_243 wl_185 vdd gnd cell_6t
Xbit_r186_c243 bl_243 br_243 wl_186 vdd gnd cell_6t
Xbit_r187_c243 bl_243 br_243 wl_187 vdd gnd cell_6t
Xbit_r188_c243 bl_243 br_243 wl_188 vdd gnd cell_6t
Xbit_r189_c243 bl_243 br_243 wl_189 vdd gnd cell_6t
Xbit_r190_c243 bl_243 br_243 wl_190 vdd gnd cell_6t
Xbit_r191_c243 bl_243 br_243 wl_191 vdd gnd cell_6t
Xbit_r192_c243 bl_243 br_243 wl_192 vdd gnd cell_6t
Xbit_r193_c243 bl_243 br_243 wl_193 vdd gnd cell_6t
Xbit_r194_c243 bl_243 br_243 wl_194 vdd gnd cell_6t
Xbit_r195_c243 bl_243 br_243 wl_195 vdd gnd cell_6t
Xbit_r196_c243 bl_243 br_243 wl_196 vdd gnd cell_6t
Xbit_r197_c243 bl_243 br_243 wl_197 vdd gnd cell_6t
Xbit_r198_c243 bl_243 br_243 wl_198 vdd gnd cell_6t
Xbit_r199_c243 bl_243 br_243 wl_199 vdd gnd cell_6t
Xbit_r200_c243 bl_243 br_243 wl_200 vdd gnd cell_6t
Xbit_r201_c243 bl_243 br_243 wl_201 vdd gnd cell_6t
Xbit_r202_c243 bl_243 br_243 wl_202 vdd gnd cell_6t
Xbit_r203_c243 bl_243 br_243 wl_203 vdd gnd cell_6t
Xbit_r204_c243 bl_243 br_243 wl_204 vdd gnd cell_6t
Xbit_r205_c243 bl_243 br_243 wl_205 vdd gnd cell_6t
Xbit_r206_c243 bl_243 br_243 wl_206 vdd gnd cell_6t
Xbit_r207_c243 bl_243 br_243 wl_207 vdd gnd cell_6t
Xbit_r208_c243 bl_243 br_243 wl_208 vdd gnd cell_6t
Xbit_r209_c243 bl_243 br_243 wl_209 vdd gnd cell_6t
Xbit_r210_c243 bl_243 br_243 wl_210 vdd gnd cell_6t
Xbit_r211_c243 bl_243 br_243 wl_211 vdd gnd cell_6t
Xbit_r212_c243 bl_243 br_243 wl_212 vdd gnd cell_6t
Xbit_r213_c243 bl_243 br_243 wl_213 vdd gnd cell_6t
Xbit_r214_c243 bl_243 br_243 wl_214 vdd gnd cell_6t
Xbit_r215_c243 bl_243 br_243 wl_215 vdd gnd cell_6t
Xbit_r216_c243 bl_243 br_243 wl_216 vdd gnd cell_6t
Xbit_r217_c243 bl_243 br_243 wl_217 vdd gnd cell_6t
Xbit_r218_c243 bl_243 br_243 wl_218 vdd gnd cell_6t
Xbit_r219_c243 bl_243 br_243 wl_219 vdd gnd cell_6t
Xbit_r220_c243 bl_243 br_243 wl_220 vdd gnd cell_6t
Xbit_r221_c243 bl_243 br_243 wl_221 vdd gnd cell_6t
Xbit_r222_c243 bl_243 br_243 wl_222 vdd gnd cell_6t
Xbit_r223_c243 bl_243 br_243 wl_223 vdd gnd cell_6t
Xbit_r224_c243 bl_243 br_243 wl_224 vdd gnd cell_6t
Xbit_r225_c243 bl_243 br_243 wl_225 vdd gnd cell_6t
Xbit_r226_c243 bl_243 br_243 wl_226 vdd gnd cell_6t
Xbit_r227_c243 bl_243 br_243 wl_227 vdd gnd cell_6t
Xbit_r228_c243 bl_243 br_243 wl_228 vdd gnd cell_6t
Xbit_r229_c243 bl_243 br_243 wl_229 vdd gnd cell_6t
Xbit_r230_c243 bl_243 br_243 wl_230 vdd gnd cell_6t
Xbit_r231_c243 bl_243 br_243 wl_231 vdd gnd cell_6t
Xbit_r232_c243 bl_243 br_243 wl_232 vdd gnd cell_6t
Xbit_r233_c243 bl_243 br_243 wl_233 vdd gnd cell_6t
Xbit_r234_c243 bl_243 br_243 wl_234 vdd gnd cell_6t
Xbit_r235_c243 bl_243 br_243 wl_235 vdd gnd cell_6t
Xbit_r236_c243 bl_243 br_243 wl_236 vdd gnd cell_6t
Xbit_r237_c243 bl_243 br_243 wl_237 vdd gnd cell_6t
Xbit_r238_c243 bl_243 br_243 wl_238 vdd gnd cell_6t
Xbit_r239_c243 bl_243 br_243 wl_239 vdd gnd cell_6t
Xbit_r240_c243 bl_243 br_243 wl_240 vdd gnd cell_6t
Xbit_r241_c243 bl_243 br_243 wl_241 vdd gnd cell_6t
Xbit_r242_c243 bl_243 br_243 wl_242 vdd gnd cell_6t
Xbit_r243_c243 bl_243 br_243 wl_243 vdd gnd cell_6t
Xbit_r244_c243 bl_243 br_243 wl_244 vdd gnd cell_6t
Xbit_r245_c243 bl_243 br_243 wl_245 vdd gnd cell_6t
Xbit_r246_c243 bl_243 br_243 wl_246 vdd gnd cell_6t
Xbit_r247_c243 bl_243 br_243 wl_247 vdd gnd cell_6t
Xbit_r248_c243 bl_243 br_243 wl_248 vdd gnd cell_6t
Xbit_r249_c243 bl_243 br_243 wl_249 vdd gnd cell_6t
Xbit_r250_c243 bl_243 br_243 wl_250 vdd gnd cell_6t
Xbit_r251_c243 bl_243 br_243 wl_251 vdd gnd cell_6t
Xbit_r252_c243 bl_243 br_243 wl_252 vdd gnd cell_6t
Xbit_r253_c243 bl_243 br_243 wl_253 vdd gnd cell_6t
Xbit_r254_c243 bl_243 br_243 wl_254 vdd gnd cell_6t
Xbit_r255_c243 bl_243 br_243 wl_255 vdd gnd cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd cell_6t
Xbit_r1_c244 bl_244 br_244 wl_1 vdd gnd cell_6t
Xbit_r2_c244 bl_244 br_244 wl_2 vdd gnd cell_6t
Xbit_r3_c244 bl_244 br_244 wl_3 vdd gnd cell_6t
Xbit_r4_c244 bl_244 br_244 wl_4 vdd gnd cell_6t
Xbit_r5_c244 bl_244 br_244 wl_5 vdd gnd cell_6t
Xbit_r6_c244 bl_244 br_244 wl_6 vdd gnd cell_6t
Xbit_r7_c244 bl_244 br_244 wl_7 vdd gnd cell_6t
Xbit_r8_c244 bl_244 br_244 wl_8 vdd gnd cell_6t
Xbit_r9_c244 bl_244 br_244 wl_9 vdd gnd cell_6t
Xbit_r10_c244 bl_244 br_244 wl_10 vdd gnd cell_6t
Xbit_r11_c244 bl_244 br_244 wl_11 vdd gnd cell_6t
Xbit_r12_c244 bl_244 br_244 wl_12 vdd gnd cell_6t
Xbit_r13_c244 bl_244 br_244 wl_13 vdd gnd cell_6t
Xbit_r14_c244 bl_244 br_244 wl_14 vdd gnd cell_6t
Xbit_r15_c244 bl_244 br_244 wl_15 vdd gnd cell_6t
Xbit_r16_c244 bl_244 br_244 wl_16 vdd gnd cell_6t
Xbit_r17_c244 bl_244 br_244 wl_17 vdd gnd cell_6t
Xbit_r18_c244 bl_244 br_244 wl_18 vdd gnd cell_6t
Xbit_r19_c244 bl_244 br_244 wl_19 vdd gnd cell_6t
Xbit_r20_c244 bl_244 br_244 wl_20 vdd gnd cell_6t
Xbit_r21_c244 bl_244 br_244 wl_21 vdd gnd cell_6t
Xbit_r22_c244 bl_244 br_244 wl_22 vdd gnd cell_6t
Xbit_r23_c244 bl_244 br_244 wl_23 vdd gnd cell_6t
Xbit_r24_c244 bl_244 br_244 wl_24 vdd gnd cell_6t
Xbit_r25_c244 bl_244 br_244 wl_25 vdd gnd cell_6t
Xbit_r26_c244 bl_244 br_244 wl_26 vdd gnd cell_6t
Xbit_r27_c244 bl_244 br_244 wl_27 vdd gnd cell_6t
Xbit_r28_c244 bl_244 br_244 wl_28 vdd gnd cell_6t
Xbit_r29_c244 bl_244 br_244 wl_29 vdd gnd cell_6t
Xbit_r30_c244 bl_244 br_244 wl_30 vdd gnd cell_6t
Xbit_r31_c244 bl_244 br_244 wl_31 vdd gnd cell_6t
Xbit_r32_c244 bl_244 br_244 wl_32 vdd gnd cell_6t
Xbit_r33_c244 bl_244 br_244 wl_33 vdd gnd cell_6t
Xbit_r34_c244 bl_244 br_244 wl_34 vdd gnd cell_6t
Xbit_r35_c244 bl_244 br_244 wl_35 vdd gnd cell_6t
Xbit_r36_c244 bl_244 br_244 wl_36 vdd gnd cell_6t
Xbit_r37_c244 bl_244 br_244 wl_37 vdd gnd cell_6t
Xbit_r38_c244 bl_244 br_244 wl_38 vdd gnd cell_6t
Xbit_r39_c244 bl_244 br_244 wl_39 vdd gnd cell_6t
Xbit_r40_c244 bl_244 br_244 wl_40 vdd gnd cell_6t
Xbit_r41_c244 bl_244 br_244 wl_41 vdd gnd cell_6t
Xbit_r42_c244 bl_244 br_244 wl_42 vdd gnd cell_6t
Xbit_r43_c244 bl_244 br_244 wl_43 vdd gnd cell_6t
Xbit_r44_c244 bl_244 br_244 wl_44 vdd gnd cell_6t
Xbit_r45_c244 bl_244 br_244 wl_45 vdd gnd cell_6t
Xbit_r46_c244 bl_244 br_244 wl_46 vdd gnd cell_6t
Xbit_r47_c244 bl_244 br_244 wl_47 vdd gnd cell_6t
Xbit_r48_c244 bl_244 br_244 wl_48 vdd gnd cell_6t
Xbit_r49_c244 bl_244 br_244 wl_49 vdd gnd cell_6t
Xbit_r50_c244 bl_244 br_244 wl_50 vdd gnd cell_6t
Xbit_r51_c244 bl_244 br_244 wl_51 vdd gnd cell_6t
Xbit_r52_c244 bl_244 br_244 wl_52 vdd gnd cell_6t
Xbit_r53_c244 bl_244 br_244 wl_53 vdd gnd cell_6t
Xbit_r54_c244 bl_244 br_244 wl_54 vdd gnd cell_6t
Xbit_r55_c244 bl_244 br_244 wl_55 vdd gnd cell_6t
Xbit_r56_c244 bl_244 br_244 wl_56 vdd gnd cell_6t
Xbit_r57_c244 bl_244 br_244 wl_57 vdd gnd cell_6t
Xbit_r58_c244 bl_244 br_244 wl_58 vdd gnd cell_6t
Xbit_r59_c244 bl_244 br_244 wl_59 vdd gnd cell_6t
Xbit_r60_c244 bl_244 br_244 wl_60 vdd gnd cell_6t
Xbit_r61_c244 bl_244 br_244 wl_61 vdd gnd cell_6t
Xbit_r62_c244 bl_244 br_244 wl_62 vdd gnd cell_6t
Xbit_r63_c244 bl_244 br_244 wl_63 vdd gnd cell_6t
Xbit_r64_c244 bl_244 br_244 wl_64 vdd gnd cell_6t
Xbit_r65_c244 bl_244 br_244 wl_65 vdd gnd cell_6t
Xbit_r66_c244 bl_244 br_244 wl_66 vdd gnd cell_6t
Xbit_r67_c244 bl_244 br_244 wl_67 vdd gnd cell_6t
Xbit_r68_c244 bl_244 br_244 wl_68 vdd gnd cell_6t
Xbit_r69_c244 bl_244 br_244 wl_69 vdd gnd cell_6t
Xbit_r70_c244 bl_244 br_244 wl_70 vdd gnd cell_6t
Xbit_r71_c244 bl_244 br_244 wl_71 vdd gnd cell_6t
Xbit_r72_c244 bl_244 br_244 wl_72 vdd gnd cell_6t
Xbit_r73_c244 bl_244 br_244 wl_73 vdd gnd cell_6t
Xbit_r74_c244 bl_244 br_244 wl_74 vdd gnd cell_6t
Xbit_r75_c244 bl_244 br_244 wl_75 vdd gnd cell_6t
Xbit_r76_c244 bl_244 br_244 wl_76 vdd gnd cell_6t
Xbit_r77_c244 bl_244 br_244 wl_77 vdd gnd cell_6t
Xbit_r78_c244 bl_244 br_244 wl_78 vdd gnd cell_6t
Xbit_r79_c244 bl_244 br_244 wl_79 vdd gnd cell_6t
Xbit_r80_c244 bl_244 br_244 wl_80 vdd gnd cell_6t
Xbit_r81_c244 bl_244 br_244 wl_81 vdd gnd cell_6t
Xbit_r82_c244 bl_244 br_244 wl_82 vdd gnd cell_6t
Xbit_r83_c244 bl_244 br_244 wl_83 vdd gnd cell_6t
Xbit_r84_c244 bl_244 br_244 wl_84 vdd gnd cell_6t
Xbit_r85_c244 bl_244 br_244 wl_85 vdd gnd cell_6t
Xbit_r86_c244 bl_244 br_244 wl_86 vdd gnd cell_6t
Xbit_r87_c244 bl_244 br_244 wl_87 vdd gnd cell_6t
Xbit_r88_c244 bl_244 br_244 wl_88 vdd gnd cell_6t
Xbit_r89_c244 bl_244 br_244 wl_89 vdd gnd cell_6t
Xbit_r90_c244 bl_244 br_244 wl_90 vdd gnd cell_6t
Xbit_r91_c244 bl_244 br_244 wl_91 vdd gnd cell_6t
Xbit_r92_c244 bl_244 br_244 wl_92 vdd gnd cell_6t
Xbit_r93_c244 bl_244 br_244 wl_93 vdd gnd cell_6t
Xbit_r94_c244 bl_244 br_244 wl_94 vdd gnd cell_6t
Xbit_r95_c244 bl_244 br_244 wl_95 vdd gnd cell_6t
Xbit_r96_c244 bl_244 br_244 wl_96 vdd gnd cell_6t
Xbit_r97_c244 bl_244 br_244 wl_97 vdd gnd cell_6t
Xbit_r98_c244 bl_244 br_244 wl_98 vdd gnd cell_6t
Xbit_r99_c244 bl_244 br_244 wl_99 vdd gnd cell_6t
Xbit_r100_c244 bl_244 br_244 wl_100 vdd gnd cell_6t
Xbit_r101_c244 bl_244 br_244 wl_101 vdd gnd cell_6t
Xbit_r102_c244 bl_244 br_244 wl_102 vdd gnd cell_6t
Xbit_r103_c244 bl_244 br_244 wl_103 vdd gnd cell_6t
Xbit_r104_c244 bl_244 br_244 wl_104 vdd gnd cell_6t
Xbit_r105_c244 bl_244 br_244 wl_105 vdd gnd cell_6t
Xbit_r106_c244 bl_244 br_244 wl_106 vdd gnd cell_6t
Xbit_r107_c244 bl_244 br_244 wl_107 vdd gnd cell_6t
Xbit_r108_c244 bl_244 br_244 wl_108 vdd gnd cell_6t
Xbit_r109_c244 bl_244 br_244 wl_109 vdd gnd cell_6t
Xbit_r110_c244 bl_244 br_244 wl_110 vdd gnd cell_6t
Xbit_r111_c244 bl_244 br_244 wl_111 vdd gnd cell_6t
Xbit_r112_c244 bl_244 br_244 wl_112 vdd gnd cell_6t
Xbit_r113_c244 bl_244 br_244 wl_113 vdd gnd cell_6t
Xbit_r114_c244 bl_244 br_244 wl_114 vdd gnd cell_6t
Xbit_r115_c244 bl_244 br_244 wl_115 vdd gnd cell_6t
Xbit_r116_c244 bl_244 br_244 wl_116 vdd gnd cell_6t
Xbit_r117_c244 bl_244 br_244 wl_117 vdd gnd cell_6t
Xbit_r118_c244 bl_244 br_244 wl_118 vdd gnd cell_6t
Xbit_r119_c244 bl_244 br_244 wl_119 vdd gnd cell_6t
Xbit_r120_c244 bl_244 br_244 wl_120 vdd gnd cell_6t
Xbit_r121_c244 bl_244 br_244 wl_121 vdd gnd cell_6t
Xbit_r122_c244 bl_244 br_244 wl_122 vdd gnd cell_6t
Xbit_r123_c244 bl_244 br_244 wl_123 vdd gnd cell_6t
Xbit_r124_c244 bl_244 br_244 wl_124 vdd gnd cell_6t
Xbit_r125_c244 bl_244 br_244 wl_125 vdd gnd cell_6t
Xbit_r126_c244 bl_244 br_244 wl_126 vdd gnd cell_6t
Xbit_r127_c244 bl_244 br_244 wl_127 vdd gnd cell_6t
Xbit_r128_c244 bl_244 br_244 wl_128 vdd gnd cell_6t
Xbit_r129_c244 bl_244 br_244 wl_129 vdd gnd cell_6t
Xbit_r130_c244 bl_244 br_244 wl_130 vdd gnd cell_6t
Xbit_r131_c244 bl_244 br_244 wl_131 vdd gnd cell_6t
Xbit_r132_c244 bl_244 br_244 wl_132 vdd gnd cell_6t
Xbit_r133_c244 bl_244 br_244 wl_133 vdd gnd cell_6t
Xbit_r134_c244 bl_244 br_244 wl_134 vdd gnd cell_6t
Xbit_r135_c244 bl_244 br_244 wl_135 vdd gnd cell_6t
Xbit_r136_c244 bl_244 br_244 wl_136 vdd gnd cell_6t
Xbit_r137_c244 bl_244 br_244 wl_137 vdd gnd cell_6t
Xbit_r138_c244 bl_244 br_244 wl_138 vdd gnd cell_6t
Xbit_r139_c244 bl_244 br_244 wl_139 vdd gnd cell_6t
Xbit_r140_c244 bl_244 br_244 wl_140 vdd gnd cell_6t
Xbit_r141_c244 bl_244 br_244 wl_141 vdd gnd cell_6t
Xbit_r142_c244 bl_244 br_244 wl_142 vdd gnd cell_6t
Xbit_r143_c244 bl_244 br_244 wl_143 vdd gnd cell_6t
Xbit_r144_c244 bl_244 br_244 wl_144 vdd gnd cell_6t
Xbit_r145_c244 bl_244 br_244 wl_145 vdd gnd cell_6t
Xbit_r146_c244 bl_244 br_244 wl_146 vdd gnd cell_6t
Xbit_r147_c244 bl_244 br_244 wl_147 vdd gnd cell_6t
Xbit_r148_c244 bl_244 br_244 wl_148 vdd gnd cell_6t
Xbit_r149_c244 bl_244 br_244 wl_149 vdd gnd cell_6t
Xbit_r150_c244 bl_244 br_244 wl_150 vdd gnd cell_6t
Xbit_r151_c244 bl_244 br_244 wl_151 vdd gnd cell_6t
Xbit_r152_c244 bl_244 br_244 wl_152 vdd gnd cell_6t
Xbit_r153_c244 bl_244 br_244 wl_153 vdd gnd cell_6t
Xbit_r154_c244 bl_244 br_244 wl_154 vdd gnd cell_6t
Xbit_r155_c244 bl_244 br_244 wl_155 vdd gnd cell_6t
Xbit_r156_c244 bl_244 br_244 wl_156 vdd gnd cell_6t
Xbit_r157_c244 bl_244 br_244 wl_157 vdd gnd cell_6t
Xbit_r158_c244 bl_244 br_244 wl_158 vdd gnd cell_6t
Xbit_r159_c244 bl_244 br_244 wl_159 vdd gnd cell_6t
Xbit_r160_c244 bl_244 br_244 wl_160 vdd gnd cell_6t
Xbit_r161_c244 bl_244 br_244 wl_161 vdd gnd cell_6t
Xbit_r162_c244 bl_244 br_244 wl_162 vdd gnd cell_6t
Xbit_r163_c244 bl_244 br_244 wl_163 vdd gnd cell_6t
Xbit_r164_c244 bl_244 br_244 wl_164 vdd gnd cell_6t
Xbit_r165_c244 bl_244 br_244 wl_165 vdd gnd cell_6t
Xbit_r166_c244 bl_244 br_244 wl_166 vdd gnd cell_6t
Xbit_r167_c244 bl_244 br_244 wl_167 vdd gnd cell_6t
Xbit_r168_c244 bl_244 br_244 wl_168 vdd gnd cell_6t
Xbit_r169_c244 bl_244 br_244 wl_169 vdd gnd cell_6t
Xbit_r170_c244 bl_244 br_244 wl_170 vdd gnd cell_6t
Xbit_r171_c244 bl_244 br_244 wl_171 vdd gnd cell_6t
Xbit_r172_c244 bl_244 br_244 wl_172 vdd gnd cell_6t
Xbit_r173_c244 bl_244 br_244 wl_173 vdd gnd cell_6t
Xbit_r174_c244 bl_244 br_244 wl_174 vdd gnd cell_6t
Xbit_r175_c244 bl_244 br_244 wl_175 vdd gnd cell_6t
Xbit_r176_c244 bl_244 br_244 wl_176 vdd gnd cell_6t
Xbit_r177_c244 bl_244 br_244 wl_177 vdd gnd cell_6t
Xbit_r178_c244 bl_244 br_244 wl_178 vdd gnd cell_6t
Xbit_r179_c244 bl_244 br_244 wl_179 vdd gnd cell_6t
Xbit_r180_c244 bl_244 br_244 wl_180 vdd gnd cell_6t
Xbit_r181_c244 bl_244 br_244 wl_181 vdd gnd cell_6t
Xbit_r182_c244 bl_244 br_244 wl_182 vdd gnd cell_6t
Xbit_r183_c244 bl_244 br_244 wl_183 vdd gnd cell_6t
Xbit_r184_c244 bl_244 br_244 wl_184 vdd gnd cell_6t
Xbit_r185_c244 bl_244 br_244 wl_185 vdd gnd cell_6t
Xbit_r186_c244 bl_244 br_244 wl_186 vdd gnd cell_6t
Xbit_r187_c244 bl_244 br_244 wl_187 vdd gnd cell_6t
Xbit_r188_c244 bl_244 br_244 wl_188 vdd gnd cell_6t
Xbit_r189_c244 bl_244 br_244 wl_189 vdd gnd cell_6t
Xbit_r190_c244 bl_244 br_244 wl_190 vdd gnd cell_6t
Xbit_r191_c244 bl_244 br_244 wl_191 vdd gnd cell_6t
Xbit_r192_c244 bl_244 br_244 wl_192 vdd gnd cell_6t
Xbit_r193_c244 bl_244 br_244 wl_193 vdd gnd cell_6t
Xbit_r194_c244 bl_244 br_244 wl_194 vdd gnd cell_6t
Xbit_r195_c244 bl_244 br_244 wl_195 vdd gnd cell_6t
Xbit_r196_c244 bl_244 br_244 wl_196 vdd gnd cell_6t
Xbit_r197_c244 bl_244 br_244 wl_197 vdd gnd cell_6t
Xbit_r198_c244 bl_244 br_244 wl_198 vdd gnd cell_6t
Xbit_r199_c244 bl_244 br_244 wl_199 vdd gnd cell_6t
Xbit_r200_c244 bl_244 br_244 wl_200 vdd gnd cell_6t
Xbit_r201_c244 bl_244 br_244 wl_201 vdd gnd cell_6t
Xbit_r202_c244 bl_244 br_244 wl_202 vdd gnd cell_6t
Xbit_r203_c244 bl_244 br_244 wl_203 vdd gnd cell_6t
Xbit_r204_c244 bl_244 br_244 wl_204 vdd gnd cell_6t
Xbit_r205_c244 bl_244 br_244 wl_205 vdd gnd cell_6t
Xbit_r206_c244 bl_244 br_244 wl_206 vdd gnd cell_6t
Xbit_r207_c244 bl_244 br_244 wl_207 vdd gnd cell_6t
Xbit_r208_c244 bl_244 br_244 wl_208 vdd gnd cell_6t
Xbit_r209_c244 bl_244 br_244 wl_209 vdd gnd cell_6t
Xbit_r210_c244 bl_244 br_244 wl_210 vdd gnd cell_6t
Xbit_r211_c244 bl_244 br_244 wl_211 vdd gnd cell_6t
Xbit_r212_c244 bl_244 br_244 wl_212 vdd gnd cell_6t
Xbit_r213_c244 bl_244 br_244 wl_213 vdd gnd cell_6t
Xbit_r214_c244 bl_244 br_244 wl_214 vdd gnd cell_6t
Xbit_r215_c244 bl_244 br_244 wl_215 vdd gnd cell_6t
Xbit_r216_c244 bl_244 br_244 wl_216 vdd gnd cell_6t
Xbit_r217_c244 bl_244 br_244 wl_217 vdd gnd cell_6t
Xbit_r218_c244 bl_244 br_244 wl_218 vdd gnd cell_6t
Xbit_r219_c244 bl_244 br_244 wl_219 vdd gnd cell_6t
Xbit_r220_c244 bl_244 br_244 wl_220 vdd gnd cell_6t
Xbit_r221_c244 bl_244 br_244 wl_221 vdd gnd cell_6t
Xbit_r222_c244 bl_244 br_244 wl_222 vdd gnd cell_6t
Xbit_r223_c244 bl_244 br_244 wl_223 vdd gnd cell_6t
Xbit_r224_c244 bl_244 br_244 wl_224 vdd gnd cell_6t
Xbit_r225_c244 bl_244 br_244 wl_225 vdd gnd cell_6t
Xbit_r226_c244 bl_244 br_244 wl_226 vdd gnd cell_6t
Xbit_r227_c244 bl_244 br_244 wl_227 vdd gnd cell_6t
Xbit_r228_c244 bl_244 br_244 wl_228 vdd gnd cell_6t
Xbit_r229_c244 bl_244 br_244 wl_229 vdd gnd cell_6t
Xbit_r230_c244 bl_244 br_244 wl_230 vdd gnd cell_6t
Xbit_r231_c244 bl_244 br_244 wl_231 vdd gnd cell_6t
Xbit_r232_c244 bl_244 br_244 wl_232 vdd gnd cell_6t
Xbit_r233_c244 bl_244 br_244 wl_233 vdd gnd cell_6t
Xbit_r234_c244 bl_244 br_244 wl_234 vdd gnd cell_6t
Xbit_r235_c244 bl_244 br_244 wl_235 vdd gnd cell_6t
Xbit_r236_c244 bl_244 br_244 wl_236 vdd gnd cell_6t
Xbit_r237_c244 bl_244 br_244 wl_237 vdd gnd cell_6t
Xbit_r238_c244 bl_244 br_244 wl_238 vdd gnd cell_6t
Xbit_r239_c244 bl_244 br_244 wl_239 vdd gnd cell_6t
Xbit_r240_c244 bl_244 br_244 wl_240 vdd gnd cell_6t
Xbit_r241_c244 bl_244 br_244 wl_241 vdd gnd cell_6t
Xbit_r242_c244 bl_244 br_244 wl_242 vdd gnd cell_6t
Xbit_r243_c244 bl_244 br_244 wl_243 vdd gnd cell_6t
Xbit_r244_c244 bl_244 br_244 wl_244 vdd gnd cell_6t
Xbit_r245_c244 bl_244 br_244 wl_245 vdd gnd cell_6t
Xbit_r246_c244 bl_244 br_244 wl_246 vdd gnd cell_6t
Xbit_r247_c244 bl_244 br_244 wl_247 vdd gnd cell_6t
Xbit_r248_c244 bl_244 br_244 wl_248 vdd gnd cell_6t
Xbit_r249_c244 bl_244 br_244 wl_249 vdd gnd cell_6t
Xbit_r250_c244 bl_244 br_244 wl_250 vdd gnd cell_6t
Xbit_r251_c244 bl_244 br_244 wl_251 vdd gnd cell_6t
Xbit_r252_c244 bl_244 br_244 wl_252 vdd gnd cell_6t
Xbit_r253_c244 bl_244 br_244 wl_253 vdd gnd cell_6t
Xbit_r254_c244 bl_244 br_244 wl_254 vdd gnd cell_6t
Xbit_r255_c244 bl_244 br_244 wl_255 vdd gnd cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd cell_6t
Xbit_r1_c245 bl_245 br_245 wl_1 vdd gnd cell_6t
Xbit_r2_c245 bl_245 br_245 wl_2 vdd gnd cell_6t
Xbit_r3_c245 bl_245 br_245 wl_3 vdd gnd cell_6t
Xbit_r4_c245 bl_245 br_245 wl_4 vdd gnd cell_6t
Xbit_r5_c245 bl_245 br_245 wl_5 vdd gnd cell_6t
Xbit_r6_c245 bl_245 br_245 wl_6 vdd gnd cell_6t
Xbit_r7_c245 bl_245 br_245 wl_7 vdd gnd cell_6t
Xbit_r8_c245 bl_245 br_245 wl_8 vdd gnd cell_6t
Xbit_r9_c245 bl_245 br_245 wl_9 vdd gnd cell_6t
Xbit_r10_c245 bl_245 br_245 wl_10 vdd gnd cell_6t
Xbit_r11_c245 bl_245 br_245 wl_11 vdd gnd cell_6t
Xbit_r12_c245 bl_245 br_245 wl_12 vdd gnd cell_6t
Xbit_r13_c245 bl_245 br_245 wl_13 vdd gnd cell_6t
Xbit_r14_c245 bl_245 br_245 wl_14 vdd gnd cell_6t
Xbit_r15_c245 bl_245 br_245 wl_15 vdd gnd cell_6t
Xbit_r16_c245 bl_245 br_245 wl_16 vdd gnd cell_6t
Xbit_r17_c245 bl_245 br_245 wl_17 vdd gnd cell_6t
Xbit_r18_c245 bl_245 br_245 wl_18 vdd gnd cell_6t
Xbit_r19_c245 bl_245 br_245 wl_19 vdd gnd cell_6t
Xbit_r20_c245 bl_245 br_245 wl_20 vdd gnd cell_6t
Xbit_r21_c245 bl_245 br_245 wl_21 vdd gnd cell_6t
Xbit_r22_c245 bl_245 br_245 wl_22 vdd gnd cell_6t
Xbit_r23_c245 bl_245 br_245 wl_23 vdd gnd cell_6t
Xbit_r24_c245 bl_245 br_245 wl_24 vdd gnd cell_6t
Xbit_r25_c245 bl_245 br_245 wl_25 vdd gnd cell_6t
Xbit_r26_c245 bl_245 br_245 wl_26 vdd gnd cell_6t
Xbit_r27_c245 bl_245 br_245 wl_27 vdd gnd cell_6t
Xbit_r28_c245 bl_245 br_245 wl_28 vdd gnd cell_6t
Xbit_r29_c245 bl_245 br_245 wl_29 vdd gnd cell_6t
Xbit_r30_c245 bl_245 br_245 wl_30 vdd gnd cell_6t
Xbit_r31_c245 bl_245 br_245 wl_31 vdd gnd cell_6t
Xbit_r32_c245 bl_245 br_245 wl_32 vdd gnd cell_6t
Xbit_r33_c245 bl_245 br_245 wl_33 vdd gnd cell_6t
Xbit_r34_c245 bl_245 br_245 wl_34 vdd gnd cell_6t
Xbit_r35_c245 bl_245 br_245 wl_35 vdd gnd cell_6t
Xbit_r36_c245 bl_245 br_245 wl_36 vdd gnd cell_6t
Xbit_r37_c245 bl_245 br_245 wl_37 vdd gnd cell_6t
Xbit_r38_c245 bl_245 br_245 wl_38 vdd gnd cell_6t
Xbit_r39_c245 bl_245 br_245 wl_39 vdd gnd cell_6t
Xbit_r40_c245 bl_245 br_245 wl_40 vdd gnd cell_6t
Xbit_r41_c245 bl_245 br_245 wl_41 vdd gnd cell_6t
Xbit_r42_c245 bl_245 br_245 wl_42 vdd gnd cell_6t
Xbit_r43_c245 bl_245 br_245 wl_43 vdd gnd cell_6t
Xbit_r44_c245 bl_245 br_245 wl_44 vdd gnd cell_6t
Xbit_r45_c245 bl_245 br_245 wl_45 vdd gnd cell_6t
Xbit_r46_c245 bl_245 br_245 wl_46 vdd gnd cell_6t
Xbit_r47_c245 bl_245 br_245 wl_47 vdd gnd cell_6t
Xbit_r48_c245 bl_245 br_245 wl_48 vdd gnd cell_6t
Xbit_r49_c245 bl_245 br_245 wl_49 vdd gnd cell_6t
Xbit_r50_c245 bl_245 br_245 wl_50 vdd gnd cell_6t
Xbit_r51_c245 bl_245 br_245 wl_51 vdd gnd cell_6t
Xbit_r52_c245 bl_245 br_245 wl_52 vdd gnd cell_6t
Xbit_r53_c245 bl_245 br_245 wl_53 vdd gnd cell_6t
Xbit_r54_c245 bl_245 br_245 wl_54 vdd gnd cell_6t
Xbit_r55_c245 bl_245 br_245 wl_55 vdd gnd cell_6t
Xbit_r56_c245 bl_245 br_245 wl_56 vdd gnd cell_6t
Xbit_r57_c245 bl_245 br_245 wl_57 vdd gnd cell_6t
Xbit_r58_c245 bl_245 br_245 wl_58 vdd gnd cell_6t
Xbit_r59_c245 bl_245 br_245 wl_59 vdd gnd cell_6t
Xbit_r60_c245 bl_245 br_245 wl_60 vdd gnd cell_6t
Xbit_r61_c245 bl_245 br_245 wl_61 vdd gnd cell_6t
Xbit_r62_c245 bl_245 br_245 wl_62 vdd gnd cell_6t
Xbit_r63_c245 bl_245 br_245 wl_63 vdd gnd cell_6t
Xbit_r64_c245 bl_245 br_245 wl_64 vdd gnd cell_6t
Xbit_r65_c245 bl_245 br_245 wl_65 vdd gnd cell_6t
Xbit_r66_c245 bl_245 br_245 wl_66 vdd gnd cell_6t
Xbit_r67_c245 bl_245 br_245 wl_67 vdd gnd cell_6t
Xbit_r68_c245 bl_245 br_245 wl_68 vdd gnd cell_6t
Xbit_r69_c245 bl_245 br_245 wl_69 vdd gnd cell_6t
Xbit_r70_c245 bl_245 br_245 wl_70 vdd gnd cell_6t
Xbit_r71_c245 bl_245 br_245 wl_71 vdd gnd cell_6t
Xbit_r72_c245 bl_245 br_245 wl_72 vdd gnd cell_6t
Xbit_r73_c245 bl_245 br_245 wl_73 vdd gnd cell_6t
Xbit_r74_c245 bl_245 br_245 wl_74 vdd gnd cell_6t
Xbit_r75_c245 bl_245 br_245 wl_75 vdd gnd cell_6t
Xbit_r76_c245 bl_245 br_245 wl_76 vdd gnd cell_6t
Xbit_r77_c245 bl_245 br_245 wl_77 vdd gnd cell_6t
Xbit_r78_c245 bl_245 br_245 wl_78 vdd gnd cell_6t
Xbit_r79_c245 bl_245 br_245 wl_79 vdd gnd cell_6t
Xbit_r80_c245 bl_245 br_245 wl_80 vdd gnd cell_6t
Xbit_r81_c245 bl_245 br_245 wl_81 vdd gnd cell_6t
Xbit_r82_c245 bl_245 br_245 wl_82 vdd gnd cell_6t
Xbit_r83_c245 bl_245 br_245 wl_83 vdd gnd cell_6t
Xbit_r84_c245 bl_245 br_245 wl_84 vdd gnd cell_6t
Xbit_r85_c245 bl_245 br_245 wl_85 vdd gnd cell_6t
Xbit_r86_c245 bl_245 br_245 wl_86 vdd gnd cell_6t
Xbit_r87_c245 bl_245 br_245 wl_87 vdd gnd cell_6t
Xbit_r88_c245 bl_245 br_245 wl_88 vdd gnd cell_6t
Xbit_r89_c245 bl_245 br_245 wl_89 vdd gnd cell_6t
Xbit_r90_c245 bl_245 br_245 wl_90 vdd gnd cell_6t
Xbit_r91_c245 bl_245 br_245 wl_91 vdd gnd cell_6t
Xbit_r92_c245 bl_245 br_245 wl_92 vdd gnd cell_6t
Xbit_r93_c245 bl_245 br_245 wl_93 vdd gnd cell_6t
Xbit_r94_c245 bl_245 br_245 wl_94 vdd gnd cell_6t
Xbit_r95_c245 bl_245 br_245 wl_95 vdd gnd cell_6t
Xbit_r96_c245 bl_245 br_245 wl_96 vdd gnd cell_6t
Xbit_r97_c245 bl_245 br_245 wl_97 vdd gnd cell_6t
Xbit_r98_c245 bl_245 br_245 wl_98 vdd gnd cell_6t
Xbit_r99_c245 bl_245 br_245 wl_99 vdd gnd cell_6t
Xbit_r100_c245 bl_245 br_245 wl_100 vdd gnd cell_6t
Xbit_r101_c245 bl_245 br_245 wl_101 vdd gnd cell_6t
Xbit_r102_c245 bl_245 br_245 wl_102 vdd gnd cell_6t
Xbit_r103_c245 bl_245 br_245 wl_103 vdd gnd cell_6t
Xbit_r104_c245 bl_245 br_245 wl_104 vdd gnd cell_6t
Xbit_r105_c245 bl_245 br_245 wl_105 vdd gnd cell_6t
Xbit_r106_c245 bl_245 br_245 wl_106 vdd gnd cell_6t
Xbit_r107_c245 bl_245 br_245 wl_107 vdd gnd cell_6t
Xbit_r108_c245 bl_245 br_245 wl_108 vdd gnd cell_6t
Xbit_r109_c245 bl_245 br_245 wl_109 vdd gnd cell_6t
Xbit_r110_c245 bl_245 br_245 wl_110 vdd gnd cell_6t
Xbit_r111_c245 bl_245 br_245 wl_111 vdd gnd cell_6t
Xbit_r112_c245 bl_245 br_245 wl_112 vdd gnd cell_6t
Xbit_r113_c245 bl_245 br_245 wl_113 vdd gnd cell_6t
Xbit_r114_c245 bl_245 br_245 wl_114 vdd gnd cell_6t
Xbit_r115_c245 bl_245 br_245 wl_115 vdd gnd cell_6t
Xbit_r116_c245 bl_245 br_245 wl_116 vdd gnd cell_6t
Xbit_r117_c245 bl_245 br_245 wl_117 vdd gnd cell_6t
Xbit_r118_c245 bl_245 br_245 wl_118 vdd gnd cell_6t
Xbit_r119_c245 bl_245 br_245 wl_119 vdd gnd cell_6t
Xbit_r120_c245 bl_245 br_245 wl_120 vdd gnd cell_6t
Xbit_r121_c245 bl_245 br_245 wl_121 vdd gnd cell_6t
Xbit_r122_c245 bl_245 br_245 wl_122 vdd gnd cell_6t
Xbit_r123_c245 bl_245 br_245 wl_123 vdd gnd cell_6t
Xbit_r124_c245 bl_245 br_245 wl_124 vdd gnd cell_6t
Xbit_r125_c245 bl_245 br_245 wl_125 vdd gnd cell_6t
Xbit_r126_c245 bl_245 br_245 wl_126 vdd gnd cell_6t
Xbit_r127_c245 bl_245 br_245 wl_127 vdd gnd cell_6t
Xbit_r128_c245 bl_245 br_245 wl_128 vdd gnd cell_6t
Xbit_r129_c245 bl_245 br_245 wl_129 vdd gnd cell_6t
Xbit_r130_c245 bl_245 br_245 wl_130 vdd gnd cell_6t
Xbit_r131_c245 bl_245 br_245 wl_131 vdd gnd cell_6t
Xbit_r132_c245 bl_245 br_245 wl_132 vdd gnd cell_6t
Xbit_r133_c245 bl_245 br_245 wl_133 vdd gnd cell_6t
Xbit_r134_c245 bl_245 br_245 wl_134 vdd gnd cell_6t
Xbit_r135_c245 bl_245 br_245 wl_135 vdd gnd cell_6t
Xbit_r136_c245 bl_245 br_245 wl_136 vdd gnd cell_6t
Xbit_r137_c245 bl_245 br_245 wl_137 vdd gnd cell_6t
Xbit_r138_c245 bl_245 br_245 wl_138 vdd gnd cell_6t
Xbit_r139_c245 bl_245 br_245 wl_139 vdd gnd cell_6t
Xbit_r140_c245 bl_245 br_245 wl_140 vdd gnd cell_6t
Xbit_r141_c245 bl_245 br_245 wl_141 vdd gnd cell_6t
Xbit_r142_c245 bl_245 br_245 wl_142 vdd gnd cell_6t
Xbit_r143_c245 bl_245 br_245 wl_143 vdd gnd cell_6t
Xbit_r144_c245 bl_245 br_245 wl_144 vdd gnd cell_6t
Xbit_r145_c245 bl_245 br_245 wl_145 vdd gnd cell_6t
Xbit_r146_c245 bl_245 br_245 wl_146 vdd gnd cell_6t
Xbit_r147_c245 bl_245 br_245 wl_147 vdd gnd cell_6t
Xbit_r148_c245 bl_245 br_245 wl_148 vdd gnd cell_6t
Xbit_r149_c245 bl_245 br_245 wl_149 vdd gnd cell_6t
Xbit_r150_c245 bl_245 br_245 wl_150 vdd gnd cell_6t
Xbit_r151_c245 bl_245 br_245 wl_151 vdd gnd cell_6t
Xbit_r152_c245 bl_245 br_245 wl_152 vdd gnd cell_6t
Xbit_r153_c245 bl_245 br_245 wl_153 vdd gnd cell_6t
Xbit_r154_c245 bl_245 br_245 wl_154 vdd gnd cell_6t
Xbit_r155_c245 bl_245 br_245 wl_155 vdd gnd cell_6t
Xbit_r156_c245 bl_245 br_245 wl_156 vdd gnd cell_6t
Xbit_r157_c245 bl_245 br_245 wl_157 vdd gnd cell_6t
Xbit_r158_c245 bl_245 br_245 wl_158 vdd gnd cell_6t
Xbit_r159_c245 bl_245 br_245 wl_159 vdd gnd cell_6t
Xbit_r160_c245 bl_245 br_245 wl_160 vdd gnd cell_6t
Xbit_r161_c245 bl_245 br_245 wl_161 vdd gnd cell_6t
Xbit_r162_c245 bl_245 br_245 wl_162 vdd gnd cell_6t
Xbit_r163_c245 bl_245 br_245 wl_163 vdd gnd cell_6t
Xbit_r164_c245 bl_245 br_245 wl_164 vdd gnd cell_6t
Xbit_r165_c245 bl_245 br_245 wl_165 vdd gnd cell_6t
Xbit_r166_c245 bl_245 br_245 wl_166 vdd gnd cell_6t
Xbit_r167_c245 bl_245 br_245 wl_167 vdd gnd cell_6t
Xbit_r168_c245 bl_245 br_245 wl_168 vdd gnd cell_6t
Xbit_r169_c245 bl_245 br_245 wl_169 vdd gnd cell_6t
Xbit_r170_c245 bl_245 br_245 wl_170 vdd gnd cell_6t
Xbit_r171_c245 bl_245 br_245 wl_171 vdd gnd cell_6t
Xbit_r172_c245 bl_245 br_245 wl_172 vdd gnd cell_6t
Xbit_r173_c245 bl_245 br_245 wl_173 vdd gnd cell_6t
Xbit_r174_c245 bl_245 br_245 wl_174 vdd gnd cell_6t
Xbit_r175_c245 bl_245 br_245 wl_175 vdd gnd cell_6t
Xbit_r176_c245 bl_245 br_245 wl_176 vdd gnd cell_6t
Xbit_r177_c245 bl_245 br_245 wl_177 vdd gnd cell_6t
Xbit_r178_c245 bl_245 br_245 wl_178 vdd gnd cell_6t
Xbit_r179_c245 bl_245 br_245 wl_179 vdd gnd cell_6t
Xbit_r180_c245 bl_245 br_245 wl_180 vdd gnd cell_6t
Xbit_r181_c245 bl_245 br_245 wl_181 vdd gnd cell_6t
Xbit_r182_c245 bl_245 br_245 wl_182 vdd gnd cell_6t
Xbit_r183_c245 bl_245 br_245 wl_183 vdd gnd cell_6t
Xbit_r184_c245 bl_245 br_245 wl_184 vdd gnd cell_6t
Xbit_r185_c245 bl_245 br_245 wl_185 vdd gnd cell_6t
Xbit_r186_c245 bl_245 br_245 wl_186 vdd gnd cell_6t
Xbit_r187_c245 bl_245 br_245 wl_187 vdd gnd cell_6t
Xbit_r188_c245 bl_245 br_245 wl_188 vdd gnd cell_6t
Xbit_r189_c245 bl_245 br_245 wl_189 vdd gnd cell_6t
Xbit_r190_c245 bl_245 br_245 wl_190 vdd gnd cell_6t
Xbit_r191_c245 bl_245 br_245 wl_191 vdd gnd cell_6t
Xbit_r192_c245 bl_245 br_245 wl_192 vdd gnd cell_6t
Xbit_r193_c245 bl_245 br_245 wl_193 vdd gnd cell_6t
Xbit_r194_c245 bl_245 br_245 wl_194 vdd gnd cell_6t
Xbit_r195_c245 bl_245 br_245 wl_195 vdd gnd cell_6t
Xbit_r196_c245 bl_245 br_245 wl_196 vdd gnd cell_6t
Xbit_r197_c245 bl_245 br_245 wl_197 vdd gnd cell_6t
Xbit_r198_c245 bl_245 br_245 wl_198 vdd gnd cell_6t
Xbit_r199_c245 bl_245 br_245 wl_199 vdd gnd cell_6t
Xbit_r200_c245 bl_245 br_245 wl_200 vdd gnd cell_6t
Xbit_r201_c245 bl_245 br_245 wl_201 vdd gnd cell_6t
Xbit_r202_c245 bl_245 br_245 wl_202 vdd gnd cell_6t
Xbit_r203_c245 bl_245 br_245 wl_203 vdd gnd cell_6t
Xbit_r204_c245 bl_245 br_245 wl_204 vdd gnd cell_6t
Xbit_r205_c245 bl_245 br_245 wl_205 vdd gnd cell_6t
Xbit_r206_c245 bl_245 br_245 wl_206 vdd gnd cell_6t
Xbit_r207_c245 bl_245 br_245 wl_207 vdd gnd cell_6t
Xbit_r208_c245 bl_245 br_245 wl_208 vdd gnd cell_6t
Xbit_r209_c245 bl_245 br_245 wl_209 vdd gnd cell_6t
Xbit_r210_c245 bl_245 br_245 wl_210 vdd gnd cell_6t
Xbit_r211_c245 bl_245 br_245 wl_211 vdd gnd cell_6t
Xbit_r212_c245 bl_245 br_245 wl_212 vdd gnd cell_6t
Xbit_r213_c245 bl_245 br_245 wl_213 vdd gnd cell_6t
Xbit_r214_c245 bl_245 br_245 wl_214 vdd gnd cell_6t
Xbit_r215_c245 bl_245 br_245 wl_215 vdd gnd cell_6t
Xbit_r216_c245 bl_245 br_245 wl_216 vdd gnd cell_6t
Xbit_r217_c245 bl_245 br_245 wl_217 vdd gnd cell_6t
Xbit_r218_c245 bl_245 br_245 wl_218 vdd gnd cell_6t
Xbit_r219_c245 bl_245 br_245 wl_219 vdd gnd cell_6t
Xbit_r220_c245 bl_245 br_245 wl_220 vdd gnd cell_6t
Xbit_r221_c245 bl_245 br_245 wl_221 vdd gnd cell_6t
Xbit_r222_c245 bl_245 br_245 wl_222 vdd gnd cell_6t
Xbit_r223_c245 bl_245 br_245 wl_223 vdd gnd cell_6t
Xbit_r224_c245 bl_245 br_245 wl_224 vdd gnd cell_6t
Xbit_r225_c245 bl_245 br_245 wl_225 vdd gnd cell_6t
Xbit_r226_c245 bl_245 br_245 wl_226 vdd gnd cell_6t
Xbit_r227_c245 bl_245 br_245 wl_227 vdd gnd cell_6t
Xbit_r228_c245 bl_245 br_245 wl_228 vdd gnd cell_6t
Xbit_r229_c245 bl_245 br_245 wl_229 vdd gnd cell_6t
Xbit_r230_c245 bl_245 br_245 wl_230 vdd gnd cell_6t
Xbit_r231_c245 bl_245 br_245 wl_231 vdd gnd cell_6t
Xbit_r232_c245 bl_245 br_245 wl_232 vdd gnd cell_6t
Xbit_r233_c245 bl_245 br_245 wl_233 vdd gnd cell_6t
Xbit_r234_c245 bl_245 br_245 wl_234 vdd gnd cell_6t
Xbit_r235_c245 bl_245 br_245 wl_235 vdd gnd cell_6t
Xbit_r236_c245 bl_245 br_245 wl_236 vdd gnd cell_6t
Xbit_r237_c245 bl_245 br_245 wl_237 vdd gnd cell_6t
Xbit_r238_c245 bl_245 br_245 wl_238 vdd gnd cell_6t
Xbit_r239_c245 bl_245 br_245 wl_239 vdd gnd cell_6t
Xbit_r240_c245 bl_245 br_245 wl_240 vdd gnd cell_6t
Xbit_r241_c245 bl_245 br_245 wl_241 vdd gnd cell_6t
Xbit_r242_c245 bl_245 br_245 wl_242 vdd gnd cell_6t
Xbit_r243_c245 bl_245 br_245 wl_243 vdd gnd cell_6t
Xbit_r244_c245 bl_245 br_245 wl_244 vdd gnd cell_6t
Xbit_r245_c245 bl_245 br_245 wl_245 vdd gnd cell_6t
Xbit_r246_c245 bl_245 br_245 wl_246 vdd gnd cell_6t
Xbit_r247_c245 bl_245 br_245 wl_247 vdd gnd cell_6t
Xbit_r248_c245 bl_245 br_245 wl_248 vdd gnd cell_6t
Xbit_r249_c245 bl_245 br_245 wl_249 vdd gnd cell_6t
Xbit_r250_c245 bl_245 br_245 wl_250 vdd gnd cell_6t
Xbit_r251_c245 bl_245 br_245 wl_251 vdd gnd cell_6t
Xbit_r252_c245 bl_245 br_245 wl_252 vdd gnd cell_6t
Xbit_r253_c245 bl_245 br_245 wl_253 vdd gnd cell_6t
Xbit_r254_c245 bl_245 br_245 wl_254 vdd gnd cell_6t
Xbit_r255_c245 bl_245 br_245 wl_255 vdd gnd cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd cell_6t
Xbit_r1_c246 bl_246 br_246 wl_1 vdd gnd cell_6t
Xbit_r2_c246 bl_246 br_246 wl_2 vdd gnd cell_6t
Xbit_r3_c246 bl_246 br_246 wl_3 vdd gnd cell_6t
Xbit_r4_c246 bl_246 br_246 wl_4 vdd gnd cell_6t
Xbit_r5_c246 bl_246 br_246 wl_5 vdd gnd cell_6t
Xbit_r6_c246 bl_246 br_246 wl_6 vdd gnd cell_6t
Xbit_r7_c246 bl_246 br_246 wl_7 vdd gnd cell_6t
Xbit_r8_c246 bl_246 br_246 wl_8 vdd gnd cell_6t
Xbit_r9_c246 bl_246 br_246 wl_9 vdd gnd cell_6t
Xbit_r10_c246 bl_246 br_246 wl_10 vdd gnd cell_6t
Xbit_r11_c246 bl_246 br_246 wl_11 vdd gnd cell_6t
Xbit_r12_c246 bl_246 br_246 wl_12 vdd gnd cell_6t
Xbit_r13_c246 bl_246 br_246 wl_13 vdd gnd cell_6t
Xbit_r14_c246 bl_246 br_246 wl_14 vdd gnd cell_6t
Xbit_r15_c246 bl_246 br_246 wl_15 vdd gnd cell_6t
Xbit_r16_c246 bl_246 br_246 wl_16 vdd gnd cell_6t
Xbit_r17_c246 bl_246 br_246 wl_17 vdd gnd cell_6t
Xbit_r18_c246 bl_246 br_246 wl_18 vdd gnd cell_6t
Xbit_r19_c246 bl_246 br_246 wl_19 vdd gnd cell_6t
Xbit_r20_c246 bl_246 br_246 wl_20 vdd gnd cell_6t
Xbit_r21_c246 bl_246 br_246 wl_21 vdd gnd cell_6t
Xbit_r22_c246 bl_246 br_246 wl_22 vdd gnd cell_6t
Xbit_r23_c246 bl_246 br_246 wl_23 vdd gnd cell_6t
Xbit_r24_c246 bl_246 br_246 wl_24 vdd gnd cell_6t
Xbit_r25_c246 bl_246 br_246 wl_25 vdd gnd cell_6t
Xbit_r26_c246 bl_246 br_246 wl_26 vdd gnd cell_6t
Xbit_r27_c246 bl_246 br_246 wl_27 vdd gnd cell_6t
Xbit_r28_c246 bl_246 br_246 wl_28 vdd gnd cell_6t
Xbit_r29_c246 bl_246 br_246 wl_29 vdd gnd cell_6t
Xbit_r30_c246 bl_246 br_246 wl_30 vdd gnd cell_6t
Xbit_r31_c246 bl_246 br_246 wl_31 vdd gnd cell_6t
Xbit_r32_c246 bl_246 br_246 wl_32 vdd gnd cell_6t
Xbit_r33_c246 bl_246 br_246 wl_33 vdd gnd cell_6t
Xbit_r34_c246 bl_246 br_246 wl_34 vdd gnd cell_6t
Xbit_r35_c246 bl_246 br_246 wl_35 vdd gnd cell_6t
Xbit_r36_c246 bl_246 br_246 wl_36 vdd gnd cell_6t
Xbit_r37_c246 bl_246 br_246 wl_37 vdd gnd cell_6t
Xbit_r38_c246 bl_246 br_246 wl_38 vdd gnd cell_6t
Xbit_r39_c246 bl_246 br_246 wl_39 vdd gnd cell_6t
Xbit_r40_c246 bl_246 br_246 wl_40 vdd gnd cell_6t
Xbit_r41_c246 bl_246 br_246 wl_41 vdd gnd cell_6t
Xbit_r42_c246 bl_246 br_246 wl_42 vdd gnd cell_6t
Xbit_r43_c246 bl_246 br_246 wl_43 vdd gnd cell_6t
Xbit_r44_c246 bl_246 br_246 wl_44 vdd gnd cell_6t
Xbit_r45_c246 bl_246 br_246 wl_45 vdd gnd cell_6t
Xbit_r46_c246 bl_246 br_246 wl_46 vdd gnd cell_6t
Xbit_r47_c246 bl_246 br_246 wl_47 vdd gnd cell_6t
Xbit_r48_c246 bl_246 br_246 wl_48 vdd gnd cell_6t
Xbit_r49_c246 bl_246 br_246 wl_49 vdd gnd cell_6t
Xbit_r50_c246 bl_246 br_246 wl_50 vdd gnd cell_6t
Xbit_r51_c246 bl_246 br_246 wl_51 vdd gnd cell_6t
Xbit_r52_c246 bl_246 br_246 wl_52 vdd gnd cell_6t
Xbit_r53_c246 bl_246 br_246 wl_53 vdd gnd cell_6t
Xbit_r54_c246 bl_246 br_246 wl_54 vdd gnd cell_6t
Xbit_r55_c246 bl_246 br_246 wl_55 vdd gnd cell_6t
Xbit_r56_c246 bl_246 br_246 wl_56 vdd gnd cell_6t
Xbit_r57_c246 bl_246 br_246 wl_57 vdd gnd cell_6t
Xbit_r58_c246 bl_246 br_246 wl_58 vdd gnd cell_6t
Xbit_r59_c246 bl_246 br_246 wl_59 vdd gnd cell_6t
Xbit_r60_c246 bl_246 br_246 wl_60 vdd gnd cell_6t
Xbit_r61_c246 bl_246 br_246 wl_61 vdd gnd cell_6t
Xbit_r62_c246 bl_246 br_246 wl_62 vdd gnd cell_6t
Xbit_r63_c246 bl_246 br_246 wl_63 vdd gnd cell_6t
Xbit_r64_c246 bl_246 br_246 wl_64 vdd gnd cell_6t
Xbit_r65_c246 bl_246 br_246 wl_65 vdd gnd cell_6t
Xbit_r66_c246 bl_246 br_246 wl_66 vdd gnd cell_6t
Xbit_r67_c246 bl_246 br_246 wl_67 vdd gnd cell_6t
Xbit_r68_c246 bl_246 br_246 wl_68 vdd gnd cell_6t
Xbit_r69_c246 bl_246 br_246 wl_69 vdd gnd cell_6t
Xbit_r70_c246 bl_246 br_246 wl_70 vdd gnd cell_6t
Xbit_r71_c246 bl_246 br_246 wl_71 vdd gnd cell_6t
Xbit_r72_c246 bl_246 br_246 wl_72 vdd gnd cell_6t
Xbit_r73_c246 bl_246 br_246 wl_73 vdd gnd cell_6t
Xbit_r74_c246 bl_246 br_246 wl_74 vdd gnd cell_6t
Xbit_r75_c246 bl_246 br_246 wl_75 vdd gnd cell_6t
Xbit_r76_c246 bl_246 br_246 wl_76 vdd gnd cell_6t
Xbit_r77_c246 bl_246 br_246 wl_77 vdd gnd cell_6t
Xbit_r78_c246 bl_246 br_246 wl_78 vdd gnd cell_6t
Xbit_r79_c246 bl_246 br_246 wl_79 vdd gnd cell_6t
Xbit_r80_c246 bl_246 br_246 wl_80 vdd gnd cell_6t
Xbit_r81_c246 bl_246 br_246 wl_81 vdd gnd cell_6t
Xbit_r82_c246 bl_246 br_246 wl_82 vdd gnd cell_6t
Xbit_r83_c246 bl_246 br_246 wl_83 vdd gnd cell_6t
Xbit_r84_c246 bl_246 br_246 wl_84 vdd gnd cell_6t
Xbit_r85_c246 bl_246 br_246 wl_85 vdd gnd cell_6t
Xbit_r86_c246 bl_246 br_246 wl_86 vdd gnd cell_6t
Xbit_r87_c246 bl_246 br_246 wl_87 vdd gnd cell_6t
Xbit_r88_c246 bl_246 br_246 wl_88 vdd gnd cell_6t
Xbit_r89_c246 bl_246 br_246 wl_89 vdd gnd cell_6t
Xbit_r90_c246 bl_246 br_246 wl_90 vdd gnd cell_6t
Xbit_r91_c246 bl_246 br_246 wl_91 vdd gnd cell_6t
Xbit_r92_c246 bl_246 br_246 wl_92 vdd gnd cell_6t
Xbit_r93_c246 bl_246 br_246 wl_93 vdd gnd cell_6t
Xbit_r94_c246 bl_246 br_246 wl_94 vdd gnd cell_6t
Xbit_r95_c246 bl_246 br_246 wl_95 vdd gnd cell_6t
Xbit_r96_c246 bl_246 br_246 wl_96 vdd gnd cell_6t
Xbit_r97_c246 bl_246 br_246 wl_97 vdd gnd cell_6t
Xbit_r98_c246 bl_246 br_246 wl_98 vdd gnd cell_6t
Xbit_r99_c246 bl_246 br_246 wl_99 vdd gnd cell_6t
Xbit_r100_c246 bl_246 br_246 wl_100 vdd gnd cell_6t
Xbit_r101_c246 bl_246 br_246 wl_101 vdd gnd cell_6t
Xbit_r102_c246 bl_246 br_246 wl_102 vdd gnd cell_6t
Xbit_r103_c246 bl_246 br_246 wl_103 vdd gnd cell_6t
Xbit_r104_c246 bl_246 br_246 wl_104 vdd gnd cell_6t
Xbit_r105_c246 bl_246 br_246 wl_105 vdd gnd cell_6t
Xbit_r106_c246 bl_246 br_246 wl_106 vdd gnd cell_6t
Xbit_r107_c246 bl_246 br_246 wl_107 vdd gnd cell_6t
Xbit_r108_c246 bl_246 br_246 wl_108 vdd gnd cell_6t
Xbit_r109_c246 bl_246 br_246 wl_109 vdd gnd cell_6t
Xbit_r110_c246 bl_246 br_246 wl_110 vdd gnd cell_6t
Xbit_r111_c246 bl_246 br_246 wl_111 vdd gnd cell_6t
Xbit_r112_c246 bl_246 br_246 wl_112 vdd gnd cell_6t
Xbit_r113_c246 bl_246 br_246 wl_113 vdd gnd cell_6t
Xbit_r114_c246 bl_246 br_246 wl_114 vdd gnd cell_6t
Xbit_r115_c246 bl_246 br_246 wl_115 vdd gnd cell_6t
Xbit_r116_c246 bl_246 br_246 wl_116 vdd gnd cell_6t
Xbit_r117_c246 bl_246 br_246 wl_117 vdd gnd cell_6t
Xbit_r118_c246 bl_246 br_246 wl_118 vdd gnd cell_6t
Xbit_r119_c246 bl_246 br_246 wl_119 vdd gnd cell_6t
Xbit_r120_c246 bl_246 br_246 wl_120 vdd gnd cell_6t
Xbit_r121_c246 bl_246 br_246 wl_121 vdd gnd cell_6t
Xbit_r122_c246 bl_246 br_246 wl_122 vdd gnd cell_6t
Xbit_r123_c246 bl_246 br_246 wl_123 vdd gnd cell_6t
Xbit_r124_c246 bl_246 br_246 wl_124 vdd gnd cell_6t
Xbit_r125_c246 bl_246 br_246 wl_125 vdd gnd cell_6t
Xbit_r126_c246 bl_246 br_246 wl_126 vdd gnd cell_6t
Xbit_r127_c246 bl_246 br_246 wl_127 vdd gnd cell_6t
Xbit_r128_c246 bl_246 br_246 wl_128 vdd gnd cell_6t
Xbit_r129_c246 bl_246 br_246 wl_129 vdd gnd cell_6t
Xbit_r130_c246 bl_246 br_246 wl_130 vdd gnd cell_6t
Xbit_r131_c246 bl_246 br_246 wl_131 vdd gnd cell_6t
Xbit_r132_c246 bl_246 br_246 wl_132 vdd gnd cell_6t
Xbit_r133_c246 bl_246 br_246 wl_133 vdd gnd cell_6t
Xbit_r134_c246 bl_246 br_246 wl_134 vdd gnd cell_6t
Xbit_r135_c246 bl_246 br_246 wl_135 vdd gnd cell_6t
Xbit_r136_c246 bl_246 br_246 wl_136 vdd gnd cell_6t
Xbit_r137_c246 bl_246 br_246 wl_137 vdd gnd cell_6t
Xbit_r138_c246 bl_246 br_246 wl_138 vdd gnd cell_6t
Xbit_r139_c246 bl_246 br_246 wl_139 vdd gnd cell_6t
Xbit_r140_c246 bl_246 br_246 wl_140 vdd gnd cell_6t
Xbit_r141_c246 bl_246 br_246 wl_141 vdd gnd cell_6t
Xbit_r142_c246 bl_246 br_246 wl_142 vdd gnd cell_6t
Xbit_r143_c246 bl_246 br_246 wl_143 vdd gnd cell_6t
Xbit_r144_c246 bl_246 br_246 wl_144 vdd gnd cell_6t
Xbit_r145_c246 bl_246 br_246 wl_145 vdd gnd cell_6t
Xbit_r146_c246 bl_246 br_246 wl_146 vdd gnd cell_6t
Xbit_r147_c246 bl_246 br_246 wl_147 vdd gnd cell_6t
Xbit_r148_c246 bl_246 br_246 wl_148 vdd gnd cell_6t
Xbit_r149_c246 bl_246 br_246 wl_149 vdd gnd cell_6t
Xbit_r150_c246 bl_246 br_246 wl_150 vdd gnd cell_6t
Xbit_r151_c246 bl_246 br_246 wl_151 vdd gnd cell_6t
Xbit_r152_c246 bl_246 br_246 wl_152 vdd gnd cell_6t
Xbit_r153_c246 bl_246 br_246 wl_153 vdd gnd cell_6t
Xbit_r154_c246 bl_246 br_246 wl_154 vdd gnd cell_6t
Xbit_r155_c246 bl_246 br_246 wl_155 vdd gnd cell_6t
Xbit_r156_c246 bl_246 br_246 wl_156 vdd gnd cell_6t
Xbit_r157_c246 bl_246 br_246 wl_157 vdd gnd cell_6t
Xbit_r158_c246 bl_246 br_246 wl_158 vdd gnd cell_6t
Xbit_r159_c246 bl_246 br_246 wl_159 vdd gnd cell_6t
Xbit_r160_c246 bl_246 br_246 wl_160 vdd gnd cell_6t
Xbit_r161_c246 bl_246 br_246 wl_161 vdd gnd cell_6t
Xbit_r162_c246 bl_246 br_246 wl_162 vdd gnd cell_6t
Xbit_r163_c246 bl_246 br_246 wl_163 vdd gnd cell_6t
Xbit_r164_c246 bl_246 br_246 wl_164 vdd gnd cell_6t
Xbit_r165_c246 bl_246 br_246 wl_165 vdd gnd cell_6t
Xbit_r166_c246 bl_246 br_246 wl_166 vdd gnd cell_6t
Xbit_r167_c246 bl_246 br_246 wl_167 vdd gnd cell_6t
Xbit_r168_c246 bl_246 br_246 wl_168 vdd gnd cell_6t
Xbit_r169_c246 bl_246 br_246 wl_169 vdd gnd cell_6t
Xbit_r170_c246 bl_246 br_246 wl_170 vdd gnd cell_6t
Xbit_r171_c246 bl_246 br_246 wl_171 vdd gnd cell_6t
Xbit_r172_c246 bl_246 br_246 wl_172 vdd gnd cell_6t
Xbit_r173_c246 bl_246 br_246 wl_173 vdd gnd cell_6t
Xbit_r174_c246 bl_246 br_246 wl_174 vdd gnd cell_6t
Xbit_r175_c246 bl_246 br_246 wl_175 vdd gnd cell_6t
Xbit_r176_c246 bl_246 br_246 wl_176 vdd gnd cell_6t
Xbit_r177_c246 bl_246 br_246 wl_177 vdd gnd cell_6t
Xbit_r178_c246 bl_246 br_246 wl_178 vdd gnd cell_6t
Xbit_r179_c246 bl_246 br_246 wl_179 vdd gnd cell_6t
Xbit_r180_c246 bl_246 br_246 wl_180 vdd gnd cell_6t
Xbit_r181_c246 bl_246 br_246 wl_181 vdd gnd cell_6t
Xbit_r182_c246 bl_246 br_246 wl_182 vdd gnd cell_6t
Xbit_r183_c246 bl_246 br_246 wl_183 vdd gnd cell_6t
Xbit_r184_c246 bl_246 br_246 wl_184 vdd gnd cell_6t
Xbit_r185_c246 bl_246 br_246 wl_185 vdd gnd cell_6t
Xbit_r186_c246 bl_246 br_246 wl_186 vdd gnd cell_6t
Xbit_r187_c246 bl_246 br_246 wl_187 vdd gnd cell_6t
Xbit_r188_c246 bl_246 br_246 wl_188 vdd gnd cell_6t
Xbit_r189_c246 bl_246 br_246 wl_189 vdd gnd cell_6t
Xbit_r190_c246 bl_246 br_246 wl_190 vdd gnd cell_6t
Xbit_r191_c246 bl_246 br_246 wl_191 vdd gnd cell_6t
Xbit_r192_c246 bl_246 br_246 wl_192 vdd gnd cell_6t
Xbit_r193_c246 bl_246 br_246 wl_193 vdd gnd cell_6t
Xbit_r194_c246 bl_246 br_246 wl_194 vdd gnd cell_6t
Xbit_r195_c246 bl_246 br_246 wl_195 vdd gnd cell_6t
Xbit_r196_c246 bl_246 br_246 wl_196 vdd gnd cell_6t
Xbit_r197_c246 bl_246 br_246 wl_197 vdd gnd cell_6t
Xbit_r198_c246 bl_246 br_246 wl_198 vdd gnd cell_6t
Xbit_r199_c246 bl_246 br_246 wl_199 vdd gnd cell_6t
Xbit_r200_c246 bl_246 br_246 wl_200 vdd gnd cell_6t
Xbit_r201_c246 bl_246 br_246 wl_201 vdd gnd cell_6t
Xbit_r202_c246 bl_246 br_246 wl_202 vdd gnd cell_6t
Xbit_r203_c246 bl_246 br_246 wl_203 vdd gnd cell_6t
Xbit_r204_c246 bl_246 br_246 wl_204 vdd gnd cell_6t
Xbit_r205_c246 bl_246 br_246 wl_205 vdd gnd cell_6t
Xbit_r206_c246 bl_246 br_246 wl_206 vdd gnd cell_6t
Xbit_r207_c246 bl_246 br_246 wl_207 vdd gnd cell_6t
Xbit_r208_c246 bl_246 br_246 wl_208 vdd gnd cell_6t
Xbit_r209_c246 bl_246 br_246 wl_209 vdd gnd cell_6t
Xbit_r210_c246 bl_246 br_246 wl_210 vdd gnd cell_6t
Xbit_r211_c246 bl_246 br_246 wl_211 vdd gnd cell_6t
Xbit_r212_c246 bl_246 br_246 wl_212 vdd gnd cell_6t
Xbit_r213_c246 bl_246 br_246 wl_213 vdd gnd cell_6t
Xbit_r214_c246 bl_246 br_246 wl_214 vdd gnd cell_6t
Xbit_r215_c246 bl_246 br_246 wl_215 vdd gnd cell_6t
Xbit_r216_c246 bl_246 br_246 wl_216 vdd gnd cell_6t
Xbit_r217_c246 bl_246 br_246 wl_217 vdd gnd cell_6t
Xbit_r218_c246 bl_246 br_246 wl_218 vdd gnd cell_6t
Xbit_r219_c246 bl_246 br_246 wl_219 vdd gnd cell_6t
Xbit_r220_c246 bl_246 br_246 wl_220 vdd gnd cell_6t
Xbit_r221_c246 bl_246 br_246 wl_221 vdd gnd cell_6t
Xbit_r222_c246 bl_246 br_246 wl_222 vdd gnd cell_6t
Xbit_r223_c246 bl_246 br_246 wl_223 vdd gnd cell_6t
Xbit_r224_c246 bl_246 br_246 wl_224 vdd gnd cell_6t
Xbit_r225_c246 bl_246 br_246 wl_225 vdd gnd cell_6t
Xbit_r226_c246 bl_246 br_246 wl_226 vdd gnd cell_6t
Xbit_r227_c246 bl_246 br_246 wl_227 vdd gnd cell_6t
Xbit_r228_c246 bl_246 br_246 wl_228 vdd gnd cell_6t
Xbit_r229_c246 bl_246 br_246 wl_229 vdd gnd cell_6t
Xbit_r230_c246 bl_246 br_246 wl_230 vdd gnd cell_6t
Xbit_r231_c246 bl_246 br_246 wl_231 vdd gnd cell_6t
Xbit_r232_c246 bl_246 br_246 wl_232 vdd gnd cell_6t
Xbit_r233_c246 bl_246 br_246 wl_233 vdd gnd cell_6t
Xbit_r234_c246 bl_246 br_246 wl_234 vdd gnd cell_6t
Xbit_r235_c246 bl_246 br_246 wl_235 vdd gnd cell_6t
Xbit_r236_c246 bl_246 br_246 wl_236 vdd gnd cell_6t
Xbit_r237_c246 bl_246 br_246 wl_237 vdd gnd cell_6t
Xbit_r238_c246 bl_246 br_246 wl_238 vdd gnd cell_6t
Xbit_r239_c246 bl_246 br_246 wl_239 vdd gnd cell_6t
Xbit_r240_c246 bl_246 br_246 wl_240 vdd gnd cell_6t
Xbit_r241_c246 bl_246 br_246 wl_241 vdd gnd cell_6t
Xbit_r242_c246 bl_246 br_246 wl_242 vdd gnd cell_6t
Xbit_r243_c246 bl_246 br_246 wl_243 vdd gnd cell_6t
Xbit_r244_c246 bl_246 br_246 wl_244 vdd gnd cell_6t
Xbit_r245_c246 bl_246 br_246 wl_245 vdd gnd cell_6t
Xbit_r246_c246 bl_246 br_246 wl_246 vdd gnd cell_6t
Xbit_r247_c246 bl_246 br_246 wl_247 vdd gnd cell_6t
Xbit_r248_c246 bl_246 br_246 wl_248 vdd gnd cell_6t
Xbit_r249_c246 bl_246 br_246 wl_249 vdd gnd cell_6t
Xbit_r250_c246 bl_246 br_246 wl_250 vdd gnd cell_6t
Xbit_r251_c246 bl_246 br_246 wl_251 vdd gnd cell_6t
Xbit_r252_c246 bl_246 br_246 wl_252 vdd gnd cell_6t
Xbit_r253_c246 bl_246 br_246 wl_253 vdd gnd cell_6t
Xbit_r254_c246 bl_246 br_246 wl_254 vdd gnd cell_6t
Xbit_r255_c246 bl_246 br_246 wl_255 vdd gnd cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd cell_6t
Xbit_r1_c247 bl_247 br_247 wl_1 vdd gnd cell_6t
Xbit_r2_c247 bl_247 br_247 wl_2 vdd gnd cell_6t
Xbit_r3_c247 bl_247 br_247 wl_3 vdd gnd cell_6t
Xbit_r4_c247 bl_247 br_247 wl_4 vdd gnd cell_6t
Xbit_r5_c247 bl_247 br_247 wl_5 vdd gnd cell_6t
Xbit_r6_c247 bl_247 br_247 wl_6 vdd gnd cell_6t
Xbit_r7_c247 bl_247 br_247 wl_7 vdd gnd cell_6t
Xbit_r8_c247 bl_247 br_247 wl_8 vdd gnd cell_6t
Xbit_r9_c247 bl_247 br_247 wl_9 vdd gnd cell_6t
Xbit_r10_c247 bl_247 br_247 wl_10 vdd gnd cell_6t
Xbit_r11_c247 bl_247 br_247 wl_11 vdd gnd cell_6t
Xbit_r12_c247 bl_247 br_247 wl_12 vdd gnd cell_6t
Xbit_r13_c247 bl_247 br_247 wl_13 vdd gnd cell_6t
Xbit_r14_c247 bl_247 br_247 wl_14 vdd gnd cell_6t
Xbit_r15_c247 bl_247 br_247 wl_15 vdd gnd cell_6t
Xbit_r16_c247 bl_247 br_247 wl_16 vdd gnd cell_6t
Xbit_r17_c247 bl_247 br_247 wl_17 vdd gnd cell_6t
Xbit_r18_c247 bl_247 br_247 wl_18 vdd gnd cell_6t
Xbit_r19_c247 bl_247 br_247 wl_19 vdd gnd cell_6t
Xbit_r20_c247 bl_247 br_247 wl_20 vdd gnd cell_6t
Xbit_r21_c247 bl_247 br_247 wl_21 vdd gnd cell_6t
Xbit_r22_c247 bl_247 br_247 wl_22 vdd gnd cell_6t
Xbit_r23_c247 bl_247 br_247 wl_23 vdd gnd cell_6t
Xbit_r24_c247 bl_247 br_247 wl_24 vdd gnd cell_6t
Xbit_r25_c247 bl_247 br_247 wl_25 vdd gnd cell_6t
Xbit_r26_c247 bl_247 br_247 wl_26 vdd gnd cell_6t
Xbit_r27_c247 bl_247 br_247 wl_27 vdd gnd cell_6t
Xbit_r28_c247 bl_247 br_247 wl_28 vdd gnd cell_6t
Xbit_r29_c247 bl_247 br_247 wl_29 vdd gnd cell_6t
Xbit_r30_c247 bl_247 br_247 wl_30 vdd gnd cell_6t
Xbit_r31_c247 bl_247 br_247 wl_31 vdd gnd cell_6t
Xbit_r32_c247 bl_247 br_247 wl_32 vdd gnd cell_6t
Xbit_r33_c247 bl_247 br_247 wl_33 vdd gnd cell_6t
Xbit_r34_c247 bl_247 br_247 wl_34 vdd gnd cell_6t
Xbit_r35_c247 bl_247 br_247 wl_35 vdd gnd cell_6t
Xbit_r36_c247 bl_247 br_247 wl_36 vdd gnd cell_6t
Xbit_r37_c247 bl_247 br_247 wl_37 vdd gnd cell_6t
Xbit_r38_c247 bl_247 br_247 wl_38 vdd gnd cell_6t
Xbit_r39_c247 bl_247 br_247 wl_39 vdd gnd cell_6t
Xbit_r40_c247 bl_247 br_247 wl_40 vdd gnd cell_6t
Xbit_r41_c247 bl_247 br_247 wl_41 vdd gnd cell_6t
Xbit_r42_c247 bl_247 br_247 wl_42 vdd gnd cell_6t
Xbit_r43_c247 bl_247 br_247 wl_43 vdd gnd cell_6t
Xbit_r44_c247 bl_247 br_247 wl_44 vdd gnd cell_6t
Xbit_r45_c247 bl_247 br_247 wl_45 vdd gnd cell_6t
Xbit_r46_c247 bl_247 br_247 wl_46 vdd gnd cell_6t
Xbit_r47_c247 bl_247 br_247 wl_47 vdd gnd cell_6t
Xbit_r48_c247 bl_247 br_247 wl_48 vdd gnd cell_6t
Xbit_r49_c247 bl_247 br_247 wl_49 vdd gnd cell_6t
Xbit_r50_c247 bl_247 br_247 wl_50 vdd gnd cell_6t
Xbit_r51_c247 bl_247 br_247 wl_51 vdd gnd cell_6t
Xbit_r52_c247 bl_247 br_247 wl_52 vdd gnd cell_6t
Xbit_r53_c247 bl_247 br_247 wl_53 vdd gnd cell_6t
Xbit_r54_c247 bl_247 br_247 wl_54 vdd gnd cell_6t
Xbit_r55_c247 bl_247 br_247 wl_55 vdd gnd cell_6t
Xbit_r56_c247 bl_247 br_247 wl_56 vdd gnd cell_6t
Xbit_r57_c247 bl_247 br_247 wl_57 vdd gnd cell_6t
Xbit_r58_c247 bl_247 br_247 wl_58 vdd gnd cell_6t
Xbit_r59_c247 bl_247 br_247 wl_59 vdd gnd cell_6t
Xbit_r60_c247 bl_247 br_247 wl_60 vdd gnd cell_6t
Xbit_r61_c247 bl_247 br_247 wl_61 vdd gnd cell_6t
Xbit_r62_c247 bl_247 br_247 wl_62 vdd gnd cell_6t
Xbit_r63_c247 bl_247 br_247 wl_63 vdd gnd cell_6t
Xbit_r64_c247 bl_247 br_247 wl_64 vdd gnd cell_6t
Xbit_r65_c247 bl_247 br_247 wl_65 vdd gnd cell_6t
Xbit_r66_c247 bl_247 br_247 wl_66 vdd gnd cell_6t
Xbit_r67_c247 bl_247 br_247 wl_67 vdd gnd cell_6t
Xbit_r68_c247 bl_247 br_247 wl_68 vdd gnd cell_6t
Xbit_r69_c247 bl_247 br_247 wl_69 vdd gnd cell_6t
Xbit_r70_c247 bl_247 br_247 wl_70 vdd gnd cell_6t
Xbit_r71_c247 bl_247 br_247 wl_71 vdd gnd cell_6t
Xbit_r72_c247 bl_247 br_247 wl_72 vdd gnd cell_6t
Xbit_r73_c247 bl_247 br_247 wl_73 vdd gnd cell_6t
Xbit_r74_c247 bl_247 br_247 wl_74 vdd gnd cell_6t
Xbit_r75_c247 bl_247 br_247 wl_75 vdd gnd cell_6t
Xbit_r76_c247 bl_247 br_247 wl_76 vdd gnd cell_6t
Xbit_r77_c247 bl_247 br_247 wl_77 vdd gnd cell_6t
Xbit_r78_c247 bl_247 br_247 wl_78 vdd gnd cell_6t
Xbit_r79_c247 bl_247 br_247 wl_79 vdd gnd cell_6t
Xbit_r80_c247 bl_247 br_247 wl_80 vdd gnd cell_6t
Xbit_r81_c247 bl_247 br_247 wl_81 vdd gnd cell_6t
Xbit_r82_c247 bl_247 br_247 wl_82 vdd gnd cell_6t
Xbit_r83_c247 bl_247 br_247 wl_83 vdd gnd cell_6t
Xbit_r84_c247 bl_247 br_247 wl_84 vdd gnd cell_6t
Xbit_r85_c247 bl_247 br_247 wl_85 vdd gnd cell_6t
Xbit_r86_c247 bl_247 br_247 wl_86 vdd gnd cell_6t
Xbit_r87_c247 bl_247 br_247 wl_87 vdd gnd cell_6t
Xbit_r88_c247 bl_247 br_247 wl_88 vdd gnd cell_6t
Xbit_r89_c247 bl_247 br_247 wl_89 vdd gnd cell_6t
Xbit_r90_c247 bl_247 br_247 wl_90 vdd gnd cell_6t
Xbit_r91_c247 bl_247 br_247 wl_91 vdd gnd cell_6t
Xbit_r92_c247 bl_247 br_247 wl_92 vdd gnd cell_6t
Xbit_r93_c247 bl_247 br_247 wl_93 vdd gnd cell_6t
Xbit_r94_c247 bl_247 br_247 wl_94 vdd gnd cell_6t
Xbit_r95_c247 bl_247 br_247 wl_95 vdd gnd cell_6t
Xbit_r96_c247 bl_247 br_247 wl_96 vdd gnd cell_6t
Xbit_r97_c247 bl_247 br_247 wl_97 vdd gnd cell_6t
Xbit_r98_c247 bl_247 br_247 wl_98 vdd gnd cell_6t
Xbit_r99_c247 bl_247 br_247 wl_99 vdd gnd cell_6t
Xbit_r100_c247 bl_247 br_247 wl_100 vdd gnd cell_6t
Xbit_r101_c247 bl_247 br_247 wl_101 vdd gnd cell_6t
Xbit_r102_c247 bl_247 br_247 wl_102 vdd gnd cell_6t
Xbit_r103_c247 bl_247 br_247 wl_103 vdd gnd cell_6t
Xbit_r104_c247 bl_247 br_247 wl_104 vdd gnd cell_6t
Xbit_r105_c247 bl_247 br_247 wl_105 vdd gnd cell_6t
Xbit_r106_c247 bl_247 br_247 wl_106 vdd gnd cell_6t
Xbit_r107_c247 bl_247 br_247 wl_107 vdd gnd cell_6t
Xbit_r108_c247 bl_247 br_247 wl_108 vdd gnd cell_6t
Xbit_r109_c247 bl_247 br_247 wl_109 vdd gnd cell_6t
Xbit_r110_c247 bl_247 br_247 wl_110 vdd gnd cell_6t
Xbit_r111_c247 bl_247 br_247 wl_111 vdd gnd cell_6t
Xbit_r112_c247 bl_247 br_247 wl_112 vdd gnd cell_6t
Xbit_r113_c247 bl_247 br_247 wl_113 vdd gnd cell_6t
Xbit_r114_c247 bl_247 br_247 wl_114 vdd gnd cell_6t
Xbit_r115_c247 bl_247 br_247 wl_115 vdd gnd cell_6t
Xbit_r116_c247 bl_247 br_247 wl_116 vdd gnd cell_6t
Xbit_r117_c247 bl_247 br_247 wl_117 vdd gnd cell_6t
Xbit_r118_c247 bl_247 br_247 wl_118 vdd gnd cell_6t
Xbit_r119_c247 bl_247 br_247 wl_119 vdd gnd cell_6t
Xbit_r120_c247 bl_247 br_247 wl_120 vdd gnd cell_6t
Xbit_r121_c247 bl_247 br_247 wl_121 vdd gnd cell_6t
Xbit_r122_c247 bl_247 br_247 wl_122 vdd gnd cell_6t
Xbit_r123_c247 bl_247 br_247 wl_123 vdd gnd cell_6t
Xbit_r124_c247 bl_247 br_247 wl_124 vdd gnd cell_6t
Xbit_r125_c247 bl_247 br_247 wl_125 vdd gnd cell_6t
Xbit_r126_c247 bl_247 br_247 wl_126 vdd gnd cell_6t
Xbit_r127_c247 bl_247 br_247 wl_127 vdd gnd cell_6t
Xbit_r128_c247 bl_247 br_247 wl_128 vdd gnd cell_6t
Xbit_r129_c247 bl_247 br_247 wl_129 vdd gnd cell_6t
Xbit_r130_c247 bl_247 br_247 wl_130 vdd gnd cell_6t
Xbit_r131_c247 bl_247 br_247 wl_131 vdd gnd cell_6t
Xbit_r132_c247 bl_247 br_247 wl_132 vdd gnd cell_6t
Xbit_r133_c247 bl_247 br_247 wl_133 vdd gnd cell_6t
Xbit_r134_c247 bl_247 br_247 wl_134 vdd gnd cell_6t
Xbit_r135_c247 bl_247 br_247 wl_135 vdd gnd cell_6t
Xbit_r136_c247 bl_247 br_247 wl_136 vdd gnd cell_6t
Xbit_r137_c247 bl_247 br_247 wl_137 vdd gnd cell_6t
Xbit_r138_c247 bl_247 br_247 wl_138 vdd gnd cell_6t
Xbit_r139_c247 bl_247 br_247 wl_139 vdd gnd cell_6t
Xbit_r140_c247 bl_247 br_247 wl_140 vdd gnd cell_6t
Xbit_r141_c247 bl_247 br_247 wl_141 vdd gnd cell_6t
Xbit_r142_c247 bl_247 br_247 wl_142 vdd gnd cell_6t
Xbit_r143_c247 bl_247 br_247 wl_143 vdd gnd cell_6t
Xbit_r144_c247 bl_247 br_247 wl_144 vdd gnd cell_6t
Xbit_r145_c247 bl_247 br_247 wl_145 vdd gnd cell_6t
Xbit_r146_c247 bl_247 br_247 wl_146 vdd gnd cell_6t
Xbit_r147_c247 bl_247 br_247 wl_147 vdd gnd cell_6t
Xbit_r148_c247 bl_247 br_247 wl_148 vdd gnd cell_6t
Xbit_r149_c247 bl_247 br_247 wl_149 vdd gnd cell_6t
Xbit_r150_c247 bl_247 br_247 wl_150 vdd gnd cell_6t
Xbit_r151_c247 bl_247 br_247 wl_151 vdd gnd cell_6t
Xbit_r152_c247 bl_247 br_247 wl_152 vdd gnd cell_6t
Xbit_r153_c247 bl_247 br_247 wl_153 vdd gnd cell_6t
Xbit_r154_c247 bl_247 br_247 wl_154 vdd gnd cell_6t
Xbit_r155_c247 bl_247 br_247 wl_155 vdd gnd cell_6t
Xbit_r156_c247 bl_247 br_247 wl_156 vdd gnd cell_6t
Xbit_r157_c247 bl_247 br_247 wl_157 vdd gnd cell_6t
Xbit_r158_c247 bl_247 br_247 wl_158 vdd gnd cell_6t
Xbit_r159_c247 bl_247 br_247 wl_159 vdd gnd cell_6t
Xbit_r160_c247 bl_247 br_247 wl_160 vdd gnd cell_6t
Xbit_r161_c247 bl_247 br_247 wl_161 vdd gnd cell_6t
Xbit_r162_c247 bl_247 br_247 wl_162 vdd gnd cell_6t
Xbit_r163_c247 bl_247 br_247 wl_163 vdd gnd cell_6t
Xbit_r164_c247 bl_247 br_247 wl_164 vdd gnd cell_6t
Xbit_r165_c247 bl_247 br_247 wl_165 vdd gnd cell_6t
Xbit_r166_c247 bl_247 br_247 wl_166 vdd gnd cell_6t
Xbit_r167_c247 bl_247 br_247 wl_167 vdd gnd cell_6t
Xbit_r168_c247 bl_247 br_247 wl_168 vdd gnd cell_6t
Xbit_r169_c247 bl_247 br_247 wl_169 vdd gnd cell_6t
Xbit_r170_c247 bl_247 br_247 wl_170 vdd gnd cell_6t
Xbit_r171_c247 bl_247 br_247 wl_171 vdd gnd cell_6t
Xbit_r172_c247 bl_247 br_247 wl_172 vdd gnd cell_6t
Xbit_r173_c247 bl_247 br_247 wl_173 vdd gnd cell_6t
Xbit_r174_c247 bl_247 br_247 wl_174 vdd gnd cell_6t
Xbit_r175_c247 bl_247 br_247 wl_175 vdd gnd cell_6t
Xbit_r176_c247 bl_247 br_247 wl_176 vdd gnd cell_6t
Xbit_r177_c247 bl_247 br_247 wl_177 vdd gnd cell_6t
Xbit_r178_c247 bl_247 br_247 wl_178 vdd gnd cell_6t
Xbit_r179_c247 bl_247 br_247 wl_179 vdd gnd cell_6t
Xbit_r180_c247 bl_247 br_247 wl_180 vdd gnd cell_6t
Xbit_r181_c247 bl_247 br_247 wl_181 vdd gnd cell_6t
Xbit_r182_c247 bl_247 br_247 wl_182 vdd gnd cell_6t
Xbit_r183_c247 bl_247 br_247 wl_183 vdd gnd cell_6t
Xbit_r184_c247 bl_247 br_247 wl_184 vdd gnd cell_6t
Xbit_r185_c247 bl_247 br_247 wl_185 vdd gnd cell_6t
Xbit_r186_c247 bl_247 br_247 wl_186 vdd gnd cell_6t
Xbit_r187_c247 bl_247 br_247 wl_187 vdd gnd cell_6t
Xbit_r188_c247 bl_247 br_247 wl_188 vdd gnd cell_6t
Xbit_r189_c247 bl_247 br_247 wl_189 vdd gnd cell_6t
Xbit_r190_c247 bl_247 br_247 wl_190 vdd gnd cell_6t
Xbit_r191_c247 bl_247 br_247 wl_191 vdd gnd cell_6t
Xbit_r192_c247 bl_247 br_247 wl_192 vdd gnd cell_6t
Xbit_r193_c247 bl_247 br_247 wl_193 vdd gnd cell_6t
Xbit_r194_c247 bl_247 br_247 wl_194 vdd gnd cell_6t
Xbit_r195_c247 bl_247 br_247 wl_195 vdd gnd cell_6t
Xbit_r196_c247 bl_247 br_247 wl_196 vdd gnd cell_6t
Xbit_r197_c247 bl_247 br_247 wl_197 vdd gnd cell_6t
Xbit_r198_c247 bl_247 br_247 wl_198 vdd gnd cell_6t
Xbit_r199_c247 bl_247 br_247 wl_199 vdd gnd cell_6t
Xbit_r200_c247 bl_247 br_247 wl_200 vdd gnd cell_6t
Xbit_r201_c247 bl_247 br_247 wl_201 vdd gnd cell_6t
Xbit_r202_c247 bl_247 br_247 wl_202 vdd gnd cell_6t
Xbit_r203_c247 bl_247 br_247 wl_203 vdd gnd cell_6t
Xbit_r204_c247 bl_247 br_247 wl_204 vdd gnd cell_6t
Xbit_r205_c247 bl_247 br_247 wl_205 vdd gnd cell_6t
Xbit_r206_c247 bl_247 br_247 wl_206 vdd gnd cell_6t
Xbit_r207_c247 bl_247 br_247 wl_207 vdd gnd cell_6t
Xbit_r208_c247 bl_247 br_247 wl_208 vdd gnd cell_6t
Xbit_r209_c247 bl_247 br_247 wl_209 vdd gnd cell_6t
Xbit_r210_c247 bl_247 br_247 wl_210 vdd gnd cell_6t
Xbit_r211_c247 bl_247 br_247 wl_211 vdd gnd cell_6t
Xbit_r212_c247 bl_247 br_247 wl_212 vdd gnd cell_6t
Xbit_r213_c247 bl_247 br_247 wl_213 vdd gnd cell_6t
Xbit_r214_c247 bl_247 br_247 wl_214 vdd gnd cell_6t
Xbit_r215_c247 bl_247 br_247 wl_215 vdd gnd cell_6t
Xbit_r216_c247 bl_247 br_247 wl_216 vdd gnd cell_6t
Xbit_r217_c247 bl_247 br_247 wl_217 vdd gnd cell_6t
Xbit_r218_c247 bl_247 br_247 wl_218 vdd gnd cell_6t
Xbit_r219_c247 bl_247 br_247 wl_219 vdd gnd cell_6t
Xbit_r220_c247 bl_247 br_247 wl_220 vdd gnd cell_6t
Xbit_r221_c247 bl_247 br_247 wl_221 vdd gnd cell_6t
Xbit_r222_c247 bl_247 br_247 wl_222 vdd gnd cell_6t
Xbit_r223_c247 bl_247 br_247 wl_223 vdd gnd cell_6t
Xbit_r224_c247 bl_247 br_247 wl_224 vdd gnd cell_6t
Xbit_r225_c247 bl_247 br_247 wl_225 vdd gnd cell_6t
Xbit_r226_c247 bl_247 br_247 wl_226 vdd gnd cell_6t
Xbit_r227_c247 bl_247 br_247 wl_227 vdd gnd cell_6t
Xbit_r228_c247 bl_247 br_247 wl_228 vdd gnd cell_6t
Xbit_r229_c247 bl_247 br_247 wl_229 vdd gnd cell_6t
Xbit_r230_c247 bl_247 br_247 wl_230 vdd gnd cell_6t
Xbit_r231_c247 bl_247 br_247 wl_231 vdd gnd cell_6t
Xbit_r232_c247 bl_247 br_247 wl_232 vdd gnd cell_6t
Xbit_r233_c247 bl_247 br_247 wl_233 vdd gnd cell_6t
Xbit_r234_c247 bl_247 br_247 wl_234 vdd gnd cell_6t
Xbit_r235_c247 bl_247 br_247 wl_235 vdd gnd cell_6t
Xbit_r236_c247 bl_247 br_247 wl_236 vdd gnd cell_6t
Xbit_r237_c247 bl_247 br_247 wl_237 vdd gnd cell_6t
Xbit_r238_c247 bl_247 br_247 wl_238 vdd gnd cell_6t
Xbit_r239_c247 bl_247 br_247 wl_239 vdd gnd cell_6t
Xbit_r240_c247 bl_247 br_247 wl_240 vdd gnd cell_6t
Xbit_r241_c247 bl_247 br_247 wl_241 vdd gnd cell_6t
Xbit_r242_c247 bl_247 br_247 wl_242 vdd gnd cell_6t
Xbit_r243_c247 bl_247 br_247 wl_243 vdd gnd cell_6t
Xbit_r244_c247 bl_247 br_247 wl_244 vdd gnd cell_6t
Xbit_r245_c247 bl_247 br_247 wl_245 vdd gnd cell_6t
Xbit_r246_c247 bl_247 br_247 wl_246 vdd gnd cell_6t
Xbit_r247_c247 bl_247 br_247 wl_247 vdd gnd cell_6t
Xbit_r248_c247 bl_247 br_247 wl_248 vdd gnd cell_6t
Xbit_r249_c247 bl_247 br_247 wl_249 vdd gnd cell_6t
Xbit_r250_c247 bl_247 br_247 wl_250 vdd gnd cell_6t
Xbit_r251_c247 bl_247 br_247 wl_251 vdd gnd cell_6t
Xbit_r252_c247 bl_247 br_247 wl_252 vdd gnd cell_6t
Xbit_r253_c247 bl_247 br_247 wl_253 vdd gnd cell_6t
Xbit_r254_c247 bl_247 br_247 wl_254 vdd gnd cell_6t
Xbit_r255_c247 bl_247 br_247 wl_255 vdd gnd cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd cell_6t
Xbit_r1_c248 bl_248 br_248 wl_1 vdd gnd cell_6t
Xbit_r2_c248 bl_248 br_248 wl_2 vdd gnd cell_6t
Xbit_r3_c248 bl_248 br_248 wl_3 vdd gnd cell_6t
Xbit_r4_c248 bl_248 br_248 wl_4 vdd gnd cell_6t
Xbit_r5_c248 bl_248 br_248 wl_5 vdd gnd cell_6t
Xbit_r6_c248 bl_248 br_248 wl_6 vdd gnd cell_6t
Xbit_r7_c248 bl_248 br_248 wl_7 vdd gnd cell_6t
Xbit_r8_c248 bl_248 br_248 wl_8 vdd gnd cell_6t
Xbit_r9_c248 bl_248 br_248 wl_9 vdd gnd cell_6t
Xbit_r10_c248 bl_248 br_248 wl_10 vdd gnd cell_6t
Xbit_r11_c248 bl_248 br_248 wl_11 vdd gnd cell_6t
Xbit_r12_c248 bl_248 br_248 wl_12 vdd gnd cell_6t
Xbit_r13_c248 bl_248 br_248 wl_13 vdd gnd cell_6t
Xbit_r14_c248 bl_248 br_248 wl_14 vdd gnd cell_6t
Xbit_r15_c248 bl_248 br_248 wl_15 vdd gnd cell_6t
Xbit_r16_c248 bl_248 br_248 wl_16 vdd gnd cell_6t
Xbit_r17_c248 bl_248 br_248 wl_17 vdd gnd cell_6t
Xbit_r18_c248 bl_248 br_248 wl_18 vdd gnd cell_6t
Xbit_r19_c248 bl_248 br_248 wl_19 vdd gnd cell_6t
Xbit_r20_c248 bl_248 br_248 wl_20 vdd gnd cell_6t
Xbit_r21_c248 bl_248 br_248 wl_21 vdd gnd cell_6t
Xbit_r22_c248 bl_248 br_248 wl_22 vdd gnd cell_6t
Xbit_r23_c248 bl_248 br_248 wl_23 vdd gnd cell_6t
Xbit_r24_c248 bl_248 br_248 wl_24 vdd gnd cell_6t
Xbit_r25_c248 bl_248 br_248 wl_25 vdd gnd cell_6t
Xbit_r26_c248 bl_248 br_248 wl_26 vdd gnd cell_6t
Xbit_r27_c248 bl_248 br_248 wl_27 vdd gnd cell_6t
Xbit_r28_c248 bl_248 br_248 wl_28 vdd gnd cell_6t
Xbit_r29_c248 bl_248 br_248 wl_29 vdd gnd cell_6t
Xbit_r30_c248 bl_248 br_248 wl_30 vdd gnd cell_6t
Xbit_r31_c248 bl_248 br_248 wl_31 vdd gnd cell_6t
Xbit_r32_c248 bl_248 br_248 wl_32 vdd gnd cell_6t
Xbit_r33_c248 bl_248 br_248 wl_33 vdd gnd cell_6t
Xbit_r34_c248 bl_248 br_248 wl_34 vdd gnd cell_6t
Xbit_r35_c248 bl_248 br_248 wl_35 vdd gnd cell_6t
Xbit_r36_c248 bl_248 br_248 wl_36 vdd gnd cell_6t
Xbit_r37_c248 bl_248 br_248 wl_37 vdd gnd cell_6t
Xbit_r38_c248 bl_248 br_248 wl_38 vdd gnd cell_6t
Xbit_r39_c248 bl_248 br_248 wl_39 vdd gnd cell_6t
Xbit_r40_c248 bl_248 br_248 wl_40 vdd gnd cell_6t
Xbit_r41_c248 bl_248 br_248 wl_41 vdd gnd cell_6t
Xbit_r42_c248 bl_248 br_248 wl_42 vdd gnd cell_6t
Xbit_r43_c248 bl_248 br_248 wl_43 vdd gnd cell_6t
Xbit_r44_c248 bl_248 br_248 wl_44 vdd gnd cell_6t
Xbit_r45_c248 bl_248 br_248 wl_45 vdd gnd cell_6t
Xbit_r46_c248 bl_248 br_248 wl_46 vdd gnd cell_6t
Xbit_r47_c248 bl_248 br_248 wl_47 vdd gnd cell_6t
Xbit_r48_c248 bl_248 br_248 wl_48 vdd gnd cell_6t
Xbit_r49_c248 bl_248 br_248 wl_49 vdd gnd cell_6t
Xbit_r50_c248 bl_248 br_248 wl_50 vdd gnd cell_6t
Xbit_r51_c248 bl_248 br_248 wl_51 vdd gnd cell_6t
Xbit_r52_c248 bl_248 br_248 wl_52 vdd gnd cell_6t
Xbit_r53_c248 bl_248 br_248 wl_53 vdd gnd cell_6t
Xbit_r54_c248 bl_248 br_248 wl_54 vdd gnd cell_6t
Xbit_r55_c248 bl_248 br_248 wl_55 vdd gnd cell_6t
Xbit_r56_c248 bl_248 br_248 wl_56 vdd gnd cell_6t
Xbit_r57_c248 bl_248 br_248 wl_57 vdd gnd cell_6t
Xbit_r58_c248 bl_248 br_248 wl_58 vdd gnd cell_6t
Xbit_r59_c248 bl_248 br_248 wl_59 vdd gnd cell_6t
Xbit_r60_c248 bl_248 br_248 wl_60 vdd gnd cell_6t
Xbit_r61_c248 bl_248 br_248 wl_61 vdd gnd cell_6t
Xbit_r62_c248 bl_248 br_248 wl_62 vdd gnd cell_6t
Xbit_r63_c248 bl_248 br_248 wl_63 vdd gnd cell_6t
Xbit_r64_c248 bl_248 br_248 wl_64 vdd gnd cell_6t
Xbit_r65_c248 bl_248 br_248 wl_65 vdd gnd cell_6t
Xbit_r66_c248 bl_248 br_248 wl_66 vdd gnd cell_6t
Xbit_r67_c248 bl_248 br_248 wl_67 vdd gnd cell_6t
Xbit_r68_c248 bl_248 br_248 wl_68 vdd gnd cell_6t
Xbit_r69_c248 bl_248 br_248 wl_69 vdd gnd cell_6t
Xbit_r70_c248 bl_248 br_248 wl_70 vdd gnd cell_6t
Xbit_r71_c248 bl_248 br_248 wl_71 vdd gnd cell_6t
Xbit_r72_c248 bl_248 br_248 wl_72 vdd gnd cell_6t
Xbit_r73_c248 bl_248 br_248 wl_73 vdd gnd cell_6t
Xbit_r74_c248 bl_248 br_248 wl_74 vdd gnd cell_6t
Xbit_r75_c248 bl_248 br_248 wl_75 vdd gnd cell_6t
Xbit_r76_c248 bl_248 br_248 wl_76 vdd gnd cell_6t
Xbit_r77_c248 bl_248 br_248 wl_77 vdd gnd cell_6t
Xbit_r78_c248 bl_248 br_248 wl_78 vdd gnd cell_6t
Xbit_r79_c248 bl_248 br_248 wl_79 vdd gnd cell_6t
Xbit_r80_c248 bl_248 br_248 wl_80 vdd gnd cell_6t
Xbit_r81_c248 bl_248 br_248 wl_81 vdd gnd cell_6t
Xbit_r82_c248 bl_248 br_248 wl_82 vdd gnd cell_6t
Xbit_r83_c248 bl_248 br_248 wl_83 vdd gnd cell_6t
Xbit_r84_c248 bl_248 br_248 wl_84 vdd gnd cell_6t
Xbit_r85_c248 bl_248 br_248 wl_85 vdd gnd cell_6t
Xbit_r86_c248 bl_248 br_248 wl_86 vdd gnd cell_6t
Xbit_r87_c248 bl_248 br_248 wl_87 vdd gnd cell_6t
Xbit_r88_c248 bl_248 br_248 wl_88 vdd gnd cell_6t
Xbit_r89_c248 bl_248 br_248 wl_89 vdd gnd cell_6t
Xbit_r90_c248 bl_248 br_248 wl_90 vdd gnd cell_6t
Xbit_r91_c248 bl_248 br_248 wl_91 vdd gnd cell_6t
Xbit_r92_c248 bl_248 br_248 wl_92 vdd gnd cell_6t
Xbit_r93_c248 bl_248 br_248 wl_93 vdd gnd cell_6t
Xbit_r94_c248 bl_248 br_248 wl_94 vdd gnd cell_6t
Xbit_r95_c248 bl_248 br_248 wl_95 vdd gnd cell_6t
Xbit_r96_c248 bl_248 br_248 wl_96 vdd gnd cell_6t
Xbit_r97_c248 bl_248 br_248 wl_97 vdd gnd cell_6t
Xbit_r98_c248 bl_248 br_248 wl_98 vdd gnd cell_6t
Xbit_r99_c248 bl_248 br_248 wl_99 vdd gnd cell_6t
Xbit_r100_c248 bl_248 br_248 wl_100 vdd gnd cell_6t
Xbit_r101_c248 bl_248 br_248 wl_101 vdd gnd cell_6t
Xbit_r102_c248 bl_248 br_248 wl_102 vdd gnd cell_6t
Xbit_r103_c248 bl_248 br_248 wl_103 vdd gnd cell_6t
Xbit_r104_c248 bl_248 br_248 wl_104 vdd gnd cell_6t
Xbit_r105_c248 bl_248 br_248 wl_105 vdd gnd cell_6t
Xbit_r106_c248 bl_248 br_248 wl_106 vdd gnd cell_6t
Xbit_r107_c248 bl_248 br_248 wl_107 vdd gnd cell_6t
Xbit_r108_c248 bl_248 br_248 wl_108 vdd gnd cell_6t
Xbit_r109_c248 bl_248 br_248 wl_109 vdd gnd cell_6t
Xbit_r110_c248 bl_248 br_248 wl_110 vdd gnd cell_6t
Xbit_r111_c248 bl_248 br_248 wl_111 vdd gnd cell_6t
Xbit_r112_c248 bl_248 br_248 wl_112 vdd gnd cell_6t
Xbit_r113_c248 bl_248 br_248 wl_113 vdd gnd cell_6t
Xbit_r114_c248 bl_248 br_248 wl_114 vdd gnd cell_6t
Xbit_r115_c248 bl_248 br_248 wl_115 vdd gnd cell_6t
Xbit_r116_c248 bl_248 br_248 wl_116 vdd gnd cell_6t
Xbit_r117_c248 bl_248 br_248 wl_117 vdd gnd cell_6t
Xbit_r118_c248 bl_248 br_248 wl_118 vdd gnd cell_6t
Xbit_r119_c248 bl_248 br_248 wl_119 vdd gnd cell_6t
Xbit_r120_c248 bl_248 br_248 wl_120 vdd gnd cell_6t
Xbit_r121_c248 bl_248 br_248 wl_121 vdd gnd cell_6t
Xbit_r122_c248 bl_248 br_248 wl_122 vdd gnd cell_6t
Xbit_r123_c248 bl_248 br_248 wl_123 vdd gnd cell_6t
Xbit_r124_c248 bl_248 br_248 wl_124 vdd gnd cell_6t
Xbit_r125_c248 bl_248 br_248 wl_125 vdd gnd cell_6t
Xbit_r126_c248 bl_248 br_248 wl_126 vdd gnd cell_6t
Xbit_r127_c248 bl_248 br_248 wl_127 vdd gnd cell_6t
Xbit_r128_c248 bl_248 br_248 wl_128 vdd gnd cell_6t
Xbit_r129_c248 bl_248 br_248 wl_129 vdd gnd cell_6t
Xbit_r130_c248 bl_248 br_248 wl_130 vdd gnd cell_6t
Xbit_r131_c248 bl_248 br_248 wl_131 vdd gnd cell_6t
Xbit_r132_c248 bl_248 br_248 wl_132 vdd gnd cell_6t
Xbit_r133_c248 bl_248 br_248 wl_133 vdd gnd cell_6t
Xbit_r134_c248 bl_248 br_248 wl_134 vdd gnd cell_6t
Xbit_r135_c248 bl_248 br_248 wl_135 vdd gnd cell_6t
Xbit_r136_c248 bl_248 br_248 wl_136 vdd gnd cell_6t
Xbit_r137_c248 bl_248 br_248 wl_137 vdd gnd cell_6t
Xbit_r138_c248 bl_248 br_248 wl_138 vdd gnd cell_6t
Xbit_r139_c248 bl_248 br_248 wl_139 vdd gnd cell_6t
Xbit_r140_c248 bl_248 br_248 wl_140 vdd gnd cell_6t
Xbit_r141_c248 bl_248 br_248 wl_141 vdd gnd cell_6t
Xbit_r142_c248 bl_248 br_248 wl_142 vdd gnd cell_6t
Xbit_r143_c248 bl_248 br_248 wl_143 vdd gnd cell_6t
Xbit_r144_c248 bl_248 br_248 wl_144 vdd gnd cell_6t
Xbit_r145_c248 bl_248 br_248 wl_145 vdd gnd cell_6t
Xbit_r146_c248 bl_248 br_248 wl_146 vdd gnd cell_6t
Xbit_r147_c248 bl_248 br_248 wl_147 vdd gnd cell_6t
Xbit_r148_c248 bl_248 br_248 wl_148 vdd gnd cell_6t
Xbit_r149_c248 bl_248 br_248 wl_149 vdd gnd cell_6t
Xbit_r150_c248 bl_248 br_248 wl_150 vdd gnd cell_6t
Xbit_r151_c248 bl_248 br_248 wl_151 vdd gnd cell_6t
Xbit_r152_c248 bl_248 br_248 wl_152 vdd gnd cell_6t
Xbit_r153_c248 bl_248 br_248 wl_153 vdd gnd cell_6t
Xbit_r154_c248 bl_248 br_248 wl_154 vdd gnd cell_6t
Xbit_r155_c248 bl_248 br_248 wl_155 vdd gnd cell_6t
Xbit_r156_c248 bl_248 br_248 wl_156 vdd gnd cell_6t
Xbit_r157_c248 bl_248 br_248 wl_157 vdd gnd cell_6t
Xbit_r158_c248 bl_248 br_248 wl_158 vdd gnd cell_6t
Xbit_r159_c248 bl_248 br_248 wl_159 vdd gnd cell_6t
Xbit_r160_c248 bl_248 br_248 wl_160 vdd gnd cell_6t
Xbit_r161_c248 bl_248 br_248 wl_161 vdd gnd cell_6t
Xbit_r162_c248 bl_248 br_248 wl_162 vdd gnd cell_6t
Xbit_r163_c248 bl_248 br_248 wl_163 vdd gnd cell_6t
Xbit_r164_c248 bl_248 br_248 wl_164 vdd gnd cell_6t
Xbit_r165_c248 bl_248 br_248 wl_165 vdd gnd cell_6t
Xbit_r166_c248 bl_248 br_248 wl_166 vdd gnd cell_6t
Xbit_r167_c248 bl_248 br_248 wl_167 vdd gnd cell_6t
Xbit_r168_c248 bl_248 br_248 wl_168 vdd gnd cell_6t
Xbit_r169_c248 bl_248 br_248 wl_169 vdd gnd cell_6t
Xbit_r170_c248 bl_248 br_248 wl_170 vdd gnd cell_6t
Xbit_r171_c248 bl_248 br_248 wl_171 vdd gnd cell_6t
Xbit_r172_c248 bl_248 br_248 wl_172 vdd gnd cell_6t
Xbit_r173_c248 bl_248 br_248 wl_173 vdd gnd cell_6t
Xbit_r174_c248 bl_248 br_248 wl_174 vdd gnd cell_6t
Xbit_r175_c248 bl_248 br_248 wl_175 vdd gnd cell_6t
Xbit_r176_c248 bl_248 br_248 wl_176 vdd gnd cell_6t
Xbit_r177_c248 bl_248 br_248 wl_177 vdd gnd cell_6t
Xbit_r178_c248 bl_248 br_248 wl_178 vdd gnd cell_6t
Xbit_r179_c248 bl_248 br_248 wl_179 vdd gnd cell_6t
Xbit_r180_c248 bl_248 br_248 wl_180 vdd gnd cell_6t
Xbit_r181_c248 bl_248 br_248 wl_181 vdd gnd cell_6t
Xbit_r182_c248 bl_248 br_248 wl_182 vdd gnd cell_6t
Xbit_r183_c248 bl_248 br_248 wl_183 vdd gnd cell_6t
Xbit_r184_c248 bl_248 br_248 wl_184 vdd gnd cell_6t
Xbit_r185_c248 bl_248 br_248 wl_185 vdd gnd cell_6t
Xbit_r186_c248 bl_248 br_248 wl_186 vdd gnd cell_6t
Xbit_r187_c248 bl_248 br_248 wl_187 vdd gnd cell_6t
Xbit_r188_c248 bl_248 br_248 wl_188 vdd gnd cell_6t
Xbit_r189_c248 bl_248 br_248 wl_189 vdd gnd cell_6t
Xbit_r190_c248 bl_248 br_248 wl_190 vdd gnd cell_6t
Xbit_r191_c248 bl_248 br_248 wl_191 vdd gnd cell_6t
Xbit_r192_c248 bl_248 br_248 wl_192 vdd gnd cell_6t
Xbit_r193_c248 bl_248 br_248 wl_193 vdd gnd cell_6t
Xbit_r194_c248 bl_248 br_248 wl_194 vdd gnd cell_6t
Xbit_r195_c248 bl_248 br_248 wl_195 vdd gnd cell_6t
Xbit_r196_c248 bl_248 br_248 wl_196 vdd gnd cell_6t
Xbit_r197_c248 bl_248 br_248 wl_197 vdd gnd cell_6t
Xbit_r198_c248 bl_248 br_248 wl_198 vdd gnd cell_6t
Xbit_r199_c248 bl_248 br_248 wl_199 vdd gnd cell_6t
Xbit_r200_c248 bl_248 br_248 wl_200 vdd gnd cell_6t
Xbit_r201_c248 bl_248 br_248 wl_201 vdd gnd cell_6t
Xbit_r202_c248 bl_248 br_248 wl_202 vdd gnd cell_6t
Xbit_r203_c248 bl_248 br_248 wl_203 vdd gnd cell_6t
Xbit_r204_c248 bl_248 br_248 wl_204 vdd gnd cell_6t
Xbit_r205_c248 bl_248 br_248 wl_205 vdd gnd cell_6t
Xbit_r206_c248 bl_248 br_248 wl_206 vdd gnd cell_6t
Xbit_r207_c248 bl_248 br_248 wl_207 vdd gnd cell_6t
Xbit_r208_c248 bl_248 br_248 wl_208 vdd gnd cell_6t
Xbit_r209_c248 bl_248 br_248 wl_209 vdd gnd cell_6t
Xbit_r210_c248 bl_248 br_248 wl_210 vdd gnd cell_6t
Xbit_r211_c248 bl_248 br_248 wl_211 vdd gnd cell_6t
Xbit_r212_c248 bl_248 br_248 wl_212 vdd gnd cell_6t
Xbit_r213_c248 bl_248 br_248 wl_213 vdd gnd cell_6t
Xbit_r214_c248 bl_248 br_248 wl_214 vdd gnd cell_6t
Xbit_r215_c248 bl_248 br_248 wl_215 vdd gnd cell_6t
Xbit_r216_c248 bl_248 br_248 wl_216 vdd gnd cell_6t
Xbit_r217_c248 bl_248 br_248 wl_217 vdd gnd cell_6t
Xbit_r218_c248 bl_248 br_248 wl_218 vdd gnd cell_6t
Xbit_r219_c248 bl_248 br_248 wl_219 vdd gnd cell_6t
Xbit_r220_c248 bl_248 br_248 wl_220 vdd gnd cell_6t
Xbit_r221_c248 bl_248 br_248 wl_221 vdd gnd cell_6t
Xbit_r222_c248 bl_248 br_248 wl_222 vdd gnd cell_6t
Xbit_r223_c248 bl_248 br_248 wl_223 vdd gnd cell_6t
Xbit_r224_c248 bl_248 br_248 wl_224 vdd gnd cell_6t
Xbit_r225_c248 bl_248 br_248 wl_225 vdd gnd cell_6t
Xbit_r226_c248 bl_248 br_248 wl_226 vdd gnd cell_6t
Xbit_r227_c248 bl_248 br_248 wl_227 vdd gnd cell_6t
Xbit_r228_c248 bl_248 br_248 wl_228 vdd gnd cell_6t
Xbit_r229_c248 bl_248 br_248 wl_229 vdd gnd cell_6t
Xbit_r230_c248 bl_248 br_248 wl_230 vdd gnd cell_6t
Xbit_r231_c248 bl_248 br_248 wl_231 vdd gnd cell_6t
Xbit_r232_c248 bl_248 br_248 wl_232 vdd gnd cell_6t
Xbit_r233_c248 bl_248 br_248 wl_233 vdd gnd cell_6t
Xbit_r234_c248 bl_248 br_248 wl_234 vdd gnd cell_6t
Xbit_r235_c248 bl_248 br_248 wl_235 vdd gnd cell_6t
Xbit_r236_c248 bl_248 br_248 wl_236 vdd gnd cell_6t
Xbit_r237_c248 bl_248 br_248 wl_237 vdd gnd cell_6t
Xbit_r238_c248 bl_248 br_248 wl_238 vdd gnd cell_6t
Xbit_r239_c248 bl_248 br_248 wl_239 vdd gnd cell_6t
Xbit_r240_c248 bl_248 br_248 wl_240 vdd gnd cell_6t
Xbit_r241_c248 bl_248 br_248 wl_241 vdd gnd cell_6t
Xbit_r242_c248 bl_248 br_248 wl_242 vdd gnd cell_6t
Xbit_r243_c248 bl_248 br_248 wl_243 vdd gnd cell_6t
Xbit_r244_c248 bl_248 br_248 wl_244 vdd gnd cell_6t
Xbit_r245_c248 bl_248 br_248 wl_245 vdd gnd cell_6t
Xbit_r246_c248 bl_248 br_248 wl_246 vdd gnd cell_6t
Xbit_r247_c248 bl_248 br_248 wl_247 vdd gnd cell_6t
Xbit_r248_c248 bl_248 br_248 wl_248 vdd gnd cell_6t
Xbit_r249_c248 bl_248 br_248 wl_249 vdd gnd cell_6t
Xbit_r250_c248 bl_248 br_248 wl_250 vdd gnd cell_6t
Xbit_r251_c248 bl_248 br_248 wl_251 vdd gnd cell_6t
Xbit_r252_c248 bl_248 br_248 wl_252 vdd gnd cell_6t
Xbit_r253_c248 bl_248 br_248 wl_253 vdd gnd cell_6t
Xbit_r254_c248 bl_248 br_248 wl_254 vdd gnd cell_6t
Xbit_r255_c248 bl_248 br_248 wl_255 vdd gnd cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd cell_6t
Xbit_r1_c249 bl_249 br_249 wl_1 vdd gnd cell_6t
Xbit_r2_c249 bl_249 br_249 wl_2 vdd gnd cell_6t
Xbit_r3_c249 bl_249 br_249 wl_3 vdd gnd cell_6t
Xbit_r4_c249 bl_249 br_249 wl_4 vdd gnd cell_6t
Xbit_r5_c249 bl_249 br_249 wl_5 vdd gnd cell_6t
Xbit_r6_c249 bl_249 br_249 wl_6 vdd gnd cell_6t
Xbit_r7_c249 bl_249 br_249 wl_7 vdd gnd cell_6t
Xbit_r8_c249 bl_249 br_249 wl_8 vdd gnd cell_6t
Xbit_r9_c249 bl_249 br_249 wl_9 vdd gnd cell_6t
Xbit_r10_c249 bl_249 br_249 wl_10 vdd gnd cell_6t
Xbit_r11_c249 bl_249 br_249 wl_11 vdd gnd cell_6t
Xbit_r12_c249 bl_249 br_249 wl_12 vdd gnd cell_6t
Xbit_r13_c249 bl_249 br_249 wl_13 vdd gnd cell_6t
Xbit_r14_c249 bl_249 br_249 wl_14 vdd gnd cell_6t
Xbit_r15_c249 bl_249 br_249 wl_15 vdd gnd cell_6t
Xbit_r16_c249 bl_249 br_249 wl_16 vdd gnd cell_6t
Xbit_r17_c249 bl_249 br_249 wl_17 vdd gnd cell_6t
Xbit_r18_c249 bl_249 br_249 wl_18 vdd gnd cell_6t
Xbit_r19_c249 bl_249 br_249 wl_19 vdd gnd cell_6t
Xbit_r20_c249 bl_249 br_249 wl_20 vdd gnd cell_6t
Xbit_r21_c249 bl_249 br_249 wl_21 vdd gnd cell_6t
Xbit_r22_c249 bl_249 br_249 wl_22 vdd gnd cell_6t
Xbit_r23_c249 bl_249 br_249 wl_23 vdd gnd cell_6t
Xbit_r24_c249 bl_249 br_249 wl_24 vdd gnd cell_6t
Xbit_r25_c249 bl_249 br_249 wl_25 vdd gnd cell_6t
Xbit_r26_c249 bl_249 br_249 wl_26 vdd gnd cell_6t
Xbit_r27_c249 bl_249 br_249 wl_27 vdd gnd cell_6t
Xbit_r28_c249 bl_249 br_249 wl_28 vdd gnd cell_6t
Xbit_r29_c249 bl_249 br_249 wl_29 vdd gnd cell_6t
Xbit_r30_c249 bl_249 br_249 wl_30 vdd gnd cell_6t
Xbit_r31_c249 bl_249 br_249 wl_31 vdd gnd cell_6t
Xbit_r32_c249 bl_249 br_249 wl_32 vdd gnd cell_6t
Xbit_r33_c249 bl_249 br_249 wl_33 vdd gnd cell_6t
Xbit_r34_c249 bl_249 br_249 wl_34 vdd gnd cell_6t
Xbit_r35_c249 bl_249 br_249 wl_35 vdd gnd cell_6t
Xbit_r36_c249 bl_249 br_249 wl_36 vdd gnd cell_6t
Xbit_r37_c249 bl_249 br_249 wl_37 vdd gnd cell_6t
Xbit_r38_c249 bl_249 br_249 wl_38 vdd gnd cell_6t
Xbit_r39_c249 bl_249 br_249 wl_39 vdd gnd cell_6t
Xbit_r40_c249 bl_249 br_249 wl_40 vdd gnd cell_6t
Xbit_r41_c249 bl_249 br_249 wl_41 vdd gnd cell_6t
Xbit_r42_c249 bl_249 br_249 wl_42 vdd gnd cell_6t
Xbit_r43_c249 bl_249 br_249 wl_43 vdd gnd cell_6t
Xbit_r44_c249 bl_249 br_249 wl_44 vdd gnd cell_6t
Xbit_r45_c249 bl_249 br_249 wl_45 vdd gnd cell_6t
Xbit_r46_c249 bl_249 br_249 wl_46 vdd gnd cell_6t
Xbit_r47_c249 bl_249 br_249 wl_47 vdd gnd cell_6t
Xbit_r48_c249 bl_249 br_249 wl_48 vdd gnd cell_6t
Xbit_r49_c249 bl_249 br_249 wl_49 vdd gnd cell_6t
Xbit_r50_c249 bl_249 br_249 wl_50 vdd gnd cell_6t
Xbit_r51_c249 bl_249 br_249 wl_51 vdd gnd cell_6t
Xbit_r52_c249 bl_249 br_249 wl_52 vdd gnd cell_6t
Xbit_r53_c249 bl_249 br_249 wl_53 vdd gnd cell_6t
Xbit_r54_c249 bl_249 br_249 wl_54 vdd gnd cell_6t
Xbit_r55_c249 bl_249 br_249 wl_55 vdd gnd cell_6t
Xbit_r56_c249 bl_249 br_249 wl_56 vdd gnd cell_6t
Xbit_r57_c249 bl_249 br_249 wl_57 vdd gnd cell_6t
Xbit_r58_c249 bl_249 br_249 wl_58 vdd gnd cell_6t
Xbit_r59_c249 bl_249 br_249 wl_59 vdd gnd cell_6t
Xbit_r60_c249 bl_249 br_249 wl_60 vdd gnd cell_6t
Xbit_r61_c249 bl_249 br_249 wl_61 vdd gnd cell_6t
Xbit_r62_c249 bl_249 br_249 wl_62 vdd gnd cell_6t
Xbit_r63_c249 bl_249 br_249 wl_63 vdd gnd cell_6t
Xbit_r64_c249 bl_249 br_249 wl_64 vdd gnd cell_6t
Xbit_r65_c249 bl_249 br_249 wl_65 vdd gnd cell_6t
Xbit_r66_c249 bl_249 br_249 wl_66 vdd gnd cell_6t
Xbit_r67_c249 bl_249 br_249 wl_67 vdd gnd cell_6t
Xbit_r68_c249 bl_249 br_249 wl_68 vdd gnd cell_6t
Xbit_r69_c249 bl_249 br_249 wl_69 vdd gnd cell_6t
Xbit_r70_c249 bl_249 br_249 wl_70 vdd gnd cell_6t
Xbit_r71_c249 bl_249 br_249 wl_71 vdd gnd cell_6t
Xbit_r72_c249 bl_249 br_249 wl_72 vdd gnd cell_6t
Xbit_r73_c249 bl_249 br_249 wl_73 vdd gnd cell_6t
Xbit_r74_c249 bl_249 br_249 wl_74 vdd gnd cell_6t
Xbit_r75_c249 bl_249 br_249 wl_75 vdd gnd cell_6t
Xbit_r76_c249 bl_249 br_249 wl_76 vdd gnd cell_6t
Xbit_r77_c249 bl_249 br_249 wl_77 vdd gnd cell_6t
Xbit_r78_c249 bl_249 br_249 wl_78 vdd gnd cell_6t
Xbit_r79_c249 bl_249 br_249 wl_79 vdd gnd cell_6t
Xbit_r80_c249 bl_249 br_249 wl_80 vdd gnd cell_6t
Xbit_r81_c249 bl_249 br_249 wl_81 vdd gnd cell_6t
Xbit_r82_c249 bl_249 br_249 wl_82 vdd gnd cell_6t
Xbit_r83_c249 bl_249 br_249 wl_83 vdd gnd cell_6t
Xbit_r84_c249 bl_249 br_249 wl_84 vdd gnd cell_6t
Xbit_r85_c249 bl_249 br_249 wl_85 vdd gnd cell_6t
Xbit_r86_c249 bl_249 br_249 wl_86 vdd gnd cell_6t
Xbit_r87_c249 bl_249 br_249 wl_87 vdd gnd cell_6t
Xbit_r88_c249 bl_249 br_249 wl_88 vdd gnd cell_6t
Xbit_r89_c249 bl_249 br_249 wl_89 vdd gnd cell_6t
Xbit_r90_c249 bl_249 br_249 wl_90 vdd gnd cell_6t
Xbit_r91_c249 bl_249 br_249 wl_91 vdd gnd cell_6t
Xbit_r92_c249 bl_249 br_249 wl_92 vdd gnd cell_6t
Xbit_r93_c249 bl_249 br_249 wl_93 vdd gnd cell_6t
Xbit_r94_c249 bl_249 br_249 wl_94 vdd gnd cell_6t
Xbit_r95_c249 bl_249 br_249 wl_95 vdd gnd cell_6t
Xbit_r96_c249 bl_249 br_249 wl_96 vdd gnd cell_6t
Xbit_r97_c249 bl_249 br_249 wl_97 vdd gnd cell_6t
Xbit_r98_c249 bl_249 br_249 wl_98 vdd gnd cell_6t
Xbit_r99_c249 bl_249 br_249 wl_99 vdd gnd cell_6t
Xbit_r100_c249 bl_249 br_249 wl_100 vdd gnd cell_6t
Xbit_r101_c249 bl_249 br_249 wl_101 vdd gnd cell_6t
Xbit_r102_c249 bl_249 br_249 wl_102 vdd gnd cell_6t
Xbit_r103_c249 bl_249 br_249 wl_103 vdd gnd cell_6t
Xbit_r104_c249 bl_249 br_249 wl_104 vdd gnd cell_6t
Xbit_r105_c249 bl_249 br_249 wl_105 vdd gnd cell_6t
Xbit_r106_c249 bl_249 br_249 wl_106 vdd gnd cell_6t
Xbit_r107_c249 bl_249 br_249 wl_107 vdd gnd cell_6t
Xbit_r108_c249 bl_249 br_249 wl_108 vdd gnd cell_6t
Xbit_r109_c249 bl_249 br_249 wl_109 vdd gnd cell_6t
Xbit_r110_c249 bl_249 br_249 wl_110 vdd gnd cell_6t
Xbit_r111_c249 bl_249 br_249 wl_111 vdd gnd cell_6t
Xbit_r112_c249 bl_249 br_249 wl_112 vdd gnd cell_6t
Xbit_r113_c249 bl_249 br_249 wl_113 vdd gnd cell_6t
Xbit_r114_c249 bl_249 br_249 wl_114 vdd gnd cell_6t
Xbit_r115_c249 bl_249 br_249 wl_115 vdd gnd cell_6t
Xbit_r116_c249 bl_249 br_249 wl_116 vdd gnd cell_6t
Xbit_r117_c249 bl_249 br_249 wl_117 vdd gnd cell_6t
Xbit_r118_c249 bl_249 br_249 wl_118 vdd gnd cell_6t
Xbit_r119_c249 bl_249 br_249 wl_119 vdd gnd cell_6t
Xbit_r120_c249 bl_249 br_249 wl_120 vdd gnd cell_6t
Xbit_r121_c249 bl_249 br_249 wl_121 vdd gnd cell_6t
Xbit_r122_c249 bl_249 br_249 wl_122 vdd gnd cell_6t
Xbit_r123_c249 bl_249 br_249 wl_123 vdd gnd cell_6t
Xbit_r124_c249 bl_249 br_249 wl_124 vdd gnd cell_6t
Xbit_r125_c249 bl_249 br_249 wl_125 vdd gnd cell_6t
Xbit_r126_c249 bl_249 br_249 wl_126 vdd gnd cell_6t
Xbit_r127_c249 bl_249 br_249 wl_127 vdd gnd cell_6t
Xbit_r128_c249 bl_249 br_249 wl_128 vdd gnd cell_6t
Xbit_r129_c249 bl_249 br_249 wl_129 vdd gnd cell_6t
Xbit_r130_c249 bl_249 br_249 wl_130 vdd gnd cell_6t
Xbit_r131_c249 bl_249 br_249 wl_131 vdd gnd cell_6t
Xbit_r132_c249 bl_249 br_249 wl_132 vdd gnd cell_6t
Xbit_r133_c249 bl_249 br_249 wl_133 vdd gnd cell_6t
Xbit_r134_c249 bl_249 br_249 wl_134 vdd gnd cell_6t
Xbit_r135_c249 bl_249 br_249 wl_135 vdd gnd cell_6t
Xbit_r136_c249 bl_249 br_249 wl_136 vdd gnd cell_6t
Xbit_r137_c249 bl_249 br_249 wl_137 vdd gnd cell_6t
Xbit_r138_c249 bl_249 br_249 wl_138 vdd gnd cell_6t
Xbit_r139_c249 bl_249 br_249 wl_139 vdd gnd cell_6t
Xbit_r140_c249 bl_249 br_249 wl_140 vdd gnd cell_6t
Xbit_r141_c249 bl_249 br_249 wl_141 vdd gnd cell_6t
Xbit_r142_c249 bl_249 br_249 wl_142 vdd gnd cell_6t
Xbit_r143_c249 bl_249 br_249 wl_143 vdd gnd cell_6t
Xbit_r144_c249 bl_249 br_249 wl_144 vdd gnd cell_6t
Xbit_r145_c249 bl_249 br_249 wl_145 vdd gnd cell_6t
Xbit_r146_c249 bl_249 br_249 wl_146 vdd gnd cell_6t
Xbit_r147_c249 bl_249 br_249 wl_147 vdd gnd cell_6t
Xbit_r148_c249 bl_249 br_249 wl_148 vdd gnd cell_6t
Xbit_r149_c249 bl_249 br_249 wl_149 vdd gnd cell_6t
Xbit_r150_c249 bl_249 br_249 wl_150 vdd gnd cell_6t
Xbit_r151_c249 bl_249 br_249 wl_151 vdd gnd cell_6t
Xbit_r152_c249 bl_249 br_249 wl_152 vdd gnd cell_6t
Xbit_r153_c249 bl_249 br_249 wl_153 vdd gnd cell_6t
Xbit_r154_c249 bl_249 br_249 wl_154 vdd gnd cell_6t
Xbit_r155_c249 bl_249 br_249 wl_155 vdd gnd cell_6t
Xbit_r156_c249 bl_249 br_249 wl_156 vdd gnd cell_6t
Xbit_r157_c249 bl_249 br_249 wl_157 vdd gnd cell_6t
Xbit_r158_c249 bl_249 br_249 wl_158 vdd gnd cell_6t
Xbit_r159_c249 bl_249 br_249 wl_159 vdd gnd cell_6t
Xbit_r160_c249 bl_249 br_249 wl_160 vdd gnd cell_6t
Xbit_r161_c249 bl_249 br_249 wl_161 vdd gnd cell_6t
Xbit_r162_c249 bl_249 br_249 wl_162 vdd gnd cell_6t
Xbit_r163_c249 bl_249 br_249 wl_163 vdd gnd cell_6t
Xbit_r164_c249 bl_249 br_249 wl_164 vdd gnd cell_6t
Xbit_r165_c249 bl_249 br_249 wl_165 vdd gnd cell_6t
Xbit_r166_c249 bl_249 br_249 wl_166 vdd gnd cell_6t
Xbit_r167_c249 bl_249 br_249 wl_167 vdd gnd cell_6t
Xbit_r168_c249 bl_249 br_249 wl_168 vdd gnd cell_6t
Xbit_r169_c249 bl_249 br_249 wl_169 vdd gnd cell_6t
Xbit_r170_c249 bl_249 br_249 wl_170 vdd gnd cell_6t
Xbit_r171_c249 bl_249 br_249 wl_171 vdd gnd cell_6t
Xbit_r172_c249 bl_249 br_249 wl_172 vdd gnd cell_6t
Xbit_r173_c249 bl_249 br_249 wl_173 vdd gnd cell_6t
Xbit_r174_c249 bl_249 br_249 wl_174 vdd gnd cell_6t
Xbit_r175_c249 bl_249 br_249 wl_175 vdd gnd cell_6t
Xbit_r176_c249 bl_249 br_249 wl_176 vdd gnd cell_6t
Xbit_r177_c249 bl_249 br_249 wl_177 vdd gnd cell_6t
Xbit_r178_c249 bl_249 br_249 wl_178 vdd gnd cell_6t
Xbit_r179_c249 bl_249 br_249 wl_179 vdd gnd cell_6t
Xbit_r180_c249 bl_249 br_249 wl_180 vdd gnd cell_6t
Xbit_r181_c249 bl_249 br_249 wl_181 vdd gnd cell_6t
Xbit_r182_c249 bl_249 br_249 wl_182 vdd gnd cell_6t
Xbit_r183_c249 bl_249 br_249 wl_183 vdd gnd cell_6t
Xbit_r184_c249 bl_249 br_249 wl_184 vdd gnd cell_6t
Xbit_r185_c249 bl_249 br_249 wl_185 vdd gnd cell_6t
Xbit_r186_c249 bl_249 br_249 wl_186 vdd gnd cell_6t
Xbit_r187_c249 bl_249 br_249 wl_187 vdd gnd cell_6t
Xbit_r188_c249 bl_249 br_249 wl_188 vdd gnd cell_6t
Xbit_r189_c249 bl_249 br_249 wl_189 vdd gnd cell_6t
Xbit_r190_c249 bl_249 br_249 wl_190 vdd gnd cell_6t
Xbit_r191_c249 bl_249 br_249 wl_191 vdd gnd cell_6t
Xbit_r192_c249 bl_249 br_249 wl_192 vdd gnd cell_6t
Xbit_r193_c249 bl_249 br_249 wl_193 vdd gnd cell_6t
Xbit_r194_c249 bl_249 br_249 wl_194 vdd gnd cell_6t
Xbit_r195_c249 bl_249 br_249 wl_195 vdd gnd cell_6t
Xbit_r196_c249 bl_249 br_249 wl_196 vdd gnd cell_6t
Xbit_r197_c249 bl_249 br_249 wl_197 vdd gnd cell_6t
Xbit_r198_c249 bl_249 br_249 wl_198 vdd gnd cell_6t
Xbit_r199_c249 bl_249 br_249 wl_199 vdd gnd cell_6t
Xbit_r200_c249 bl_249 br_249 wl_200 vdd gnd cell_6t
Xbit_r201_c249 bl_249 br_249 wl_201 vdd gnd cell_6t
Xbit_r202_c249 bl_249 br_249 wl_202 vdd gnd cell_6t
Xbit_r203_c249 bl_249 br_249 wl_203 vdd gnd cell_6t
Xbit_r204_c249 bl_249 br_249 wl_204 vdd gnd cell_6t
Xbit_r205_c249 bl_249 br_249 wl_205 vdd gnd cell_6t
Xbit_r206_c249 bl_249 br_249 wl_206 vdd gnd cell_6t
Xbit_r207_c249 bl_249 br_249 wl_207 vdd gnd cell_6t
Xbit_r208_c249 bl_249 br_249 wl_208 vdd gnd cell_6t
Xbit_r209_c249 bl_249 br_249 wl_209 vdd gnd cell_6t
Xbit_r210_c249 bl_249 br_249 wl_210 vdd gnd cell_6t
Xbit_r211_c249 bl_249 br_249 wl_211 vdd gnd cell_6t
Xbit_r212_c249 bl_249 br_249 wl_212 vdd gnd cell_6t
Xbit_r213_c249 bl_249 br_249 wl_213 vdd gnd cell_6t
Xbit_r214_c249 bl_249 br_249 wl_214 vdd gnd cell_6t
Xbit_r215_c249 bl_249 br_249 wl_215 vdd gnd cell_6t
Xbit_r216_c249 bl_249 br_249 wl_216 vdd gnd cell_6t
Xbit_r217_c249 bl_249 br_249 wl_217 vdd gnd cell_6t
Xbit_r218_c249 bl_249 br_249 wl_218 vdd gnd cell_6t
Xbit_r219_c249 bl_249 br_249 wl_219 vdd gnd cell_6t
Xbit_r220_c249 bl_249 br_249 wl_220 vdd gnd cell_6t
Xbit_r221_c249 bl_249 br_249 wl_221 vdd gnd cell_6t
Xbit_r222_c249 bl_249 br_249 wl_222 vdd gnd cell_6t
Xbit_r223_c249 bl_249 br_249 wl_223 vdd gnd cell_6t
Xbit_r224_c249 bl_249 br_249 wl_224 vdd gnd cell_6t
Xbit_r225_c249 bl_249 br_249 wl_225 vdd gnd cell_6t
Xbit_r226_c249 bl_249 br_249 wl_226 vdd gnd cell_6t
Xbit_r227_c249 bl_249 br_249 wl_227 vdd gnd cell_6t
Xbit_r228_c249 bl_249 br_249 wl_228 vdd gnd cell_6t
Xbit_r229_c249 bl_249 br_249 wl_229 vdd gnd cell_6t
Xbit_r230_c249 bl_249 br_249 wl_230 vdd gnd cell_6t
Xbit_r231_c249 bl_249 br_249 wl_231 vdd gnd cell_6t
Xbit_r232_c249 bl_249 br_249 wl_232 vdd gnd cell_6t
Xbit_r233_c249 bl_249 br_249 wl_233 vdd gnd cell_6t
Xbit_r234_c249 bl_249 br_249 wl_234 vdd gnd cell_6t
Xbit_r235_c249 bl_249 br_249 wl_235 vdd gnd cell_6t
Xbit_r236_c249 bl_249 br_249 wl_236 vdd gnd cell_6t
Xbit_r237_c249 bl_249 br_249 wl_237 vdd gnd cell_6t
Xbit_r238_c249 bl_249 br_249 wl_238 vdd gnd cell_6t
Xbit_r239_c249 bl_249 br_249 wl_239 vdd gnd cell_6t
Xbit_r240_c249 bl_249 br_249 wl_240 vdd gnd cell_6t
Xbit_r241_c249 bl_249 br_249 wl_241 vdd gnd cell_6t
Xbit_r242_c249 bl_249 br_249 wl_242 vdd gnd cell_6t
Xbit_r243_c249 bl_249 br_249 wl_243 vdd gnd cell_6t
Xbit_r244_c249 bl_249 br_249 wl_244 vdd gnd cell_6t
Xbit_r245_c249 bl_249 br_249 wl_245 vdd gnd cell_6t
Xbit_r246_c249 bl_249 br_249 wl_246 vdd gnd cell_6t
Xbit_r247_c249 bl_249 br_249 wl_247 vdd gnd cell_6t
Xbit_r248_c249 bl_249 br_249 wl_248 vdd gnd cell_6t
Xbit_r249_c249 bl_249 br_249 wl_249 vdd gnd cell_6t
Xbit_r250_c249 bl_249 br_249 wl_250 vdd gnd cell_6t
Xbit_r251_c249 bl_249 br_249 wl_251 vdd gnd cell_6t
Xbit_r252_c249 bl_249 br_249 wl_252 vdd gnd cell_6t
Xbit_r253_c249 bl_249 br_249 wl_253 vdd gnd cell_6t
Xbit_r254_c249 bl_249 br_249 wl_254 vdd gnd cell_6t
Xbit_r255_c249 bl_249 br_249 wl_255 vdd gnd cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd cell_6t
Xbit_r1_c250 bl_250 br_250 wl_1 vdd gnd cell_6t
Xbit_r2_c250 bl_250 br_250 wl_2 vdd gnd cell_6t
Xbit_r3_c250 bl_250 br_250 wl_3 vdd gnd cell_6t
Xbit_r4_c250 bl_250 br_250 wl_4 vdd gnd cell_6t
Xbit_r5_c250 bl_250 br_250 wl_5 vdd gnd cell_6t
Xbit_r6_c250 bl_250 br_250 wl_6 vdd gnd cell_6t
Xbit_r7_c250 bl_250 br_250 wl_7 vdd gnd cell_6t
Xbit_r8_c250 bl_250 br_250 wl_8 vdd gnd cell_6t
Xbit_r9_c250 bl_250 br_250 wl_9 vdd gnd cell_6t
Xbit_r10_c250 bl_250 br_250 wl_10 vdd gnd cell_6t
Xbit_r11_c250 bl_250 br_250 wl_11 vdd gnd cell_6t
Xbit_r12_c250 bl_250 br_250 wl_12 vdd gnd cell_6t
Xbit_r13_c250 bl_250 br_250 wl_13 vdd gnd cell_6t
Xbit_r14_c250 bl_250 br_250 wl_14 vdd gnd cell_6t
Xbit_r15_c250 bl_250 br_250 wl_15 vdd gnd cell_6t
Xbit_r16_c250 bl_250 br_250 wl_16 vdd gnd cell_6t
Xbit_r17_c250 bl_250 br_250 wl_17 vdd gnd cell_6t
Xbit_r18_c250 bl_250 br_250 wl_18 vdd gnd cell_6t
Xbit_r19_c250 bl_250 br_250 wl_19 vdd gnd cell_6t
Xbit_r20_c250 bl_250 br_250 wl_20 vdd gnd cell_6t
Xbit_r21_c250 bl_250 br_250 wl_21 vdd gnd cell_6t
Xbit_r22_c250 bl_250 br_250 wl_22 vdd gnd cell_6t
Xbit_r23_c250 bl_250 br_250 wl_23 vdd gnd cell_6t
Xbit_r24_c250 bl_250 br_250 wl_24 vdd gnd cell_6t
Xbit_r25_c250 bl_250 br_250 wl_25 vdd gnd cell_6t
Xbit_r26_c250 bl_250 br_250 wl_26 vdd gnd cell_6t
Xbit_r27_c250 bl_250 br_250 wl_27 vdd gnd cell_6t
Xbit_r28_c250 bl_250 br_250 wl_28 vdd gnd cell_6t
Xbit_r29_c250 bl_250 br_250 wl_29 vdd gnd cell_6t
Xbit_r30_c250 bl_250 br_250 wl_30 vdd gnd cell_6t
Xbit_r31_c250 bl_250 br_250 wl_31 vdd gnd cell_6t
Xbit_r32_c250 bl_250 br_250 wl_32 vdd gnd cell_6t
Xbit_r33_c250 bl_250 br_250 wl_33 vdd gnd cell_6t
Xbit_r34_c250 bl_250 br_250 wl_34 vdd gnd cell_6t
Xbit_r35_c250 bl_250 br_250 wl_35 vdd gnd cell_6t
Xbit_r36_c250 bl_250 br_250 wl_36 vdd gnd cell_6t
Xbit_r37_c250 bl_250 br_250 wl_37 vdd gnd cell_6t
Xbit_r38_c250 bl_250 br_250 wl_38 vdd gnd cell_6t
Xbit_r39_c250 bl_250 br_250 wl_39 vdd gnd cell_6t
Xbit_r40_c250 bl_250 br_250 wl_40 vdd gnd cell_6t
Xbit_r41_c250 bl_250 br_250 wl_41 vdd gnd cell_6t
Xbit_r42_c250 bl_250 br_250 wl_42 vdd gnd cell_6t
Xbit_r43_c250 bl_250 br_250 wl_43 vdd gnd cell_6t
Xbit_r44_c250 bl_250 br_250 wl_44 vdd gnd cell_6t
Xbit_r45_c250 bl_250 br_250 wl_45 vdd gnd cell_6t
Xbit_r46_c250 bl_250 br_250 wl_46 vdd gnd cell_6t
Xbit_r47_c250 bl_250 br_250 wl_47 vdd gnd cell_6t
Xbit_r48_c250 bl_250 br_250 wl_48 vdd gnd cell_6t
Xbit_r49_c250 bl_250 br_250 wl_49 vdd gnd cell_6t
Xbit_r50_c250 bl_250 br_250 wl_50 vdd gnd cell_6t
Xbit_r51_c250 bl_250 br_250 wl_51 vdd gnd cell_6t
Xbit_r52_c250 bl_250 br_250 wl_52 vdd gnd cell_6t
Xbit_r53_c250 bl_250 br_250 wl_53 vdd gnd cell_6t
Xbit_r54_c250 bl_250 br_250 wl_54 vdd gnd cell_6t
Xbit_r55_c250 bl_250 br_250 wl_55 vdd gnd cell_6t
Xbit_r56_c250 bl_250 br_250 wl_56 vdd gnd cell_6t
Xbit_r57_c250 bl_250 br_250 wl_57 vdd gnd cell_6t
Xbit_r58_c250 bl_250 br_250 wl_58 vdd gnd cell_6t
Xbit_r59_c250 bl_250 br_250 wl_59 vdd gnd cell_6t
Xbit_r60_c250 bl_250 br_250 wl_60 vdd gnd cell_6t
Xbit_r61_c250 bl_250 br_250 wl_61 vdd gnd cell_6t
Xbit_r62_c250 bl_250 br_250 wl_62 vdd gnd cell_6t
Xbit_r63_c250 bl_250 br_250 wl_63 vdd gnd cell_6t
Xbit_r64_c250 bl_250 br_250 wl_64 vdd gnd cell_6t
Xbit_r65_c250 bl_250 br_250 wl_65 vdd gnd cell_6t
Xbit_r66_c250 bl_250 br_250 wl_66 vdd gnd cell_6t
Xbit_r67_c250 bl_250 br_250 wl_67 vdd gnd cell_6t
Xbit_r68_c250 bl_250 br_250 wl_68 vdd gnd cell_6t
Xbit_r69_c250 bl_250 br_250 wl_69 vdd gnd cell_6t
Xbit_r70_c250 bl_250 br_250 wl_70 vdd gnd cell_6t
Xbit_r71_c250 bl_250 br_250 wl_71 vdd gnd cell_6t
Xbit_r72_c250 bl_250 br_250 wl_72 vdd gnd cell_6t
Xbit_r73_c250 bl_250 br_250 wl_73 vdd gnd cell_6t
Xbit_r74_c250 bl_250 br_250 wl_74 vdd gnd cell_6t
Xbit_r75_c250 bl_250 br_250 wl_75 vdd gnd cell_6t
Xbit_r76_c250 bl_250 br_250 wl_76 vdd gnd cell_6t
Xbit_r77_c250 bl_250 br_250 wl_77 vdd gnd cell_6t
Xbit_r78_c250 bl_250 br_250 wl_78 vdd gnd cell_6t
Xbit_r79_c250 bl_250 br_250 wl_79 vdd gnd cell_6t
Xbit_r80_c250 bl_250 br_250 wl_80 vdd gnd cell_6t
Xbit_r81_c250 bl_250 br_250 wl_81 vdd gnd cell_6t
Xbit_r82_c250 bl_250 br_250 wl_82 vdd gnd cell_6t
Xbit_r83_c250 bl_250 br_250 wl_83 vdd gnd cell_6t
Xbit_r84_c250 bl_250 br_250 wl_84 vdd gnd cell_6t
Xbit_r85_c250 bl_250 br_250 wl_85 vdd gnd cell_6t
Xbit_r86_c250 bl_250 br_250 wl_86 vdd gnd cell_6t
Xbit_r87_c250 bl_250 br_250 wl_87 vdd gnd cell_6t
Xbit_r88_c250 bl_250 br_250 wl_88 vdd gnd cell_6t
Xbit_r89_c250 bl_250 br_250 wl_89 vdd gnd cell_6t
Xbit_r90_c250 bl_250 br_250 wl_90 vdd gnd cell_6t
Xbit_r91_c250 bl_250 br_250 wl_91 vdd gnd cell_6t
Xbit_r92_c250 bl_250 br_250 wl_92 vdd gnd cell_6t
Xbit_r93_c250 bl_250 br_250 wl_93 vdd gnd cell_6t
Xbit_r94_c250 bl_250 br_250 wl_94 vdd gnd cell_6t
Xbit_r95_c250 bl_250 br_250 wl_95 vdd gnd cell_6t
Xbit_r96_c250 bl_250 br_250 wl_96 vdd gnd cell_6t
Xbit_r97_c250 bl_250 br_250 wl_97 vdd gnd cell_6t
Xbit_r98_c250 bl_250 br_250 wl_98 vdd gnd cell_6t
Xbit_r99_c250 bl_250 br_250 wl_99 vdd gnd cell_6t
Xbit_r100_c250 bl_250 br_250 wl_100 vdd gnd cell_6t
Xbit_r101_c250 bl_250 br_250 wl_101 vdd gnd cell_6t
Xbit_r102_c250 bl_250 br_250 wl_102 vdd gnd cell_6t
Xbit_r103_c250 bl_250 br_250 wl_103 vdd gnd cell_6t
Xbit_r104_c250 bl_250 br_250 wl_104 vdd gnd cell_6t
Xbit_r105_c250 bl_250 br_250 wl_105 vdd gnd cell_6t
Xbit_r106_c250 bl_250 br_250 wl_106 vdd gnd cell_6t
Xbit_r107_c250 bl_250 br_250 wl_107 vdd gnd cell_6t
Xbit_r108_c250 bl_250 br_250 wl_108 vdd gnd cell_6t
Xbit_r109_c250 bl_250 br_250 wl_109 vdd gnd cell_6t
Xbit_r110_c250 bl_250 br_250 wl_110 vdd gnd cell_6t
Xbit_r111_c250 bl_250 br_250 wl_111 vdd gnd cell_6t
Xbit_r112_c250 bl_250 br_250 wl_112 vdd gnd cell_6t
Xbit_r113_c250 bl_250 br_250 wl_113 vdd gnd cell_6t
Xbit_r114_c250 bl_250 br_250 wl_114 vdd gnd cell_6t
Xbit_r115_c250 bl_250 br_250 wl_115 vdd gnd cell_6t
Xbit_r116_c250 bl_250 br_250 wl_116 vdd gnd cell_6t
Xbit_r117_c250 bl_250 br_250 wl_117 vdd gnd cell_6t
Xbit_r118_c250 bl_250 br_250 wl_118 vdd gnd cell_6t
Xbit_r119_c250 bl_250 br_250 wl_119 vdd gnd cell_6t
Xbit_r120_c250 bl_250 br_250 wl_120 vdd gnd cell_6t
Xbit_r121_c250 bl_250 br_250 wl_121 vdd gnd cell_6t
Xbit_r122_c250 bl_250 br_250 wl_122 vdd gnd cell_6t
Xbit_r123_c250 bl_250 br_250 wl_123 vdd gnd cell_6t
Xbit_r124_c250 bl_250 br_250 wl_124 vdd gnd cell_6t
Xbit_r125_c250 bl_250 br_250 wl_125 vdd gnd cell_6t
Xbit_r126_c250 bl_250 br_250 wl_126 vdd gnd cell_6t
Xbit_r127_c250 bl_250 br_250 wl_127 vdd gnd cell_6t
Xbit_r128_c250 bl_250 br_250 wl_128 vdd gnd cell_6t
Xbit_r129_c250 bl_250 br_250 wl_129 vdd gnd cell_6t
Xbit_r130_c250 bl_250 br_250 wl_130 vdd gnd cell_6t
Xbit_r131_c250 bl_250 br_250 wl_131 vdd gnd cell_6t
Xbit_r132_c250 bl_250 br_250 wl_132 vdd gnd cell_6t
Xbit_r133_c250 bl_250 br_250 wl_133 vdd gnd cell_6t
Xbit_r134_c250 bl_250 br_250 wl_134 vdd gnd cell_6t
Xbit_r135_c250 bl_250 br_250 wl_135 vdd gnd cell_6t
Xbit_r136_c250 bl_250 br_250 wl_136 vdd gnd cell_6t
Xbit_r137_c250 bl_250 br_250 wl_137 vdd gnd cell_6t
Xbit_r138_c250 bl_250 br_250 wl_138 vdd gnd cell_6t
Xbit_r139_c250 bl_250 br_250 wl_139 vdd gnd cell_6t
Xbit_r140_c250 bl_250 br_250 wl_140 vdd gnd cell_6t
Xbit_r141_c250 bl_250 br_250 wl_141 vdd gnd cell_6t
Xbit_r142_c250 bl_250 br_250 wl_142 vdd gnd cell_6t
Xbit_r143_c250 bl_250 br_250 wl_143 vdd gnd cell_6t
Xbit_r144_c250 bl_250 br_250 wl_144 vdd gnd cell_6t
Xbit_r145_c250 bl_250 br_250 wl_145 vdd gnd cell_6t
Xbit_r146_c250 bl_250 br_250 wl_146 vdd gnd cell_6t
Xbit_r147_c250 bl_250 br_250 wl_147 vdd gnd cell_6t
Xbit_r148_c250 bl_250 br_250 wl_148 vdd gnd cell_6t
Xbit_r149_c250 bl_250 br_250 wl_149 vdd gnd cell_6t
Xbit_r150_c250 bl_250 br_250 wl_150 vdd gnd cell_6t
Xbit_r151_c250 bl_250 br_250 wl_151 vdd gnd cell_6t
Xbit_r152_c250 bl_250 br_250 wl_152 vdd gnd cell_6t
Xbit_r153_c250 bl_250 br_250 wl_153 vdd gnd cell_6t
Xbit_r154_c250 bl_250 br_250 wl_154 vdd gnd cell_6t
Xbit_r155_c250 bl_250 br_250 wl_155 vdd gnd cell_6t
Xbit_r156_c250 bl_250 br_250 wl_156 vdd gnd cell_6t
Xbit_r157_c250 bl_250 br_250 wl_157 vdd gnd cell_6t
Xbit_r158_c250 bl_250 br_250 wl_158 vdd gnd cell_6t
Xbit_r159_c250 bl_250 br_250 wl_159 vdd gnd cell_6t
Xbit_r160_c250 bl_250 br_250 wl_160 vdd gnd cell_6t
Xbit_r161_c250 bl_250 br_250 wl_161 vdd gnd cell_6t
Xbit_r162_c250 bl_250 br_250 wl_162 vdd gnd cell_6t
Xbit_r163_c250 bl_250 br_250 wl_163 vdd gnd cell_6t
Xbit_r164_c250 bl_250 br_250 wl_164 vdd gnd cell_6t
Xbit_r165_c250 bl_250 br_250 wl_165 vdd gnd cell_6t
Xbit_r166_c250 bl_250 br_250 wl_166 vdd gnd cell_6t
Xbit_r167_c250 bl_250 br_250 wl_167 vdd gnd cell_6t
Xbit_r168_c250 bl_250 br_250 wl_168 vdd gnd cell_6t
Xbit_r169_c250 bl_250 br_250 wl_169 vdd gnd cell_6t
Xbit_r170_c250 bl_250 br_250 wl_170 vdd gnd cell_6t
Xbit_r171_c250 bl_250 br_250 wl_171 vdd gnd cell_6t
Xbit_r172_c250 bl_250 br_250 wl_172 vdd gnd cell_6t
Xbit_r173_c250 bl_250 br_250 wl_173 vdd gnd cell_6t
Xbit_r174_c250 bl_250 br_250 wl_174 vdd gnd cell_6t
Xbit_r175_c250 bl_250 br_250 wl_175 vdd gnd cell_6t
Xbit_r176_c250 bl_250 br_250 wl_176 vdd gnd cell_6t
Xbit_r177_c250 bl_250 br_250 wl_177 vdd gnd cell_6t
Xbit_r178_c250 bl_250 br_250 wl_178 vdd gnd cell_6t
Xbit_r179_c250 bl_250 br_250 wl_179 vdd gnd cell_6t
Xbit_r180_c250 bl_250 br_250 wl_180 vdd gnd cell_6t
Xbit_r181_c250 bl_250 br_250 wl_181 vdd gnd cell_6t
Xbit_r182_c250 bl_250 br_250 wl_182 vdd gnd cell_6t
Xbit_r183_c250 bl_250 br_250 wl_183 vdd gnd cell_6t
Xbit_r184_c250 bl_250 br_250 wl_184 vdd gnd cell_6t
Xbit_r185_c250 bl_250 br_250 wl_185 vdd gnd cell_6t
Xbit_r186_c250 bl_250 br_250 wl_186 vdd gnd cell_6t
Xbit_r187_c250 bl_250 br_250 wl_187 vdd gnd cell_6t
Xbit_r188_c250 bl_250 br_250 wl_188 vdd gnd cell_6t
Xbit_r189_c250 bl_250 br_250 wl_189 vdd gnd cell_6t
Xbit_r190_c250 bl_250 br_250 wl_190 vdd gnd cell_6t
Xbit_r191_c250 bl_250 br_250 wl_191 vdd gnd cell_6t
Xbit_r192_c250 bl_250 br_250 wl_192 vdd gnd cell_6t
Xbit_r193_c250 bl_250 br_250 wl_193 vdd gnd cell_6t
Xbit_r194_c250 bl_250 br_250 wl_194 vdd gnd cell_6t
Xbit_r195_c250 bl_250 br_250 wl_195 vdd gnd cell_6t
Xbit_r196_c250 bl_250 br_250 wl_196 vdd gnd cell_6t
Xbit_r197_c250 bl_250 br_250 wl_197 vdd gnd cell_6t
Xbit_r198_c250 bl_250 br_250 wl_198 vdd gnd cell_6t
Xbit_r199_c250 bl_250 br_250 wl_199 vdd gnd cell_6t
Xbit_r200_c250 bl_250 br_250 wl_200 vdd gnd cell_6t
Xbit_r201_c250 bl_250 br_250 wl_201 vdd gnd cell_6t
Xbit_r202_c250 bl_250 br_250 wl_202 vdd gnd cell_6t
Xbit_r203_c250 bl_250 br_250 wl_203 vdd gnd cell_6t
Xbit_r204_c250 bl_250 br_250 wl_204 vdd gnd cell_6t
Xbit_r205_c250 bl_250 br_250 wl_205 vdd gnd cell_6t
Xbit_r206_c250 bl_250 br_250 wl_206 vdd gnd cell_6t
Xbit_r207_c250 bl_250 br_250 wl_207 vdd gnd cell_6t
Xbit_r208_c250 bl_250 br_250 wl_208 vdd gnd cell_6t
Xbit_r209_c250 bl_250 br_250 wl_209 vdd gnd cell_6t
Xbit_r210_c250 bl_250 br_250 wl_210 vdd gnd cell_6t
Xbit_r211_c250 bl_250 br_250 wl_211 vdd gnd cell_6t
Xbit_r212_c250 bl_250 br_250 wl_212 vdd gnd cell_6t
Xbit_r213_c250 bl_250 br_250 wl_213 vdd gnd cell_6t
Xbit_r214_c250 bl_250 br_250 wl_214 vdd gnd cell_6t
Xbit_r215_c250 bl_250 br_250 wl_215 vdd gnd cell_6t
Xbit_r216_c250 bl_250 br_250 wl_216 vdd gnd cell_6t
Xbit_r217_c250 bl_250 br_250 wl_217 vdd gnd cell_6t
Xbit_r218_c250 bl_250 br_250 wl_218 vdd gnd cell_6t
Xbit_r219_c250 bl_250 br_250 wl_219 vdd gnd cell_6t
Xbit_r220_c250 bl_250 br_250 wl_220 vdd gnd cell_6t
Xbit_r221_c250 bl_250 br_250 wl_221 vdd gnd cell_6t
Xbit_r222_c250 bl_250 br_250 wl_222 vdd gnd cell_6t
Xbit_r223_c250 bl_250 br_250 wl_223 vdd gnd cell_6t
Xbit_r224_c250 bl_250 br_250 wl_224 vdd gnd cell_6t
Xbit_r225_c250 bl_250 br_250 wl_225 vdd gnd cell_6t
Xbit_r226_c250 bl_250 br_250 wl_226 vdd gnd cell_6t
Xbit_r227_c250 bl_250 br_250 wl_227 vdd gnd cell_6t
Xbit_r228_c250 bl_250 br_250 wl_228 vdd gnd cell_6t
Xbit_r229_c250 bl_250 br_250 wl_229 vdd gnd cell_6t
Xbit_r230_c250 bl_250 br_250 wl_230 vdd gnd cell_6t
Xbit_r231_c250 bl_250 br_250 wl_231 vdd gnd cell_6t
Xbit_r232_c250 bl_250 br_250 wl_232 vdd gnd cell_6t
Xbit_r233_c250 bl_250 br_250 wl_233 vdd gnd cell_6t
Xbit_r234_c250 bl_250 br_250 wl_234 vdd gnd cell_6t
Xbit_r235_c250 bl_250 br_250 wl_235 vdd gnd cell_6t
Xbit_r236_c250 bl_250 br_250 wl_236 vdd gnd cell_6t
Xbit_r237_c250 bl_250 br_250 wl_237 vdd gnd cell_6t
Xbit_r238_c250 bl_250 br_250 wl_238 vdd gnd cell_6t
Xbit_r239_c250 bl_250 br_250 wl_239 vdd gnd cell_6t
Xbit_r240_c250 bl_250 br_250 wl_240 vdd gnd cell_6t
Xbit_r241_c250 bl_250 br_250 wl_241 vdd gnd cell_6t
Xbit_r242_c250 bl_250 br_250 wl_242 vdd gnd cell_6t
Xbit_r243_c250 bl_250 br_250 wl_243 vdd gnd cell_6t
Xbit_r244_c250 bl_250 br_250 wl_244 vdd gnd cell_6t
Xbit_r245_c250 bl_250 br_250 wl_245 vdd gnd cell_6t
Xbit_r246_c250 bl_250 br_250 wl_246 vdd gnd cell_6t
Xbit_r247_c250 bl_250 br_250 wl_247 vdd gnd cell_6t
Xbit_r248_c250 bl_250 br_250 wl_248 vdd gnd cell_6t
Xbit_r249_c250 bl_250 br_250 wl_249 vdd gnd cell_6t
Xbit_r250_c250 bl_250 br_250 wl_250 vdd gnd cell_6t
Xbit_r251_c250 bl_250 br_250 wl_251 vdd gnd cell_6t
Xbit_r252_c250 bl_250 br_250 wl_252 vdd gnd cell_6t
Xbit_r253_c250 bl_250 br_250 wl_253 vdd gnd cell_6t
Xbit_r254_c250 bl_250 br_250 wl_254 vdd gnd cell_6t
Xbit_r255_c250 bl_250 br_250 wl_255 vdd gnd cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd cell_6t
Xbit_r1_c251 bl_251 br_251 wl_1 vdd gnd cell_6t
Xbit_r2_c251 bl_251 br_251 wl_2 vdd gnd cell_6t
Xbit_r3_c251 bl_251 br_251 wl_3 vdd gnd cell_6t
Xbit_r4_c251 bl_251 br_251 wl_4 vdd gnd cell_6t
Xbit_r5_c251 bl_251 br_251 wl_5 vdd gnd cell_6t
Xbit_r6_c251 bl_251 br_251 wl_6 vdd gnd cell_6t
Xbit_r7_c251 bl_251 br_251 wl_7 vdd gnd cell_6t
Xbit_r8_c251 bl_251 br_251 wl_8 vdd gnd cell_6t
Xbit_r9_c251 bl_251 br_251 wl_9 vdd gnd cell_6t
Xbit_r10_c251 bl_251 br_251 wl_10 vdd gnd cell_6t
Xbit_r11_c251 bl_251 br_251 wl_11 vdd gnd cell_6t
Xbit_r12_c251 bl_251 br_251 wl_12 vdd gnd cell_6t
Xbit_r13_c251 bl_251 br_251 wl_13 vdd gnd cell_6t
Xbit_r14_c251 bl_251 br_251 wl_14 vdd gnd cell_6t
Xbit_r15_c251 bl_251 br_251 wl_15 vdd gnd cell_6t
Xbit_r16_c251 bl_251 br_251 wl_16 vdd gnd cell_6t
Xbit_r17_c251 bl_251 br_251 wl_17 vdd gnd cell_6t
Xbit_r18_c251 bl_251 br_251 wl_18 vdd gnd cell_6t
Xbit_r19_c251 bl_251 br_251 wl_19 vdd gnd cell_6t
Xbit_r20_c251 bl_251 br_251 wl_20 vdd gnd cell_6t
Xbit_r21_c251 bl_251 br_251 wl_21 vdd gnd cell_6t
Xbit_r22_c251 bl_251 br_251 wl_22 vdd gnd cell_6t
Xbit_r23_c251 bl_251 br_251 wl_23 vdd gnd cell_6t
Xbit_r24_c251 bl_251 br_251 wl_24 vdd gnd cell_6t
Xbit_r25_c251 bl_251 br_251 wl_25 vdd gnd cell_6t
Xbit_r26_c251 bl_251 br_251 wl_26 vdd gnd cell_6t
Xbit_r27_c251 bl_251 br_251 wl_27 vdd gnd cell_6t
Xbit_r28_c251 bl_251 br_251 wl_28 vdd gnd cell_6t
Xbit_r29_c251 bl_251 br_251 wl_29 vdd gnd cell_6t
Xbit_r30_c251 bl_251 br_251 wl_30 vdd gnd cell_6t
Xbit_r31_c251 bl_251 br_251 wl_31 vdd gnd cell_6t
Xbit_r32_c251 bl_251 br_251 wl_32 vdd gnd cell_6t
Xbit_r33_c251 bl_251 br_251 wl_33 vdd gnd cell_6t
Xbit_r34_c251 bl_251 br_251 wl_34 vdd gnd cell_6t
Xbit_r35_c251 bl_251 br_251 wl_35 vdd gnd cell_6t
Xbit_r36_c251 bl_251 br_251 wl_36 vdd gnd cell_6t
Xbit_r37_c251 bl_251 br_251 wl_37 vdd gnd cell_6t
Xbit_r38_c251 bl_251 br_251 wl_38 vdd gnd cell_6t
Xbit_r39_c251 bl_251 br_251 wl_39 vdd gnd cell_6t
Xbit_r40_c251 bl_251 br_251 wl_40 vdd gnd cell_6t
Xbit_r41_c251 bl_251 br_251 wl_41 vdd gnd cell_6t
Xbit_r42_c251 bl_251 br_251 wl_42 vdd gnd cell_6t
Xbit_r43_c251 bl_251 br_251 wl_43 vdd gnd cell_6t
Xbit_r44_c251 bl_251 br_251 wl_44 vdd gnd cell_6t
Xbit_r45_c251 bl_251 br_251 wl_45 vdd gnd cell_6t
Xbit_r46_c251 bl_251 br_251 wl_46 vdd gnd cell_6t
Xbit_r47_c251 bl_251 br_251 wl_47 vdd gnd cell_6t
Xbit_r48_c251 bl_251 br_251 wl_48 vdd gnd cell_6t
Xbit_r49_c251 bl_251 br_251 wl_49 vdd gnd cell_6t
Xbit_r50_c251 bl_251 br_251 wl_50 vdd gnd cell_6t
Xbit_r51_c251 bl_251 br_251 wl_51 vdd gnd cell_6t
Xbit_r52_c251 bl_251 br_251 wl_52 vdd gnd cell_6t
Xbit_r53_c251 bl_251 br_251 wl_53 vdd gnd cell_6t
Xbit_r54_c251 bl_251 br_251 wl_54 vdd gnd cell_6t
Xbit_r55_c251 bl_251 br_251 wl_55 vdd gnd cell_6t
Xbit_r56_c251 bl_251 br_251 wl_56 vdd gnd cell_6t
Xbit_r57_c251 bl_251 br_251 wl_57 vdd gnd cell_6t
Xbit_r58_c251 bl_251 br_251 wl_58 vdd gnd cell_6t
Xbit_r59_c251 bl_251 br_251 wl_59 vdd gnd cell_6t
Xbit_r60_c251 bl_251 br_251 wl_60 vdd gnd cell_6t
Xbit_r61_c251 bl_251 br_251 wl_61 vdd gnd cell_6t
Xbit_r62_c251 bl_251 br_251 wl_62 vdd gnd cell_6t
Xbit_r63_c251 bl_251 br_251 wl_63 vdd gnd cell_6t
Xbit_r64_c251 bl_251 br_251 wl_64 vdd gnd cell_6t
Xbit_r65_c251 bl_251 br_251 wl_65 vdd gnd cell_6t
Xbit_r66_c251 bl_251 br_251 wl_66 vdd gnd cell_6t
Xbit_r67_c251 bl_251 br_251 wl_67 vdd gnd cell_6t
Xbit_r68_c251 bl_251 br_251 wl_68 vdd gnd cell_6t
Xbit_r69_c251 bl_251 br_251 wl_69 vdd gnd cell_6t
Xbit_r70_c251 bl_251 br_251 wl_70 vdd gnd cell_6t
Xbit_r71_c251 bl_251 br_251 wl_71 vdd gnd cell_6t
Xbit_r72_c251 bl_251 br_251 wl_72 vdd gnd cell_6t
Xbit_r73_c251 bl_251 br_251 wl_73 vdd gnd cell_6t
Xbit_r74_c251 bl_251 br_251 wl_74 vdd gnd cell_6t
Xbit_r75_c251 bl_251 br_251 wl_75 vdd gnd cell_6t
Xbit_r76_c251 bl_251 br_251 wl_76 vdd gnd cell_6t
Xbit_r77_c251 bl_251 br_251 wl_77 vdd gnd cell_6t
Xbit_r78_c251 bl_251 br_251 wl_78 vdd gnd cell_6t
Xbit_r79_c251 bl_251 br_251 wl_79 vdd gnd cell_6t
Xbit_r80_c251 bl_251 br_251 wl_80 vdd gnd cell_6t
Xbit_r81_c251 bl_251 br_251 wl_81 vdd gnd cell_6t
Xbit_r82_c251 bl_251 br_251 wl_82 vdd gnd cell_6t
Xbit_r83_c251 bl_251 br_251 wl_83 vdd gnd cell_6t
Xbit_r84_c251 bl_251 br_251 wl_84 vdd gnd cell_6t
Xbit_r85_c251 bl_251 br_251 wl_85 vdd gnd cell_6t
Xbit_r86_c251 bl_251 br_251 wl_86 vdd gnd cell_6t
Xbit_r87_c251 bl_251 br_251 wl_87 vdd gnd cell_6t
Xbit_r88_c251 bl_251 br_251 wl_88 vdd gnd cell_6t
Xbit_r89_c251 bl_251 br_251 wl_89 vdd gnd cell_6t
Xbit_r90_c251 bl_251 br_251 wl_90 vdd gnd cell_6t
Xbit_r91_c251 bl_251 br_251 wl_91 vdd gnd cell_6t
Xbit_r92_c251 bl_251 br_251 wl_92 vdd gnd cell_6t
Xbit_r93_c251 bl_251 br_251 wl_93 vdd gnd cell_6t
Xbit_r94_c251 bl_251 br_251 wl_94 vdd gnd cell_6t
Xbit_r95_c251 bl_251 br_251 wl_95 vdd gnd cell_6t
Xbit_r96_c251 bl_251 br_251 wl_96 vdd gnd cell_6t
Xbit_r97_c251 bl_251 br_251 wl_97 vdd gnd cell_6t
Xbit_r98_c251 bl_251 br_251 wl_98 vdd gnd cell_6t
Xbit_r99_c251 bl_251 br_251 wl_99 vdd gnd cell_6t
Xbit_r100_c251 bl_251 br_251 wl_100 vdd gnd cell_6t
Xbit_r101_c251 bl_251 br_251 wl_101 vdd gnd cell_6t
Xbit_r102_c251 bl_251 br_251 wl_102 vdd gnd cell_6t
Xbit_r103_c251 bl_251 br_251 wl_103 vdd gnd cell_6t
Xbit_r104_c251 bl_251 br_251 wl_104 vdd gnd cell_6t
Xbit_r105_c251 bl_251 br_251 wl_105 vdd gnd cell_6t
Xbit_r106_c251 bl_251 br_251 wl_106 vdd gnd cell_6t
Xbit_r107_c251 bl_251 br_251 wl_107 vdd gnd cell_6t
Xbit_r108_c251 bl_251 br_251 wl_108 vdd gnd cell_6t
Xbit_r109_c251 bl_251 br_251 wl_109 vdd gnd cell_6t
Xbit_r110_c251 bl_251 br_251 wl_110 vdd gnd cell_6t
Xbit_r111_c251 bl_251 br_251 wl_111 vdd gnd cell_6t
Xbit_r112_c251 bl_251 br_251 wl_112 vdd gnd cell_6t
Xbit_r113_c251 bl_251 br_251 wl_113 vdd gnd cell_6t
Xbit_r114_c251 bl_251 br_251 wl_114 vdd gnd cell_6t
Xbit_r115_c251 bl_251 br_251 wl_115 vdd gnd cell_6t
Xbit_r116_c251 bl_251 br_251 wl_116 vdd gnd cell_6t
Xbit_r117_c251 bl_251 br_251 wl_117 vdd gnd cell_6t
Xbit_r118_c251 bl_251 br_251 wl_118 vdd gnd cell_6t
Xbit_r119_c251 bl_251 br_251 wl_119 vdd gnd cell_6t
Xbit_r120_c251 bl_251 br_251 wl_120 vdd gnd cell_6t
Xbit_r121_c251 bl_251 br_251 wl_121 vdd gnd cell_6t
Xbit_r122_c251 bl_251 br_251 wl_122 vdd gnd cell_6t
Xbit_r123_c251 bl_251 br_251 wl_123 vdd gnd cell_6t
Xbit_r124_c251 bl_251 br_251 wl_124 vdd gnd cell_6t
Xbit_r125_c251 bl_251 br_251 wl_125 vdd gnd cell_6t
Xbit_r126_c251 bl_251 br_251 wl_126 vdd gnd cell_6t
Xbit_r127_c251 bl_251 br_251 wl_127 vdd gnd cell_6t
Xbit_r128_c251 bl_251 br_251 wl_128 vdd gnd cell_6t
Xbit_r129_c251 bl_251 br_251 wl_129 vdd gnd cell_6t
Xbit_r130_c251 bl_251 br_251 wl_130 vdd gnd cell_6t
Xbit_r131_c251 bl_251 br_251 wl_131 vdd gnd cell_6t
Xbit_r132_c251 bl_251 br_251 wl_132 vdd gnd cell_6t
Xbit_r133_c251 bl_251 br_251 wl_133 vdd gnd cell_6t
Xbit_r134_c251 bl_251 br_251 wl_134 vdd gnd cell_6t
Xbit_r135_c251 bl_251 br_251 wl_135 vdd gnd cell_6t
Xbit_r136_c251 bl_251 br_251 wl_136 vdd gnd cell_6t
Xbit_r137_c251 bl_251 br_251 wl_137 vdd gnd cell_6t
Xbit_r138_c251 bl_251 br_251 wl_138 vdd gnd cell_6t
Xbit_r139_c251 bl_251 br_251 wl_139 vdd gnd cell_6t
Xbit_r140_c251 bl_251 br_251 wl_140 vdd gnd cell_6t
Xbit_r141_c251 bl_251 br_251 wl_141 vdd gnd cell_6t
Xbit_r142_c251 bl_251 br_251 wl_142 vdd gnd cell_6t
Xbit_r143_c251 bl_251 br_251 wl_143 vdd gnd cell_6t
Xbit_r144_c251 bl_251 br_251 wl_144 vdd gnd cell_6t
Xbit_r145_c251 bl_251 br_251 wl_145 vdd gnd cell_6t
Xbit_r146_c251 bl_251 br_251 wl_146 vdd gnd cell_6t
Xbit_r147_c251 bl_251 br_251 wl_147 vdd gnd cell_6t
Xbit_r148_c251 bl_251 br_251 wl_148 vdd gnd cell_6t
Xbit_r149_c251 bl_251 br_251 wl_149 vdd gnd cell_6t
Xbit_r150_c251 bl_251 br_251 wl_150 vdd gnd cell_6t
Xbit_r151_c251 bl_251 br_251 wl_151 vdd gnd cell_6t
Xbit_r152_c251 bl_251 br_251 wl_152 vdd gnd cell_6t
Xbit_r153_c251 bl_251 br_251 wl_153 vdd gnd cell_6t
Xbit_r154_c251 bl_251 br_251 wl_154 vdd gnd cell_6t
Xbit_r155_c251 bl_251 br_251 wl_155 vdd gnd cell_6t
Xbit_r156_c251 bl_251 br_251 wl_156 vdd gnd cell_6t
Xbit_r157_c251 bl_251 br_251 wl_157 vdd gnd cell_6t
Xbit_r158_c251 bl_251 br_251 wl_158 vdd gnd cell_6t
Xbit_r159_c251 bl_251 br_251 wl_159 vdd gnd cell_6t
Xbit_r160_c251 bl_251 br_251 wl_160 vdd gnd cell_6t
Xbit_r161_c251 bl_251 br_251 wl_161 vdd gnd cell_6t
Xbit_r162_c251 bl_251 br_251 wl_162 vdd gnd cell_6t
Xbit_r163_c251 bl_251 br_251 wl_163 vdd gnd cell_6t
Xbit_r164_c251 bl_251 br_251 wl_164 vdd gnd cell_6t
Xbit_r165_c251 bl_251 br_251 wl_165 vdd gnd cell_6t
Xbit_r166_c251 bl_251 br_251 wl_166 vdd gnd cell_6t
Xbit_r167_c251 bl_251 br_251 wl_167 vdd gnd cell_6t
Xbit_r168_c251 bl_251 br_251 wl_168 vdd gnd cell_6t
Xbit_r169_c251 bl_251 br_251 wl_169 vdd gnd cell_6t
Xbit_r170_c251 bl_251 br_251 wl_170 vdd gnd cell_6t
Xbit_r171_c251 bl_251 br_251 wl_171 vdd gnd cell_6t
Xbit_r172_c251 bl_251 br_251 wl_172 vdd gnd cell_6t
Xbit_r173_c251 bl_251 br_251 wl_173 vdd gnd cell_6t
Xbit_r174_c251 bl_251 br_251 wl_174 vdd gnd cell_6t
Xbit_r175_c251 bl_251 br_251 wl_175 vdd gnd cell_6t
Xbit_r176_c251 bl_251 br_251 wl_176 vdd gnd cell_6t
Xbit_r177_c251 bl_251 br_251 wl_177 vdd gnd cell_6t
Xbit_r178_c251 bl_251 br_251 wl_178 vdd gnd cell_6t
Xbit_r179_c251 bl_251 br_251 wl_179 vdd gnd cell_6t
Xbit_r180_c251 bl_251 br_251 wl_180 vdd gnd cell_6t
Xbit_r181_c251 bl_251 br_251 wl_181 vdd gnd cell_6t
Xbit_r182_c251 bl_251 br_251 wl_182 vdd gnd cell_6t
Xbit_r183_c251 bl_251 br_251 wl_183 vdd gnd cell_6t
Xbit_r184_c251 bl_251 br_251 wl_184 vdd gnd cell_6t
Xbit_r185_c251 bl_251 br_251 wl_185 vdd gnd cell_6t
Xbit_r186_c251 bl_251 br_251 wl_186 vdd gnd cell_6t
Xbit_r187_c251 bl_251 br_251 wl_187 vdd gnd cell_6t
Xbit_r188_c251 bl_251 br_251 wl_188 vdd gnd cell_6t
Xbit_r189_c251 bl_251 br_251 wl_189 vdd gnd cell_6t
Xbit_r190_c251 bl_251 br_251 wl_190 vdd gnd cell_6t
Xbit_r191_c251 bl_251 br_251 wl_191 vdd gnd cell_6t
Xbit_r192_c251 bl_251 br_251 wl_192 vdd gnd cell_6t
Xbit_r193_c251 bl_251 br_251 wl_193 vdd gnd cell_6t
Xbit_r194_c251 bl_251 br_251 wl_194 vdd gnd cell_6t
Xbit_r195_c251 bl_251 br_251 wl_195 vdd gnd cell_6t
Xbit_r196_c251 bl_251 br_251 wl_196 vdd gnd cell_6t
Xbit_r197_c251 bl_251 br_251 wl_197 vdd gnd cell_6t
Xbit_r198_c251 bl_251 br_251 wl_198 vdd gnd cell_6t
Xbit_r199_c251 bl_251 br_251 wl_199 vdd gnd cell_6t
Xbit_r200_c251 bl_251 br_251 wl_200 vdd gnd cell_6t
Xbit_r201_c251 bl_251 br_251 wl_201 vdd gnd cell_6t
Xbit_r202_c251 bl_251 br_251 wl_202 vdd gnd cell_6t
Xbit_r203_c251 bl_251 br_251 wl_203 vdd gnd cell_6t
Xbit_r204_c251 bl_251 br_251 wl_204 vdd gnd cell_6t
Xbit_r205_c251 bl_251 br_251 wl_205 vdd gnd cell_6t
Xbit_r206_c251 bl_251 br_251 wl_206 vdd gnd cell_6t
Xbit_r207_c251 bl_251 br_251 wl_207 vdd gnd cell_6t
Xbit_r208_c251 bl_251 br_251 wl_208 vdd gnd cell_6t
Xbit_r209_c251 bl_251 br_251 wl_209 vdd gnd cell_6t
Xbit_r210_c251 bl_251 br_251 wl_210 vdd gnd cell_6t
Xbit_r211_c251 bl_251 br_251 wl_211 vdd gnd cell_6t
Xbit_r212_c251 bl_251 br_251 wl_212 vdd gnd cell_6t
Xbit_r213_c251 bl_251 br_251 wl_213 vdd gnd cell_6t
Xbit_r214_c251 bl_251 br_251 wl_214 vdd gnd cell_6t
Xbit_r215_c251 bl_251 br_251 wl_215 vdd gnd cell_6t
Xbit_r216_c251 bl_251 br_251 wl_216 vdd gnd cell_6t
Xbit_r217_c251 bl_251 br_251 wl_217 vdd gnd cell_6t
Xbit_r218_c251 bl_251 br_251 wl_218 vdd gnd cell_6t
Xbit_r219_c251 bl_251 br_251 wl_219 vdd gnd cell_6t
Xbit_r220_c251 bl_251 br_251 wl_220 vdd gnd cell_6t
Xbit_r221_c251 bl_251 br_251 wl_221 vdd gnd cell_6t
Xbit_r222_c251 bl_251 br_251 wl_222 vdd gnd cell_6t
Xbit_r223_c251 bl_251 br_251 wl_223 vdd gnd cell_6t
Xbit_r224_c251 bl_251 br_251 wl_224 vdd gnd cell_6t
Xbit_r225_c251 bl_251 br_251 wl_225 vdd gnd cell_6t
Xbit_r226_c251 bl_251 br_251 wl_226 vdd gnd cell_6t
Xbit_r227_c251 bl_251 br_251 wl_227 vdd gnd cell_6t
Xbit_r228_c251 bl_251 br_251 wl_228 vdd gnd cell_6t
Xbit_r229_c251 bl_251 br_251 wl_229 vdd gnd cell_6t
Xbit_r230_c251 bl_251 br_251 wl_230 vdd gnd cell_6t
Xbit_r231_c251 bl_251 br_251 wl_231 vdd gnd cell_6t
Xbit_r232_c251 bl_251 br_251 wl_232 vdd gnd cell_6t
Xbit_r233_c251 bl_251 br_251 wl_233 vdd gnd cell_6t
Xbit_r234_c251 bl_251 br_251 wl_234 vdd gnd cell_6t
Xbit_r235_c251 bl_251 br_251 wl_235 vdd gnd cell_6t
Xbit_r236_c251 bl_251 br_251 wl_236 vdd gnd cell_6t
Xbit_r237_c251 bl_251 br_251 wl_237 vdd gnd cell_6t
Xbit_r238_c251 bl_251 br_251 wl_238 vdd gnd cell_6t
Xbit_r239_c251 bl_251 br_251 wl_239 vdd gnd cell_6t
Xbit_r240_c251 bl_251 br_251 wl_240 vdd gnd cell_6t
Xbit_r241_c251 bl_251 br_251 wl_241 vdd gnd cell_6t
Xbit_r242_c251 bl_251 br_251 wl_242 vdd gnd cell_6t
Xbit_r243_c251 bl_251 br_251 wl_243 vdd gnd cell_6t
Xbit_r244_c251 bl_251 br_251 wl_244 vdd gnd cell_6t
Xbit_r245_c251 bl_251 br_251 wl_245 vdd gnd cell_6t
Xbit_r246_c251 bl_251 br_251 wl_246 vdd gnd cell_6t
Xbit_r247_c251 bl_251 br_251 wl_247 vdd gnd cell_6t
Xbit_r248_c251 bl_251 br_251 wl_248 vdd gnd cell_6t
Xbit_r249_c251 bl_251 br_251 wl_249 vdd gnd cell_6t
Xbit_r250_c251 bl_251 br_251 wl_250 vdd gnd cell_6t
Xbit_r251_c251 bl_251 br_251 wl_251 vdd gnd cell_6t
Xbit_r252_c251 bl_251 br_251 wl_252 vdd gnd cell_6t
Xbit_r253_c251 bl_251 br_251 wl_253 vdd gnd cell_6t
Xbit_r254_c251 bl_251 br_251 wl_254 vdd gnd cell_6t
Xbit_r255_c251 bl_251 br_251 wl_255 vdd gnd cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd cell_6t
Xbit_r1_c252 bl_252 br_252 wl_1 vdd gnd cell_6t
Xbit_r2_c252 bl_252 br_252 wl_2 vdd gnd cell_6t
Xbit_r3_c252 bl_252 br_252 wl_3 vdd gnd cell_6t
Xbit_r4_c252 bl_252 br_252 wl_4 vdd gnd cell_6t
Xbit_r5_c252 bl_252 br_252 wl_5 vdd gnd cell_6t
Xbit_r6_c252 bl_252 br_252 wl_6 vdd gnd cell_6t
Xbit_r7_c252 bl_252 br_252 wl_7 vdd gnd cell_6t
Xbit_r8_c252 bl_252 br_252 wl_8 vdd gnd cell_6t
Xbit_r9_c252 bl_252 br_252 wl_9 vdd gnd cell_6t
Xbit_r10_c252 bl_252 br_252 wl_10 vdd gnd cell_6t
Xbit_r11_c252 bl_252 br_252 wl_11 vdd gnd cell_6t
Xbit_r12_c252 bl_252 br_252 wl_12 vdd gnd cell_6t
Xbit_r13_c252 bl_252 br_252 wl_13 vdd gnd cell_6t
Xbit_r14_c252 bl_252 br_252 wl_14 vdd gnd cell_6t
Xbit_r15_c252 bl_252 br_252 wl_15 vdd gnd cell_6t
Xbit_r16_c252 bl_252 br_252 wl_16 vdd gnd cell_6t
Xbit_r17_c252 bl_252 br_252 wl_17 vdd gnd cell_6t
Xbit_r18_c252 bl_252 br_252 wl_18 vdd gnd cell_6t
Xbit_r19_c252 bl_252 br_252 wl_19 vdd gnd cell_6t
Xbit_r20_c252 bl_252 br_252 wl_20 vdd gnd cell_6t
Xbit_r21_c252 bl_252 br_252 wl_21 vdd gnd cell_6t
Xbit_r22_c252 bl_252 br_252 wl_22 vdd gnd cell_6t
Xbit_r23_c252 bl_252 br_252 wl_23 vdd gnd cell_6t
Xbit_r24_c252 bl_252 br_252 wl_24 vdd gnd cell_6t
Xbit_r25_c252 bl_252 br_252 wl_25 vdd gnd cell_6t
Xbit_r26_c252 bl_252 br_252 wl_26 vdd gnd cell_6t
Xbit_r27_c252 bl_252 br_252 wl_27 vdd gnd cell_6t
Xbit_r28_c252 bl_252 br_252 wl_28 vdd gnd cell_6t
Xbit_r29_c252 bl_252 br_252 wl_29 vdd gnd cell_6t
Xbit_r30_c252 bl_252 br_252 wl_30 vdd gnd cell_6t
Xbit_r31_c252 bl_252 br_252 wl_31 vdd gnd cell_6t
Xbit_r32_c252 bl_252 br_252 wl_32 vdd gnd cell_6t
Xbit_r33_c252 bl_252 br_252 wl_33 vdd gnd cell_6t
Xbit_r34_c252 bl_252 br_252 wl_34 vdd gnd cell_6t
Xbit_r35_c252 bl_252 br_252 wl_35 vdd gnd cell_6t
Xbit_r36_c252 bl_252 br_252 wl_36 vdd gnd cell_6t
Xbit_r37_c252 bl_252 br_252 wl_37 vdd gnd cell_6t
Xbit_r38_c252 bl_252 br_252 wl_38 vdd gnd cell_6t
Xbit_r39_c252 bl_252 br_252 wl_39 vdd gnd cell_6t
Xbit_r40_c252 bl_252 br_252 wl_40 vdd gnd cell_6t
Xbit_r41_c252 bl_252 br_252 wl_41 vdd gnd cell_6t
Xbit_r42_c252 bl_252 br_252 wl_42 vdd gnd cell_6t
Xbit_r43_c252 bl_252 br_252 wl_43 vdd gnd cell_6t
Xbit_r44_c252 bl_252 br_252 wl_44 vdd gnd cell_6t
Xbit_r45_c252 bl_252 br_252 wl_45 vdd gnd cell_6t
Xbit_r46_c252 bl_252 br_252 wl_46 vdd gnd cell_6t
Xbit_r47_c252 bl_252 br_252 wl_47 vdd gnd cell_6t
Xbit_r48_c252 bl_252 br_252 wl_48 vdd gnd cell_6t
Xbit_r49_c252 bl_252 br_252 wl_49 vdd gnd cell_6t
Xbit_r50_c252 bl_252 br_252 wl_50 vdd gnd cell_6t
Xbit_r51_c252 bl_252 br_252 wl_51 vdd gnd cell_6t
Xbit_r52_c252 bl_252 br_252 wl_52 vdd gnd cell_6t
Xbit_r53_c252 bl_252 br_252 wl_53 vdd gnd cell_6t
Xbit_r54_c252 bl_252 br_252 wl_54 vdd gnd cell_6t
Xbit_r55_c252 bl_252 br_252 wl_55 vdd gnd cell_6t
Xbit_r56_c252 bl_252 br_252 wl_56 vdd gnd cell_6t
Xbit_r57_c252 bl_252 br_252 wl_57 vdd gnd cell_6t
Xbit_r58_c252 bl_252 br_252 wl_58 vdd gnd cell_6t
Xbit_r59_c252 bl_252 br_252 wl_59 vdd gnd cell_6t
Xbit_r60_c252 bl_252 br_252 wl_60 vdd gnd cell_6t
Xbit_r61_c252 bl_252 br_252 wl_61 vdd gnd cell_6t
Xbit_r62_c252 bl_252 br_252 wl_62 vdd gnd cell_6t
Xbit_r63_c252 bl_252 br_252 wl_63 vdd gnd cell_6t
Xbit_r64_c252 bl_252 br_252 wl_64 vdd gnd cell_6t
Xbit_r65_c252 bl_252 br_252 wl_65 vdd gnd cell_6t
Xbit_r66_c252 bl_252 br_252 wl_66 vdd gnd cell_6t
Xbit_r67_c252 bl_252 br_252 wl_67 vdd gnd cell_6t
Xbit_r68_c252 bl_252 br_252 wl_68 vdd gnd cell_6t
Xbit_r69_c252 bl_252 br_252 wl_69 vdd gnd cell_6t
Xbit_r70_c252 bl_252 br_252 wl_70 vdd gnd cell_6t
Xbit_r71_c252 bl_252 br_252 wl_71 vdd gnd cell_6t
Xbit_r72_c252 bl_252 br_252 wl_72 vdd gnd cell_6t
Xbit_r73_c252 bl_252 br_252 wl_73 vdd gnd cell_6t
Xbit_r74_c252 bl_252 br_252 wl_74 vdd gnd cell_6t
Xbit_r75_c252 bl_252 br_252 wl_75 vdd gnd cell_6t
Xbit_r76_c252 bl_252 br_252 wl_76 vdd gnd cell_6t
Xbit_r77_c252 bl_252 br_252 wl_77 vdd gnd cell_6t
Xbit_r78_c252 bl_252 br_252 wl_78 vdd gnd cell_6t
Xbit_r79_c252 bl_252 br_252 wl_79 vdd gnd cell_6t
Xbit_r80_c252 bl_252 br_252 wl_80 vdd gnd cell_6t
Xbit_r81_c252 bl_252 br_252 wl_81 vdd gnd cell_6t
Xbit_r82_c252 bl_252 br_252 wl_82 vdd gnd cell_6t
Xbit_r83_c252 bl_252 br_252 wl_83 vdd gnd cell_6t
Xbit_r84_c252 bl_252 br_252 wl_84 vdd gnd cell_6t
Xbit_r85_c252 bl_252 br_252 wl_85 vdd gnd cell_6t
Xbit_r86_c252 bl_252 br_252 wl_86 vdd gnd cell_6t
Xbit_r87_c252 bl_252 br_252 wl_87 vdd gnd cell_6t
Xbit_r88_c252 bl_252 br_252 wl_88 vdd gnd cell_6t
Xbit_r89_c252 bl_252 br_252 wl_89 vdd gnd cell_6t
Xbit_r90_c252 bl_252 br_252 wl_90 vdd gnd cell_6t
Xbit_r91_c252 bl_252 br_252 wl_91 vdd gnd cell_6t
Xbit_r92_c252 bl_252 br_252 wl_92 vdd gnd cell_6t
Xbit_r93_c252 bl_252 br_252 wl_93 vdd gnd cell_6t
Xbit_r94_c252 bl_252 br_252 wl_94 vdd gnd cell_6t
Xbit_r95_c252 bl_252 br_252 wl_95 vdd gnd cell_6t
Xbit_r96_c252 bl_252 br_252 wl_96 vdd gnd cell_6t
Xbit_r97_c252 bl_252 br_252 wl_97 vdd gnd cell_6t
Xbit_r98_c252 bl_252 br_252 wl_98 vdd gnd cell_6t
Xbit_r99_c252 bl_252 br_252 wl_99 vdd gnd cell_6t
Xbit_r100_c252 bl_252 br_252 wl_100 vdd gnd cell_6t
Xbit_r101_c252 bl_252 br_252 wl_101 vdd gnd cell_6t
Xbit_r102_c252 bl_252 br_252 wl_102 vdd gnd cell_6t
Xbit_r103_c252 bl_252 br_252 wl_103 vdd gnd cell_6t
Xbit_r104_c252 bl_252 br_252 wl_104 vdd gnd cell_6t
Xbit_r105_c252 bl_252 br_252 wl_105 vdd gnd cell_6t
Xbit_r106_c252 bl_252 br_252 wl_106 vdd gnd cell_6t
Xbit_r107_c252 bl_252 br_252 wl_107 vdd gnd cell_6t
Xbit_r108_c252 bl_252 br_252 wl_108 vdd gnd cell_6t
Xbit_r109_c252 bl_252 br_252 wl_109 vdd gnd cell_6t
Xbit_r110_c252 bl_252 br_252 wl_110 vdd gnd cell_6t
Xbit_r111_c252 bl_252 br_252 wl_111 vdd gnd cell_6t
Xbit_r112_c252 bl_252 br_252 wl_112 vdd gnd cell_6t
Xbit_r113_c252 bl_252 br_252 wl_113 vdd gnd cell_6t
Xbit_r114_c252 bl_252 br_252 wl_114 vdd gnd cell_6t
Xbit_r115_c252 bl_252 br_252 wl_115 vdd gnd cell_6t
Xbit_r116_c252 bl_252 br_252 wl_116 vdd gnd cell_6t
Xbit_r117_c252 bl_252 br_252 wl_117 vdd gnd cell_6t
Xbit_r118_c252 bl_252 br_252 wl_118 vdd gnd cell_6t
Xbit_r119_c252 bl_252 br_252 wl_119 vdd gnd cell_6t
Xbit_r120_c252 bl_252 br_252 wl_120 vdd gnd cell_6t
Xbit_r121_c252 bl_252 br_252 wl_121 vdd gnd cell_6t
Xbit_r122_c252 bl_252 br_252 wl_122 vdd gnd cell_6t
Xbit_r123_c252 bl_252 br_252 wl_123 vdd gnd cell_6t
Xbit_r124_c252 bl_252 br_252 wl_124 vdd gnd cell_6t
Xbit_r125_c252 bl_252 br_252 wl_125 vdd gnd cell_6t
Xbit_r126_c252 bl_252 br_252 wl_126 vdd gnd cell_6t
Xbit_r127_c252 bl_252 br_252 wl_127 vdd gnd cell_6t
Xbit_r128_c252 bl_252 br_252 wl_128 vdd gnd cell_6t
Xbit_r129_c252 bl_252 br_252 wl_129 vdd gnd cell_6t
Xbit_r130_c252 bl_252 br_252 wl_130 vdd gnd cell_6t
Xbit_r131_c252 bl_252 br_252 wl_131 vdd gnd cell_6t
Xbit_r132_c252 bl_252 br_252 wl_132 vdd gnd cell_6t
Xbit_r133_c252 bl_252 br_252 wl_133 vdd gnd cell_6t
Xbit_r134_c252 bl_252 br_252 wl_134 vdd gnd cell_6t
Xbit_r135_c252 bl_252 br_252 wl_135 vdd gnd cell_6t
Xbit_r136_c252 bl_252 br_252 wl_136 vdd gnd cell_6t
Xbit_r137_c252 bl_252 br_252 wl_137 vdd gnd cell_6t
Xbit_r138_c252 bl_252 br_252 wl_138 vdd gnd cell_6t
Xbit_r139_c252 bl_252 br_252 wl_139 vdd gnd cell_6t
Xbit_r140_c252 bl_252 br_252 wl_140 vdd gnd cell_6t
Xbit_r141_c252 bl_252 br_252 wl_141 vdd gnd cell_6t
Xbit_r142_c252 bl_252 br_252 wl_142 vdd gnd cell_6t
Xbit_r143_c252 bl_252 br_252 wl_143 vdd gnd cell_6t
Xbit_r144_c252 bl_252 br_252 wl_144 vdd gnd cell_6t
Xbit_r145_c252 bl_252 br_252 wl_145 vdd gnd cell_6t
Xbit_r146_c252 bl_252 br_252 wl_146 vdd gnd cell_6t
Xbit_r147_c252 bl_252 br_252 wl_147 vdd gnd cell_6t
Xbit_r148_c252 bl_252 br_252 wl_148 vdd gnd cell_6t
Xbit_r149_c252 bl_252 br_252 wl_149 vdd gnd cell_6t
Xbit_r150_c252 bl_252 br_252 wl_150 vdd gnd cell_6t
Xbit_r151_c252 bl_252 br_252 wl_151 vdd gnd cell_6t
Xbit_r152_c252 bl_252 br_252 wl_152 vdd gnd cell_6t
Xbit_r153_c252 bl_252 br_252 wl_153 vdd gnd cell_6t
Xbit_r154_c252 bl_252 br_252 wl_154 vdd gnd cell_6t
Xbit_r155_c252 bl_252 br_252 wl_155 vdd gnd cell_6t
Xbit_r156_c252 bl_252 br_252 wl_156 vdd gnd cell_6t
Xbit_r157_c252 bl_252 br_252 wl_157 vdd gnd cell_6t
Xbit_r158_c252 bl_252 br_252 wl_158 vdd gnd cell_6t
Xbit_r159_c252 bl_252 br_252 wl_159 vdd gnd cell_6t
Xbit_r160_c252 bl_252 br_252 wl_160 vdd gnd cell_6t
Xbit_r161_c252 bl_252 br_252 wl_161 vdd gnd cell_6t
Xbit_r162_c252 bl_252 br_252 wl_162 vdd gnd cell_6t
Xbit_r163_c252 bl_252 br_252 wl_163 vdd gnd cell_6t
Xbit_r164_c252 bl_252 br_252 wl_164 vdd gnd cell_6t
Xbit_r165_c252 bl_252 br_252 wl_165 vdd gnd cell_6t
Xbit_r166_c252 bl_252 br_252 wl_166 vdd gnd cell_6t
Xbit_r167_c252 bl_252 br_252 wl_167 vdd gnd cell_6t
Xbit_r168_c252 bl_252 br_252 wl_168 vdd gnd cell_6t
Xbit_r169_c252 bl_252 br_252 wl_169 vdd gnd cell_6t
Xbit_r170_c252 bl_252 br_252 wl_170 vdd gnd cell_6t
Xbit_r171_c252 bl_252 br_252 wl_171 vdd gnd cell_6t
Xbit_r172_c252 bl_252 br_252 wl_172 vdd gnd cell_6t
Xbit_r173_c252 bl_252 br_252 wl_173 vdd gnd cell_6t
Xbit_r174_c252 bl_252 br_252 wl_174 vdd gnd cell_6t
Xbit_r175_c252 bl_252 br_252 wl_175 vdd gnd cell_6t
Xbit_r176_c252 bl_252 br_252 wl_176 vdd gnd cell_6t
Xbit_r177_c252 bl_252 br_252 wl_177 vdd gnd cell_6t
Xbit_r178_c252 bl_252 br_252 wl_178 vdd gnd cell_6t
Xbit_r179_c252 bl_252 br_252 wl_179 vdd gnd cell_6t
Xbit_r180_c252 bl_252 br_252 wl_180 vdd gnd cell_6t
Xbit_r181_c252 bl_252 br_252 wl_181 vdd gnd cell_6t
Xbit_r182_c252 bl_252 br_252 wl_182 vdd gnd cell_6t
Xbit_r183_c252 bl_252 br_252 wl_183 vdd gnd cell_6t
Xbit_r184_c252 bl_252 br_252 wl_184 vdd gnd cell_6t
Xbit_r185_c252 bl_252 br_252 wl_185 vdd gnd cell_6t
Xbit_r186_c252 bl_252 br_252 wl_186 vdd gnd cell_6t
Xbit_r187_c252 bl_252 br_252 wl_187 vdd gnd cell_6t
Xbit_r188_c252 bl_252 br_252 wl_188 vdd gnd cell_6t
Xbit_r189_c252 bl_252 br_252 wl_189 vdd gnd cell_6t
Xbit_r190_c252 bl_252 br_252 wl_190 vdd gnd cell_6t
Xbit_r191_c252 bl_252 br_252 wl_191 vdd gnd cell_6t
Xbit_r192_c252 bl_252 br_252 wl_192 vdd gnd cell_6t
Xbit_r193_c252 bl_252 br_252 wl_193 vdd gnd cell_6t
Xbit_r194_c252 bl_252 br_252 wl_194 vdd gnd cell_6t
Xbit_r195_c252 bl_252 br_252 wl_195 vdd gnd cell_6t
Xbit_r196_c252 bl_252 br_252 wl_196 vdd gnd cell_6t
Xbit_r197_c252 bl_252 br_252 wl_197 vdd gnd cell_6t
Xbit_r198_c252 bl_252 br_252 wl_198 vdd gnd cell_6t
Xbit_r199_c252 bl_252 br_252 wl_199 vdd gnd cell_6t
Xbit_r200_c252 bl_252 br_252 wl_200 vdd gnd cell_6t
Xbit_r201_c252 bl_252 br_252 wl_201 vdd gnd cell_6t
Xbit_r202_c252 bl_252 br_252 wl_202 vdd gnd cell_6t
Xbit_r203_c252 bl_252 br_252 wl_203 vdd gnd cell_6t
Xbit_r204_c252 bl_252 br_252 wl_204 vdd gnd cell_6t
Xbit_r205_c252 bl_252 br_252 wl_205 vdd gnd cell_6t
Xbit_r206_c252 bl_252 br_252 wl_206 vdd gnd cell_6t
Xbit_r207_c252 bl_252 br_252 wl_207 vdd gnd cell_6t
Xbit_r208_c252 bl_252 br_252 wl_208 vdd gnd cell_6t
Xbit_r209_c252 bl_252 br_252 wl_209 vdd gnd cell_6t
Xbit_r210_c252 bl_252 br_252 wl_210 vdd gnd cell_6t
Xbit_r211_c252 bl_252 br_252 wl_211 vdd gnd cell_6t
Xbit_r212_c252 bl_252 br_252 wl_212 vdd gnd cell_6t
Xbit_r213_c252 bl_252 br_252 wl_213 vdd gnd cell_6t
Xbit_r214_c252 bl_252 br_252 wl_214 vdd gnd cell_6t
Xbit_r215_c252 bl_252 br_252 wl_215 vdd gnd cell_6t
Xbit_r216_c252 bl_252 br_252 wl_216 vdd gnd cell_6t
Xbit_r217_c252 bl_252 br_252 wl_217 vdd gnd cell_6t
Xbit_r218_c252 bl_252 br_252 wl_218 vdd gnd cell_6t
Xbit_r219_c252 bl_252 br_252 wl_219 vdd gnd cell_6t
Xbit_r220_c252 bl_252 br_252 wl_220 vdd gnd cell_6t
Xbit_r221_c252 bl_252 br_252 wl_221 vdd gnd cell_6t
Xbit_r222_c252 bl_252 br_252 wl_222 vdd gnd cell_6t
Xbit_r223_c252 bl_252 br_252 wl_223 vdd gnd cell_6t
Xbit_r224_c252 bl_252 br_252 wl_224 vdd gnd cell_6t
Xbit_r225_c252 bl_252 br_252 wl_225 vdd gnd cell_6t
Xbit_r226_c252 bl_252 br_252 wl_226 vdd gnd cell_6t
Xbit_r227_c252 bl_252 br_252 wl_227 vdd gnd cell_6t
Xbit_r228_c252 bl_252 br_252 wl_228 vdd gnd cell_6t
Xbit_r229_c252 bl_252 br_252 wl_229 vdd gnd cell_6t
Xbit_r230_c252 bl_252 br_252 wl_230 vdd gnd cell_6t
Xbit_r231_c252 bl_252 br_252 wl_231 vdd gnd cell_6t
Xbit_r232_c252 bl_252 br_252 wl_232 vdd gnd cell_6t
Xbit_r233_c252 bl_252 br_252 wl_233 vdd gnd cell_6t
Xbit_r234_c252 bl_252 br_252 wl_234 vdd gnd cell_6t
Xbit_r235_c252 bl_252 br_252 wl_235 vdd gnd cell_6t
Xbit_r236_c252 bl_252 br_252 wl_236 vdd gnd cell_6t
Xbit_r237_c252 bl_252 br_252 wl_237 vdd gnd cell_6t
Xbit_r238_c252 bl_252 br_252 wl_238 vdd gnd cell_6t
Xbit_r239_c252 bl_252 br_252 wl_239 vdd gnd cell_6t
Xbit_r240_c252 bl_252 br_252 wl_240 vdd gnd cell_6t
Xbit_r241_c252 bl_252 br_252 wl_241 vdd gnd cell_6t
Xbit_r242_c252 bl_252 br_252 wl_242 vdd gnd cell_6t
Xbit_r243_c252 bl_252 br_252 wl_243 vdd gnd cell_6t
Xbit_r244_c252 bl_252 br_252 wl_244 vdd gnd cell_6t
Xbit_r245_c252 bl_252 br_252 wl_245 vdd gnd cell_6t
Xbit_r246_c252 bl_252 br_252 wl_246 vdd gnd cell_6t
Xbit_r247_c252 bl_252 br_252 wl_247 vdd gnd cell_6t
Xbit_r248_c252 bl_252 br_252 wl_248 vdd gnd cell_6t
Xbit_r249_c252 bl_252 br_252 wl_249 vdd gnd cell_6t
Xbit_r250_c252 bl_252 br_252 wl_250 vdd gnd cell_6t
Xbit_r251_c252 bl_252 br_252 wl_251 vdd gnd cell_6t
Xbit_r252_c252 bl_252 br_252 wl_252 vdd gnd cell_6t
Xbit_r253_c252 bl_252 br_252 wl_253 vdd gnd cell_6t
Xbit_r254_c252 bl_252 br_252 wl_254 vdd gnd cell_6t
Xbit_r255_c252 bl_252 br_252 wl_255 vdd gnd cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd cell_6t
Xbit_r1_c253 bl_253 br_253 wl_1 vdd gnd cell_6t
Xbit_r2_c253 bl_253 br_253 wl_2 vdd gnd cell_6t
Xbit_r3_c253 bl_253 br_253 wl_3 vdd gnd cell_6t
Xbit_r4_c253 bl_253 br_253 wl_4 vdd gnd cell_6t
Xbit_r5_c253 bl_253 br_253 wl_5 vdd gnd cell_6t
Xbit_r6_c253 bl_253 br_253 wl_6 vdd gnd cell_6t
Xbit_r7_c253 bl_253 br_253 wl_7 vdd gnd cell_6t
Xbit_r8_c253 bl_253 br_253 wl_8 vdd gnd cell_6t
Xbit_r9_c253 bl_253 br_253 wl_9 vdd gnd cell_6t
Xbit_r10_c253 bl_253 br_253 wl_10 vdd gnd cell_6t
Xbit_r11_c253 bl_253 br_253 wl_11 vdd gnd cell_6t
Xbit_r12_c253 bl_253 br_253 wl_12 vdd gnd cell_6t
Xbit_r13_c253 bl_253 br_253 wl_13 vdd gnd cell_6t
Xbit_r14_c253 bl_253 br_253 wl_14 vdd gnd cell_6t
Xbit_r15_c253 bl_253 br_253 wl_15 vdd gnd cell_6t
Xbit_r16_c253 bl_253 br_253 wl_16 vdd gnd cell_6t
Xbit_r17_c253 bl_253 br_253 wl_17 vdd gnd cell_6t
Xbit_r18_c253 bl_253 br_253 wl_18 vdd gnd cell_6t
Xbit_r19_c253 bl_253 br_253 wl_19 vdd gnd cell_6t
Xbit_r20_c253 bl_253 br_253 wl_20 vdd gnd cell_6t
Xbit_r21_c253 bl_253 br_253 wl_21 vdd gnd cell_6t
Xbit_r22_c253 bl_253 br_253 wl_22 vdd gnd cell_6t
Xbit_r23_c253 bl_253 br_253 wl_23 vdd gnd cell_6t
Xbit_r24_c253 bl_253 br_253 wl_24 vdd gnd cell_6t
Xbit_r25_c253 bl_253 br_253 wl_25 vdd gnd cell_6t
Xbit_r26_c253 bl_253 br_253 wl_26 vdd gnd cell_6t
Xbit_r27_c253 bl_253 br_253 wl_27 vdd gnd cell_6t
Xbit_r28_c253 bl_253 br_253 wl_28 vdd gnd cell_6t
Xbit_r29_c253 bl_253 br_253 wl_29 vdd gnd cell_6t
Xbit_r30_c253 bl_253 br_253 wl_30 vdd gnd cell_6t
Xbit_r31_c253 bl_253 br_253 wl_31 vdd gnd cell_6t
Xbit_r32_c253 bl_253 br_253 wl_32 vdd gnd cell_6t
Xbit_r33_c253 bl_253 br_253 wl_33 vdd gnd cell_6t
Xbit_r34_c253 bl_253 br_253 wl_34 vdd gnd cell_6t
Xbit_r35_c253 bl_253 br_253 wl_35 vdd gnd cell_6t
Xbit_r36_c253 bl_253 br_253 wl_36 vdd gnd cell_6t
Xbit_r37_c253 bl_253 br_253 wl_37 vdd gnd cell_6t
Xbit_r38_c253 bl_253 br_253 wl_38 vdd gnd cell_6t
Xbit_r39_c253 bl_253 br_253 wl_39 vdd gnd cell_6t
Xbit_r40_c253 bl_253 br_253 wl_40 vdd gnd cell_6t
Xbit_r41_c253 bl_253 br_253 wl_41 vdd gnd cell_6t
Xbit_r42_c253 bl_253 br_253 wl_42 vdd gnd cell_6t
Xbit_r43_c253 bl_253 br_253 wl_43 vdd gnd cell_6t
Xbit_r44_c253 bl_253 br_253 wl_44 vdd gnd cell_6t
Xbit_r45_c253 bl_253 br_253 wl_45 vdd gnd cell_6t
Xbit_r46_c253 bl_253 br_253 wl_46 vdd gnd cell_6t
Xbit_r47_c253 bl_253 br_253 wl_47 vdd gnd cell_6t
Xbit_r48_c253 bl_253 br_253 wl_48 vdd gnd cell_6t
Xbit_r49_c253 bl_253 br_253 wl_49 vdd gnd cell_6t
Xbit_r50_c253 bl_253 br_253 wl_50 vdd gnd cell_6t
Xbit_r51_c253 bl_253 br_253 wl_51 vdd gnd cell_6t
Xbit_r52_c253 bl_253 br_253 wl_52 vdd gnd cell_6t
Xbit_r53_c253 bl_253 br_253 wl_53 vdd gnd cell_6t
Xbit_r54_c253 bl_253 br_253 wl_54 vdd gnd cell_6t
Xbit_r55_c253 bl_253 br_253 wl_55 vdd gnd cell_6t
Xbit_r56_c253 bl_253 br_253 wl_56 vdd gnd cell_6t
Xbit_r57_c253 bl_253 br_253 wl_57 vdd gnd cell_6t
Xbit_r58_c253 bl_253 br_253 wl_58 vdd gnd cell_6t
Xbit_r59_c253 bl_253 br_253 wl_59 vdd gnd cell_6t
Xbit_r60_c253 bl_253 br_253 wl_60 vdd gnd cell_6t
Xbit_r61_c253 bl_253 br_253 wl_61 vdd gnd cell_6t
Xbit_r62_c253 bl_253 br_253 wl_62 vdd gnd cell_6t
Xbit_r63_c253 bl_253 br_253 wl_63 vdd gnd cell_6t
Xbit_r64_c253 bl_253 br_253 wl_64 vdd gnd cell_6t
Xbit_r65_c253 bl_253 br_253 wl_65 vdd gnd cell_6t
Xbit_r66_c253 bl_253 br_253 wl_66 vdd gnd cell_6t
Xbit_r67_c253 bl_253 br_253 wl_67 vdd gnd cell_6t
Xbit_r68_c253 bl_253 br_253 wl_68 vdd gnd cell_6t
Xbit_r69_c253 bl_253 br_253 wl_69 vdd gnd cell_6t
Xbit_r70_c253 bl_253 br_253 wl_70 vdd gnd cell_6t
Xbit_r71_c253 bl_253 br_253 wl_71 vdd gnd cell_6t
Xbit_r72_c253 bl_253 br_253 wl_72 vdd gnd cell_6t
Xbit_r73_c253 bl_253 br_253 wl_73 vdd gnd cell_6t
Xbit_r74_c253 bl_253 br_253 wl_74 vdd gnd cell_6t
Xbit_r75_c253 bl_253 br_253 wl_75 vdd gnd cell_6t
Xbit_r76_c253 bl_253 br_253 wl_76 vdd gnd cell_6t
Xbit_r77_c253 bl_253 br_253 wl_77 vdd gnd cell_6t
Xbit_r78_c253 bl_253 br_253 wl_78 vdd gnd cell_6t
Xbit_r79_c253 bl_253 br_253 wl_79 vdd gnd cell_6t
Xbit_r80_c253 bl_253 br_253 wl_80 vdd gnd cell_6t
Xbit_r81_c253 bl_253 br_253 wl_81 vdd gnd cell_6t
Xbit_r82_c253 bl_253 br_253 wl_82 vdd gnd cell_6t
Xbit_r83_c253 bl_253 br_253 wl_83 vdd gnd cell_6t
Xbit_r84_c253 bl_253 br_253 wl_84 vdd gnd cell_6t
Xbit_r85_c253 bl_253 br_253 wl_85 vdd gnd cell_6t
Xbit_r86_c253 bl_253 br_253 wl_86 vdd gnd cell_6t
Xbit_r87_c253 bl_253 br_253 wl_87 vdd gnd cell_6t
Xbit_r88_c253 bl_253 br_253 wl_88 vdd gnd cell_6t
Xbit_r89_c253 bl_253 br_253 wl_89 vdd gnd cell_6t
Xbit_r90_c253 bl_253 br_253 wl_90 vdd gnd cell_6t
Xbit_r91_c253 bl_253 br_253 wl_91 vdd gnd cell_6t
Xbit_r92_c253 bl_253 br_253 wl_92 vdd gnd cell_6t
Xbit_r93_c253 bl_253 br_253 wl_93 vdd gnd cell_6t
Xbit_r94_c253 bl_253 br_253 wl_94 vdd gnd cell_6t
Xbit_r95_c253 bl_253 br_253 wl_95 vdd gnd cell_6t
Xbit_r96_c253 bl_253 br_253 wl_96 vdd gnd cell_6t
Xbit_r97_c253 bl_253 br_253 wl_97 vdd gnd cell_6t
Xbit_r98_c253 bl_253 br_253 wl_98 vdd gnd cell_6t
Xbit_r99_c253 bl_253 br_253 wl_99 vdd gnd cell_6t
Xbit_r100_c253 bl_253 br_253 wl_100 vdd gnd cell_6t
Xbit_r101_c253 bl_253 br_253 wl_101 vdd gnd cell_6t
Xbit_r102_c253 bl_253 br_253 wl_102 vdd gnd cell_6t
Xbit_r103_c253 bl_253 br_253 wl_103 vdd gnd cell_6t
Xbit_r104_c253 bl_253 br_253 wl_104 vdd gnd cell_6t
Xbit_r105_c253 bl_253 br_253 wl_105 vdd gnd cell_6t
Xbit_r106_c253 bl_253 br_253 wl_106 vdd gnd cell_6t
Xbit_r107_c253 bl_253 br_253 wl_107 vdd gnd cell_6t
Xbit_r108_c253 bl_253 br_253 wl_108 vdd gnd cell_6t
Xbit_r109_c253 bl_253 br_253 wl_109 vdd gnd cell_6t
Xbit_r110_c253 bl_253 br_253 wl_110 vdd gnd cell_6t
Xbit_r111_c253 bl_253 br_253 wl_111 vdd gnd cell_6t
Xbit_r112_c253 bl_253 br_253 wl_112 vdd gnd cell_6t
Xbit_r113_c253 bl_253 br_253 wl_113 vdd gnd cell_6t
Xbit_r114_c253 bl_253 br_253 wl_114 vdd gnd cell_6t
Xbit_r115_c253 bl_253 br_253 wl_115 vdd gnd cell_6t
Xbit_r116_c253 bl_253 br_253 wl_116 vdd gnd cell_6t
Xbit_r117_c253 bl_253 br_253 wl_117 vdd gnd cell_6t
Xbit_r118_c253 bl_253 br_253 wl_118 vdd gnd cell_6t
Xbit_r119_c253 bl_253 br_253 wl_119 vdd gnd cell_6t
Xbit_r120_c253 bl_253 br_253 wl_120 vdd gnd cell_6t
Xbit_r121_c253 bl_253 br_253 wl_121 vdd gnd cell_6t
Xbit_r122_c253 bl_253 br_253 wl_122 vdd gnd cell_6t
Xbit_r123_c253 bl_253 br_253 wl_123 vdd gnd cell_6t
Xbit_r124_c253 bl_253 br_253 wl_124 vdd gnd cell_6t
Xbit_r125_c253 bl_253 br_253 wl_125 vdd gnd cell_6t
Xbit_r126_c253 bl_253 br_253 wl_126 vdd gnd cell_6t
Xbit_r127_c253 bl_253 br_253 wl_127 vdd gnd cell_6t
Xbit_r128_c253 bl_253 br_253 wl_128 vdd gnd cell_6t
Xbit_r129_c253 bl_253 br_253 wl_129 vdd gnd cell_6t
Xbit_r130_c253 bl_253 br_253 wl_130 vdd gnd cell_6t
Xbit_r131_c253 bl_253 br_253 wl_131 vdd gnd cell_6t
Xbit_r132_c253 bl_253 br_253 wl_132 vdd gnd cell_6t
Xbit_r133_c253 bl_253 br_253 wl_133 vdd gnd cell_6t
Xbit_r134_c253 bl_253 br_253 wl_134 vdd gnd cell_6t
Xbit_r135_c253 bl_253 br_253 wl_135 vdd gnd cell_6t
Xbit_r136_c253 bl_253 br_253 wl_136 vdd gnd cell_6t
Xbit_r137_c253 bl_253 br_253 wl_137 vdd gnd cell_6t
Xbit_r138_c253 bl_253 br_253 wl_138 vdd gnd cell_6t
Xbit_r139_c253 bl_253 br_253 wl_139 vdd gnd cell_6t
Xbit_r140_c253 bl_253 br_253 wl_140 vdd gnd cell_6t
Xbit_r141_c253 bl_253 br_253 wl_141 vdd gnd cell_6t
Xbit_r142_c253 bl_253 br_253 wl_142 vdd gnd cell_6t
Xbit_r143_c253 bl_253 br_253 wl_143 vdd gnd cell_6t
Xbit_r144_c253 bl_253 br_253 wl_144 vdd gnd cell_6t
Xbit_r145_c253 bl_253 br_253 wl_145 vdd gnd cell_6t
Xbit_r146_c253 bl_253 br_253 wl_146 vdd gnd cell_6t
Xbit_r147_c253 bl_253 br_253 wl_147 vdd gnd cell_6t
Xbit_r148_c253 bl_253 br_253 wl_148 vdd gnd cell_6t
Xbit_r149_c253 bl_253 br_253 wl_149 vdd gnd cell_6t
Xbit_r150_c253 bl_253 br_253 wl_150 vdd gnd cell_6t
Xbit_r151_c253 bl_253 br_253 wl_151 vdd gnd cell_6t
Xbit_r152_c253 bl_253 br_253 wl_152 vdd gnd cell_6t
Xbit_r153_c253 bl_253 br_253 wl_153 vdd gnd cell_6t
Xbit_r154_c253 bl_253 br_253 wl_154 vdd gnd cell_6t
Xbit_r155_c253 bl_253 br_253 wl_155 vdd gnd cell_6t
Xbit_r156_c253 bl_253 br_253 wl_156 vdd gnd cell_6t
Xbit_r157_c253 bl_253 br_253 wl_157 vdd gnd cell_6t
Xbit_r158_c253 bl_253 br_253 wl_158 vdd gnd cell_6t
Xbit_r159_c253 bl_253 br_253 wl_159 vdd gnd cell_6t
Xbit_r160_c253 bl_253 br_253 wl_160 vdd gnd cell_6t
Xbit_r161_c253 bl_253 br_253 wl_161 vdd gnd cell_6t
Xbit_r162_c253 bl_253 br_253 wl_162 vdd gnd cell_6t
Xbit_r163_c253 bl_253 br_253 wl_163 vdd gnd cell_6t
Xbit_r164_c253 bl_253 br_253 wl_164 vdd gnd cell_6t
Xbit_r165_c253 bl_253 br_253 wl_165 vdd gnd cell_6t
Xbit_r166_c253 bl_253 br_253 wl_166 vdd gnd cell_6t
Xbit_r167_c253 bl_253 br_253 wl_167 vdd gnd cell_6t
Xbit_r168_c253 bl_253 br_253 wl_168 vdd gnd cell_6t
Xbit_r169_c253 bl_253 br_253 wl_169 vdd gnd cell_6t
Xbit_r170_c253 bl_253 br_253 wl_170 vdd gnd cell_6t
Xbit_r171_c253 bl_253 br_253 wl_171 vdd gnd cell_6t
Xbit_r172_c253 bl_253 br_253 wl_172 vdd gnd cell_6t
Xbit_r173_c253 bl_253 br_253 wl_173 vdd gnd cell_6t
Xbit_r174_c253 bl_253 br_253 wl_174 vdd gnd cell_6t
Xbit_r175_c253 bl_253 br_253 wl_175 vdd gnd cell_6t
Xbit_r176_c253 bl_253 br_253 wl_176 vdd gnd cell_6t
Xbit_r177_c253 bl_253 br_253 wl_177 vdd gnd cell_6t
Xbit_r178_c253 bl_253 br_253 wl_178 vdd gnd cell_6t
Xbit_r179_c253 bl_253 br_253 wl_179 vdd gnd cell_6t
Xbit_r180_c253 bl_253 br_253 wl_180 vdd gnd cell_6t
Xbit_r181_c253 bl_253 br_253 wl_181 vdd gnd cell_6t
Xbit_r182_c253 bl_253 br_253 wl_182 vdd gnd cell_6t
Xbit_r183_c253 bl_253 br_253 wl_183 vdd gnd cell_6t
Xbit_r184_c253 bl_253 br_253 wl_184 vdd gnd cell_6t
Xbit_r185_c253 bl_253 br_253 wl_185 vdd gnd cell_6t
Xbit_r186_c253 bl_253 br_253 wl_186 vdd gnd cell_6t
Xbit_r187_c253 bl_253 br_253 wl_187 vdd gnd cell_6t
Xbit_r188_c253 bl_253 br_253 wl_188 vdd gnd cell_6t
Xbit_r189_c253 bl_253 br_253 wl_189 vdd gnd cell_6t
Xbit_r190_c253 bl_253 br_253 wl_190 vdd gnd cell_6t
Xbit_r191_c253 bl_253 br_253 wl_191 vdd gnd cell_6t
Xbit_r192_c253 bl_253 br_253 wl_192 vdd gnd cell_6t
Xbit_r193_c253 bl_253 br_253 wl_193 vdd gnd cell_6t
Xbit_r194_c253 bl_253 br_253 wl_194 vdd gnd cell_6t
Xbit_r195_c253 bl_253 br_253 wl_195 vdd gnd cell_6t
Xbit_r196_c253 bl_253 br_253 wl_196 vdd gnd cell_6t
Xbit_r197_c253 bl_253 br_253 wl_197 vdd gnd cell_6t
Xbit_r198_c253 bl_253 br_253 wl_198 vdd gnd cell_6t
Xbit_r199_c253 bl_253 br_253 wl_199 vdd gnd cell_6t
Xbit_r200_c253 bl_253 br_253 wl_200 vdd gnd cell_6t
Xbit_r201_c253 bl_253 br_253 wl_201 vdd gnd cell_6t
Xbit_r202_c253 bl_253 br_253 wl_202 vdd gnd cell_6t
Xbit_r203_c253 bl_253 br_253 wl_203 vdd gnd cell_6t
Xbit_r204_c253 bl_253 br_253 wl_204 vdd gnd cell_6t
Xbit_r205_c253 bl_253 br_253 wl_205 vdd gnd cell_6t
Xbit_r206_c253 bl_253 br_253 wl_206 vdd gnd cell_6t
Xbit_r207_c253 bl_253 br_253 wl_207 vdd gnd cell_6t
Xbit_r208_c253 bl_253 br_253 wl_208 vdd gnd cell_6t
Xbit_r209_c253 bl_253 br_253 wl_209 vdd gnd cell_6t
Xbit_r210_c253 bl_253 br_253 wl_210 vdd gnd cell_6t
Xbit_r211_c253 bl_253 br_253 wl_211 vdd gnd cell_6t
Xbit_r212_c253 bl_253 br_253 wl_212 vdd gnd cell_6t
Xbit_r213_c253 bl_253 br_253 wl_213 vdd gnd cell_6t
Xbit_r214_c253 bl_253 br_253 wl_214 vdd gnd cell_6t
Xbit_r215_c253 bl_253 br_253 wl_215 vdd gnd cell_6t
Xbit_r216_c253 bl_253 br_253 wl_216 vdd gnd cell_6t
Xbit_r217_c253 bl_253 br_253 wl_217 vdd gnd cell_6t
Xbit_r218_c253 bl_253 br_253 wl_218 vdd gnd cell_6t
Xbit_r219_c253 bl_253 br_253 wl_219 vdd gnd cell_6t
Xbit_r220_c253 bl_253 br_253 wl_220 vdd gnd cell_6t
Xbit_r221_c253 bl_253 br_253 wl_221 vdd gnd cell_6t
Xbit_r222_c253 bl_253 br_253 wl_222 vdd gnd cell_6t
Xbit_r223_c253 bl_253 br_253 wl_223 vdd gnd cell_6t
Xbit_r224_c253 bl_253 br_253 wl_224 vdd gnd cell_6t
Xbit_r225_c253 bl_253 br_253 wl_225 vdd gnd cell_6t
Xbit_r226_c253 bl_253 br_253 wl_226 vdd gnd cell_6t
Xbit_r227_c253 bl_253 br_253 wl_227 vdd gnd cell_6t
Xbit_r228_c253 bl_253 br_253 wl_228 vdd gnd cell_6t
Xbit_r229_c253 bl_253 br_253 wl_229 vdd gnd cell_6t
Xbit_r230_c253 bl_253 br_253 wl_230 vdd gnd cell_6t
Xbit_r231_c253 bl_253 br_253 wl_231 vdd gnd cell_6t
Xbit_r232_c253 bl_253 br_253 wl_232 vdd gnd cell_6t
Xbit_r233_c253 bl_253 br_253 wl_233 vdd gnd cell_6t
Xbit_r234_c253 bl_253 br_253 wl_234 vdd gnd cell_6t
Xbit_r235_c253 bl_253 br_253 wl_235 vdd gnd cell_6t
Xbit_r236_c253 bl_253 br_253 wl_236 vdd gnd cell_6t
Xbit_r237_c253 bl_253 br_253 wl_237 vdd gnd cell_6t
Xbit_r238_c253 bl_253 br_253 wl_238 vdd gnd cell_6t
Xbit_r239_c253 bl_253 br_253 wl_239 vdd gnd cell_6t
Xbit_r240_c253 bl_253 br_253 wl_240 vdd gnd cell_6t
Xbit_r241_c253 bl_253 br_253 wl_241 vdd gnd cell_6t
Xbit_r242_c253 bl_253 br_253 wl_242 vdd gnd cell_6t
Xbit_r243_c253 bl_253 br_253 wl_243 vdd gnd cell_6t
Xbit_r244_c253 bl_253 br_253 wl_244 vdd gnd cell_6t
Xbit_r245_c253 bl_253 br_253 wl_245 vdd gnd cell_6t
Xbit_r246_c253 bl_253 br_253 wl_246 vdd gnd cell_6t
Xbit_r247_c253 bl_253 br_253 wl_247 vdd gnd cell_6t
Xbit_r248_c253 bl_253 br_253 wl_248 vdd gnd cell_6t
Xbit_r249_c253 bl_253 br_253 wl_249 vdd gnd cell_6t
Xbit_r250_c253 bl_253 br_253 wl_250 vdd gnd cell_6t
Xbit_r251_c253 bl_253 br_253 wl_251 vdd gnd cell_6t
Xbit_r252_c253 bl_253 br_253 wl_252 vdd gnd cell_6t
Xbit_r253_c253 bl_253 br_253 wl_253 vdd gnd cell_6t
Xbit_r254_c253 bl_253 br_253 wl_254 vdd gnd cell_6t
Xbit_r255_c253 bl_253 br_253 wl_255 vdd gnd cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd cell_6t
Xbit_r1_c254 bl_254 br_254 wl_1 vdd gnd cell_6t
Xbit_r2_c254 bl_254 br_254 wl_2 vdd gnd cell_6t
Xbit_r3_c254 bl_254 br_254 wl_3 vdd gnd cell_6t
Xbit_r4_c254 bl_254 br_254 wl_4 vdd gnd cell_6t
Xbit_r5_c254 bl_254 br_254 wl_5 vdd gnd cell_6t
Xbit_r6_c254 bl_254 br_254 wl_6 vdd gnd cell_6t
Xbit_r7_c254 bl_254 br_254 wl_7 vdd gnd cell_6t
Xbit_r8_c254 bl_254 br_254 wl_8 vdd gnd cell_6t
Xbit_r9_c254 bl_254 br_254 wl_9 vdd gnd cell_6t
Xbit_r10_c254 bl_254 br_254 wl_10 vdd gnd cell_6t
Xbit_r11_c254 bl_254 br_254 wl_11 vdd gnd cell_6t
Xbit_r12_c254 bl_254 br_254 wl_12 vdd gnd cell_6t
Xbit_r13_c254 bl_254 br_254 wl_13 vdd gnd cell_6t
Xbit_r14_c254 bl_254 br_254 wl_14 vdd gnd cell_6t
Xbit_r15_c254 bl_254 br_254 wl_15 vdd gnd cell_6t
Xbit_r16_c254 bl_254 br_254 wl_16 vdd gnd cell_6t
Xbit_r17_c254 bl_254 br_254 wl_17 vdd gnd cell_6t
Xbit_r18_c254 bl_254 br_254 wl_18 vdd gnd cell_6t
Xbit_r19_c254 bl_254 br_254 wl_19 vdd gnd cell_6t
Xbit_r20_c254 bl_254 br_254 wl_20 vdd gnd cell_6t
Xbit_r21_c254 bl_254 br_254 wl_21 vdd gnd cell_6t
Xbit_r22_c254 bl_254 br_254 wl_22 vdd gnd cell_6t
Xbit_r23_c254 bl_254 br_254 wl_23 vdd gnd cell_6t
Xbit_r24_c254 bl_254 br_254 wl_24 vdd gnd cell_6t
Xbit_r25_c254 bl_254 br_254 wl_25 vdd gnd cell_6t
Xbit_r26_c254 bl_254 br_254 wl_26 vdd gnd cell_6t
Xbit_r27_c254 bl_254 br_254 wl_27 vdd gnd cell_6t
Xbit_r28_c254 bl_254 br_254 wl_28 vdd gnd cell_6t
Xbit_r29_c254 bl_254 br_254 wl_29 vdd gnd cell_6t
Xbit_r30_c254 bl_254 br_254 wl_30 vdd gnd cell_6t
Xbit_r31_c254 bl_254 br_254 wl_31 vdd gnd cell_6t
Xbit_r32_c254 bl_254 br_254 wl_32 vdd gnd cell_6t
Xbit_r33_c254 bl_254 br_254 wl_33 vdd gnd cell_6t
Xbit_r34_c254 bl_254 br_254 wl_34 vdd gnd cell_6t
Xbit_r35_c254 bl_254 br_254 wl_35 vdd gnd cell_6t
Xbit_r36_c254 bl_254 br_254 wl_36 vdd gnd cell_6t
Xbit_r37_c254 bl_254 br_254 wl_37 vdd gnd cell_6t
Xbit_r38_c254 bl_254 br_254 wl_38 vdd gnd cell_6t
Xbit_r39_c254 bl_254 br_254 wl_39 vdd gnd cell_6t
Xbit_r40_c254 bl_254 br_254 wl_40 vdd gnd cell_6t
Xbit_r41_c254 bl_254 br_254 wl_41 vdd gnd cell_6t
Xbit_r42_c254 bl_254 br_254 wl_42 vdd gnd cell_6t
Xbit_r43_c254 bl_254 br_254 wl_43 vdd gnd cell_6t
Xbit_r44_c254 bl_254 br_254 wl_44 vdd gnd cell_6t
Xbit_r45_c254 bl_254 br_254 wl_45 vdd gnd cell_6t
Xbit_r46_c254 bl_254 br_254 wl_46 vdd gnd cell_6t
Xbit_r47_c254 bl_254 br_254 wl_47 vdd gnd cell_6t
Xbit_r48_c254 bl_254 br_254 wl_48 vdd gnd cell_6t
Xbit_r49_c254 bl_254 br_254 wl_49 vdd gnd cell_6t
Xbit_r50_c254 bl_254 br_254 wl_50 vdd gnd cell_6t
Xbit_r51_c254 bl_254 br_254 wl_51 vdd gnd cell_6t
Xbit_r52_c254 bl_254 br_254 wl_52 vdd gnd cell_6t
Xbit_r53_c254 bl_254 br_254 wl_53 vdd gnd cell_6t
Xbit_r54_c254 bl_254 br_254 wl_54 vdd gnd cell_6t
Xbit_r55_c254 bl_254 br_254 wl_55 vdd gnd cell_6t
Xbit_r56_c254 bl_254 br_254 wl_56 vdd gnd cell_6t
Xbit_r57_c254 bl_254 br_254 wl_57 vdd gnd cell_6t
Xbit_r58_c254 bl_254 br_254 wl_58 vdd gnd cell_6t
Xbit_r59_c254 bl_254 br_254 wl_59 vdd gnd cell_6t
Xbit_r60_c254 bl_254 br_254 wl_60 vdd gnd cell_6t
Xbit_r61_c254 bl_254 br_254 wl_61 vdd gnd cell_6t
Xbit_r62_c254 bl_254 br_254 wl_62 vdd gnd cell_6t
Xbit_r63_c254 bl_254 br_254 wl_63 vdd gnd cell_6t
Xbit_r64_c254 bl_254 br_254 wl_64 vdd gnd cell_6t
Xbit_r65_c254 bl_254 br_254 wl_65 vdd gnd cell_6t
Xbit_r66_c254 bl_254 br_254 wl_66 vdd gnd cell_6t
Xbit_r67_c254 bl_254 br_254 wl_67 vdd gnd cell_6t
Xbit_r68_c254 bl_254 br_254 wl_68 vdd gnd cell_6t
Xbit_r69_c254 bl_254 br_254 wl_69 vdd gnd cell_6t
Xbit_r70_c254 bl_254 br_254 wl_70 vdd gnd cell_6t
Xbit_r71_c254 bl_254 br_254 wl_71 vdd gnd cell_6t
Xbit_r72_c254 bl_254 br_254 wl_72 vdd gnd cell_6t
Xbit_r73_c254 bl_254 br_254 wl_73 vdd gnd cell_6t
Xbit_r74_c254 bl_254 br_254 wl_74 vdd gnd cell_6t
Xbit_r75_c254 bl_254 br_254 wl_75 vdd gnd cell_6t
Xbit_r76_c254 bl_254 br_254 wl_76 vdd gnd cell_6t
Xbit_r77_c254 bl_254 br_254 wl_77 vdd gnd cell_6t
Xbit_r78_c254 bl_254 br_254 wl_78 vdd gnd cell_6t
Xbit_r79_c254 bl_254 br_254 wl_79 vdd gnd cell_6t
Xbit_r80_c254 bl_254 br_254 wl_80 vdd gnd cell_6t
Xbit_r81_c254 bl_254 br_254 wl_81 vdd gnd cell_6t
Xbit_r82_c254 bl_254 br_254 wl_82 vdd gnd cell_6t
Xbit_r83_c254 bl_254 br_254 wl_83 vdd gnd cell_6t
Xbit_r84_c254 bl_254 br_254 wl_84 vdd gnd cell_6t
Xbit_r85_c254 bl_254 br_254 wl_85 vdd gnd cell_6t
Xbit_r86_c254 bl_254 br_254 wl_86 vdd gnd cell_6t
Xbit_r87_c254 bl_254 br_254 wl_87 vdd gnd cell_6t
Xbit_r88_c254 bl_254 br_254 wl_88 vdd gnd cell_6t
Xbit_r89_c254 bl_254 br_254 wl_89 vdd gnd cell_6t
Xbit_r90_c254 bl_254 br_254 wl_90 vdd gnd cell_6t
Xbit_r91_c254 bl_254 br_254 wl_91 vdd gnd cell_6t
Xbit_r92_c254 bl_254 br_254 wl_92 vdd gnd cell_6t
Xbit_r93_c254 bl_254 br_254 wl_93 vdd gnd cell_6t
Xbit_r94_c254 bl_254 br_254 wl_94 vdd gnd cell_6t
Xbit_r95_c254 bl_254 br_254 wl_95 vdd gnd cell_6t
Xbit_r96_c254 bl_254 br_254 wl_96 vdd gnd cell_6t
Xbit_r97_c254 bl_254 br_254 wl_97 vdd gnd cell_6t
Xbit_r98_c254 bl_254 br_254 wl_98 vdd gnd cell_6t
Xbit_r99_c254 bl_254 br_254 wl_99 vdd gnd cell_6t
Xbit_r100_c254 bl_254 br_254 wl_100 vdd gnd cell_6t
Xbit_r101_c254 bl_254 br_254 wl_101 vdd gnd cell_6t
Xbit_r102_c254 bl_254 br_254 wl_102 vdd gnd cell_6t
Xbit_r103_c254 bl_254 br_254 wl_103 vdd gnd cell_6t
Xbit_r104_c254 bl_254 br_254 wl_104 vdd gnd cell_6t
Xbit_r105_c254 bl_254 br_254 wl_105 vdd gnd cell_6t
Xbit_r106_c254 bl_254 br_254 wl_106 vdd gnd cell_6t
Xbit_r107_c254 bl_254 br_254 wl_107 vdd gnd cell_6t
Xbit_r108_c254 bl_254 br_254 wl_108 vdd gnd cell_6t
Xbit_r109_c254 bl_254 br_254 wl_109 vdd gnd cell_6t
Xbit_r110_c254 bl_254 br_254 wl_110 vdd gnd cell_6t
Xbit_r111_c254 bl_254 br_254 wl_111 vdd gnd cell_6t
Xbit_r112_c254 bl_254 br_254 wl_112 vdd gnd cell_6t
Xbit_r113_c254 bl_254 br_254 wl_113 vdd gnd cell_6t
Xbit_r114_c254 bl_254 br_254 wl_114 vdd gnd cell_6t
Xbit_r115_c254 bl_254 br_254 wl_115 vdd gnd cell_6t
Xbit_r116_c254 bl_254 br_254 wl_116 vdd gnd cell_6t
Xbit_r117_c254 bl_254 br_254 wl_117 vdd gnd cell_6t
Xbit_r118_c254 bl_254 br_254 wl_118 vdd gnd cell_6t
Xbit_r119_c254 bl_254 br_254 wl_119 vdd gnd cell_6t
Xbit_r120_c254 bl_254 br_254 wl_120 vdd gnd cell_6t
Xbit_r121_c254 bl_254 br_254 wl_121 vdd gnd cell_6t
Xbit_r122_c254 bl_254 br_254 wl_122 vdd gnd cell_6t
Xbit_r123_c254 bl_254 br_254 wl_123 vdd gnd cell_6t
Xbit_r124_c254 bl_254 br_254 wl_124 vdd gnd cell_6t
Xbit_r125_c254 bl_254 br_254 wl_125 vdd gnd cell_6t
Xbit_r126_c254 bl_254 br_254 wl_126 vdd gnd cell_6t
Xbit_r127_c254 bl_254 br_254 wl_127 vdd gnd cell_6t
Xbit_r128_c254 bl_254 br_254 wl_128 vdd gnd cell_6t
Xbit_r129_c254 bl_254 br_254 wl_129 vdd gnd cell_6t
Xbit_r130_c254 bl_254 br_254 wl_130 vdd gnd cell_6t
Xbit_r131_c254 bl_254 br_254 wl_131 vdd gnd cell_6t
Xbit_r132_c254 bl_254 br_254 wl_132 vdd gnd cell_6t
Xbit_r133_c254 bl_254 br_254 wl_133 vdd gnd cell_6t
Xbit_r134_c254 bl_254 br_254 wl_134 vdd gnd cell_6t
Xbit_r135_c254 bl_254 br_254 wl_135 vdd gnd cell_6t
Xbit_r136_c254 bl_254 br_254 wl_136 vdd gnd cell_6t
Xbit_r137_c254 bl_254 br_254 wl_137 vdd gnd cell_6t
Xbit_r138_c254 bl_254 br_254 wl_138 vdd gnd cell_6t
Xbit_r139_c254 bl_254 br_254 wl_139 vdd gnd cell_6t
Xbit_r140_c254 bl_254 br_254 wl_140 vdd gnd cell_6t
Xbit_r141_c254 bl_254 br_254 wl_141 vdd gnd cell_6t
Xbit_r142_c254 bl_254 br_254 wl_142 vdd gnd cell_6t
Xbit_r143_c254 bl_254 br_254 wl_143 vdd gnd cell_6t
Xbit_r144_c254 bl_254 br_254 wl_144 vdd gnd cell_6t
Xbit_r145_c254 bl_254 br_254 wl_145 vdd gnd cell_6t
Xbit_r146_c254 bl_254 br_254 wl_146 vdd gnd cell_6t
Xbit_r147_c254 bl_254 br_254 wl_147 vdd gnd cell_6t
Xbit_r148_c254 bl_254 br_254 wl_148 vdd gnd cell_6t
Xbit_r149_c254 bl_254 br_254 wl_149 vdd gnd cell_6t
Xbit_r150_c254 bl_254 br_254 wl_150 vdd gnd cell_6t
Xbit_r151_c254 bl_254 br_254 wl_151 vdd gnd cell_6t
Xbit_r152_c254 bl_254 br_254 wl_152 vdd gnd cell_6t
Xbit_r153_c254 bl_254 br_254 wl_153 vdd gnd cell_6t
Xbit_r154_c254 bl_254 br_254 wl_154 vdd gnd cell_6t
Xbit_r155_c254 bl_254 br_254 wl_155 vdd gnd cell_6t
Xbit_r156_c254 bl_254 br_254 wl_156 vdd gnd cell_6t
Xbit_r157_c254 bl_254 br_254 wl_157 vdd gnd cell_6t
Xbit_r158_c254 bl_254 br_254 wl_158 vdd gnd cell_6t
Xbit_r159_c254 bl_254 br_254 wl_159 vdd gnd cell_6t
Xbit_r160_c254 bl_254 br_254 wl_160 vdd gnd cell_6t
Xbit_r161_c254 bl_254 br_254 wl_161 vdd gnd cell_6t
Xbit_r162_c254 bl_254 br_254 wl_162 vdd gnd cell_6t
Xbit_r163_c254 bl_254 br_254 wl_163 vdd gnd cell_6t
Xbit_r164_c254 bl_254 br_254 wl_164 vdd gnd cell_6t
Xbit_r165_c254 bl_254 br_254 wl_165 vdd gnd cell_6t
Xbit_r166_c254 bl_254 br_254 wl_166 vdd gnd cell_6t
Xbit_r167_c254 bl_254 br_254 wl_167 vdd gnd cell_6t
Xbit_r168_c254 bl_254 br_254 wl_168 vdd gnd cell_6t
Xbit_r169_c254 bl_254 br_254 wl_169 vdd gnd cell_6t
Xbit_r170_c254 bl_254 br_254 wl_170 vdd gnd cell_6t
Xbit_r171_c254 bl_254 br_254 wl_171 vdd gnd cell_6t
Xbit_r172_c254 bl_254 br_254 wl_172 vdd gnd cell_6t
Xbit_r173_c254 bl_254 br_254 wl_173 vdd gnd cell_6t
Xbit_r174_c254 bl_254 br_254 wl_174 vdd gnd cell_6t
Xbit_r175_c254 bl_254 br_254 wl_175 vdd gnd cell_6t
Xbit_r176_c254 bl_254 br_254 wl_176 vdd gnd cell_6t
Xbit_r177_c254 bl_254 br_254 wl_177 vdd gnd cell_6t
Xbit_r178_c254 bl_254 br_254 wl_178 vdd gnd cell_6t
Xbit_r179_c254 bl_254 br_254 wl_179 vdd gnd cell_6t
Xbit_r180_c254 bl_254 br_254 wl_180 vdd gnd cell_6t
Xbit_r181_c254 bl_254 br_254 wl_181 vdd gnd cell_6t
Xbit_r182_c254 bl_254 br_254 wl_182 vdd gnd cell_6t
Xbit_r183_c254 bl_254 br_254 wl_183 vdd gnd cell_6t
Xbit_r184_c254 bl_254 br_254 wl_184 vdd gnd cell_6t
Xbit_r185_c254 bl_254 br_254 wl_185 vdd gnd cell_6t
Xbit_r186_c254 bl_254 br_254 wl_186 vdd gnd cell_6t
Xbit_r187_c254 bl_254 br_254 wl_187 vdd gnd cell_6t
Xbit_r188_c254 bl_254 br_254 wl_188 vdd gnd cell_6t
Xbit_r189_c254 bl_254 br_254 wl_189 vdd gnd cell_6t
Xbit_r190_c254 bl_254 br_254 wl_190 vdd gnd cell_6t
Xbit_r191_c254 bl_254 br_254 wl_191 vdd gnd cell_6t
Xbit_r192_c254 bl_254 br_254 wl_192 vdd gnd cell_6t
Xbit_r193_c254 bl_254 br_254 wl_193 vdd gnd cell_6t
Xbit_r194_c254 bl_254 br_254 wl_194 vdd gnd cell_6t
Xbit_r195_c254 bl_254 br_254 wl_195 vdd gnd cell_6t
Xbit_r196_c254 bl_254 br_254 wl_196 vdd gnd cell_6t
Xbit_r197_c254 bl_254 br_254 wl_197 vdd gnd cell_6t
Xbit_r198_c254 bl_254 br_254 wl_198 vdd gnd cell_6t
Xbit_r199_c254 bl_254 br_254 wl_199 vdd gnd cell_6t
Xbit_r200_c254 bl_254 br_254 wl_200 vdd gnd cell_6t
Xbit_r201_c254 bl_254 br_254 wl_201 vdd gnd cell_6t
Xbit_r202_c254 bl_254 br_254 wl_202 vdd gnd cell_6t
Xbit_r203_c254 bl_254 br_254 wl_203 vdd gnd cell_6t
Xbit_r204_c254 bl_254 br_254 wl_204 vdd gnd cell_6t
Xbit_r205_c254 bl_254 br_254 wl_205 vdd gnd cell_6t
Xbit_r206_c254 bl_254 br_254 wl_206 vdd gnd cell_6t
Xbit_r207_c254 bl_254 br_254 wl_207 vdd gnd cell_6t
Xbit_r208_c254 bl_254 br_254 wl_208 vdd gnd cell_6t
Xbit_r209_c254 bl_254 br_254 wl_209 vdd gnd cell_6t
Xbit_r210_c254 bl_254 br_254 wl_210 vdd gnd cell_6t
Xbit_r211_c254 bl_254 br_254 wl_211 vdd gnd cell_6t
Xbit_r212_c254 bl_254 br_254 wl_212 vdd gnd cell_6t
Xbit_r213_c254 bl_254 br_254 wl_213 vdd gnd cell_6t
Xbit_r214_c254 bl_254 br_254 wl_214 vdd gnd cell_6t
Xbit_r215_c254 bl_254 br_254 wl_215 vdd gnd cell_6t
Xbit_r216_c254 bl_254 br_254 wl_216 vdd gnd cell_6t
Xbit_r217_c254 bl_254 br_254 wl_217 vdd gnd cell_6t
Xbit_r218_c254 bl_254 br_254 wl_218 vdd gnd cell_6t
Xbit_r219_c254 bl_254 br_254 wl_219 vdd gnd cell_6t
Xbit_r220_c254 bl_254 br_254 wl_220 vdd gnd cell_6t
Xbit_r221_c254 bl_254 br_254 wl_221 vdd gnd cell_6t
Xbit_r222_c254 bl_254 br_254 wl_222 vdd gnd cell_6t
Xbit_r223_c254 bl_254 br_254 wl_223 vdd gnd cell_6t
Xbit_r224_c254 bl_254 br_254 wl_224 vdd gnd cell_6t
Xbit_r225_c254 bl_254 br_254 wl_225 vdd gnd cell_6t
Xbit_r226_c254 bl_254 br_254 wl_226 vdd gnd cell_6t
Xbit_r227_c254 bl_254 br_254 wl_227 vdd gnd cell_6t
Xbit_r228_c254 bl_254 br_254 wl_228 vdd gnd cell_6t
Xbit_r229_c254 bl_254 br_254 wl_229 vdd gnd cell_6t
Xbit_r230_c254 bl_254 br_254 wl_230 vdd gnd cell_6t
Xbit_r231_c254 bl_254 br_254 wl_231 vdd gnd cell_6t
Xbit_r232_c254 bl_254 br_254 wl_232 vdd gnd cell_6t
Xbit_r233_c254 bl_254 br_254 wl_233 vdd gnd cell_6t
Xbit_r234_c254 bl_254 br_254 wl_234 vdd gnd cell_6t
Xbit_r235_c254 bl_254 br_254 wl_235 vdd gnd cell_6t
Xbit_r236_c254 bl_254 br_254 wl_236 vdd gnd cell_6t
Xbit_r237_c254 bl_254 br_254 wl_237 vdd gnd cell_6t
Xbit_r238_c254 bl_254 br_254 wl_238 vdd gnd cell_6t
Xbit_r239_c254 bl_254 br_254 wl_239 vdd gnd cell_6t
Xbit_r240_c254 bl_254 br_254 wl_240 vdd gnd cell_6t
Xbit_r241_c254 bl_254 br_254 wl_241 vdd gnd cell_6t
Xbit_r242_c254 bl_254 br_254 wl_242 vdd gnd cell_6t
Xbit_r243_c254 bl_254 br_254 wl_243 vdd gnd cell_6t
Xbit_r244_c254 bl_254 br_254 wl_244 vdd gnd cell_6t
Xbit_r245_c254 bl_254 br_254 wl_245 vdd gnd cell_6t
Xbit_r246_c254 bl_254 br_254 wl_246 vdd gnd cell_6t
Xbit_r247_c254 bl_254 br_254 wl_247 vdd gnd cell_6t
Xbit_r248_c254 bl_254 br_254 wl_248 vdd gnd cell_6t
Xbit_r249_c254 bl_254 br_254 wl_249 vdd gnd cell_6t
Xbit_r250_c254 bl_254 br_254 wl_250 vdd gnd cell_6t
Xbit_r251_c254 bl_254 br_254 wl_251 vdd gnd cell_6t
Xbit_r252_c254 bl_254 br_254 wl_252 vdd gnd cell_6t
Xbit_r253_c254 bl_254 br_254 wl_253 vdd gnd cell_6t
Xbit_r254_c254 bl_254 br_254 wl_254 vdd gnd cell_6t
Xbit_r255_c254 bl_254 br_254 wl_255 vdd gnd cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd cell_6t
Xbit_r1_c255 bl_255 br_255 wl_1 vdd gnd cell_6t
Xbit_r2_c255 bl_255 br_255 wl_2 vdd gnd cell_6t
Xbit_r3_c255 bl_255 br_255 wl_3 vdd gnd cell_6t
Xbit_r4_c255 bl_255 br_255 wl_4 vdd gnd cell_6t
Xbit_r5_c255 bl_255 br_255 wl_5 vdd gnd cell_6t
Xbit_r6_c255 bl_255 br_255 wl_6 vdd gnd cell_6t
Xbit_r7_c255 bl_255 br_255 wl_7 vdd gnd cell_6t
Xbit_r8_c255 bl_255 br_255 wl_8 vdd gnd cell_6t
Xbit_r9_c255 bl_255 br_255 wl_9 vdd gnd cell_6t
Xbit_r10_c255 bl_255 br_255 wl_10 vdd gnd cell_6t
Xbit_r11_c255 bl_255 br_255 wl_11 vdd gnd cell_6t
Xbit_r12_c255 bl_255 br_255 wl_12 vdd gnd cell_6t
Xbit_r13_c255 bl_255 br_255 wl_13 vdd gnd cell_6t
Xbit_r14_c255 bl_255 br_255 wl_14 vdd gnd cell_6t
Xbit_r15_c255 bl_255 br_255 wl_15 vdd gnd cell_6t
Xbit_r16_c255 bl_255 br_255 wl_16 vdd gnd cell_6t
Xbit_r17_c255 bl_255 br_255 wl_17 vdd gnd cell_6t
Xbit_r18_c255 bl_255 br_255 wl_18 vdd gnd cell_6t
Xbit_r19_c255 bl_255 br_255 wl_19 vdd gnd cell_6t
Xbit_r20_c255 bl_255 br_255 wl_20 vdd gnd cell_6t
Xbit_r21_c255 bl_255 br_255 wl_21 vdd gnd cell_6t
Xbit_r22_c255 bl_255 br_255 wl_22 vdd gnd cell_6t
Xbit_r23_c255 bl_255 br_255 wl_23 vdd gnd cell_6t
Xbit_r24_c255 bl_255 br_255 wl_24 vdd gnd cell_6t
Xbit_r25_c255 bl_255 br_255 wl_25 vdd gnd cell_6t
Xbit_r26_c255 bl_255 br_255 wl_26 vdd gnd cell_6t
Xbit_r27_c255 bl_255 br_255 wl_27 vdd gnd cell_6t
Xbit_r28_c255 bl_255 br_255 wl_28 vdd gnd cell_6t
Xbit_r29_c255 bl_255 br_255 wl_29 vdd gnd cell_6t
Xbit_r30_c255 bl_255 br_255 wl_30 vdd gnd cell_6t
Xbit_r31_c255 bl_255 br_255 wl_31 vdd gnd cell_6t
Xbit_r32_c255 bl_255 br_255 wl_32 vdd gnd cell_6t
Xbit_r33_c255 bl_255 br_255 wl_33 vdd gnd cell_6t
Xbit_r34_c255 bl_255 br_255 wl_34 vdd gnd cell_6t
Xbit_r35_c255 bl_255 br_255 wl_35 vdd gnd cell_6t
Xbit_r36_c255 bl_255 br_255 wl_36 vdd gnd cell_6t
Xbit_r37_c255 bl_255 br_255 wl_37 vdd gnd cell_6t
Xbit_r38_c255 bl_255 br_255 wl_38 vdd gnd cell_6t
Xbit_r39_c255 bl_255 br_255 wl_39 vdd gnd cell_6t
Xbit_r40_c255 bl_255 br_255 wl_40 vdd gnd cell_6t
Xbit_r41_c255 bl_255 br_255 wl_41 vdd gnd cell_6t
Xbit_r42_c255 bl_255 br_255 wl_42 vdd gnd cell_6t
Xbit_r43_c255 bl_255 br_255 wl_43 vdd gnd cell_6t
Xbit_r44_c255 bl_255 br_255 wl_44 vdd gnd cell_6t
Xbit_r45_c255 bl_255 br_255 wl_45 vdd gnd cell_6t
Xbit_r46_c255 bl_255 br_255 wl_46 vdd gnd cell_6t
Xbit_r47_c255 bl_255 br_255 wl_47 vdd gnd cell_6t
Xbit_r48_c255 bl_255 br_255 wl_48 vdd gnd cell_6t
Xbit_r49_c255 bl_255 br_255 wl_49 vdd gnd cell_6t
Xbit_r50_c255 bl_255 br_255 wl_50 vdd gnd cell_6t
Xbit_r51_c255 bl_255 br_255 wl_51 vdd gnd cell_6t
Xbit_r52_c255 bl_255 br_255 wl_52 vdd gnd cell_6t
Xbit_r53_c255 bl_255 br_255 wl_53 vdd gnd cell_6t
Xbit_r54_c255 bl_255 br_255 wl_54 vdd gnd cell_6t
Xbit_r55_c255 bl_255 br_255 wl_55 vdd gnd cell_6t
Xbit_r56_c255 bl_255 br_255 wl_56 vdd gnd cell_6t
Xbit_r57_c255 bl_255 br_255 wl_57 vdd gnd cell_6t
Xbit_r58_c255 bl_255 br_255 wl_58 vdd gnd cell_6t
Xbit_r59_c255 bl_255 br_255 wl_59 vdd gnd cell_6t
Xbit_r60_c255 bl_255 br_255 wl_60 vdd gnd cell_6t
Xbit_r61_c255 bl_255 br_255 wl_61 vdd gnd cell_6t
Xbit_r62_c255 bl_255 br_255 wl_62 vdd gnd cell_6t
Xbit_r63_c255 bl_255 br_255 wl_63 vdd gnd cell_6t
Xbit_r64_c255 bl_255 br_255 wl_64 vdd gnd cell_6t
Xbit_r65_c255 bl_255 br_255 wl_65 vdd gnd cell_6t
Xbit_r66_c255 bl_255 br_255 wl_66 vdd gnd cell_6t
Xbit_r67_c255 bl_255 br_255 wl_67 vdd gnd cell_6t
Xbit_r68_c255 bl_255 br_255 wl_68 vdd gnd cell_6t
Xbit_r69_c255 bl_255 br_255 wl_69 vdd gnd cell_6t
Xbit_r70_c255 bl_255 br_255 wl_70 vdd gnd cell_6t
Xbit_r71_c255 bl_255 br_255 wl_71 vdd gnd cell_6t
Xbit_r72_c255 bl_255 br_255 wl_72 vdd gnd cell_6t
Xbit_r73_c255 bl_255 br_255 wl_73 vdd gnd cell_6t
Xbit_r74_c255 bl_255 br_255 wl_74 vdd gnd cell_6t
Xbit_r75_c255 bl_255 br_255 wl_75 vdd gnd cell_6t
Xbit_r76_c255 bl_255 br_255 wl_76 vdd gnd cell_6t
Xbit_r77_c255 bl_255 br_255 wl_77 vdd gnd cell_6t
Xbit_r78_c255 bl_255 br_255 wl_78 vdd gnd cell_6t
Xbit_r79_c255 bl_255 br_255 wl_79 vdd gnd cell_6t
Xbit_r80_c255 bl_255 br_255 wl_80 vdd gnd cell_6t
Xbit_r81_c255 bl_255 br_255 wl_81 vdd gnd cell_6t
Xbit_r82_c255 bl_255 br_255 wl_82 vdd gnd cell_6t
Xbit_r83_c255 bl_255 br_255 wl_83 vdd gnd cell_6t
Xbit_r84_c255 bl_255 br_255 wl_84 vdd gnd cell_6t
Xbit_r85_c255 bl_255 br_255 wl_85 vdd gnd cell_6t
Xbit_r86_c255 bl_255 br_255 wl_86 vdd gnd cell_6t
Xbit_r87_c255 bl_255 br_255 wl_87 vdd gnd cell_6t
Xbit_r88_c255 bl_255 br_255 wl_88 vdd gnd cell_6t
Xbit_r89_c255 bl_255 br_255 wl_89 vdd gnd cell_6t
Xbit_r90_c255 bl_255 br_255 wl_90 vdd gnd cell_6t
Xbit_r91_c255 bl_255 br_255 wl_91 vdd gnd cell_6t
Xbit_r92_c255 bl_255 br_255 wl_92 vdd gnd cell_6t
Xbit_r93_c255 bl_255 br_255 wl_93 vdd gnd cell_6t
Xbit_r94_c255 bl_255 br_255 wl_94 vdd gnd cell_6t
Xbit_r95_c255 bl_255 br_255 wl_95 vdd gnd cell_6t
Xbit_r96_c255 bl_255 br_255 wl_96 vdd gnd cell_6t
Xbit_r97_c255 bl_255 br_255 wl_97 vdd gnd cell_6t
Xbit_r98_c255 bl_255 br_255 wl_98 vdd gnd cell_6t
Xbit_r99_c255 bl_255 br_255 wl_99 vdd gnd cell_6t
Xbit_r100_c255 bl_255 br_255 wl_100 vdd gnd cell_6t
Xbit_r101_c255 bl_255 br_255 wl_101 vdd gnd cell_6t
Xbit_r102_c255 bl_255 br_255 wl_102 vdd gnd cell_6t
Xbit_r103_c255 bl_255 br_255 wl_103 vdd gnd cell_6t
Xbit_r104_c255 bl_255 br_255 wl_104 vdd gnd cell_6t
Xbit_r105_c255 bl_255 br_255 wl_105 vdd gnd cell_6t
Xbit_r106_c255 bl_255 br_255 wl_106 vdd gnd cell_6t
Xbit_r107_c255 bl_255 br_255 wl_107 vdd gnd cell_6t
Xbit_r108_c255 bl_255 br_255 wl_108 vdd gnd cell_6t
Xbit_r109_c255 bl_255 br_255 wl_109 vdd gnd cell_6t
Xbit_r110_c255 bl_255 br_255 wl_110 vdd gnd cell_6t
Xbit_r111_c255 bl_255 br_255 wl_111 vdd gnd cell_6t
Xbit_r112_c255 bl_255 br_255 wl_112 vdd gnd cell_6t
Xbit_r113_c255 bl_255 br_255 wl_113 vdd gnd cell_6t
Xbit_r114_c255 bl_255 br_255 wl_114 vdd gnd cell_6t
Xbit_r115_c255 bl_255 br_255 wl_115 vdd gnd cell_6t
Xbit_r116_c255 bl_255 br_255 wl_116 vdd gnd cell_6t
Xbit_r117_c255 bl_255 br_255 wl_117 vdd gnd cell_6t
Xbit_r118_c255 bl_255 br_255 wl_118 vdd gnd cell_6t
Xbit_r119_c255 bl_255 br_255 wl_119 vdd gnd cell_6t
Xbit_r120_c255 bl_255 br_255 wl_120 vdd gnd cell_6t
Xbit_r121_c255 bl_255 br_255 wl_121 vdd gnd cell_6t
Xbit_r122_c255 bl_255 br_255 wl_122 vdd gnd cell_6t
Xbit_r123_c255 bl_255 br_255 wl_123 vdd gnd cell_6t
Xbit_r124_c255 bl_255 br_255 wl_124 vdd gnd cell_6t
Xbit_r125_c255 bl_255 br_255 wl_125 vdd gnd cell_6t
Xbit_r126_c255 bl_255 br_255 wl_126 vdd gnd cell_6t
Xbit_r127_c255 bl_255 br_255 wl_127 vdd gnd cell_6t
Xbit_r128_c255 bl_255 br_255 wl_128 vdd gnd cell_6t
Xbit_r129_c255 bl_255 br_255 wl_129 vdd gnd cell_6t
Xbit_r130_c255 bl_255 br_255 wl_130 vdd gnd cell_6t
Xbit_r131_c255 bl_255 br_255 wl_131 vdd gnd cell_6t
Xbit_r132_c255 bl_255 br_255 wl_132 vdd gnd cell_6t
Xbit_r133_c255 bl_255 br_255 wl_133 vdd gnd cell_6t
Xbit_r134_c255 bl_255 br_255 wl_134 vdd gnd cell_6t
Xbit_r135_c255 bl_255 br_255 wl_135 vdd gnd cell_6t
Xbit_r136_c255 bl_255 br_255 wl_136 vdd gnd cell_6t
Xbit_r137_c255 bl_255 br_255 wl_137 vdd gnd cell_6t
Xbit_r138_c255 bl_255 br_255 wl_138 vdd gnd cell_6t
Xbit_r139_c255 bl_255 br_255 wl_139 vdd gnd cell_6t
Xbit_r140_c255 bl_255 br_255 wl_140 vdd gnd cell_6t
Xbit_r141_c255 bl_255 br_255 wl_141 vdd gnd cell_6t
Xbit_r142_c255 bl_255 br_255 wl_142 vdd gnd cell_6t
Xbit_r143_c255 bl_255 br_255 wl_143 vdd gnd cell_6t
Xbit_r144_c255 bl_255 br_255 wl_144 vdd gnd cell_6t
Xbit_r145_c255 bl_255 br_255 wl_145 vdd gnd cell_6t
Xbit_r146_c255 bl_255 br_255 wl_146 vdd gnd cell_6t
Xbit_r147_c255 bl_255 br_255 wl_147 vdd gnd cell_6t
Xbit_r148_c255 bl_255 br_255 wl_148 vdd gnd cell_6t
Xbit_r149_c255 bl_255 br_255 wl_149 vdd gnd cell_6t
Xbit_r150_c255 bl_255 br_255 wl_150 vdd gnd cell_6t
Xbit_r151_c255 bl_255 br_255 wl_151 vdd gnd cell_6t
Xbit_r152_c255 bl_255 br_255 wl_152 vdd gnd cell_6t
Xbit_r153_c255 bl_255 br_255 wl_153 vdd gnd cell_6t
Xbit_r154_c255 bl_255 br_255 wl_154 vdd gnd cell_6t
Xbit_r155_c255 bl_255 br_255 wl_155 vdd gnd cell_6t
Xbit_r156_c255 bl_255 br_255 wl_156 vdd gnd cell_6t
Xbit_r157_c255 bl_255 br_255 wl_157 vdd gnd cell_6t
Xbit_r158_c255 bl_255 br_255 wl_158 vdd gnd cell_6t
Xbit_r159_c255 bl_255 br_255 wl_159 vdd gnd cell_6t
Xbit_r160_c255 bl_255 br_255 wl_160 vdd gnd cell_6t
Xbit_r161_c255 bl_255 br_255 wl_161 vdd gnd cell_6t
Xbit_r162_c255 bl_255 br_255 wl_162 vdd gnd cell_6t
Xbit_r163_c255 bl_255 br_255 wl_163 vdd gnd cell_6t
Xbit_r164_c255 bl_255 br_255 wl_164 vdd gnd cell_6t
Xbit_r165_c255 bl_255 br_255 wl_165 vdd gnd cell_6t
Xbit_r166_c255 bl_255 br_255 wl_166 vdd gnd cell_6t
Xbit_r167_c255 bl_255 br_255 wl_167 vdd gnd cell_6t
Xbit_r168_c255 bl_255 br_255 wl_168 vdd gnd cell_6t
Xbit_r169_c255 bl_255 br_255 wl_169 vdd gnd cell_6t
Xbit_r170_c255 bl_255 br_255 wl_170 vdd gnd cell_6t
Xbit_r171_c255 bl_255 br_255 wl_171 vdd gnd cell_6t
Xbit_r172_c255 bl_255 br_255 wl_172 vdd gnd cell_6t
Xbit_r173_c255 bl_255 br_255 wl_173 vdd gnd cell_6t
Xbit_r174_c255 bl_255 br_255 wl_174 vdd gnd cell_6t
Xbit_r175_c255 bl_255 br_255 wl_175 vdd gnd cell_6t
Xbit_r176_c255 bl_255 br_255 wl_176 vdd gnd cell_6t
Xbit_r177_c255 bl_255 br_255 wl_177 vdd gnd cell_6t
Xbit_r178_c255 bl_255 br_255 wl_178 vdd gnd cell_6t
Xbit_r179_c255 bl_255 br_255 wl_179 vdd gnd cell_6t
Xbit_r180_c255 bl_255 br_255 wl_180 vdd gnd cell_6t
Xbit_r181_c255 bl_255 br_255 wl_181 vdd gnd cell_6t
Xbit_r182_c255 bl_255 br_255 wl_182 vdd gnd cell_6t
Xbit_r183_c255 bl_255 br_255 wl_183 vdd gnd cell_6t
Xbit_r184_c255 bl_255 br_255 wl_184 vdd gnd cell_6t
Xbit_r185_c255 bl_255 br_255 wl_185 vdd gnd cell_6t
Xbit_r186_c255 bl_255 br_255 wl_186 vdd gnd cell_6t
Xbit_r187_c255 bl_255 br_255 wl_187 vdd gnd cell_6t
Xbit_r188_c255 bl_255 br_255 wl_188 vdd gnd cell_6t
Xbit_r189_c255 bl_255 br_255 wl_189 vdd gnd cell_6t
Xbit_r190_c255 bl_255 br_255 wl_190 vdd gnd cell_6t
Xbit_r191_c255 bl_255 br_255 wl_191 vdd gnd cell_6t
Xbit_r192_c255 bl_255 br_255 wl_192 vdd gnd cell_6t
Xbit_r193_c255 bl_255 br_255 wl_193 vdd gnd cell_6t
Xbit_r194_c255 bl_255 br_255 wl_194 vdd gnd cell_6t
Xbit_r195_c255 bl_255 br_255 wl_195 vdd gnd cell_6t
Xbit_r196_c255 bl_255 br_255 wl_196 vdd gnd cell_6t
Xbit_r197_c255 bl_255 br_255 wl_197 vdd gnd cell_6t
Xbit_r198_c255 bl_255 br_255 wl_198 vdd gnd cell_6t
Xbit_r199_c255 bl_255 br_255 wl_199 vdd gnd cell_6t
Xbit_r200_c255 bl_255 br_255 wl_200 vdd gnd cell_6t
Xbit_r201_c255 bl_255 br_255 wl_201 vdd gnd cell_6t
Xbit_r202_c255 bl_255 br_255 wl_202 vdd gnd cell_6t
Xbit_r203_c255 bl_255 br_255 wl_203 vdd gnd cell_6t
Xbit_r204_c255 bl_255 br_255 wl_204 vdd gnd cell_6t
Xbit_r205_c255 bl_255 br_255 wl_205 vdd gnd cell_6t
Xbit_r206_c255 bl_255 br_255 wl_206 vdd gnd cell_6t
Xbit_r207_c255 bl_255 br_255 wl_207 vdd gnd cell_6t
Xbit_r208_c255 bl_255 br_255 wl_208 vdd gnd cell_6t
Xbit_r209_c255 bl_255 br_255 wl_209 vdd gnd cell_6t
Xbit_r210_c255 bl_255 br_255 wl_210 vdd gnd cell_6t
Xbit_r211_c255 bl_255 br_255 wl_211 vdd gnd cell_6t
Xbit_r212_c255 bl_255 br_255 wl_212 vdd gnd cell_6t
Xbit_r213_c255 bl_255 br_255 wl_213 vdd gnd cell_6t
Xbit_r214_c255 bl_255 br_255 wl_214 vdd gnd cell_6t
Xbit_r215_c255 bl_255 br_255 wl_215 vdd gnd cell_6t
Xbit_r216_c255 bl_255 br_255 wl_216 vdd gnd cell_6t
Xbit_r217_c255 bl_255 br_255 wl_217 vdd gnd cell_6t
Xbit_r218_c255 bl_255 br_255 wl_218 vdd gnd cell_6t
Xbit_r219_c255 bl_255 br_255 wl_219 vdd gnd cell_6t
Xbit_r220_c255 bl_255 br_255 wl_220 vdd gnd cell_6t
Xbit_r221_c255 bl_255 br_255 wl_221 vdd gnd cell_6t
Xbit_r222_c255 bl_255 br_255 wl_222 vdd gnd cell_6t
Xbit_r223_c255 bl_255 br_255 wl_223 vdd gnd cell_6t
Xbit_r224_c255 bl_255 br_255 wl_224 vdd gnd cell_6t
Xbit_r225_c255 bl_255 br_255 wl_225 vdd gnd cell_6t
Xbit_r226_c255 bl_255 br_255 wl_226 vdd gnd cell_6t
Xbit_r227_c255 bl_255 br_255 wl_227 vdd gnd cell_6t
Xbit_r228_c255 bl_255 br_255 wl_228 vdd gnd cell_6t
Xbit_r229_c255 bl_255 br_255 wl_229 vdd gnd cell_6t
Xbit_r230_c255 bl_255 br_255 wl_230 vdd gnd cell_6t
Xbit_r231_c255 bl_255 br_255 wl_231 vdd gnd cell_6t
Xbit_r232_c255 bl_255 br_255 wl_232 vdd gnd cell_6t
Xbit_r233_c255 bl_255 br_255 wl_233 vdd gnd cell_6t
Xbit_r234_c255 bl_255 br_255 wl_234 vdd gnd cell_6t
Xbit_r235_c255 bl_255 br_255 wl_235 vdd gnd cell_6t
Xbit_r236_c255 bl_255 br_255 wl_236 vdd gnd cell_6t
Xbit_r237_c255 bl_255 br_255 wl_237 vdd gnd cell_6t
Xbit_r238_c255 bl_255 br_255 wl_238 vdd gnd cell_6t
Xbit_r239_c255 bl_255 br_255 wl_239 vdd gnd cell_6t
Xbit_r240_c255 bl_255 br_255 wl_240 vdd gnd cell_6t
Xbit_r241_c255 bl_255 br_255 wl_241 vdd gnd cell_6t
Xbit_r242_c255 bl_255 br_255 wl_242 vdd gnd cell_6t
Xbit_r243_c255 bl_255 br_255 wl_243 vdd gnd cell_6t
Xbit_r244_c255 bl_255 br_255 wl_244 vdd gnd cell_6t
Xbit_r245_c255 bl_255 br_255 wl_245 vdd gnd cell_6t
Xbit_r246_c255 bl_255 br_255 wl_246 vdd gnd cell_6t
Xbit_r247_c255 bl_255 br_255 wl_247 vdd gnd cell_6t
Xbit_r248_c255 bl_255 br_255 wl_248 vdd gnd cell_6t
Xbit_r249_c255 bl_255 br_255 wl_249 vdd gnd cell_6t
Xbit_r250_c255 bl_255 br_255 wl_250 vdd gnd cell_6t
Xbit_r251_c255 bl_255 br_255 wl_251 vdd gnd cell_6t
Xbit_r252_c255 bl_255 br_255 wl_252 vdd gnd cell_6t
Xbit_r253_c255 bl_255 br_255 wl_253 vdd gnd cell_6t
Xbit_r254_c255 bl_255 br_255 wl_254 vdd gnd cell_6t
Xbit_r255_c255 bl_255 br_255 wl_255 vdd gnd cell_6t
.ENDS bitcell_array_0

.SUBCKT replica_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 vdd Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 vdd Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q vdd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q vdd vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl vdd gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT dummy_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl_noconn wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br_noconn wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT replica_column_0 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 wl_256 wl_257 wl_258 vdd gnd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* INPUT : wl_131 
* INPUT : wl_132 
* INPUT : wl_133 
* INPUT : wl_134 
* INPUT : wl_135 
* INPUT : wl_136 
* INPUT : wl_137 
* INPUT : wl_138 
* INPUT : wl_139 
* INPUT : wl_140 
* INPUT : wl_141 
* INPUT : wl_142 
* INPUT : wl_143 
* INPUT : wl_144 
* INPUT : wl_145 
* INPUT : wl_146 
* INPUT : wl_147 
* INPUT : wl_148 
* INPUT : wl_149 
* INPUT : wl_150 
* INPUT : wl_151 
* INPUT : wl_152 
* INPUT : wl_153 
* INPUT : wl_154 
* INPUT : wl_155 
* INPUT : wl_156 
* INPUT : wl_157 
* INPUT : wl_158 
* INPUT : wl_159 
* INPUT : wl_160 
* INPUT : wl_161 
* INPUT : wl_162 
* INPUT : wl_163 
* INPUT : wl_164 
* INPUT : wl_165 
* INPUT : wl_166 
* INPUT : wl_167 
* INPUT : wl_168 
* INPUT : wl_169 
* INPUT : wl_170 
* INPUT : wl_171 
* INPUT : wl_172 
* INPUT : wl_173 
* INPUT : wl_174 
* INPUT : wl_175 
* INPUT : wl_176 
* INPUT : wl_177 
* INPUT : wl_178 
* INPUT : wl_179 
* INPUT : wl_180 
* INPUT : wl_181 
* INPUT : wl_182 
* INPUT : wl_183 
* INPUT : wl_184 
* INPUT : wl_185 
* INPUT : wl_186 
* INPUT : wl_187 
* INPUT : wl_188 
* INPUT : wl_189 
* INPUT : wl_190 
* INPUT : wl_191 
* INPUT : wl_192 
* INPUT : wl_193 
* INPUT : wl_194 
* INPUT : wl_195 
* INPUT : wl_196 
* INPUT : wl_197 
* INPUT : wl_198 
* INPUT : wl_199 
* INPUT : wl_200 
* INPUT : wl_201 
* INPUT : wl_202 
* INPUT : wl_203 
* INPUT : wl_204 
* INPUT : wl_205 
* INPUT : wl_206 
* INPUT : wl_207 
* INPUT : wl_208 
* INPUT : wl_209 
* INPUT : wl_210 
* INPUT : wl_211 
* INPUT : wl_212 
* INPUT : wl_213 
* INPUT : wl_214 
* INPUT : wl_215 
* INPUT : wl_216 
* INPUT : wl_217 
* INPUT : wl_218 
* INPUT : wl_219 
* INPUT : wl_220 
* INPUT : wl_221 
* INPUT : wl_222 
* INPUT : wl_223 
* INPUT : wl_224 
* INPUT : wl_225 
* INPUT : wl_226 
* INPUT : wl_227 
* INPUT : wl_228 
* INPUT : wl_229 
* INPUT : wl_230 
* INPUT : wl_231 
* INPUT : wl_232 
* INPUT : wl_233 
* INPUT : wl_234 
* INPUT : wl_235 
* INPUT : wl_236 
* INPUT : wl_237 
* INPUT : wl_238 
* INPUT : wl_239 
* INPUT : wl_240 
* INPUT : wl_241 
* INPUT : wl_242 
* INPUT : wl_243 
* INPUT : wl_244 
* INPUT : wl_245 
* INPUT : wl_246 
* INPUT : wl_247 
* INPUT : wl_248 
* INPUT : wl_249 
* INPUT : wl_250 
* INPUT : wl_251 
* INPUT : wl_252 
* INPUT : wl_253 
* INPUT : wl_254 
* INPUT : wl_255 
* INPUT : wl_256 
* INPUT : wl_257 
* INPUT : wl_258 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xrbc_1 bl_0 br_0 wl_1 vdd gnd replica_cell_6t
Xrbc_2 bl_0 br_0 wl_2 vdd gnd replica_cell_6t
Xrbc_3 bl_0 br_0 wl_3 vdd gnd replica_cell_6t
Xrbc_4 bl_0 br_0 wl_4 vdd gnd replica_cell_6t
Xrbc_5 bl_0 br_0 wl_5 vdd gnd replica_cell_6t
Xrbc_6 bl_0 br_0 wl_6 vdd gnd replica_cell_6t
Xrbc_7 bl_0 br_0 wl_7 vdd gnd replica_cell_6t
Xrbc_8 bl_0 br_0 wl_8 vdd gnd replica_cell_6t
Xrbc_9 bl_0 br_0 wl_9 vdd gnd replica_cell_6t
Xrbc_10 bl_0 br_0 wl_10 vdd gnd replica_cell_6t
Xrbc_11 bl_0 br_0 wl_11 vdd gnd replica_cell_6t
Xrbc_12 bl_0 br_0 wl_12 vdd gnd replica_cell_6t
Xrbc_13 bl_0 br_0 wl_13 vdd gnd replica_cell_6t
Xrbc_14 bl_0 br_0 wl_14 vdd gnd replica_cell_6t
Xrbc_15 bl_0 br_0 wl_15 vdd gnd replica_cell_6t
Xrbc_16 bl_0 br_0 wl_16 vdd gnd replica_cell_6t
Xrbc_17 bl_0 br_0 wl_17 vdd gnd replica_cell_6t
Xrbc_18 bl_0 br_0 wl_18 vdd gnd replica_cell_6t
Xrbc_19 bl_0 br_0 wl_19 vdd gnd replica_cell_6t
Xrbc_20 bl_0 br_0 wl_20 vdd gnd replica_cell_6t
Xrbc_21 bl_0 br_0 wl_21 vdd gnd replica_cell_6t
Xrbc_22 bl_0 br_0 wl_22 vdd gnd replica_cell_6t
Xrbc_23 bl_0 br_0 wl_23 vdd gnd replica_cell_6t
Xrbc_24 bl_0 br_0 wl_24 vdd gnd replica_cell_6t
Xrbc_25 bl_0 br_0 wl_25 vdd gnd replica_cell_6t
Xrbc_26 bl_0 br_0 wl_26 vdd gnd replica_cell_6t
Xrbc_27 bl_0 br_0 wl_27 vdd gnd replica_cell_6t
Xrbc_28 bl_0 br_0 wl_28 vdd gnd replica_cell_6t
Xrbc_29 bl_0 br_0 wl_29 vdd gnd replica_cell_6t
Xrbc_30 bl_0 br_0 wl_30 vdd gnd replica_cell_6t
Xrbc_31 bl_0 br_0 wl_31 vdd gnd replica_cell_6t
Xrbc_32 bl_0 br_0 wl_32 vdd gnd replica_cell_6t
Xrbc_33 bl_0 br_0 wl_33 vdd gnd replica_cell_6t
Xrbc_34 bl_0 br_0 wl_34 vdd gnd replica_cell_6t
Xrbc_35 bl_0 br_0 wl_35 vdd gnd replica_cell_6t
Xrbc_36 bl_0 br_0 wl_36 vdd gnd replica_cell_6t
Xrbc_37 bl_0 br_0 wl_37 vdd gnd replica_cell_6t
Xrbc_38 bl_0 br_0 wl_38 vdd gnd replica_cell_6t
Xrbc_39 bl_0 br_0 wl_39 vdd gnd replica_cell_6t
Xrbc_40 bl_0 br_0 wl_40 vdd gnd replica_cell_6t
Xrbc_41 bl_0 br_0 wl_41 vdd gnd replica_cell_6t
Xrbc_42 bl_0 br_0 wl_42 vdd gnd replica_cell_6t
Xrbc_43 bl_0 br_0 wl_43 vdd gnd replica_cell_6t
Xrbc_44 bl_0 br_0 wl_44 vdd gnd replica_cell_6t
Xrbc_45 bl_0 br_0 wl_45 vdd gnd replica_cell_6t
Xrbc_46 bl_0 br_0 wl_46 vdd gnd replica_cell_6t
Xrbc_47 bl_0 br_0 wl_47 vdd gnd replica_cell_6t
Xrbc_48 bl_0 br_0 wl_48 vdd gnd replica_cell_6t
Xrbc_49 bl_0 br_0 wl_49 vdd gnd replica_cell_6t
Xrbc_50 bl_0 br_0 wl_50 vdd gnd replica_cell_6t
Xrbc_51 bl_0 br_0 wl_51 vdd gnd replica_cell_6t
Xrbc_52 bl_0 br_0 wl_52 vdd gnd replica_cell_6t
Xrbc_53 bl_0 br_0 wl_53 vdd gnd replica_cell_6t
Xrbc_54 bl_0 br_0 wl_54 vdd gnd replica_cell_6t
Xrbc_55 bl_0 br_0 wl_55 vdd gnd replica_cell_6t
Xrbc_56 bl_0 br_0 wl_56 vdd gnd replica_cell_6t
Xrbc_57 bl_0 br_0 wl_57 vdd gnd replica_cell_6t
Xrbc_58 bl_0 br_0 wl_58 vdd gnd replica_cell_6t
Xrbc_59 bl_0 br_0 wl_59 vdd gnd replica_cell_6t
Xrbc_60 bl_0 br_0 wl_60 vdd gnd replica_cell_6t
Xrbc_61 bl_0 br_0 wl_61 vdd gnd replica_cell_6t
Xrbc_62 bl_0 br_0 wl_62 vdd gnd replica_cell_6t
Xrbc_63 bl_0 br_0 wl_63 vdd gnd replica_cell_6t
Xrbc_64 bl_0 br_0 wl_64 vdd gnd replica_cell_6t
Xrbc_65 bl_0 br_0 wl_65 vdd gnd replica_cell_6t
Xrbc_66 bl_0 br_0 wl_66 vdd gnd replica_cell_6t
Xrbc_67 bl_0 br_0 wl_67 vdd gnd replica_cell_6t
Xrbc_68 bl_0 br_0 wl_68 vdd gnd replica_cell_6t
Xrbc_69 bl_0 br_0 wl_69 vdd gnd replica_cell_6t
Xrbc_70 bl_0 br_0 wl_70 vdd gnd replica_cell_6t
Xrbc_71 bl_0 br_0 wl_71 vdd gnd replica_cell_6t
Xrbc_72 bl_0 br_0 wl_72 vdd gnd replica_cell_6t
Xrbc_73 bl_0 br_0 wl_73 vdd gnd replica_cell_6t
Xrbc_74 bl_0 br_0 wl_74 vdd gnd replica_cell_6t
Xrbc_75 bl_0 br_0 wl_75 vdd gnd replica_cell_6t
Xrbc_76 bl_0 br_0 wl_76 vdd gnd replica_cell_6t
Xrbc_77 bl_0 br_0 wl_77 vdd gnd replica_cell_6t
Xrbc_78 bl_0 br_0 wl_78 vdd gnd replica_cell_6t
Xrbc_79 bl_0 br_0 wl_79 vdd gnd replica_cell_6t
Xrbc_80 bl_0 br_0 wl_80 vdd gnd replica_cell_6t
Xrbc_81 bl_0 br_0 wl_81 vdd gnd replica_cell_6t
Xrbc_82 bl_0 br_0 wl_82 vdd gnd replica_cell_6t
Xrbc_83 bl_0 br_0 wl_83 vdd gnd replica_cell_6t
Xrbc_84 bl_0 br_0 wl_84 vdd gnd replica_cell_6t
Xrbc_85 bl_0 br_0 wl_85 vdd gnd replica_cell_6t
Xrbc_86 bl_0 br_0 wl_86 vdd gnd replica_cell_6t
Xrbc_87 bl_0 br_0 wl_87 vdd gnd replica_cell_6t
Xrbc_88 bl_0 br_0 wl_88 vdd gnd replica_cell_6t
Xrbc_89 bl_0 br_0 wl_89 vdd gnd replica_cell_6t
Xrbc_90 bl_0 br_0 wl_90 vdd gnd replica_cell_6t
Xrbc_91 bl_0 br_0 wl_91 vdd gnd replica_cell_6t
Xrbc_92 bl_0 br_0 wl_92 vdd gnd replica_cell_6t
Xrbc_93 bl_0 br_0 wl_93 vdd gnd replica_cell_6t
Xrbc_94 bl_0 br_0 wl_94 vdd gnd replica_cell_6t
Xrbc_95 bl_0 br_0 wl_95 vdd gnd replica_cell_6t
Xrbc_96 bl_0 br_0 wl_96 vdd gnd replica_cell_6t
Xrbc_97 bl_0 br_0 wl_97 vdd gnd replica_cell_6t
Xrbc_98 bl_0 br_0 wl_98 vdd gnd replica_cell_6t
Xrbc_99 bl_0 br_0 wl_99 vdd gnd replica_cell_6t
Xrbc_100 bl_0 br_0 wl_100 vdd gnd replica_cell_6t
Xrbc_101 bl_0 br_0 wl_101 vdd gnd replica_cell_6t
Xrbc_102 bl_0 br_0 wl_102 vdd gnd replica_cell_6t
Xrbc_103 bl_0 br_0 wl_103 vdd gnd replica_cell_6t
Xrbc_104 bl_0 br_0 wl_104 vdd gnd replica_cell_6t
Xrbc_105 bl_0 br_0 wl_105 vdd gnd replica_cell_6t
Xrbc_106 bl_0 br_0 wl_106 vdd gnd replica_cell_6t
Xrbc_107 bl_0 br_0 wl_107 vdd gnd replica_cell_6t
Xrbc_108 bl_0 br_0 wl_108 vdd gnd replica_cell_6t
Xrbc_109 bl_0 br_0 wl_109 vdd gnd replica_cell_6t
Xrbc_110 bl_0 br_0 wl_110 vdd gnd replica_cell_6t
Xrbc_111 bl_0 br_0 wl_111 vdd gnd replica_cell_6t
Xrbc_112 bl_0 br_0 wl_112 vdd gnd replica_cell_6t
Xrbc_113 bl_0 br_0 wl_113 vdd gnd replica_cell_6t
Xrbc_114 bl_0 br_0 wl_114 vdd gnd replica_cell_6t
Xrbc_115 bl_0 br_0 wl_115 vdd gnd replica_cell_6t
Xrbc_116 bl_0 br_0 wl_116 vdd gnd replica_cell_6t
Xrbc_117 bl_0 br_0 wl_117 vdd gnd replica_cell_6t
Xrbc_118 bl_0 br_0 wl_118 vdd gnd replica_cell_6t
Xrbc_119 bl_0 br_0 wl_119 vdd gnd replica_cell_6t
Xrbc_120 bl_0 br_0 wl_120 vdd gnd replica_cell_6t
Xrbc_121 bl_0 br_0 wl_121 vdd gnd replica_cell_6t
Xrbc_122 bl_0 br_0 wl_122 vdd gnd replica_cell_6t
Xrbc_123 bl_0 br_0 wl_123 vdd gnd replica_cell_6t
Xrbc_124 bl_0 br_0 wl_124 vdd gnd replica_cell_6t
Xrbc_125 bl_0 br_0 wl_125 vdd gnd replica_cell_6t
Xrbc_126 bl_0 br_0 wl_126 vdd gnd replica_cell_6t
Xrbc_127 bl_0 br_0 wl_127 vdd gnd replica_cell_6t
Xrbc_128 bl_0 br_0 wl_128 vdd gnd replica_cell_6t
Xrbc_129 bl_0 br_0 wl_129 vdd gnd replica_cell_6t
Xrbc_130 bl_0 br_0 wl_130 vdd gnd replica_cell_6t
Xrbc_131 bl_0 br_0 wl_131 vdd gnd replica_cell_6t
Xrbc_132 bl_0 br_0 wl_132 vdd gnd replica_cell_6t
Xrbc_133 bl_0 br_0 wl_133 vdd gnd replica_cell_6t
Xrbc_134 bl_0 br_0 wl_134 vdd gnd replica_cell_6t
Xrbc_135 bl_0 br_0 wl_135 vdd gnd replica_cell_6t
Xrbc_136 bl_0 br_0 wl_136 vdd gnd replica_cell_6t
Xrbc_137 bl_0 br_0 wl_137 vdd gnd replica_cell_6t
Xrbc_138 bl_0 br_0 wl_138 vdd gnd replica_cell_6t
Xrbc_139 bl_0 br_0 wl_139 vdd gnd replica_cell_6t
Xrbc_140 bl_0 br_0 wl_140 vdd gnd replica_cell_6t
Xrbc_141 bl_0 br_0 wl_141 vdd gnd replica_cell_6t
Xrbc_142 bl_0 br_0 wl_142 vdd gnd replica_cell_6t
Xrbc_143 bl_0 br_0 wl_143 vdd gnd replica_cell_6t
Xrbc_144 bl_0 br_0 wl_144 vdd gnd replica_cell_6t
Xrbc_145 bl_0 br_0 wl_145 vdd gnd replica_cell_6t
Xrbc_146 bl_0 br_0 wl_146 vdd gnd replica_cell_6t
Xrbc_147 bl_0 br_0 wl_147 vdd gnd replica_cell_6t
Xrbc_148 bl_0 br_0 wl_148 vdd gnd replica_cell_6t
Xrbc_149 bl_0 br_0 wl_149 vdd gnd replica_cell_6t
Xrbc_150 bl_0 br_0 wl_150 vdd gnd replica_cell_6t
Xrbc_151 bl_0 br_0 wl_151 vdd gnd replica_cell_6t
Xrbc_152 bl_0 br_0 wl_152 vdd gnd replica_cell_6t
Xrbc_153 bl_0 br_0 wl_153 vdd gnd replica_cell_6t
Xrbc_154 bl_0 br_0 wl_154 vdd gnd replica_cell_6t
Xrbc_155 bl_0 br_0 wl_155 vdd gnd replica_cell_6t
Xrbc_156 bl_0 br_0 wl_156 vdd gnd replica_cell_6t
Xrbc_157 bl_0 br_0 wl_157 vdd gnd replica_cell_6t
Xrbc_158 bl_0 br_0 wl_158 vdd gnd replica_cell_6t
Xrbc_159 bl_0 br_0 wl_159 vdd gnd replica_cell_6t
Xrbc_160 bl_0 br_0 wl_160 vdd gnd replica_cell_6t
Xrbc_161 bl_0 br_0 wl_161 vdd gnd replica_cell_6t
Xrbc_162 bl_0 br_0 wl_162 vdd gnd replica_cell_6t
Xrbc_163 bl_0 br_0 wl_163 vdd gnd replica_cell_6t
Xrbc_164 bl_0 br_0 wl_164 vdd gnd replica_cell_6t
Xrbc_165 bl_0 br_0 wl_165 vdd gnd replica_cell_6t
Xrbc_166 bl_0 br_0 wl_166 vdd gnd replica_cell_6t
Xrbc_167 bl_0 br_0 wl_167 vdd gnd replica_cell_6t
Xrbc_168 bl_0 br_0 wl_168 vdd gnd replica_cell_6t
Xrbc_169 bl_0 br_0 wl_169 vdd gnd replica_cell_6t
Xrbc_170 bl_0 br_0 wl_170 vdd gnd replica_cell_6t
Xrbc_171 bl_0 br_0 wl_171 vdd gnd replica_cell_6t
Xrbc_172 bl_0 br_0 wl_172 vdd gnd replica_cell_6t
Xrbc_173 bl_0 br_0 wl_173 vdd gnd replica_cell_6t
Xrbc_174 bl_0 br_0 wl_174 vdd gnd replica_cell_6t
Xrbc_175 bl_0 br_0 wl_175 vdd gnd replica_cell_6t
Xrbc_176 bl_0 br_0 wl_176 vdd gnd replica_cell_6t
Xrbc_177 bl_0 br_0 wl_177 vdd gnd replica_cell_6t
Xrbc_178 bl_0 br_0 wl_178 vdd gnd replica_cell_6t
Xrbc_179 bl_0 br_0 wl_179 vdd gnd replica_cell_6t
Xrbc_180 bl_0 br_0 wl_180 vdd gnd replica_cell_6t
Xrbc_181 bl_0 br_0 wl_181 vdd gnd replica_cell_6t
Xrbc_182 bl_0 br_0 wl_182 vdd gnd replica_cell_6t
Xrbc_183 bl_0 br_0 wl_183 vdd gnd replica_cell_6t
Xrbc_184 bl_0 br_0 wl_184 vdd gnd replica_cell_6t
Xrbc_185 bl_0 br_0 wl_185 vdd gnd replica_cell_6t
Xrbc_186 bl_0 br_0 wl_186 vdd gnd replica_cell_6t
Xrbc_187 bl_0 br_0 wl_187 vdd gnd replica_cell_6t
Xrbc_188 bl_0 br_0 wl_188 vdd gnd replica_cell_6t
Xrbc_189 bl_0 br_0 wl_189 vdd gnd replica_cell_6t
Xrbc_190 bl_0 br_0 wl_190 vdd gnd replica_cell_6t
Xrbc_191 bl_0 br_0 wl_191 vdd gnd replica_cell_6t
Xrbc_192 bl_0 br_0 wl_192 vdd gnd replica_cell_6t
Xrbc_193 bl_0 br_0 wl_193 vdd gnd replica_cell_6t
Xrbc_194 bl_0 br_0 wl_194 vdd gnd replica_cell_6t
Xrbc_195 bl_0 br_0 wl_195 vdd gnd replica_cell_6t
Xrbc_196 bl_0 br_0 wl_196 vdd gnd replica_cell_6t
Xrbc_197 bl_0 br_0 wl_197 vdd gnd replica_cell_6t
Xrbc_198 bl_0 br_0 wl_198 vdd gnd replica_cell_6t
Xrbc_199 bl_0 br_0 wl_199 vdd gnd replica_cell_6t
Xrbc_200 bl_0 br_0 wl_200 vdd gnd replica_cell_6t
Xrbc_201 bl_0 br_0 wl_201 vdd gnd replica_cell_6t
Xrbc_202 bl_0 br_0 wl_202 vdd gnd replica_cell_6t
Xrbc_203 bl_0 br_0 wl_203 vdd gnd replica_cell_6t
Xrbc_204 bl_0 br_0 wl_204 vdd gnd replica_cell_6t
Xrbc_205 bl_0 br_0 wl_205 vdd gnd replica_cell_6t
Xrbc_206 bl_0 br_0 wl_206 vdd gnd replica_cell_6t
Xrbc_207 bl_0 br_0 wl_207 vdd gnd replica_cell_6t
Xrbc_208 bl_0 br_0 wl_208 vdd gnd replica_cell_6t
Xrbc_209 bl_0 br_0 wl_209 vdd gnd replica_cell_6t
Xrbc_210 bl_0 br_0 wl_210 vdd gnd replica_cell_6t
Xrbc_211 bl_0 br_0 wl_211 vdd gnd replica_cell_6t
Xrbc_212 bl_0 br_0 wl_212 vdd gnd replica_cell_6t
Xrbc_213 bl_0 br_0 wl_213 vdd gnd replica_cell_6t
Xrbc_214 bl_0 br_0 wl_214 vdd gnd replica_cell_6t
Xrbc_215 bl_0 br_0 wl_215 vdd gnd replica_cell_6t
Xrbc_216 bl_0 br_0 wl_216 vdd gnd replica_cell_6t
Xrbc_217 bl_0 br_0 wl_217 vdd gnd replica_cell_6t
Xrbc_218 bl_0 br_0 wl_218 vdd gnd replica_cell_6t
Xrbc_219 bl_0 br_0 wl_219 vdd gnd replica_cell_6t
Xrbc_220 bl_0 br_0 wl_220 vdd gnd replica_cell_6t
Xrbc_221 bl_0 br_0 wl_221 vdd gnd replica_cell_6t
Xrbc_222 bl_0 br_0 wl_222 vdd gnd replica_cell_6t
Xrbc_223 bl_0 br_0 wl_223 vdd gnd replica_cell_6t
Xrbc_224 bl_0 br_0 wl_224 vdd gnd replica_cell_6t
Xrbc_225 bl_0 br_0 wl_225 vdd gnd replica_cell_6t
Xrbc_226 bl_0 br_0 wl_226 vdd gnd replica_cell_6t
Xrbc_227 bl_0 br_0 wl_227 vdd gnd replica_cell_6t
Xrbc_228 bl_0 br_0 wl_228 vdd gnd replica_cell_6t
Xrbc_229 bl_0 br_0 wl_229 vdd gnd replica_cell_6t
Xrbc_230 bl_0 br_0 wl_230 vdd gnd replica_cell_6t
Xrbc_231 bl_0 br_0 wl_231 vdd gnd replica_cell_6t
Xrbc_232 bl_0 br_0 wl_232 vdd gnd replica_cell_6t
Xrbc_233 bl_0 br_0 wl_233 vdd gnd replica_cell_6t
Xrbc_234 bl_0 br_0 wl_234 vdd gnd replica_cell_6t
Xrbc_235 bl_0 br_0 wl_235 vdd gnd replica_cell_6t
Xrbc_236 bl_0 br_0 wl_236 vdd gnd replica_cell_6t
Xrbc_237 bl_0 br_0 wl_237 vdd gnd replica_cell_6t
Xrbc_238 bl_0 br_0 wl_238 vdd gnd replica_cell_6t
Xrbc_239 bl_0 br_0 wl_239 vdd gnd replica_cell_6t
Xrbc_240 bl_0 br_0 wl_240 vdd gnd replica_cell_6t
Xrbc_241 bl_0 br_0 wl_241 vdd gnd replica_cell_6t
Xrbc_242 bl_0 br_0 wl_242 vdd gnd replica_cell_6t
Xrbc_243 bl_0 br_0 wl_243 vdd gnd replica_cell_6t
Xrbc_244 bl_0 br_0 wl_244 vdd gnd replica_cell_6t
Xrbc_245 bl_0 br_0 wl_245 vdd gnd replica_cell_6t
Xrbc_246 bl_0 br_0 wl_246 vdd gnd replica_cell_6t
Xrbc_247 bl_0 br_0 wl_247 vdd gnd replica_cell_6t
Xrbc_248 bl_0 br_0 wl_248 vdd gnd replica_cell_6t
Xrbc_249 bl_0 br_0 wl_249 vdd gnd replica_cell_6t
Xrbc_250 bl_0 br_0 wl_250 vdd gnd replica_cell_6t
Xrbc_251 bl_0 br_0 wl_251 vdd gnd replica_cell_6t
Xrbc_252 bl_0 br_0 wl_252 vdd gnd replica_cell_6t
Xrbc_253 bl_0 br_0 wl_253 vdd gnd replica_cell_6t
Xrbc_254 bl_0 br_0 wl_254 vdd gnd replica_cell_6t
Xrbc_255 bl_0 br_0 wl_255 vdd gnd replica_cell_6t
Xrbc_256 bl_0 br_0 wl_256 vdd gnd replica_cell_6t
Xrbc_257 bl_0 br_0 wl_257 vdd gnd replica_cell_6t
Xrbc_258 bl_0 br_0 wl_258 vdd gnd dummy_cell_6t
.ENDS replica_column_0

.SUBCKT dummy_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd dummy_cell_6t
.ENDS dummy_array_0

.SUBCKT dummy_array_1 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 wl_256 wl_257 wl_258 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* INPUT : wl_131 
* INPUT : wl_132 
* INPUT : wl_133 
* INPUT : wl_134 
* INPUT : wl_135 
* INPUT : wl_136 
* INPUT : wl_137 
* INPUT : wl_138 
* INPUT : wl_139 
* INPUT : wl_140 
* INPUT : wl_141 
* INPUT : wl_142 
* INPUT : wl_143 
* INPUT : wl_144 
* INPUT : wl_145 
* INPUT : wl_146 
* INPUT : wl_147 
* INPUT : wl_148 
* INPUT : wl_149 
* INPUT : wl_150 
* INPUT : wl_151 
* INPUT : wl_152 
* INPUT : wl_153 
* INPUT : wl_154 
* INPUT : wl_155 
* INPUT : wl_156 
* INPUT : wl_157 
* INPUT : wl_158 
* INPUT : wl_159 
* INPUT : wl_160 
* INPUT : wl_161 
* INPUT : wl_162 
* INPUT : wl_163 
* INPUT : wl_164 
* INPUT : wl_165 
* INPUT : wl_166 
* INPUT : wl_167 
* INPUT : wl_168 
* INPUT : wl_169 
* INPUT : wl_170 
* INPUT : wl_171 
* INPUT : wl_172 
* INPUT : wl_173 
* INPUT : wl_174 
* INPUT : wl_175 
* INPUT : wl_176 
* INPUT : wl_177 
* INPUT : wl_178 
* INPUT : wl_179 
* INPUT : wl_180 
* INPUT : wl_181 
* INPUT : wl_182 
* INPUT : wl_183 
* INPUT : wl_184 
* INPUT : wl_185 
* INPUT : wl_186 
* INPUT : wl_187 
* INPUT : wl_188 
* INPUT : wl_189 
* INPUT : wl_190 
* INPUT : wl_191 
* INPUT : wl_192 
* INPUT : wl_193 
* INPUT : wl_194 
* INPUT : wl_195 
* INPUT : wl_196 
* INPUT : wl_197 
* INPUT : wl_198 
* INPUT : wl_199 
* INPUT : wl_200 
* INPUT : wl_201 
* INPUT : wl_202 
* INPUT : wl_203 
* INPUT : wl_204 
* INPUT : wl_205 
* INPUT : wl_206 
* INPUT : wl_207 
* INPUT : wl_208 
* INPUT : wl_209 
* INPUT : wl_210 
* INPUT : wl_211 
* INPUT : wl_212 
* INPUT : wl_213 
* INPUT : wl_214 
* INPUT : wl_215 
* INPUT : wl_216 
* INPUT : wl_217 
* INPUT : wl_218 
* INPUT : wl_219 
* INPUT : wl_220 
* INPUT : wl_221 
* INPUT : wl_222 
* INPUT : wl_223 
* INPUT : wl_224 
* INPUT : wl_225 
* INPUT : wl_226 
* INPUT : wl_227 
* INPUT : wl_228 
* INPUT : wl_229 
* INPUT : wl_230 
* INPUT : wl_231 
* INPUT : wl_232 
* INPUT : wl_233 
* INPUT : wl_234 
* INPUT : wl_235 
* INPUT : wl_236 
* INPUT : wl_237 
* INPUT : wl_238 
* INPUT : wl_239 
* INPUT : wl_240 
* INPUT : wl_241 
* INPUT : wl_242 
* INPUT : wl_243 
* INPUT : wl_244 
* INPUT : wl_245 
* INPUT : wl_246 
* INPUT : wl_247 
* INPUT : wl_248 
* INPUT : wl_249 
* INPUT : wl_250 
* INPUT : wl_251 
* INPUT : wl_252 
* INPUT : wl_253 
* INPUT : wl_254 
* INPUT : wl_255 
* INPUT : wl_256 
* INPUT : wl_257 
* INPUT : wl_258 
* POWER : vdd 
* GROUND: gnd 
* rows: 259 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd dummy_cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd dummy_cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd dummy_cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd dummy_cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd dummy_cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd dummy_cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd dummy_cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd dummy_cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd dummy_cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd dummy_cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd dummy_cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd dummy_cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd dummy_cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd dummy_cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd dummy_cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd dummy_cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd dummy_cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd dummy_cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd dummy_cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd dummy_cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd dummy_cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd dummy_cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd dummy_cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd dummy_cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd dummy_cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd dummy_cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd dummy_cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd dummy_cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd dummy_cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd dummy_cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd dummy_cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd dummy_cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd dummy_cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd dummy_cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd dummy_cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd dummy_cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd dummy_cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd dummy_cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd dummy_cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd dummy_cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd dummy_cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd dummy_cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd dummy_cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd dummy_cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd dummy_cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd dummy_cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd dummy_cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd dummy_cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd dummy_cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd dummy_cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd dummy_cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd dummy_cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd dummy_cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd dummy_cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd dummy_cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd dummy_cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd dummy_cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd dummy_cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd dummy_cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd dummy_cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd dummy_cell_6t
Xbit_r128_c0 bl_0 br_0 wl_128 vdd gnd dummy_cell_6t
Xbit_r129_c0 bl_0 br_0 wl_129 vdd gnd dummy_cell_6t
Xbit_r130_c0 bl_0 br_0 wl_130 vdd gnd dummy_cell_6t
Xbit_r131_c0 bl_0 br_0 wl_131 vdd gnd dummy_cell_6t
Xbit_r132_c0 bl_0 br_0 wl_132 vdd gnd dummy_cell_6t
Xbit_r133_c0 bl_0 br_0 wl_133 vdd gnd dummy_cell_6t
Xbit_r134_c0 bl_0 br_0 wl_134 vdd gnd dummy_cell_6t
Xbit_r135_c0 bl_0 br_0 wl_135 vdd gnd dummy_cell_6t
Xbit_r136_c0 bl_0 br_0 wl_136 vdd gnd dummy_cell_6t
Xbit_r137_c0 bl_0 br_0 wl_137 vdd gnd dummy_cell_6t
Xbit_r138_c0 bl_0 br_0 wl_138 vdd gnd dummy_cell_6t
Xbit_r139_c0 bl_0 br_0 wl_139 vdd gnd dummy_cell_6t
Xbit_r140_c0 bl_0 br_0 wl_140 vdd gnd dummy_cell_6t
Xbit_r141_c0 bl_0 br_0 wl_141 vdd gnd dummy_cell_6t
Xbit_r142_c0 bl_0 br_0 wl_142 vdd gnd dummy_cell_6t
Xbit_r143_c0 bl_0 br_0 wl_143 vdd gnd dummy_cell_6t
Xbit_r144_c0 bl_0 br_0 wl_144 vdd gnd dummy_cell_6t
Xbit_r145_c0 bl_0 br_0 wl_145 vdd gnd dummy_cell_6t
Xbit_r146_c0 bl_0 br_0 wl_146 vdd gnd dummy_cell_6t
Xbit_r147_c0 bl_0 br_0 wl_147 vdd gnd dummy_cell_6t
Xbit_r148_c0 bl_0 br_0 wl_148 vdd gnd dummy_cell_6t
Xbit_r149_c0 bl_0 br_0 wl_149 vdd gnd dummy_cell_6t
Xbit_r150_c0 bl_0 br_0 wl_150 vdd gnd dummy_cell_6t
Xbit_r151_c0 bl_0 br_0 wl_151 vdd gnd dummy_cell_6t
Xbit_r152_c0 bl_0 br_0 wl_152 vdd gnd dummy_cell_6t
Xbit_r153_c0 bl_0 br_0 wl_153 vdd gnd dummy_cell_6t
Xbit_r154_c0 bl_0 br_0 wl_154 vdd gnd dummy_cell_6t
Xbit_r155_c0 bl_0 br_0 wl_155 vdd gnd dummy_cell_6t
Xbit_r156_c0 bl_0 br_0 wl_156 vdd gnd dummy_cell_6t
Xbit_r157_c0 bl_0 br_0 wl_157 vdd gnd dummy_cell_6t
Xbit_r158_c0 bl_0 br_0 wl_158 vdd gnd dummy_cell_6t
Xbit_r159_c0 bl_0 br_0 wl_159 vdd gnd dummy_cell_6t
Xbit_r160_c0 bl_0 br_0 wl_160 vdd gnd dummy_cell_6t
Xbit_r161_c0 bl_0 br_0 wl_161 vdd gnd dummy_cell_6t
Xbit_r162_c0 bl_0 br_0 wl_162 vdd gnd dummy_cell_6t
Xbit_r163_c0 bl_0 br_0 wl_163 vdd gnd dummy_cell_6t
Xbit_r164_c0 bl_0 br_0 wl_164 vdd gnd dummy_cell_6t
Xbit_r165_c0 bl_0 br_0 wl_165 vdd gnd dummy_cell_6t
Xbit_r166_c0 bl_0 br_0 wl_166 vdd gnd dummy_cell_6t
Xbit_r167_c0 bl_0 br_0 wl_167 vdd gnd dummy_cell_6t
Xbit_r168_c0 bl_0 br_0 wl_168 vdd gnd dummy_cell_6t
Xbit_r169_c0 bl_0 br_0 wl_169 vdd gnd dummy_cell_6t
Xbit_r170_c0 bl_0 br_0 wl_170 vdd gnd dummy_cell_6t
Xbit_r171_c0 bl_0 br_0 wl_171 vdd gnd dummy_cell_6t
Xbit_r172_c0 bl_0 br_0 wl_172 vdd gnd dummy_cell_6t
Xbit_r173_c0 bl_0 br_0 wl_173 vdd gnd dummy_cell_6t
Xbit_r174_c0 bl_0 br_0 wl_174 vdd gnd dummy_cell_6t
Xbit_r175_c0 bl_0 br_0 wl_175 vdd gnd dummy_cell_6t
Xbit_r176_c0 bl_0 br_0 wl_176 vdd gnd dummy_cell_6t
Xbit_r177_c0 bl_0 br_0 wl_177 vdd gnd dummy_cell_6t
Xbit_r178_c0 bl_0 br_0 wl_178 vdd gnd dummy_cell_6t
Xbit_r179_c0 bl_0 br_0 wl_179 vdd gnd dummy_cell_6t
Xbit_r180_c0 bl_0 br_0 wl_180 vdd gnd dummy_cell_6t
Xbit_r181_c0 bl_0 br_0 wl_181 vdd gnd dummy_cell_6t
Xbit_r182_c0 bl_0 br_0 wl_182 vdd gnd dummy_cell_6t
Xbit_r183_c0 bl_0 br_0 wl_183 vdd gnd dummy_cell_6t
Xbit_r184_c0 bl_0 br_0 wl_184 vdd gnd dummy_cell_6t
Xbit_r185_c0 bl_0 br_0 wl_185 vdd gnd dummy_cell_6t
Xbit_r186_c0 bl_0 br_0 wl_186 vdd gnd dummy_cell_6t
Xbit_r187_c0 bl_0 br_0 wl_187 vdd gnd dummy_cell_6t
Xbit_r188_c0 bl_0 br_0 wl_188 vdd gnd dummy_cell_6t
Xbit_r189_c0 bl_0 br_0 wl_189 vdd gnd dummy_cell_6t
Xbit_r190_c0 bl_0 br_0 wl_190 vdd gnd dummy_cell_6t
Xbit_r191_c0 bl_0 br_0 wl_191 vdd gnd dummy_cell_6t
Xbit_r192_c0 bl_0 br_0 wl_192 vdd gnd dummy_cell_6t
Xbit_r193_c0 bl_0 br_0 wl_193 vdd gnd dummy_cell_6t
Xbit_r194_c0 bl_0 br_0 wl_194 vdd gnd dummy_cell_6t
Xbit_r195_c0 bl_0 br_0 wl_195 vdd gnd dummy_cell_6t
Xbit_r196_c0 bl_0 br_0 wl_196 vdd gnd dummy_cell_6t
Xbit_r197_c0 bl_0 br_0 wl_197 vdd gnd dummy_cell_6t
Xbit_r198_c0 bl_0 br_0 wl_198 vdd gnd dummy_cell_6t
Xbit_r199_c0 bl_0 br_0 wl_199 vdd gnd dummy_cell_6t
Xbit_r200_c0 bl_0 br_0 wl_200 vdd gnd dummy_cell_6t
Xbit_r201_c0 bl_0 br_0 wl_201 vdd gnd dummy_cell_6t
Xbit_r202_c0 bl_0 br_0 wl_202 vdd gnd dummy_cell_6t
Xbit_r203_c0 bl_0 br_0 wl_203 vdd gnd dummy_cell_6t
Xbit_r204_c0 bl_0 br_0 wl_204 vdd gnd dummy_cell_6t
Xbit_r205_c0 bl_0 br_0 wl_205 vdd gnd dummy_cell_6t
Xbit_r206_c0 bl_0 br_0 wl_206 vdd gnd dummy_cell_6t
Xbit_r207_c0 bl_0 br_0 wl_207 vdd gnd dummy_cell_6t
Xbit_r208_c0 bl_0 br_0 wl_208 vdd gnd dummy_cell_6t
Xbit_r209_c0 bl_0 br_0 wl_209 vdd gnd dummy_cell_6t
Xbit_r210_c0 bl_0 br_0 wl_210 vdd gnd dummy_cell_6t
Xbit_r211_c0 bl_0 br_0 wl_211 vdd gnd dummy_cell_6t
Xbit_r212_c0 bl_0 br_0 wl_212 vdd gnd dummy_cell_6t
Xbit_r213_c0 bl_0 br_0 wl_213 vdd gnd dummy_cell_6t
Xbit_r214_c0 bl_0 br_0 wl_214 vdd gnd dummy_cell_6t
Xbit_r215_c0 bl_0 br_0 wl_215 vdd gnd dummy_cell_6t
Xbit_r216_c0 bl_0 br_0 wl_216 vdd gnd dummy_cell_6t
Xbit_r217_c0 bl_0 br_0 wl_217 vdd gnd dummy_cell_6t
Xbit_r218_c0 bl_0 br_0 wl_218 vdd gnd dummy_cell_6t
Xbit_r219_c0 bl_0 br_0 wl_219 vdd gnd dummy_cell_6t
Xbit_r220_c0 bl_0 br_0 wl_220 vdd gnd dummy_cell_6t
Xbit_r221_c0 bl_0 br_0 wl_221 vdd gnd dummy_cell_6t
Xbit_r222_c0 bl_0 br_0 wl_222 vdd gnd dummy_cell_6t
Xbit_r223_c0 bl_0 br_0 wl_223 vdd gnd dummy_cell_6t
Xbit_r224_c0 bl_0 br_0 wl_224 vdd gnd dummy_cell_6t
Xbit_r225_c0 bl_0 br_0 wl_225 vdd gnd dummy_cell_6t
Xbit_r226_c0 bl_0 br_0 wl_226 vdd gnd dummy_cell_6t
Xbit_r227_c0 bl_0 br_0 wl_227 vdd gnd dummy_cell_6t
Xbit_r228_c0 bl_0 br_0 wl_228 vdd gnd dummy_cell_6t
Xbit_r229_c0 bl_0 br_0 wl_229 vdd gnd dummy_cell_6t
Xbit_r230_c0 bl_0 br_0 wl_230 vdd gnd dummy_cell_6t
Xbit_r231_c0 bl_0 br_0 wl_231 vdd gnd dummy_cell_6t
Xbit_r232_c0 bl_0 br_0 wl_232 vdd gnd dummy_cell_6t
Xbit_r233_c0 bl_0 br_0 wl_233 vdd gnd dummy_cell_6t
Xbit_r234_c0 bl_0 br_0 wl_234 vdd gnd dummy_cell_6t
Xbit_r235_c0 bl_0 br_0 wl_235 vdd gnd dummy_cell_6t
Xbit_r236_c0 bl_0 br_0 wl_236 vdd gnd dummy_cell_6t
Xbit_r237_c0 bl_0 br_0 wl_237 vdd gnd dummy_cell_6t
Xbit_r238_c0 bl_0 br_0 wl_238 vdd gnd dummy_cell_6t
Xbit_r239_c0 bl_0 br_0 wl_239 vdd gnd dummy_cell_6t
Xbit_r240_c0 bl_0 br_0 wl_240 vdd gnd dummy_cell_6t
Xbit_r241_c0 bl_0 br_0 wl_241 vdd gnd dummy_cell_6t
Xbit_r242_c0 bl_0 br_0 wl_242 vdd gnd dummy_cell_6t
Xbit_r243_c0 bl_0 br_0 wl_243 vdd gnd dummy_cell_6t
Xbit_r244_c0 bl_0 br_0 wl_244 vdd gnd dummy_cell_6t
Xbit_r245_c0 bl_0 br_0 wl_245 vdd gnd dummy_cell_6t
Xbit_r246_c0 bl_0 br_0 wl_246 vdd gnd dummy_cell_6t
Xbit_r247_c0 bl_0 br_0 wl_247 vdd gnd dummy_cell_6t
Xbit_r248_c0 bl_0 br_0 wl_248 vdd gnd dummy_cell_6t
Xbit_r249_c0 bl_0 br_0 wl_249 vdd gnd dummy_cell_6t
Xbit_r250_c0 bl_0 br_0 wl_250 vdd gnd dummy_cell_6t
Xbit_r251_c0 bl_0 br_0 wl_251 vdd gnd dummy_cell_6t
Xbit_r252_c0 bl_0 br_0 wl_252 vdd gnd dummy_cell_6t
Xbit_r253_c0 bl_0 br_0 wl_253 vdd gnd dummy_cell_6t
Xbit_r254_c0 bl_0 br_0 wl_254 vdd gnd dummy_cell_6t
Xbit_r255_c0 bl_0 br_0 wl_255 vdd gnd dummy_cell_6t
Xbit_r256_c0 bl_0 br_0 wl_256 vdd gnd dummy_cell_6t
Xbit_r257_c0 bl_0 br_0 wl_257 vdd gnd dummy_cell_6t
Xbit_r258_c0 bl_0 br_0 wl_258 vdd gnd dummy_cell_6t
.ENDS dummy_array_1

.SUBCKT dummy_array_2 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 wl_256 wl_257 wl_258 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* INPUT : wl_131 
* INPUT : wl_132 
* INPUT : wl_133 
* INPUT : wl_134 
* INPUT : wl_135 
* INPUT : wl_136 
* INPUT : wl_137 
* INPUT : wl_138 
* INPUT : wl_139 
* INPUT : wl_140 
* INPUT : wl_141 
* INPUT : wl_142 
* INPUT : wl_143 
* INPUT : wl_144 
* INPUT : wl_145 
* INPUT : wl_146 
* INPUT : wl_147 
* INPUT : wl_148 
* INPUT : wl_149 
* INPUT : wl_150 
* INPUT : wl_151 
* INPUT : wl_152 
* INPUT : wl_153 
* INPUT : wl_154 
* INPUT : wl_155 
* INPUT : wl_156 
* INPUT : wl_157 
* INPUT : wl_158 
* INPUT : wl_159 
* INPUT : wl_160 
* INPUT : wl_161 
* INPUT : wl_162 
* INPUT : wl_163 
* INPUT : wl_164 
* INPUT : wl_165 
* INPUT : wl_166 
* INPUT : wl_167 
* INPUT : wl_168 
* INPUT : wl_169 
* INPUT : wl_170 
* INPUT : wl_171 
* INPUT : wl_172 
* INPUT : wl_173 
* INPUT : wl_174 
* INPUT : wl_175 
* INPUT : wl_176 
* INPUT : wl_177 
* INPUT : wl_178 
* INPUT : wl_179 
* INPUT : wl_180 
* INPUT : wl_181 
* INPUT : wl_182 
* INPUT : wl_183 
* INPUT : wl_184 
* INPUT : wl_185 
* INPUT : wl_186 
* INPUT : wl_187 
* INPUT : wl_188 
* INPUT : wl_189 
* INPUT : wl_190 
* INPUT : wl_191 
* INPUT : wl_192 
* INPUT : wl_193 
* INPUT : wl_194 
* INPUT : wl_195 
* INPUT : wl_196 
* INPUT : wl_197 
* INPUT : wl_198 
* INPUT : wl_199 
* INPUT : wl_200 
* INPUT : wl_201 
* INPUT : wl_202 
* INPUT : wl_203 
* INPUT : wl_204 
* INPUT : wl_205 
* INPUT : wl_206 
* INPUT : wl_207 
* INPUT : wl_208 
* INPUT : wl_209 
* INPUT : wl_210 
* INPUT : wl_211 
* INPUT : wl_212 
* INPUT : wl_213 
* INPUT : wl_214 
* INPUT : wl_215 
* INPUT : wl_216 
* INPUT : wl_217 
* INPUT : wl_218 
* INPUT : wl_219 
* INPUT : wl_220 
* INPUT : wl_221 
* INPUT : wl_222 
* INPUT : wl_223 
* INPUT : wl_224 
* INPUT : wl_225 
* INPUT : wl_226 
* INPUT : wl_227 
* INPUT : wl_228 
* INPUT : wl_229 
* INPUT : wl_230 
* INPUT : wl_231 
* INPUT : wl_232 
* INPUT : wl_233 
* INPUT : wl_234 
* INPUT : wl_235 
* INPUT : wl_236 
* INPUT : wl_237 
* INPUT : wl_238 
* INPUT : wl_239 
* INPUT : wl_240 
* INPUT : wl_241 
* INPUT : wl_242 
* INPUT : wl_243 
* INPUT : wl_244 
* INPUT : wl_245 
* INPUT : wl_246 
* INPUT : wl_247 
* INPUT : wl_248 
* INPUT : wl_249 
* INPUT : wl_250 
* INPUT : wl_251 
* INPUT : wl_252 
* INPUT : wl_253 
* INPUT : wl_254 
* INPUT : wl_255 
* INPUT : wl_256 
* INPUT : wl_257 
* INPUT : wl_258 
* POWER : vdd 
* GROUND: gnd 
* rows: 259 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd dummy_cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd dummy_cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd dummy_cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd dummy_cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd dummy_cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd dummy_cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd dummy_cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd dummy_cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd dummy_cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd dummy_cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd dummy_cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd dummy_cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd dummy_cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd dummy_cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd dummy_cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd dummy_cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd dummy_cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd dummy_cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd dummy_cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd dummy_cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd dummy_cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd dummy_cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd dummy_cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd dummy_cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd dummy_cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd dummy_cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd dummy_cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd dummy_cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd dummy_cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd dummy_cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd dummy_cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd dummy_cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd dummy_cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd dummy_cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd dummy_cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd dummy_cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd dummy_cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd dummy_cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd dummy_cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd dummy_cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd dummy_cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd dummy_cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd dummy_cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd dummy_cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd dummy_cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd dummy_cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd dummy_cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd dummy_cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd dummy_cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd dummy_cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd dummy_cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd dummy_cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd dummy_cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd dummy_cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd dummy_cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd dummy_cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd dummy_cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd dummy_cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd dummy_cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd dummy_cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd dummy_cell_6t
Xbit_r128_c0 bl_0 br_0 wl_128 vdd gnd dummy_cell_6t
Xbit_r129_c0 bl_0 br_0 wl_129 vdd gnd dummy_cell_6t
Xbit_r130_c0 bl_0 br_0 wl_130 vdd gnd dummy_cell_6t
Xbit_r131_c0 bl_0 br_0 wl_131 vdd gnd dummy_cell_6t
Xbit_r132_c0 bl_0 br_0 wl_132 vdd gnd dummy_cell_6t
Xbit_r133_c0 bl_0 br_0 wl_133 vdd gnd dummy_cell_6t
Xbit_r134_c0 bl_0 br_0 wl_134 vdd gnd dummy_cell_6t
Xbit_r135_c0 bl_0 br_0 wl_135 vdd gnd dummy_cell_6t
Xbit_r136_c0 bl_0 br_0 wl_136 vdd gnd dummy_cell_6t
Xbit_r137_c0 bl_0 br_0 wl_137 vdd gnd dummy_cell_6t
Xbit_r138_c0 bl_0 br_0 wl_138 vdd gnd dummy_cell_6t
Xbit_r139_c0 bl_0 br_0 wl_139 vdd gnd dummy_cell_6t
Xbit_r140_c0 bl_0 br_0 wl_140 vdd gnd dummy_cell_6t
Xbit_r141_c0 bl_0 br_0 wl_141 vdd gnd dummy_cell_6t
Xbit_r142_c0 bl_0 br_0 wl_142 vdd gnd dummy_cell_6t
Xbit_r143_c0 bl_0 br_0 wl_143 vdd gnd dummy_cell_6t
Xbit_r144_c0 bl_0 br_0 wl_144 vdd gnd dummy_cell_6t
Xbit_r145_c0 bl_0 br_0 wl_145 vdd gnd dummy_cell_6t
Xbit_r146_c0 bl_0 br_0 wl_146 vdd gnd dummy_cell_6t
Xbit_r147_c0 bl_0 br_0 wl_147 vdd gnd dummy_cell_6t
Xbit_r148_c0 bl_0 br_0 wl_148 vdd gnd dummy_cell_6t
Xbit_r149_c0 bl_0 br_0 wl_149 vdd gnd dummy_cell_6t
Xbit_r150_c0 bl_0 br_0 wl_150 vdd gnd dummy_cell_6t
Xbit_r151_c0 bl_0 br_0 wl_151 vdd gnd dummy_cell_6t
Xbit_r152_c0 bl_0 br_0 wl_152 vdd gnd dummy_cell_6t
Xbit_r153_c0 bl_0 br_0 wl_153 vdd gnd dummy_cell_6t
Xbit_r154_c0 bl_0 br_0 wl_154 vdd gnd dummy_cell_6t
Xbit_r155_c0 bl_0 br_0 wl_155 vdd gnd dummy_cell_6t
Xbit_r156_c0 bl_0 br_0 wl_156 vdd gnd dummy_cell_6t
Xbit_r157_c0 bl_0 br_0 wl_157 vdd gnd dummy_cell_6t
Xbit_r158_c0 bl_0 br_0 wl_158 vdd gnd dummy_cell_6t
Xbit_r159_c0 bl_0 br_0 wl_159 vdd gnd dummy_cell_6t
Xbit_r160_c0 bl_0 br_0 wl_160 vdd gnd dummy_cell_6t
Xbit_r161_c0 bl_0 br_0 wl_161 vdd gnd dummy_cell_6t
Xbit_r162_c0 bl_0 br_0 wl_162 vdd gnd dummy_cell_6t
Xbit_r163_c0 bl_0 br_0 wl_163 vdd gnd dummy_cell_6t
Xbit_r164_c0 bl_0 br_0 wl_164 vdd gnd dummy_cell_6t
Xbit_r165_c0 bl_0 br_0 wl_165 vdd gnd dummy_cell_6t
Xbit_r166_c0 bl_0 br_0 wl_166 vdd gnd dummy_cell_6t
Xbit_r167_c0 bl_0 br_0 wl_167 vdd gnd dummy_cell_6t
Xbit_r168_c0 bl_0 br_0 wl_168 vdd gnd dummy_cell_6t
Xbit_r169_c0 bl_0 br_0 wl_169 vdd gnd dummy_cell_6t
Xbit_r170_c0 bl_0 br_0 wl_170 vdd gnd dummy_cell_6t
Xbit_r171_c0 bl_0 br_0 wl_171 vdd gnd dummy_cell_6t
Xbit_r172_c0 bl_0 br_0 wl_172 vdd gnd dummy_cell_6t
Xbit_r173_c0 bl_0 br_0 wl_173 vdd gnd dummy_cell_6t
Xbit_r174_c0 bl_0 br_0 wl_174 vdd gnd dummy_cell_6t
Xbit_r175_c0 bl_0 br_0 wl_175 vdd gnd dummy_cell_6t
Xbit_r176_c0 bl_0 br_0 wl_176 vdd gnd dummy_cell_6t
Xbit_r177_c0 bl_0 br_0 wl_177 vdd gnd dummy_cell_6t
Xbit_r178_c0 bl_0 br_0 wl_178 vdd gnd dummy_cell_6t
Xbit_r179_c0 bl_0 br_0 wl_179 vdd gnd dummy_cell_6t
Xbit_r180_c0 bl_0 br_0 wl_180 vdd gnd dummy_cell_6t
Xbit_r181_c0 bl_0 br_0 wl_181 vdd gnd dummy_cell_6t
Xbit_r182_c0 bl_0 br_0 wl_182 vdd gnd dummy_cell_6t
Xbit_r183_c0 bl_0 br_0 wl_183 vdd gnd dummy_cell_6t
Xbit_r184_c0 bl_0 br_0 wl_184 vdd gnd dummy_cell_6t
Xbit_r185_c0 bl_0 br_0 wl_185 vdd gnd dummy_cell_6t
Xbit_r186_c0 bl_0 br_0 wl_186 vdd gnd dummy_cell_6t
Xbit_r187_c0 bl_0 br_0 wl_187 vdd gnd dummy_cell_6t
Xbit_r188_c0 bl_0 br_0 wl_188 vdd gnd dummy_cell_6t
Xbit_r189_c0 bl_0 br_0 wl_189 vdd gnd dummy_cell_6t
Xbit_r190_c0 bl_0 br_0 wl_190 vdd gnd dummy_cell_6t
Xbit_r191_c0 bl_0 br_0 wl_191 vdd gnd dummy_cell_6t
Xbit_r192_c0 bl_0 br_0 wl_192 vdd gnd dummy_cell_6t
Xbit_r193_c0 bl_0 br_0 wl_193 vdd gnd dummy_cell_6t
Xbit_r194_c0 bl_0 br_0 wl_194 vdd gnd dummy_cell_6t
Xbit_r195_c0 bl_0 br_0 wl_195 vdd gnd dummy_cell_6t
Xbit_r196_c0 bl_0 br_0 wl_196 vdd gnd dummy_cell_6t
Xbit_r197_c0 bl_0 br_0 wl_197 vdd gnd dummy_cell_6t
Xbit_r198_c0 bl_0 br_0 wl_198 vdd gnd dummy_cell_6t
Xbit_r199_c0 bl_0 br_0 wl_199 vdd gnd dummy_cell_6t
Xbit_r200_c0 bl_0 br_0 wl_200 vdd gnd dummy_cell_6t
Xbit_r201_c0 bl_0 br_0 wl_201 vdd gnd dummy_cell_6t
Xbit_r202_c0 bl_0 br_0 wl_202 vdd gnd dummy_cell_6t
Xbit_r203_c0 bl_0 br_0 wl_203 vdd gnd dummy_cell_6t
Xbit_r204_c0 bl_0 br_0 wl_204 vdd gnd dummy_cell_6t
Xbit_r205_c0 bl_0 br_0 wl_205 vdd gnd dummy_cell_6t
Xbit_r206_c0 bl_0 br_0 wl_206 vdd gnd dummy_cell_6t
Xbit_r207_c0 bl_0 br_0 wl_207 vdd gnd dummy_cell_6t
Xbit_r208_c0 bl_0 br_0 wl_208 vdd gnd dummy_cell_6t
Xbit_r209_c0 bl_0 br_0 wl_209 vdd gnd dummy_cell_6t
Xbit_r210_c0 bl_0 br_0 wl_210 vdd gnd dummy_cell_6t
Xbit_r211_c0 bl_0 br_0 wl_211 vdd gnd dummy_cell_6t
Xbit_r212_c0 bl_0 br_0 wl_212 vdd gnd dummy_cell_6t
Xbit_r213_c0 bl_0 br_0 wl_213 vdd gnd dummy_cell_6t
Xbit_r214_c0 bl_0 br_0 wl_214 vdd gnd dummy_cell_6t
Xbit_r215_c0 bl_0 br_0 wl_215 vdd gnd dummy_cell_6t
Xbit_r216_c0 bl_0 br_0 wl_216 vdd gnd dummy_cell_6t
Xbit_r217_c0 bl_0 br_0 wl_217 vdd gnd dummy_cell_6t
Xbit_r218_c0 bl_0 br_0 wl_218 vdd gnd dummy_cell_6t
Xbit_r219_c0 bl_0 br_0 wl_219 vdd gnd dummy_cell_6t
Xbit_r220_c0 bl_0 br_0 wl_220 vdd gnd dummy_cell_6t
Xbit_r221_c0 bl_0 br_0 wl_221 vdd gnd dummy_cell_6t
Xbit_r222_c0 bl_0 br_0 wl_222 vdd gnd dummy_cell_6t
Xbit_r223_c0 bl_0 br_0 wl_223 vdd gnd dummy_cell_6t
Xbit_r224_c0 bl_0 br_0 wl_224 vdd gnd dummy_cell_6t
Xbit_r225_c0 bl_0 br_0 wl_225 vdd gnd dummy_cell_6t
Xbit_r226_c0 bl_0 br_0 wl_226 vdd gnd dummy_cell_6t
Xbit_r227_c0 bl_0 br_0 wl_227 vdd gnd dummy_cell_6t
Xbit_r228_c0 bl_0 br_0 wl_228 vdd gnd dummy_cell_6t
Xbit_r229_c0 bl_0 br_0 wl_229 vdd gnd dummy_cell_6t
Xbit_r230_c0 bl_0 br_0 wl_230 vdd gnd dummy_cell_6t
Xbit_r231_c0 bl_0 br_0 wl_231 vdd gnd dummy_cell_6t
Xbit_r232_c0 bl_0 br_0 wl_232 vdd gnd dummy_cell_6t
Xbit_r233_c0 bl_0 br_0 wl_233 vdd gnd dummy_cell_6t
Xbit_r234_c0 bl_0 br_0 wl_234 vdd gnd dummy_cell_6t
Xbit_r235_c0 bl_0 br_0 wl_235 vdd gnd dummy_cell_6t
Xbit_r236_c0 bl_0 br_0 wl_236 vdd gnd dummy_cell_6t
Xbit_r237_c0 bl_0 br_0 wl_237 vdd gnd dummy_cell_6t
Xbit_r238_c0 bl_0 br_0 wl_238 vdd gnd dummy_cell_6t
Xbit_r239_c0 bl_0 br_0 wl_239 vdd gnd dummy_cell_6t
Xbit_r240_c0 bl_0 br_0 wl_240 vdd gnd dummy_cell_6t
Xbit_r241_c0 bl_0 br_0 wl_241 vdd gnd dummy_cell_6t
Xbit_r242_c0 bl_0 br_0 wl_242 vdd gnd dummy_cell_6t
Xbit_r243_c0 bl_0 br_0 wl_243 vdd gnd dummy_cell_6t
Xbit_r244_c0 bl_0 br_0 wl_244 vdd gnd dummy_cell_6t
Xbit_r245_c0 bl_0 br_0 wl_245 vdd gnd dummy_cell_6t
Xbit_r246_c0 bl_0 br_0 wl_246 vdd gnd dummy_cell_6t
Xbit_r247_c0 bl_0 br_0 wl_247 vdd gnd dummy_cell_6t
Xbit_r248_c0 bl_0 br_0 wl_248 vdd gnd dummy_cell_6t
Xbit_r249_c0 bl_0 br_0 wl_249 vdd gnd dummy_cell_6t
Xbit_r250_c0 bl_0 br_0 wl_250 vdd gnd dummy_cell_6t
Xbit_r251_c0 bl_0 br_0 wl_251 vdd gnd dummy_cell_6t
Xbit_r252_c0 bl_0 br_0 wl_252 vdd gnd dummy_cell_6t
Xbit_r253_c0 bl_0 br_0 wl_253 vdd gnd dummy_cell_6t
Xbit_r254_c0 bl_0 br_0 wl_254 vdd gnd dummy_cell_6t
Xbit_r255_c0 bl_0 br_0 wl_255 vdd gnd dummy_cell_6t
Xbit_r256_c0 bl_0 br_0 wl_256 vdd gnd dummy_cell_6t
Xbit_r257_c0 bl_0 br_0 wl_257 vdd gnd dummy_cell_6t
Xbit_r258_c0 bl_0 br_0 wl_258 vdd gnd dummy_cell_6t
.ENDS dummy_array_2

.SUBCKT replica_bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 rbl_wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: rbl_bl_0 
* OUTPUT: rbl_br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* INPUT : wl_131 
* INPUT : wl_132 
* INPUT : wl_133 
* INPUT : wl_134 
* INPUT : wl_135 
* INPUT : wl_136 
* INPUT : wl_137 
* INPUT : wl_138 
* INPUT : wl_139 
* INPUT : wl_140 
* INPUT : wl_141 
* INPUT : wl_142 
* INPUT : wl_143 
* INPUT : wl_144 
* INPUT : wl_145 
* INPUT : wl_146 
* INPUT : wl_147 
* INPUT : wl_148 
* INPUT : wl_149 
* INPUT : wl_150 
* INPUT : wl_151 
* INPUT : wl_152 
* INPUT : wl_153 
* INPUT : wl_154 
* INPUT : wl_155 
* INPUT : wl_156 
* INPUT : wl_157 
* INPUT : wl_158 
* INPUT : wl_159 
* INPUT : wl_160 
* INPUT : wl_161 
* INPUT : wl_162 
* INPUT : wl_163 
* INPUT : wl_164 
* INPUT : wl_165 
* INPUT : wl_166 
* INPUT : wl_167 
* INPUT : wl_168 
* INPUT : wl_169 
* INPUT : wl_170 
* INPUT : wl_171 
* INPUT : wl_172 
* INPUT : wl_173 
* INPUT : wl_174 
* INPUT : wl_175 
* INPUT : wl_176 
* INPUT : wl_177 
* INPUT : wl_178 
* INPUT : wl_179 
* INPUT : wl_180 
* INPUT : wl_181 
* INPUT : wl_182 
* INPUT : wl_183 
* INPUT : wl_184 
* INPUT : wl_185 
* INPUT : wl_186 
* INPUT : wl_187 
* INPUT : wl_188 
* INPUT : wl_189 
* INPUT : wl_190 
* INPUT : wl_191 
* INPUT : wl_192 
* INPUT : wl_193 
* INPUT : wl_194 
* INPUT : wl_195 
* INPUT : wl_196 
* INPUT : wl_197 
* INPUT : wl_198 
* INPUT : wl_199 
* INPUT : wl_200 
* INPUT : wl_201 
* INPUT : wl_202 
* INPUT : wl_203 
* INPUT : wl_204 
* INPUT : wl_205 
* INPUT : wl_206 
* INPUT : wl_207 
* INPUT : wl_208 
* INPUT : wl_209 
* INPUT : wl_210 
* INPUT : wl_211 
* INPUT : wl_212 
* INPUT : wl_213 
* INPUT : wl_214 
* INPUT : wl_215 
* INPUT : wl_216 
* INPUT : wl_217 
* INPUT : wl_218 
* INPUT : wl_219 
* INPUT : wl_220 
* INPUT : wl_221 
* INPUT : wl_222 
* INPUT : wl_223 
* INPUT : wl_224 
* INPUT : wl_225 
* INPUT : wl_226 
* INPUT : wl_227 
* INPUT : wl_228 
* INPUT : wl_229 
* INPUT : wl_230 
* INPUT : wl_231 
* INPUT : wl_232 
* INPUT : wl_233 
* INPUT : wl_234 
* INPUT : wl_235 
* INPUT : wl_236 
* INPUT : wl_237 
* INPUT : wl_238 
* INPUT : wl_239 
* INPUT : wl_240 
* INPUT : wl_241 
* INPUT : wl_242 
* INPUT : wl_243 
* INPUT : wl_244 
* INPUT : wl_245 
* INPUT : wl_246 
* INPUT : wl_247 
* INPUT : wl_248 
* INPUT : wl_249 
* INPUT : wl_250 
* INPUT : wl_251 
* INPUT : wl_252 
* INPUT : wl_253 
* INPUT : wl_254 
* INPUT : wl_255 
* INPUT : rbl_wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 256 cols: 256
Xbitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 vdd gnd bitcell_array_0
Xreplica_col_0 rbl_bl_0 rbl_br_0 dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 dummy_wl_top vdd gnd replica_column_0
Xdummy_row_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_wl_0 vdd gnd dummy_array_0
Xdummy_row_bot bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_bot vdd gnd dummy_array_0
Xdummy_row_top bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_top vdd gnd dummy_array_0
Xdummy_col_left dummy_bl_left dummy_br_left dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 dummy_wl_top vdd gnd dummy_array_1
Xdummy_col_right dummy_bl_right dummy_br_right dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 dummy_wl_top vdd gnd dummy_array_2
.ENDS replica_bitcell_array_0

.SUBCKT pinv_6 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_6

* ptx M{0} {1} pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_7 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_7

* ptx M{0} {1} nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* ptx M{0} {1} pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_8 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_8

.SUBCKT pinvbuf_0 A Zb Z vdd gnd
* INOUT : A 
* INOUT : Zb 
* INOUT : Z 
* INOUT : vdd 
* INOUT : gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_6
Xbuf_inv2 zb_int z_int vdd gnd pinv_7
Xbuf_inv3 z_int Zb vdd gnd pinv_8
Xbuf_inv4 zb_int Z vdd gnd pinv_8
.ENDS pinvbuf_0

.SUBCKT bank dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 dout0_33 dout0_34 dout0_35 dout0_36 dout0_37 dout0_38 dout0_39 dout0_40 dout0_41 dout0_42 dout0_43 dout0_44 dout0_45 dout0_46 dout0_47 dout0_48 dout0_49 dout0_50 dout0_51 dout0_52 dout0_53 dout0_54 dout0_55 dout0_56 dout0_57 dout0_58 dout0_59 dout0_60 dout0_61 dout0_62 dout0_63 dout0_64 dout0_65 dout0_66 dout0_67 dout0_68 dout0_69 dout0_70 dout0_71 dout0_72 dout0_73 dout0_74 dout0_75 dout0_76 dout0_77 dout0_78 dout0_79 dout0_80 dout0_81 dout0_82 dout0_83 dout0_84 dout0_85 dout0_86 dout0_87 dout0_88 dout0_89 dout0_90 dout0_91 dout0_92 dout0_93 dout0_94 dout0_95 dout0_96 dout0_97 dout0_98 dout0_99 dout0_100 dout0_101 dout0_102 dout0_103 dout0_104 dout0_105 dout0_106 dout0_107 dout0_108 dout0_109 dout0_110 dout0_111 dout0_112 dout0_113 dout0_114 dout0_115 dout0_116 dout0_117 dout0_118 dout0_119 dout0_120 dout0_121 dout0_122 dout0_123 dout0_124 dout0_125 dout0_126 dout0_127 rbl_bl_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 din0_33 din0_34 din0_35 din0_36 din0_37 din0_38 din0_39 din0_40 din0_41 din0_42 din0_43 din0_44 din0_45 din0_46 din0_47 din0_48 din0_49 din0_50 din0_51 din0_52 din0_53 din0_54 din0_55 din0_56 din0_57 din0_58 din0_59 din0_60 din0_61 din0_62 din0_63 din0_64 din0_65 din0_66 din0_67 din0_68 din0_69 din0_70 din0_71 din0_72 din0_73 din0_74 din0_75 din0_76 din0_77 din0_78 din0_79 din0_80 din0_81 din0_82 din0_83 din0_84 din0_85 din0_86 din0_87 din0_88 din0_89 din0_90 din0_91 din0_92 din0_93 din0_94 din0_95 din0_96 din0_97 din0_98 din0_99 din0_100 din0_101 din0_102 din0_103 din0_104 din0_105 din0_106 din0_107 din0_108 din0_109 din0_110 din0_111 din0_112 din0_113 din0_114 din0_115 din0_116 din0_117 din0_118 din0_119 din0_120 din0_121 din0_122 din0_123 din0_124 din0_125 din0_126 din0_127 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: dout0_32 
* OUTPUT: dout0_33 
* OUTPUT: dout0_34 
* OUTPUT: dout0_35 
* OUTPUT: dout0_36 
* OUTPUT: dout0_37 
* OUTPUT: dout0_38 
* OUTPUT: dout0_39 
* OUTPUT: dout0_40 
* OUTPUT: dout0_41 
* OUTPUT: dout0_42 
* OUTPUT: dout0_43 
* OUTPUT: dout0_44 
* OUTPUT: dout0_45 
* OUTPUT: dout0_46 
* OUTPUT: dout0_47 
* OUTPUT: dout0_48 
* OUTPUT: dout0_49 
* OUTPUT: dout0_50 
* OUTPUT: dout0_51 
* OUTPUT: dout0_52 
* OUTPUT: dout0_53 
* OUTPUT: dout0_54 
* OUTPUT: dout0_55 
* OUTPUT: dout0_56 
* OUTPUT: dout0_57 
* OUTPUT: dout0_58 
* OUTPUT: dout0_59 
* OUTPUT: dout0_60 
* OUTPUT: dout0_61 
* OUTPUT: dout0_62 
* OUTPUT: dout0_63 
* OUTPUT: dout0_64 
* OUTPUT: dout0_65 
* OUTPUT: dout0_66 
* OUTPUT: dout0_67 
* OUTPUT: dout0_68 
* OUTPUT: dout0_69 
* OUTPUT: dout0_70 
* OUTPUT: dout0_71 
* OUTPUT: dout0_72 
* OUTPUT: dout0_73 
* OUTPUT: dout0_74 
* OUTPUT: dout0_75 
* OUTPUT: dout0_76 
* OUTPUT: dout0_77 
* OUTPUT: dout0_78 
* OUTPUT: dout0_79 
* OUTPUT: dout0_80 
* OUTPUT: dout0_81 
* OUTPUT: dout0_82 
* OUTPUT: dout0_83 
* OUTPUT: dout0_84 
* OUTPUT: dout0_85 
* OUTPUT: dout0_86 
* OUTPUT: dout0_87 
* OUTPUT: dout0_88 
* OUTPUT: dout0_89 
* OUTPUT: dout0_90 
* OUTPUT: dout0_91 
* OUTPUT: dout0_92 
* OUTPUT: dout0_93 
* OUTPUT: dout0_94 
* OUTPUT: dout0_95 
* OUTPUT: dout0_96 
* OUTPUT: dout0_97 
* OUTPUT: dout0_98 
* OUTPUT: dout0_99 
* OUTPUT: dout0_100 
* OUTPUT: dout0_101 
* OUTPUT: dout0_102 
* OUTPUT: dout0_103 
* OUTPUT: dout0_104 
* OUTPUT: dout0_105 
* OUTPUT: dout0_106 
* OUTPUT: dout0_107 
* OUTPUT: dout0_108 
* OUTPUT: dout0_109 
* OUTPUT: dout0_110 
* OUTPUT: dout0_111 
* OUTPUT: dout0_112 
* OUTPUT: dout0_113 
* OUTPUT: dout0_114 
* OUTPUT: dout0_115 
* OUTPUT: dout0_116 
* OUTPUT: dout0_117 
* OUTPUT: dout0_118 
* OUTPUT: dout0_119 
* OUTPUT: dout0_120 
* OUTPUT: dout0_121 
* OUTPUT: dout0_122 
* OUTPUT: dout0_123 
* OUTPUT: dout0_124 
* OUTPUT: dout0_125 
* OUTPUT: dout0_126 
* OUTPUT: dout0_127 
* OUTPUT: rbl_bl_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : din0_32 
* INPUT : din0_33 
* INPUT : din0_34 
* INPUT : din0_35 
* INPUT : din0_36 
* INPUT : din0_37 
* INPUT : din0_38 
* INPUT : din0_39 
* INPUT : din0_40 
* INPUT : din0_41 
* INPUT : din0_42 
* INPUT : din0_43 
* INPUT : din0_44 
* INPUT : din0_45 
* INPUT : din0_46 
* INPUT : din0_47 
* INPUT : din0_48 
* INPUT : din0_49 
* INPUT : din0_50 
* INPUT : din0_51 
* INPUT : din0_52 
* INPUT : din0_53 
* INPUT : din0_54 
* INPUT : din0_55 
* INPUT : din0_56 
* INPUT : din0_57 
* INPUT : din0_58 
* INPUT : din0_59 
* INPUT : din0_60 
* INPUT : din0_61 
* INPUT : din0_62 
* INPUT : din0_63 
* INPUT : din0_64 
* INPUT : din0_65 
* INPUT : din0_66 
* INPUT : din0_67 
* INPUT : din0_68 
* INPUT : din0_69 
* INPUT : din0_70 
* INPUT : din0_71 
* INPUT : din0_72 
* INPUT : din0_73 
* INPUT : din0_74 
* INPUT : din0_75 
* INPUT : din0_76 
* INPUT : din0_77 
* INPUT : din0_78 
* INPUT : din0_79 
* INPUT : din0_80 
* INPUT : din0_81 
* INPUT : din0_82 
* INPUT : din0_83 
* INPUT : din0_84 
* INPUT : din0_85 
* INPUT : din0_86 
* INPUT : din0_87 
* INPUT : din0_88 
* INPUT : din0_89 
* INPUT : din0_90 
* INPUT : din0_91 
* INPUT : din0_92 
* INPUT : din0_93 
* INPUT : din0_94 
* INPUT : din0_95 
* INPUT : din0_96 
* INPUT : din0_97 
* INPUT : din0_98 
* INPUT : din0_99 
* INPUT : din0_100 
* INPUT : din0_101 
* INPUT : din0_102 
* INPUT : din0_103 
* INPUT : din0_104 
* INPUT : din0_105 
* INPUT : din0_106 
* INPUT : din0_107 
* INPUT : din0_108 
* INPUT : din0_109 
* INPUT : din0_110 
* INPUT : din0_111 
* INPUT : din0_112 
* INPUT : din0_113 
* INPUT : din0_114 
* INPUT : din0_115 
* INPUT : din0_116 
* INPUT : din0_117 
* INPUT : din0_118 
* INPUT : din0_119 
* INPUT : din0_120 
* INPUT : din0_121 
* INPUT : din0_122 
* INPUT : din0_123 
* INPUT : din0_124 
* INPUT : din0_125 
* INPUT : din0_126 
* INPUT : din0_127 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr0_8 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xreplica_bitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 wl_en0 vdd gnd replica_bitcell_array_0
Xport_data0 rbl_bl_0 rbl_br_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 dout0_32 dout0_33 dout0_34 dout0_35 dout0_36 dout0_37 dout0_38 dout0_39 dout0_40 dout0_41 dout0_42 dout0_43 dout0_44 dout0_45 dout0_46 dout0_47 dout0_48 dout0_49 dout0_50 dout0_51 dout0_52 dout0_53 dout0_54 dout0_55 dout0_56 dout0_57 dout0_58 dout0_59 dout0_60 dout0_61 dout0_62 dout0_63 dout0_64 dout0_65 dout0_66 dout0_67 dout0_68 dout0_69 dout0_70 dout0_71 dout0_72 dout0_73 dout0_74 dout0_75 dout0_76 dout0_77 dout0_78 dout0_79 dout0_80 dout0_81 dout0_82 dout0_83 dout0_84 dout0_85 dout0_86 dout0_87 dout0_88 dout0_89 dout0_90 dout0_91 dout0_92 dout0_93 dout0_94 dout0_95 dout0_96 dout0_97 dout0_98 dout0_99 dout0_100 dout0_101 dout0_102 dout0_103 dout0_104 dout0_105 dout0_106 dout0_107 dout0_108 dout0_109 dout0_110 dout0_111 dout0_112 dout0_113 dout0_114 dout0_115 dout0_116 dout0_117 dout0_118 dout0_119 dout0_120 dout0_121 dout0_122 dout0_123 dout0_124 dout0_125 dout0_126 dout0_127 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 din0_32 din0_33 din0_34 din0_35 din0_36 din0_37 din0_38 din0_39 din0_40 din0_41 din0_42 din0_43 din0_44 din0_45 din0_46 din0_47 din0_48 din0_49 din0_50 din0_51 din0_52 din0_53 din0_54 din0_55 din0_56 din0_57 din0_58 din0_59 din0_60 din0_61 din0_62 din0_63 din0_64 din0_65 din0_66 din0_67 din0_68 din0_69 din0_70 din0_71 din0_72 din0_73 din0_74 din0_75 din0_76 din0_77 din0_78 din0_79 din0_80 din0_81 din0_82 din0_83 din0_84 din0_85 din0_86 din0_87 din0_88 din0_89 din0_90 din0_91 din0_92 din0_93 din0_94 din0_95 din0_96 din0_97 din0_98 din0_99 din0_100 din0_101 din0_102 din0_103 din0_104 din0_105 din0_106 din0_107 din0_108 din0_109 din0_110 din0_111 din0_112 din0_113 din0_114 din0_115 din0_116 din0_117 din0_118 din0_119 din0_120 din0_121 din0_122 din0_123 din0_124 din0_125 din0_126 din0_127 sel0_0 sel0_1 s_en0 p_en_bar0 w_en0 vdd gnd port_data_0
Xport_address0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 wl_en0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 wl_131 wl_132 wl_133 wl_134 wl_135 wl_136 wl_137 wl_138 wl_139 wl_140 wl_141 wl_142 wl_143 wl_144 wl_145 wl_146 wl_147 wl_148 wl_149 wl_150 wl_151 wl_152 wl_153 wl_154 wl_155 wl_156 wl_157 wl_158 wl_159 wl_160 wl_161 wl_162 wl_163 wl_164 wl_165 wl_166 wl_167 wl_168 wl_169 wl_170 wl_171 wl_172 wl_173 wl_174 wl_175 wl_176 wl_177 wl_178 wl_179 wl_180 wl_181 wl_182 wl_183 wl_184 wl_185 wl_186 wl_187 wl_188 wl_189 wl_190 wl_191 wl_192 wl_193 wl_194 wl_195 wl_196 wl_197 wl_198 wl_199 wl_200 wl_201 wl_202 wl_203 wl_204 wl_205 wl_206 wl_207 wl_208 wl_209 wl_210 wl_211 wl_212 wl_213 wl_214 wl_215 wl_216 wl_217 wl_218 wl_219 wl_220 wl_221 wl_222 wl_223 wl_224 wl_225 wl_226 wl_227 wl_228 wl_229 wl_230 wl_231 wl_232 wl_233 wl_234 wl_235 wl_236 wl_237 wl_238 wl_239 wl_240 wl_241 wl_242 wl_243 wl_244 wl_245 wl_246 wl_247 wl_248 wl_249 wl_250 wl_251 wl_252 wl_253 wl_254 wl_255 vdd gnd port_address_0
Xcol_address_decoder0 addr0_0 sel0_0 sel0_1 vdd gnd pinvbuf_0
.ENDS bank

.SUBCKT dff_buf_0 D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff D qint clk vdd gnd dff
Xdff_buf_inv1 qint Qb vdd gnd pinv_7
Xdff_buf_inv2 Qb Q vdd gnd pinv_8
.ENDS dff_buf_0

.SUBCKT dff_buf_array_0 din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
Xdff_r1_c0 din_1 dout_1 dout_bar_1 clk vdd gnd dff_buf_0
.ENDS dff_buf_array_0

.SUBCKT pnand2_1 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_1

.SUBCKT pdriver_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 4]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_6
Xbuf_inv3 Zb2_int Z vdd gnd pinv_8
.ENDS pdriver_1

.SUBCKT pand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_1
Xpand2_inv zb_int Z vdd gnd pdriver_1
.ENDS pand2_0

* ptx M{0} {1} nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p

.SUBCKT pinv_9 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p
.ENDS pinv_9

* ptx M{0} {1} nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT pinv_10 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_10

.SUBCKT pbuf_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_9
Xbuf_inv2 zb_int Z vdd gnd pinv_10
.ENDS pbuf_0

* ptx M{0} {1} nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_11 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_11

* ptx M{0} {1} nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_12 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_12

* ptx M{0} {1} nmos_vtg m=9 w=0.26u l=0.05u pd=0.62u ps=0.62u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=9 w=0.78u l=0.05u pd=1.66u ps=1.66u as=0.10p ad=0.10p

.SUBCKT pinv_13 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.78u l=0.05u pd=1.66u ps=1.66u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.26u l=0.05u pd=0.62u ps=0.62u as=0.03p ad=0.03p
.ENDS pinv_13

* ptx M{0} {1} nmos_vtg m=25 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=25 w=0.8425u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p

.SUBCKT pinv_14 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=25 w=0.8425u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=25 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS pinv_14

* ptx M{0} {1} nmos_vtg m=75 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=75 w=0.845u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p

.SUBCKT pinv_15 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=75 w=0.845u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=75 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_15

.SUBCKT pdriver_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 1, 1, 3, 9, 26, 78, 235]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_6
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_6
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_6
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_6
Xbuf_inv6 Zb5_int Zb6_int vdd gnd pinv_11
Xbuf_inv7 Zb6_int Zb7_int vdd gnd pinv_12
Xbuf_inv8 Zb7_int Zb8_int vdd gnd pinv_13
Xbuf_inv9 Zb8_int Zb9_int vdd gnd pinv_14
Xbuf_inv10 Zb9_int Z vdd gnd pinv_15
.ENDS pdriver_2

* ptx M{0} {1} nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p

.SUBCKT pinv_16 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS pinv_16

* ptx M{0} {1} nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p

.SUBCKT pinv_17 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_17

.SUBCKT pdriver_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_6
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_6
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_11
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_12
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_16
Xbuf_inv6 Zb5_int Z vdd gnd pinv_17
.ENDS pdriver_3

.SUBCKT pnand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_1

* ptx M{0} {1} nmos_vtg m=43 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=43 w=0.855u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT pinv_18 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=43 w=0.855u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=43 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_18

.SUBCKT pand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_18
.ENDS pand3_0

* ptx M{0} {1} nmos_vtg m=41 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=41 w=0.8425u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p

.SUBCKT pinv_19 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=41 w=0.8425u l=0.05u pd=1.79u ps=1.79u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=41 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS pinv_19

.SUBCKT pand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_19
.ENDS pand3_1

.SUBCKT pinv_20 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_20

.SUBCKT delay_chain_0 in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0 in dout_1 vdd gnd pinv_20
Xdload_0_0 dout_1 n_0_0 vdd gnd pinv_20
Xdload_0_1 dout_1 n_0_1 vdd gnd pinv_20
Xdload_0_2 dout_1 n_0_2 vdd gnd pinv_20
Xdload_0_3 dout_1 n_0_3 vdd gnd pinv_20
Xdinv1 dout_1 dout_2 vdd gnd pinv_20
Xdload_1_0 dout_2 n_1_0 vdd gnd pinv_20
Xdload_1_1 dout_2 n_1_1 vdd gnd pinv_20
Xdload_1_2 dout_2 n_1_2 vdd gnd pinv_20
Xdload_1_3 dout_2 n_1_3 vdd gnd pinv_20
Xdinv2 dout_2 dout_3 vdd gnd pinv_20
Xdload_2_0 dout_3 n_2_0 vdd gnd pinv_20
Xdload_2_1 dout_3 n_2_1 vdd gnd pinv_20
Xdload_2_2 dout_3 n_2_2 vdd gnd pinv_20
Xdload_2_3 dout_3 n_2_3 vdd gnd pinv_20
Xdinv3 dout_3 dout_4 vdd gnd pinv_20
Xdload_3_0 dout_4 n_3_0 vdd gnd pinv_20
Xdload_3_1 dout_4 n_3_1 vdd gnd pinv_20
Xdload_3_2 dout_4 n_3_2 vdd gnd pinv_20
Xdload_3_3 dout_4 n_3_3 vdd gnd pinv_20
Xdinv4 dout_4 dout_5 vdd gnd pinv_20
Xdload_4_0 dout_5 n_4_0 vdd gnd pinv_20
Xdload_4_1 dout_5 n_4_1 vdd gnd pinv_20
Xdload_4_2 dout_5 n_4_2 vdd gnd pinv_20
Xdload_4_3 dout_5 n_4_3 vdd gnd pinv_20
Xdinv5 dout_5 dout_6 vdd gnd pinv_20
Xdload_5_0 dout_6 n_5_0 vdd gnd pinv_20
Xdload_5_1 dout_6 n_5_1 vdd gnd pinv_20
Xdload_5_2 dout_6 n_5_2 vdd gnd pinv_20
Xdload_5_3 dout_6 n_5_3 vdd gnd pinv_20
Xdinv6 dout_6 dout_7 vdd gnd pinv_20
Xdload_6_0 dout_7 n_6_0 vdd gnd pinv_20
Xdload_6_1 dout_7 n_6_1 vdd gnd pinv_20
Xdload_6_2 dout_7 n_6_2 vdd gnd pinv_20
Xdload_6_3 dout_7 n_6_3 vdd gnd pinv_20
Xdinv7 dout_7 dout_8 vdd gnd pinv_20
Xdload_7_0 dout_8 n_7_0 vdd gnd pinv_20
Xdload_7_1 dout_8 n_7_1 vdd gnd pinv_20
Xdload_7_2 dout_8 n_7_2 vdd gnd pinv_20
Xdload_7_3 dout_8 n_7_3 vdd gnd pinv_20
Xdinv8 dout_8 out vdd gnd pinv_20
Xdload_8_0 out n_8_0 vdd gnd pinv_20
Xdload_8_1 out n_8_1 vdd gnd pinv_20
Xdload_8_2 out n_8_2 vdd gnd pinv_20
Xdload_8_3 out n_8_3 vdd gnd pinv_20
.ENDS delay_chain_0

.SUBCKT control_logic_rw csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 128
Xctrl_dffs csb web cs_bar cs we_bar we clk_buf vdd gnd dff_buf_array_0
Xclkbuf clk clk_buf vdd gnd pdriver_2
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_6
Xand2_gated_clk_bar cs clk_bar gated_clk_bar vdd gnd pand2_0
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_0
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_3
Xrbl_bl_delay_inv rbl_bl_delay rbl_bl_delay_bar vdd gnd pinv_6
Xw_en_and we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd pand3_0
Xbuf_s_en_and rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd pand3_1
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain_0
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_3
.ENDS control_logic_rw

.SUBCKT sram_512_128 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36] din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43] din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50] din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57] din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64] din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71] din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78] din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85] din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92] din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99] din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106] din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113] din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120] din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] csb0 web0 clk0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35] dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41] dout0[42] dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62] dout0[63] dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69] dout0[70] dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76] dout0[77] dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83] dout0[84] dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90] dout0[91] dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97] dout0[98] dout0[99] dout0[100] dout0[101] dout0[102] dout0[103] dout0[104] dout0[105] dout0[106] dout0[107] dout0[108] dout0[109] dout0[110] dout0[111] dout0[112] dout0[113] dout0[114] dout0[115] dout0[116] dout0[117] dout0[118] dout0[119] dout0[120] dout0[121] dout0[122] dout0[123] dout0[124] dout0[125] dout0[126] dout0[127] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : din0[32] 
* INPUT : din0[33] 
* INPUT : din0[34] 
* INPUT : din0[35] 
* INPUT : din0[36] 
* INPUT : din0[37] 
* INPUT : din0[38] 
* INPUT : din0[39] 
* INPUT : din0[40] 
* INPUT : din0[41] 
* INPUT : din0[42] 
* INPUT : din0[43] 
* INPUT : din0[44] 
* INPUT : din0[45] 
* INPUT : din0[46] 
* INPUT : din0[47] 
* INPUT : din0[48] 
* INPUT : din0[49] 
* INPUT : din0[50] 
* INPUT : din0[51] 
* INPUT : din0[52] 
* INPUT : din0[53] 
* INPUT : din0[54] 
* INPUT : din0[55] 
* INPUT : din0[56] 
* INPUT : din0[57] 
* INPUT : din0[58] 
* INPUT : din0[59] 
* INPUT : din0[60] 
* INPUT : din0[61] 
* INPUT : din0[62] 
* INPUT : din0[63] 
* INPUT : din0[64] 
* INPUT : din0[65] 
* INPUT : din0[66] 
* INPUT : din0[67] 
* INPUT : din0[68] 
* INPUT : din0[69] 
* INPUT : din0[70] 
* INPUT : din0[71] 
* INPUT : din0[72] 
* INPUT : din0[73] 
* INPUT : din0[74] 
* INPUT : din0[75] 
* INPUT : din0[76] 
* INPUT : din0[77] 
* INPUT : din0[78] 
* INPUT : din0[79] 
* INPUT : din0[80] 
* INPUT : din0[81] 
* INPUT : din0[82] 
* INPUT : din0[83] 
* INPUT : din0[84] 
* INPUT : din0[85] 
* INPUT : din0[86] 
* INPUT : din0[87] 
* INPUT : din0[88] 
* INPUT : din0[89] 
* INPUT : din0[90] 
* INPUT : din0[91] 
* INPUT : din0[92] 
* INPUT : din0[93] 
* INPUT : din0[94] 
* INPUT : din0[95] 
* INPUT : din0[96] 
* INPUT : din0[97] 
* INPUT : din0[98] 
* INPUT : din0[99] 
* INPUT : din0[100] 
* INPUT : din0[101] 
* INPUT : din0[102] 
* INPUT : din0[103] 
* INPUT : din0[104] 
* INPUT : din0[105] 
* INPUT : din0[106] 
* INPUT : din0[107] 
* INPUT : din0[108] 
* INPUT : din0[109] 
* INPUT : din0[110] 
* INPUT : din0[111] 
* INPUT : din0[112] 
* INPUT : din0[113] 
* INPUT : din0[114] 
* INPUT : din0[115] 
* INPUT : din0[116] 
* INPUT : din0[117] 
* INPUT : din0[118] 
* INPUT : din0[119] 
* INPUT : din0[120] 
* INPUT : din0[121] 
* INPUT : din0[122] 
* INPUT : din0[123] 
* INPUT : din0[124] 
* INPUT : din0[125] 
* INPUT : din0[126] 
* INPUT : din0[127] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr0[8] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* OUTPUT: dout0[32] 
* OUTPUT: dout0[33] 
* OUTPUT: dout0[34] 
* OUTPUT: dout0[35] 
* OUTPUT: dout0[36] 
* OUTPUT: dout0[37] 
* OUTPUT: dout0[38] 
* OUTPUT: dout0[39] 
* OUTPUT: dout0[40] 
* OUTPUT: dout0[41] 
* OUTPUT: dout0[42] 
* OUTPUT: dout0[43] 
* OUTPUT: dout0[44] 
* OUTPUT: dout0[45] 
* OUTPUT: dout0[46] 
* OUTPUT: dout0[47] 
* OUTPUT: dout0[48] 
* OUTPUT: dout0[49] 
* OUTPUT: dout0[50] 
* OUTPUT: dout0[51] 
* OUTPUT: dout0[52] 
* OUTPUT: dout0[53] 
* OUTPUT: dout0[54] 
* OUTPUT: dout0[55] 
* OUTPUT: dout0[56] 
* OUTPUT: dout0[57] 
* OUTPUT: dout0[58] 
* OUTPUT: dout0[59] 
* OUTPUT: dout0[60] 
* OUTPUT: dout0[61] 
* OUTPUT: dout0[62] 
* OUTPUT: dout0[63] 
* OUTPUT: dout0[64] 
* OUTPUT: dout0[65] 
* OUTPUT: dout0[66] 
* OUTPUT: dout0[67] 
* OUTPUT: dout0[68] 
* OUTPUT: dout0[69] 
* OUTPUT: dout0[70] 
* OUTPUT: dout0[71] 
* OUTPUT: dout0[72] 
* OUTPUT: dout0[73] 
* OUTPUT: dout0[74] 
* OUTPUT: dout0[75] 
* OUTPUT: dout0[76] 
* OUTPUT: dout0[77] 
* OUTPUT: dout0[78] 
* OUTPUT: dout0[79] 
* OUTPUT: dout0[80] 
* OUTPUT: dout0[81] 
* OUTPUT: dout0[82] 
* OUTPUT: dout0[83] 
* OUTPUT: dout0[84] 
* OUTPUT: dout0[85] 
* OUTPUT: dout0[86] 
* OUTPUT: dout0[87] 
* OUTPUT: dout0[88] 
* OUTPUT: dout0[89] 
* OUTPUT: dout0[90] 
* OUTPUT: dout0[91] 
* OUTPUT: dout0[92] 
* OUTPUT: dout0[93] 
* OUTPUT: dout0[94] 
* OUTPUT: dout0[95] 
* OUTPUT: dout0[96] 
* OUTPUT: dout0[97] 
* OUTPUT: dout0[98] 
* OUTPUT: dout0[99] 
* OUTPUT: dout0[100] 
* OUTPUT: dout0[101] 
* OUTPUT: dout0[102] 
* OUTPUT: dout0[103] 
* OUTPUT: dout0[104] 
* OUTPUT: dout0[105] 
* OUTPUT: dout0[106] 
* OUTPUT: dout0[107] 
* OUTPUT: dout0[108] 
* OUTPUT: dout0[109] 
* OUTPUT: dout0[110] 
* OUTPUT: dout0[111] 
* OUTPUT: dout0[112] 
* OUTPUT: dout0[113] 
* OUTPUT: dout0[114] 
* OUTPUT: dout0[115] 
* OUTPUT: dout0[116] 
* OUTPUT: dout0[117] 
* OUTPUT: dout0[118] 
* OUTPUT: dout0[119] 
* OUTPUT: dout0[120] 
* OUTPUT: dout0[121] 
* OUTPUT: dout0[122] 
* OUTPUT: dout0[123] 
* OUTPUT: dout0[124] 
* OUTPUT: dout0[125] 
* OUTPUT: dout0[126] 
* OUTPUT: dout0[127] 
* POWER : vdd 
* GROUND: gnd 
Xbank0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35] dout0[36] dout0[37] dout0[38] dout0[39] dout0[40] dout0[41] dout0[42] dout0[43] dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[50] dout0[51] dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59] dout0[60] dout0[61] dout0[62] dout0[63] dout0[64] dout0[65] dout0[66] dout0[67] dout0[68] dout0[69] dout0[70] dout0[71] dout0[72] dout0[73] dout0[74] dout0[75] dout0[76] dout0[77] dout0[78] dout0[79] dout0[80] dout0[81] dout0[82] dout0[83] dout0[84] dout0[85] dout0[86] dout0[87] dout0[88] dout0[89] dout0[90] dout0[91] dout0[92] dout0[93] dout0[94] dout0[95] dout0[96] dout0[97] dout0[98] dout0[99] dout0[100] dout0[101] dout0[102] dout0[103] dout0[104] dout0[105] dout0[106] dout0[107] dout0[108] dout0[109] dout0[110] dout0[111] dout0[112] dout0[113] dout0[114] dout0[115] dout0[116] dout0[117] dout0[118] dout0[119] dout0[120] dout0[121] dout0[122] dout0[123] dout0[124] dout0[125] dout0[126] dout0[127] rbl_bl0 bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] bank_din0[32] bank_din0[33] bank_din0[34] bank_din0[35] bank_din0[36] bank_din0[37] bank_din0[38] bank_din0[39] bank_din0[40] bank_din0[41] bank_din0[42] bank_din0[43] bank_din0[44] bank_din0[45] bank_din0[46] bank_din0[47] bank_din0[48] bank_din0[49] bank_din0[50] bank_din0[51] bank_din0[52] bank_din0[53] bank_din0[54] bank_din0[55] bank_din0[56] bank_din0[57] bank_din0[58] bank_din0[59] bank_din0[60] bank_din0[61] bank_din0[62] bank_din0[63] bank_din0[64] bank_din0[65] bank_din0[66] bank_din0[67] bank_din0[68] bank_din0[69] bank_din0[70] bank_din0[71] bank_din0[72] bank_din0[73] bank_din0[74] bank_din0[75] bank_din0[76] bank_din0[77] bank_din0[78] bank_din0[79] bank_din0[80] bank_din0[81] bank_din0[82] bank_din0[83] bank_din0[84] bank_din0[85] bank_din0[86] bank_din0[87] bank_din0[88] bank_din0[89] bank_din0[90] bank_din0[91] bank_din0[92] bank_din0[93] bank_din0[94] bank_din0[95] bank_din0[96] bank_din0[97] bank_din0[98] bank_din0[99] bank_din0[100] bank_din0[101] bank_din0[102] bank_din0[103] bank_din0[104] bank_din0[105] bank_din0[106] bank_din0[107] bank_din0[108] bank_din0[109] bank_din0[110] bank_din0[111] bank_din0[112] bank_din0[113] bank_din0[114] bank_din0[115] bank_din0[116] bank_din0[117] bank_din0[118] bank_din0[119] bank_din0[120] bank_din0[121] bank_din0[122] bank_din0[123] bank_din0[124] bank_din0[125] bank_din0[126] bank_din0[127] a0[0] a0[1] a0[2] a0[3] a0[4] a0[5] a0[6] a0[7] a0[8] s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd bank
Xcontrol0 csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd control_logic_rw
Xrow_address0 addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] a0[1] a0[2] a0[3] a0[4] a0[5] a0[6] a0[7] a0[8] clk_buf0 vdd gnd row_addr_dff
Xcol_address0 addr0[0] a0[0] clk_buf0 vdd gnd col_addr_dff
Xdata_dff0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] din0[32] din0[33] din0[34] din0[35] din0[36] din0[37] din0[38] din0[39] din0[40] din0[41] din0[42] din0[43] din0[44] din0[45] din0[46] din0[47] din0[48] din0[49] din0[50] din0[51] din0[52] din0[53] din0[54] din0[55] din0[56] din0[57] din0[58] din0[59] din0[60] din0[61] din0[62] din0[63] din0[64] din0[65] din0[66] din0[67] din0[68] din0[69] din0[70] din0[71] din0[72] din0[73] din0[74] din0[75] din0[76] din0[77] din0[78] din0[79] din0[80] din0[81] din0[82] din0[83] din0[84] din0[85] din0[86] din0[87] din0[88] din0[89] din0[90] din0[91] din0[92] din0[93] din0[94] din0[95] din0[96] din0[97] din0[98] din0[99] din0[100] din0[101] din0[102] din0[103] din0[104] din0[105] din0[106] din0[107] din0[108] din0[109] din0[110] din0[111] din0[112] din0[113] din0[114] din0[115] din0[116] din0[117] din0[118] din0[119] din0[120] din0[121] din0[122] din0[123] din0[124] din0[125] din0[126] din0[127] bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] bank_din0[32] bank_din0[33] bank_din0[34] bank_din0[35] bank_din0[36] bank_din0[37] bank_din0[38] bank_din0[39] bank_din0[40] bank_din0[41] bank_din0[42] bank_din0[43] bank_din0[44] bank_din0[45] bank_din0[46] bank_din0[47] bank_din0[48] bank_din0[49] bank_din0[50] bank_din0[51] bank_din0[52] bank_din0[53] bank_din0[54] bank_din0[55] bank_din0[56] bank_din0[57] bank_din0[58] bank_din0[59] bank_din0[60] bank_din0[61] bank_din0[62] bank_din0[63] bank_din0[64] bank_din0[65] bank_din0[66] bank_din0[67] bank_din0[68] bank_din0[69] bank_din0[70] bank_din0[71] bank_din0[72] bank_din0[73] bank_din0[74] bank_din0[75] bank_din0[76] bank_din0[77] bank_din0[78] bank_din0[79] bank_din0[80] bank_din0[81] bank_din0[82] bank_din0[83] bank_din0[84] bank_din0[85] bank_din0[86] bank_din0[87] bank_din0[88] bank_din0[89] bank_din0[90] bank_din0[91] bank_din0[92] bank_din0[93] bank_din0[94] bank_din0[95] bank_din0[96] bank_din0[97] bank_din0[98] bank_din0[99] bank_din0[100] bank_din0[101] bank_din0[102] bank_din0[103] bank_din0[104] bank_din0[105] bank_din0[106] bank_din0[107] bank_din0[108] bank_din0[109] bank_din0[110] bank_din0[111] bank_din0[112] bank_din0[113] bank_din0[114] bank_din0[115] bank_din0[116] bank_din0[117] bank_din0[118] bank_din0[119] bank_din0[120] bank_din0[121] bank_din0[122] bank_din0[123] bank_din0[124] bank_din0[125] bank_din0[126] bank_din0[127] clk_buf0 vdd gnd data_dff
.ENDS sram_512_128
